magic
tech sky130B
magscale 1 2
timestamp 1736855682
<< nwell >>
rect 42475 25064 42762 25065
rect 43622 25064 43857 25065
rect 39993 25010 40233 25011
rect 39990 24777 40233 25010
rect 39990 24595 40234 24777
rect 42472 24667 42762 25064
rect 43449 24671 43931 25064
rect 48988 25061 49275 25062
rect 50135 25061 50370 25062
rect 46506 25007 46746 25008
rect 39552 24271 40744 24595
rect 41877 24200 42762 24667
rect 41877 24147 42763 24200
rect 43019 24147 43931 24671
rect 46503 24774 46746 25007
rect 46503 24592 46747 24774
rect 48985 24664 49275 25061
rect 49962 24668 50444 25061
rect 62080 25060 62367 25061
rect 63227 25060 63462 25061
rect 55522 25056 55809 25057
rect 56669 25056 56904 25057
rect 53040 25002 53280 25003
rect 46065 24268 47257 24592
rect 41877 24143 42764 24147
rect 42306 23858 42764 24143
rect 43449 23888 43931 24147
rect 48390 24197 49275 24664
rect 48390 24144 49276 24197
rect 49532 24144 50444 24668
rect 53037 24769 53280 25002
rect 53037 24587 53281 24769
rect 55519 24659 55809 25056
rect 56496 24663 56978 25056
rect 59598 25006 59838 25007
rect 52599 24263 53791 24587
rect 48390 24140 49277 24144
rect 42306 23560 42790 23858
rect 43448 23564 43932 23888
rect 48819 23855 49277 24140
rect 49962 23885 50444 24144
rect 54924 24192 55809 24659
rect 54924 24139 55810 24192
rect 56066 24139 56978 24663
rect 59595 24773 59838 25006
rect 59595 24591 59839 24773
rect 62077 24663 62367 25060
rect 63054 24667 63536 25060
rect 59157 24267 60349 24591
rect 61482 24196 62367 24663
rect 61482 24143 62368 24196
rect 62624 24143 63536 24667
rect 61482 24139 62369 24143
rect 54924 24135 55811 24139
rect 48819 23557 49303 23855
rect 49961 23561 50445 23885
rect 55353 23850 55811 24135
rect 56496 23880 56978 24139
rect 55353 23552 55837 23850
rect 56495 23556 56979 23880
rect 61911 23854 62369 24139
rect 63054 23884 63536 24143
rect 61911 23556 62395 23854
rect 63053 23560 63537 23884
rect 40007 23360 40247 23361
rect 40004 23127 40247 23360
rect 46520 23357 46760 23358
rect 40004 22945 40248 23127
rect 46517 23124 46760 23357
rect 59612 23356 59852 23357
rect 53054 23352 53294 23353
rect 39566 22621 40758 22945
rect 43718 22528 43946 23018
rect 46517 22942 46761 23124
rect 53051 23119 53294 23352
rect 59609 23123 59852 23356
rect 46079 22618 47271 22942
rect 3438 22058 5215 22348
rect 6582 22058 8359 22348
rect 3437 21858 5215 22058
rect 6581 21858 8359 22058
rect 9714 22054 11491 22344
rect 12858 22054 14635 22344
rect 16060 22058 17837 22348
rect 19204 22058 20981 22348
rect 2964 21534 5656 21858
rect 6108 21534 8800 21858
rect 9713 21854 11491 22054
rect 12857 21854 14635 22054
rect 16059 21858 17837 22058
rect 19203 21858 20981 22058
rect 22336 22054 24113 22344
rect 25480 22054 27257 22344
rect 9240 21530 11932 21854
rect 12384 21530 15076 21854
rect 15586 21534 18278 21858
rect 18730 21534 21422 21858
rect 22335 21854 24113 22054
rect 25479 21854 27257 22054
rect 41029 22328 42352 22528
rect 43412 22328 44250 22528
rect 50231 22525 50459 23015
rect 53051 22937 53295 23119
rect 52613 22613 53805 22937
rect 41029 22004 44733 22328
rect 47542 22325 48865 22525
rect 49925 22325 50763 22525
rect 56765 22520 56993 23010
rect 59609 22941 59853 23123
rect 59171 22617 60363 22941
rect 63323 22524 63551 23014
rect 21862 21530 24554 21854
rect 25006 21530 27698 21854
rect 40002 21756 40242 21757
rect 39999 21523 40242 21756
rect 39999 21341 40243 21523
rect 39561 21017 40753 21341
rect 41457 21311 42295 22004
rect 43355 21311 44193 22004
rect 47542 22001 51246 22325
rect 54076 22320 55399 22520
rect 56459 22320 57297 22520
rect 60634 22324 61957 22524
rect 63017 22324 63855 22524
rect 46515 21753 46755 21754
rect 46512 21520 46755 21753
rect 46512 21338 46756 21520
rect 46074 21014 47266 21338
rect 47970 21308 48808 22001
rect 49868 21308 50706 22001
rect 54076 21996 57780 22320
rect 60634 22000 64338 22324
rect 53049 21748 53289 21749
rect 53046 21515 53289 21748
rect 53046 21333 53290 21515
rect 52608 21009 53800 21333
rect 54504 21303 55342 21996
rect 56402 21303 57240 21996
rect 59607 21752 59847 21753
rect 59604 21519 59847 21752
rect 59604 21337 59848 21519
rect 59166 21013 60358 21337
rect 61062 21307 61900 22000
rect 62960 21307 63798 22000
rect 70651 21668 70975 22109
rect 70161 19891 70975 21668
rect 70451 19890 70975 19891
rect 59168 19460 59403 19461
rect 60263 19460 60550 19461
rect 52655 19457 52890 19458
rect 53750 19457 54037 19458
rect 39563 19456 39798 19457
rect 40658 19456 40945 19457
rect 39489 19063 39971 19456
rect 39489 18539 40401 19063
rect 40658 19059 40948 19456
rect 46121 19452 46356 19453
rect 47216 19452 47503 19453
rect 43187 19402 43427 19403
rect 43187 19169 43430 19402
rect 40658 18592 41543 19059
rect 43186 18987 43430 19169
rect 46047 19059 46529 19452
rect 42676 18663 43868 18987
rect 40657 18539 41543 18592
rect 39489 18280 39971 18539
rect 40656 18535 41543 18539
rect 46047 18535 46959 19059
rect 47216 19055 47506 19452
rect 49745 19398 49985 19399
rect 49745 19165 49988 19398
rect 47216 18588 48101 19055
rect 49744 18983 49988 19165
rect 52581 19064 53063 19457
rect 49234 18659 50426 18983
rect 47215 18535 48101 18588
rect 39488 17956 39972 18280
rect 40656 18250 41114 18535
rect 46047 18276 46529 18535
rect 47214 18531 48101 18535
rect 52581 18540 53493 19064
rect 53750 19060 54040 19457
rect 56279 19403 56519 19404
rect 56279 19170 56522 19403
rect 53750 18593 54635 19060
rect 56278 18988 56522 19170
rect 59094 19067 59576 19460
rect 55768 18664 56960 18988
rect 53749 18540 54635 18593
rect 40630 17952 41114 18250
rect 46046 17952 46530 18276
rect 47214 18246 47672 18531
rect 52581 18281 53063 18540
rect 53748 18536 54635 18540
rect 59094 18543 60006 19067
rect 60263 19063 60553 19460
rect 70651 19417 70975 19890
rect 62792 19406 63032 19407
rect 62792 19173 63035 19406
rect 60263 18596 61148 19063
rect 62791 18991 63035 19173
rect 62281 18667 63473 18991
rect 60262 18543 61148 18596
rect 47188 17948 47672 18246
rect 52580 17957 53064 18281
rect 53748 18251 54206 18536
rect 59094 18284 59576 18543
rect 60261 18539 61148 18543
rect 53722 17953 54206 18251
rect 59093 17960 59577 18284
rect 60261 18254 60719 18539
rect 70651 18524 70975 18965
rect 60235 17956 60719 18254
rect 62778 17756 63018 17757
rect 56265 17753 56505 17754
rect 43173 17752 43413 17753
rect 43173 17519 43416 17752
rect 4396 16346 5310 17126
rect 5564 16348 6478 17126
rect 4396 16082 4880 16346
rect 4396 16040 4881 16082
rect 5564 16081 6048 16348
rect 6732 16346 7646 17126
rect 7900 16348 8814 17126
rect 6732 16081 7216 16346
rect 7900 16082 8384 16348
rect 9074 16346 9988 17124
rect 5564 16040 6049 16081
rect 6732 16040 7217 16081
rect 7900 16040 8386 16082
rect 4397 15758 4881 16040
rect 5565 15757 6049 16040
rect 6733 15757 7217 16040
rect 7902 15758 8386 16040
rect 9074 15762 9558 16346
rect 10242 16344 11156 17124
rect 11410 16346 12324 17124
rect 12578 16346 13492 17124
rect 13756 16675 14948 16921
rect 15204 16675 16396 16921
rect 13755 16663 14948 16675
rect 15203 16663 16396 16675
rect 16702 16673 17894 16919
rect 18150 16673 19342 16919
rect 19670 16675 20862 16921
rect 21118 16675 22310 16921
rect 39474 16920 39702 17410
rect 43172 17337 43416 17519
rect 49731 17748 49971 17749
rect 49731 17515 49974 17748
rect 56265 17520 56508 17753
rect 62778 17523 63021 17756
rect 42662 17013 43854 17337
rect 13755 16351 14947 16663
rect 15203 16351 16395 16663
rect 16701 16661 17894 16673
rect 18149 16661 19342 16673
rect 19669 16663 20862 16675
rect 21117 16663 22310 16675
rect 22616 16673 23808 16919
rect 24064 16673 25256 16919
rect 39170 16720 40008 16920
rect 41068 16720 42391 16920
rect 46032 16916 46260 17406
rect 49730 17333 49974 17515
rect 49220 17009 50412 17333
rect 52566 16921 52794 17411
rect 56264 17338 56508 17520
rect 55754 17014 56946 17338
rect 59079 16924 59307 17414
rect 62777 17341 63021 17523
rect 62267 17017 63459 17341
rect 16701 16349 17893 16661
rect 18149 16349 19341 16661
rect 19669 16351 20861 16663
rect 21117 16351 22309 16663
rect 22615 16661 23808 16673
rect 24063 16661 25256 16673
rect 22615 16349 23807 16661
rect 24063 16349 25255 16661
rect 38687 16396 42391 16720
rect 45728 16716 46566 16916
rect 47626 16716 48949 16916
rect 52262 16721 53100 16921
rect 54160 16721 55483 16921
rect 58775 16724 59613 16924
rect 60673 16724 61996 16924
rect 70161 16747 70975 18524
rect 70451 16746 70975 16747
rect 10242 16086 10726 16344
rect 11410 16086 11894 16346
rect 10242 16038 10727 16086
rect 11410 16038 11895 16086
rect 10243 15762 10727 16038
rect 11411 15762 11895 16038
rect 12578 15756 13062 16346
rect 39227 15703 40065 16396
rect 41125 15703 41963 16396
rect 45245 16392 48949 16716
rect 51779 16397 55483 16721
rect 58292 16400 61996 16724
rect 43178 16148 43418 16149
rect 43178 15915 43421 16148
rect 43177 15733 43421 15915
rect 42667 15409 43859 15733
rect 45785 15699 46623 16392
rect 47683 15699 48521 16392
rect 49736 16144 49976 16145
rect 49736 15911 49979 16144
rect 49735 15729 49979 15911
rect 49225 15405 50417 15729
rect 52319 15704 53157 16397
rect 54217 15704 55055 16397
rect 56270 16149 56510 16150
rect 56270 15916 56513 16149
rect 56269 15734 56513 15916
rect 55759 15410 56951 15734
rect 58832 15707 59670 16400
rect 60730 15707 61568 16400
rect 70651 16273 70975 16746
rect 62783 16152 63023 16153
rect 62783 15919 63026 16152
rect 62782 15737 63026 15919
rect 62272 15413 63464 15737
rect 70647 15392 70971 15833
rect 936 14920 2713 15210
rect 4080 14920 5857 15210
rect 935 14720 2713 14920
rect 4079 14720 5857 14920
rect 7212 14916 8989 15206
rect 10356 14916 12133 15206
rect 13558 14920 15335 15210
rect 16702 14920 18479 15210
rect 462 14396 3154 14720
rect 3606 14396 6298 14720
rect 7211 14716 8989 14916
rect 10355 14716 12133 14916
rect 13557 14720 15335 14920
rect 16701 14720 18479 14920
rect 19834 14916 21611 15206
rect 22978 14916 24755 15206
rect 6738 14392 9430 14716
rect 9882 14392 12574 14716
rect 13084 14396 15776 14720
rect 16228 14396 18920 14720
rect 19833 14716 21611 14916
rect 22977 14716 24755 14916
rect 19360 14392 22052 14716
rect 22504 14392 25196 14716
rect 70157 13615 70971 15392
rect 70447 13614 70971 13615
rect 30092 12789 30416 13216
rect 70647 13141 70971 13614
rect 30092 12735 31109 12789
rect 29797 12545 31109 12735
rect 936 12186 2713 12476
rect 4080 12186 5857 12476
rect 935 11986 2713 12186
rect 4079 11986 5857 12186
rect 7212 12182 8989 12472
rect 10356 12182 12133 12472
rect 13558 12186 15335 12476
rect 16702 12186 18479 12476
rect 462 11662 3154 11986
rect 3606 11662 6298 11986
rect 7211 11982 8989 12182
rect 10355 11982 12133 12182
rect 13557 11986 15335 12186
rect 16701 11986 18479 12186
rect 19834 12182 21611 12472
rect 22978 12182 24755 12472
rect 6738 11658 9430 11982
rect 9882 11658 12574 11982
rect 13084 11662 15776 11986
rect 16228 11662 18920 11986
rect 19833 11982 21611 12182
rect 22977 11982 24755 12182
rect 29605 12069 31109 12545
rect 41521 12211 42713 12457
rect 41521 12199 42714 12211
rect 19360 11658 22052 11982
rect 22504 11658 25196 11982
rect 29797 11951 31109 12069
rect 29797 11891 30416 11951
rect 30092 11411 30416 11891
rect 41522 11887 42714 12199
rect 48070 12210 49262 12456
rect 54724 12231 55916 12477
rect 54724 12219 55917 12231
rect 48070 12198 49263 12210
rect 48071 11886 49263 12198
rect 54725 11907 55917 12219
rect 63377 12064 64569 12310
rect 63377 12052 64570 12064
rect 63378 11740 64570 12052
rect 65832 11902 66329 12359
rect 70647 12248 70971 12689
rect 65186 11656 68170 11902
rect 65186 11335 68171 11656
rect 30090 10721 30414 11148
rect 30090 10667 31107 10721
rect 29795 10477 31107 10667
rect 65613 10642 66451 11335
rect 66979 11332 68171 11335
rect 47220 10601 47507 10602
rect 48367 10601 48602 10602
rect 60499 10601 60786 10602
rect 61646 10601 61881 10602
rect 29605 10001 31107 10477
rect 34857 10311 36049 10557
rect 44738 10547 44978 10548
rect 40671 10513 40958 10514
rect 41818 10513 42053 10514
rect 38189 10459 38429 10460
rect 34857 10299 36050 10311
rect 29795 9883 31107 10001
rect 34858 9987 36050 10299
rect 38186 10226 38429 10459
rect 38186 10044 38430 10226
rect 40668 10116 40958 10513
rect 41645 10120 42127 10513
rect 44735 10314 44978 10547
rect 44735 10132 44979 10314
rect 47217 10204 47507 10601
rect 48194 10208 48676 10601
rect 58017 10547 58257 10548
rect 53874 10533 54161 10534
rect 55021 10533 55256 10534
rect 51392 10479 51632 10480
rect 29795 9823 30414 9883
rect 946 9454 2723 9744
rect 4090 9454 5867 9744
rect 945 9254 2723 9454
rect 4089 9254 5867 9454
rect 7222 9450 8999 9740
rect 10366 9450 12143 9740
rect 13568 9454 15345 9744
rect 16712 9454 18489 9744
rect 472 8930 3164 9254
rect 3616 8930 6308 9254
rect 7221 9250 8999 9450
rect 10365 9250 12143 9450
rect 13567 9254 15345 9454
rect 16711 9254 18489 9454
rect 19844 9450 21621 9740
rect 22988 9450 24765 9740
rect 6748 8926 9440 9250
rect 9892 8926 12584 9250
rect 13094 8930 15786 9254
rect 16238 8930 18930 9254
rect 19843 9250 21621 9450
rect 22987 9250 24765 9450
rect 30090 9343 30414 9823
rect 37748 9720 38940 10044
rect 40073 9649 40958 10116
rect 40073 9596 40959 9649
rect 41215 9596 42127 10120
rect 44297 9808 45489 10132
rect 46622 9737 47507 10204
rect 46622 9684 47508 9737
rect 47764 9684 48676 10208
rect 51389 10246 51632 10479
rect 51389 10064 51633 10246
rect 53871 10136 54161 10533
rect 54848 10140 55330 10533
rect 50951 9740 52143 10064
rect 46622 9680 47509 9684
rect 40073 9592 40960 9596
rect 40502 9307 40960 9592
rect 41645 9337 42127 9596
rect 47051 9395 47509 9680
rect 48194 9425 48676 9684
rect 53276 9669 54161 10136
rect 53276 9616 54162 9669
rect 54418 9616 55330 10140
rect 58014 10314 58257 10547
rect 58014 10132 58258 10314
rect 60496 10204 60786 10601
rect 61473 10208 61955 10601
rect 70157 10471 70971 12248
rect 70447 10470 70971 10471
rect 57576 9808 58768 10132
rect 59901 9737 60786 10204
rect 59901 9684 60787 9737
rect 61043 9684 61955 10208
rect 70647 9997 70971 10470
rect 59901 9680 60788 9684
rect 53276 9612 54163 9616
rect 19370 8926 22062 9250
rect 22514 8926 25206 9250
rect 30092 8652 30416 9079
rect 40502 9009 40986 9307
rect 41644 9013 42128 9337
rect 47051 9097 47535 9395
rect 48193 9101 48677 9425
rect 53705 9327 54163 9612
rect 54848 9357 55330 9616
rect 60330 9395 60788 9680
rect 61473 9425 61955 9684
rect 63372 9493 64564 9739
rect 63372 9481 64565 9493
rect 53705 9029 54189 9327
rect 54847 9033 55331 9357
rect 60330 9097 60814 9395
rect 61472 9101 61956 9425
rect 63373 9169 64565 9481
rect 70651 9046 70975 9487
rect 44752 8897 44992 8898
rect 58031 8897 58271 8898
rect 38203 8809 38443 8810
rect 30092 8598 31109 8652
rect 29797 8408 31109 8598
rect 29605 7932 31109 8408
rect 38200 8576 38443 8809
rect 44749 8664 44992 8897
rect 51406 8829 51646 8830
rect 38200 8394 38444 8576
rect 44749 8482 44993 8664
rect 51403 8596 51646 8829
rect 58028 8664 58271 8897
rect 37762 8070 38954 8394
rect 41914 7977 42142 8467
rect 44311 8158 45503 8482
rect 48463 8065 48691 8555
rect 51403 8414 51647 8596
rect 50965 8090 52157 8414
rect 29797 7814 31109 7932
rect 29797 7754 30416 7814
rect 30092 7274 30416 7754
rect 34849 7726 36041 7972
rect 39225 7777 40548 7977
rect 41608 7777 42446 7977
rect 45774 7865 47097 8065
rect 48157 7865 48995 8065
rect 55117 7997 55345 8487
rect 58028 8482 58272 8664
rect 57590 8158 58782 8482
rect 61742 8065 61970 8555
rect 34849 7714 36042 7726
rect 34850 7402 36042 7714
rect 39225 7453 42929 7777
rect 45774 7541 49478 7865
rect 52428 7797 53751 7997
rect 54811 7797 55649 7997
rect 59053 7865 60376 8065
rect 61436 7865 62274 8065
rect 38198 7205 38438 7206
rect 3081 6295 3565 6847
rect 3819 6295 4303 6847
rect 4557 6295 5041 6847
rect 5295 6295 5779 6847
rect 6035 6295 6519 6847
rect 6777 6297 7261 6847
rect 7515 6301 7999 6847
rect 8253 6297 8737 6849
rect 9843 6604 10319 6794
rect 9665 6309 10509 6604
rect 11911 6602 12387 6794
rect 13980 6604 14456 6794
rect 9185 5985 10990 6309
rect 11733 6307 12577 6602
rect 13802 6309 14646 6604
rect 16048 6602 16524 6794
rect 18117 6602 18593 6792
rect 9725 5292 10563 5985
rect 11253 5983 13058 6307
rect 13322 5985 15127 6309
rect 15870 6307 16714 6602
rect 17939 6307 18783 6602
rect 20185 6600 20661 6792
rect 22254 6602 22730 6792
rect 11793 5290 12631 5983
rect 13862 5292 14700 5985
rect 15390 5983 17195 6307
rect 17459 5983 19264 6307
rect 20007 6305 20851 6600
rect 22076 6307 22920 6602
rect 24322 6600 24798 6792
rect 15930 5290 16768 5983
rect 17999 5290 18837 5983
rect 19527 5981 21332 6305
rect 21596 5983 23401 6307
rect 24144 6305 24988 6600
rect 30090 6584 30414 7011
rect 38195 6972 38438 7205
rect 38195 6790 38439 6972
rect 30090 6530 31107 6584
rect 29795 6340 31107 6530
rect 37757 6466 38949 6790
rect 39653 6760 40491 7453
rect 41551 6760 42389 7453
rect 44747 7293 44987 7294
rect 44744 7060 44987 7293
rect 44744 6878 44988 7060
rect 44306 6554 45498 6878
rect 46202 6848 47040 7541
rect 48100 6848 48938 7541
rect 52428 7473 56132 7797
rect 59053 7541 62757 7865
rect 65834 7811 66331 8268
rect 65188 7565 68172 7811
rect 51401 7225 51641 7226
rect 51398 6992 51641 7225
rect 51398 6810 51642 6992
rect 50960 6486 52152 6810
rect 52856 6780 53694 7473
rect 54754 6780 55592 7473
rect 58026 7293 58266 7294
rect 58023 7060 58266 7293
rect 58023 6878 58267 7060
rect 57585 6554 58777 6878
rect 59481 6848 60319 7541
rect 61379 6848 62217 7541
rect 65188 7244 68173 7565
rect 70161 7269 70975 9046
rect 70451 7268 70975 7269
rect 63372 6460 64564 6706
rect 65615 6551 66453 7244
rect 66981 7241 68173 7244
rect 70651 6795 70975 7268
rect 63372 6448 64565 6460
rect 20067 5288 20905 5981
rect 22136 5290 22974 5983
rect 23664 5981 25469 6305
rect 24204 5288 25042 5981
rect 29605 5864 31107 6340
rect 63373 6136 64565 6448
rect 70651 5902 70975 6343
rect 29795 5746 31107 5864
rect 29795 5686 30414 5746
rect 30090 5206 30414 5686
rect 30090 4515 30414 4942
rect 40663 4733 40950 4734
rect 41810 4733 42045 4734
rect 60491 4733 60778 4734
rect 61638 4733 61873 4734
rect 30090 4461 31107 4515
rect 29795 4271 31107 4461
rect 34830 4448 36022 4694
rect 38181 4679 38421 4680
rect 34830 4436 36023 4448
rect 29603 3795 31107 4271
rect 34831 4124 36023 4436
rect 38178 4446 38421 4679
rect 38178 4264 38422 4446
rect 40660 4336 40950 4733
rect 41637 4340 42119 4733
rect 53869 4732 54156 4733
rect 55016 4732 55251 4733
rect 47214 4731 47501 4732
rect 48361 4731 48596 4732
rect 44732 4677 44972 4678
rect 37740 3940 38932 4264
rect 40065 3869 40950 4336
rect 40065 3816 40951 3869
rect 41207 3816 42119 4340
rect 44729 4444 44972 4677
rect 44729 4262 44973 4444
rect 47211 4334 47501 4731
rect 48188 4338 48670 4731
rect 51387 4678 51627 4679
rect 44291 3938 45483 4262
rect 40065 3812 40952 3816
rect 29795 3677 31107 3795
rect 29795 3617 30414 3677
rect 30090 3137 30414 3617
rect 40494 3527 40952 3812
rect 41637 3557 42119 3816
rect 46616 3867 47501 4334
rect 46616 3814 47502 3867
rect 47758 3814 48670 4338
rect 51384 4445 51627 4678
rect 51384 4263 51628 4445
rect 53866 4335 54156 4732
rect 54843 4339 55325 4732
rect 58009 4679 58249 4680
rect 50946 3939 52138 4263
rect 46616 3810 47503 3814
rect 40494 3229 40978 3527
rect 41636 3233 42120 3557
rect 47045 3525 47503 3810
rect 48188 3555 48670 3814
rect 53271 3868 54156 4335
rect 53271 3815 54157 3868
rect 54413 3815 55325 4339
rect 58006 4446 58249 4679
rect 58006 4264 58250 4446
rect 60488 4336 60778 4733
rect 61465 4340 61947 4733
rect 63443 4540 64635 4786
rect 63443 4528 64636 4540
rect 57568 3940 58760 4264
rect 53271 3811 54158 3815
rect 47045 3227 47529 3525
rect 48187 3231 48671 3555
rect 53700 3526 54158 3811
rect 54843 3556 55325 3815
rect 59893 3869 60778 4336
rect 59893 3816 60779 3869
rect 61035 3816 61947 4340
rect 63444 4216 64636 4528
rect 65834 4316 66331 4773
rect 59893 3812 60780 3816
rect 53700 3228 54184 3526
rect 54842 3232 55326 3556
rect 60322 3527 60780 3812
rect 61465 3557 61947 3816
rect 65188 4070 68172 4316
rect 70161 4125 70975 5902
rect 70451 4124 70975 4125
rect 65188 3749 68173 4070
rect 60322 3229 60806 3527
rect 61464 3233 61948 3557
rect 65615 3056 66453 3749
rect 66981 3746 68173 3749
rect 70651 3651 70975 4124
rect 38195 3029 38435 3030
rect 58023 3029 58263 3030
rect 653 2202 2430 2492
rect 3797 2202 5574 2492
rect 6929 2206 8706 2496
rect 10073 2206 11850 2496
rect 653 2002 2431 2202
rect 3797 2002 5575 2202
rect 6929 2006 8707 2206
rect 10073 2006 11851 2206
rect 13275 2202 15052 2492
rect 16419 2202 18196 2492
rect 19551 2206 21328 2496
rect 22695 2206 24472 2496
rect 30088 2447 30412 2874
rect 38192 2796 38435 3029
rect 51401 3028 51641 3029
rect 44746 3027 44986 3028
rect 38192 2614 38436 2796
rect 44743 2794 44986 3027
rect 51398 2795 51641 3028
rect 58020 2796 58263 3029
rect 30088 2393 31105 2447
rect 212 1678 2904 2002
rect 3356 1678 6048 2002
rect 6488 1682 9180 2006
rect 9632 1682 12324 2006
rect 13275 2002 15053 2202
rect 16419 2002 18197 2202
rect 19551 2006 21329 2206
rect 22695 2006 24473 2206
rect 29793 2203 31105 2393
rect 37754 2290 38946 2614
rect 12834 1678 15526 2002
rect 15978 1678 18670 2002
rect 19110 1682 21802 2006
rect 22254 1682 24946 2006
rect 29603 1727 31105 2203
rect 41906 2197 42134 2687
rect 44743 2612 44987 2794
rect 44305 2288 45497 2612
rect 39217 1997 40540 2197
rect 41600 1997 42438 2197
rect 48457 2195 48685 2685
rect 51398 2613 51642 2795
rect 50960 2289 52152 2613
rect 55112 2196 55340 2686
rect 58020 2614 58264 2796
rect 70647 2770 70971 3211
rect 57582 2290 58774 2614
rect 61734 2197 61962 2687
rect 29793 1609 31105 1727
rect 34846 1688 36038 1934
rect 34846 1676 36039 1688
rect 29793 1549 30412 1609
rect 30088 1069 30412 1549
rect 34847 1364 36039 1676
rect 39217 1673 42921 1997
rect 45768 1995 47091 2195
rect 48151 1995 48989 2195
rect 52423 1996 53746 2196
rect 54806 1996 55644 2196
rect 59045 1997 60368 2197
rect 61428 1997 62266 2197
rect 38190 1425 38430 1426
rect 38187 1192 38430 1425
rect 38187 1010 38431 1192
rect 30090 378 30414 805
rect 37749 686 38941 1010
rect 39645 980 40483 1673
rect 41543 980 42381 1673
rect 45768 1671 49472 1995
rect 52423 1672 56127 1996
rect 59045 1673 62749 1997
rect 44741 1423 44981 1424
rect 44738 1190 44981 1423
rect 44738 1008 44982 1190
rect 44300 684 45492 1008
rect 46196 978 47034 1671
rect 48094 978 48932 1671
rect 51396 1424 51636 1425
rect 51393 1191 51636 1424
rect 51393 1009 51637 1191
rect 50955 685 52147 1009
rect 52851 979 53689 1672
rect 54749 979 55587 1672
rect 58018 1425 58258 1426
rect 58015 1192 58258 1425
rect 58015 1010 58259 1192
rect 57577 686 58769 1010
rect 59473 980 60311 1673
rect 61371 980 62209 1673
rect 63440 1470 64632 1716
rect 63440 1458 64633 1470
rect 63441 1146 64633 1458
rect 70157 993 70971 2770
rect 70447 992 70971 993
rect 70647 519 70971 992
rect 30090 324 31107 378
rect 29795 134 31107 324
rect 29603 -342 31107 134
rect 65834 -32 66331 425
rect 29795 -460 31107 -342
rect 65188 -278 68172 -32
rect 29795 -520 30414 -460
rect 30090 -1000 30414 -520
rect 65188 -599 68173 -278
rect 70647 -374 70971 67
rect 685 -1690 2462 -1400
rect 3829 -1690 5606 -1400
rect 6961 -1686 8738 -1396
rect 10105 -1686 11882 -1396
rect 685 -1890 2463 -1690
rect 3829 -1890 5607 -1690
rect 6961 -1886 8739 -1686
rect 10105 -1886 11883 -1686
rect 13307 -1690 15084 -1400
rect 16451 -1690 18228 -1400
rect 19583 -1686 21360 -1396
rect 22727 -1686 24504 -1396
rect 244 -2214 2936 -1890
rect 3388 -2214 6080 -1890
rect 6520 -2210 9212 -1886
rect 9664 -2210 12356 -1886
rect 13307 -1890 15085 -1690
rect 16451 -1890 18229 -1690
rect 19583 -1886 21361 -1686
rect 22727 -1886 24505 -1686
rect 30088 -1690 30412 -1263
rect 63447 -1375 64639 -1129
rect 65615 -1292 66453 -599
rect 66981 -602 68173 -599
rect 63447 -1387 64640 -1375
rect 30088 -1744 31105 -1690
rect 12866 -2214 15558 -1890
rect 16010 -2214 18702 -1890
rect 19142 -2210 21834 -1886
rect 22286 -2210 24978 -1886
rect 29793 -1934 31105 -1744
rect 41557 -1805 42749 -1493
rect 48111 -1800 49303 -1488
rect 29603 -2410 31105 -1934
rect 41556 -1817 42749 -1805
rect 48110 -1812 49303 -1800
rect 54760 -1812 55952 -1500
rect 63448 -1699 64640 -1387
rect 41556 -2063 42748 -1817
rect 48110 -2058 49302 -1812
rect 54759 -1824 55952 -1812
rect 54759 -2070 55951 -1824
rect 70157 -2151 70971 -374
rect 70447 -2152 70971 -2151
rect 29793 -2528 31105 -2410
rect 29793 -2588 30412 -2528
rect 30088 -3068 30412 -2588
rect 70647 -2625 70971 -2152
<< nmos >>
rect 39883 23696 39943 24096
rect 40001 23696 40061 24096
rect 40236 23896 40296 24096
rect 41881 23622 41941 23822
rect 41999 23622 42059 23822
rect 42117 23622 42177 23822
rect 43023 23626 43083 23826
rect 43141 23626 43201 23826
rect 43259 23626 43319 23826
rect 46396 23693 46456 24093
rect 46514 23693 46574 24093
rect 46749 23893 46809 24093
rect 48394 23619 48454 23819
rect 48512 23619 48572 23819
rect 48630 23619 48690 23819
rect 49536 23623 49596 23823
rect 49654 23623 49714 23823
rect 49772 23623 49832 23823
rect 52930 23688 52990 24088
rect 53048 23688 53108 24088
rect 53283 23888 53343 24088
rect 54928 23614 54988 23814
rect 55046 23614 55106 23814
rect 55164 23614 55224 23814
rect 56070 23618 56130 23818
rect 56188 23618 56248 23818
rect 56306 23618 56366 23818
rect 59488 23692 59548 24092
rect 59606 23692 59666 24092
rect 59841 23892 59901 24092
rect 61486 23618 61546 23818
rect 61604 23618 61664 23818
rect 61722 23618 61782 23818
rect 62628 23622 62688 23822
rect 62746 23622 62806 23822
rect 62864 23622 62924 23822
rect 39897 22046 39957 22446
rect 40015 22046 40075 22446
rect 40250 22246 40310 22446
rect 3926 20463 3986 20663
rect 4122 20263 4182 20663
rect 4240 20263 4300 20663
rect 4358 20263 4418 20663
rect 4476 20263 4536 20663
rect 4668 20463 4728 20663
rect 7070 20463 7130 20663
rect 7266 20263 7326 20663
rect 7384 20263 7444 20663
rect 7502 20263 7562 20663
rect 7620 20263 7680 20663
rect 7812 20463 7872 20663
rect 10202 20459 10262 20659
rect 10398 20259 10458 20659
rect 10516 20259 10576 20659
rect 10634 20259 10694 20659
rect 10752 20259 10812 20659
rect 10944 20459 11004 20659
rect 13346 20459 13406 20659
rect 13542 20259 13602 20659
rect 13660 20259 13720 20659
rect 13778 20259 13838 20659
rect 13896 20259 13956 20659
rect 14088 20459 14148 20659
rect 16548 20463 16608 20663
rect 16744 20263 16804 20663
rect 16862 20263 16922 20663
rect 16980 20263 17040 20663
rect 17098 20263 17158 20663
rect 17290 20463 17350 20663
rect 19692 20463 19752 20663
rect 19888 20263 19948 20663
rect 20006 20263 20066 20663
rect 20124 20263 20184 20663
rect 20242 20263 20302 20663
rect 20434 20463 20494 20663
rect 46410 22043 46470 22443
rect 46528 22043 46588 22443
rect 46763 22243 46823 22443
rect 22824 20459 22884 20659
rect 23020 20259 23080 20659
rect 23138 20259 23198 20659
rect 23256 20259 23316 20659
rect 23374 20259 23434 20659
rect 23566 20459 23626 20659
rect 25968 20459 26028 20659
rect 26164 20259 26224 20659
rect 26282 20259 26342 20659
rect 26400 20259 26460 20659
rect 26518 20259 26578 20659
rect 26710 20459 26770 20659
rect 39892 20442 39952 20842
rect 40010 20442 40070 20842
rect 40245 20642 40305 20842
rect 41249 20841 41309 21041
rect 41669 20641 41729 21041
rect 41787 20641 41847 21041
rect 41905 20641 41965 21041
rect 42023 20641 42083 21041
rect 42547 20841 42607 21041
rect 43147 20841 43207 21041
rect 43567 20641 43627 21041
rect 43685 20641 43745 21041
rect 43803 20641 43863 21041
rect 43921 20641 43981 21041
rect 44445 20841 44505 21041
rect 52944 22038 53004 22438
rect 53062 22038 53122 22438
rect 53297 22238 53357 22438
rect 46405 20439 46465 20839
rect 46523 20439 46583 20839
rect 46758 20639 46818 20839
rect 47762 20838 47822 21038
rect 48182 20638 48242 21038
rect 48300 20638 48360 21038
rect 48418 20638 48478 21038
rect 48536 20638 48596 21038
rect 49060 20838 49120 21038
rect 49660 20838 49720 21038
rect 50080 20638 50140 21038
rect 50198 20638 50258 21038
rect 50316 20638 50376 21038
rect 50434 20638 50494 21038
rect 50958 20838 51018 21038
rect 59502 22042 59562 22442
rect 59620 22042 59680 22442
rect 59855 22242 59915 22442
rect 52939 20434 52999 20834
rect 53057 20434 53117 20834
rect 53292 20634 53352 20834
rect 54296 20833 54356 21033
rect 54716 20633 54776 21033
rect 54834 20633 54894 21033
rect 54952 20633 55012 21033
rect 55070 20633 55130 21033
rect 55594 20833 55654 21033
rect 56194 20833 56254 21033
rect 56614 20633 56674 21033
rect 56732 20633 56792 21033
rect 56850 20633 56910 21033
rect 56968 20633 57028 21033
rect 57492 20833 57552 21033
rect 59497 20438 59557 20838
rect 59615 20438 59675 20838
rect 59850 20638 59910 20838
rect 60854 20837 60914 21037
rect 61274 20637 61334 21037
rect 61392 20637 61452 21037
rect 61510 20637 61570 21037
rect 61628 20637 61688 21037
rect 62152 20837 62212 21037
rect 62752 20837 62812 21037
rect 63172 20637 63232 21037
rect 63290 20637 63350 21037
rect 63408 20637 63468 21037
rect 63526 20637 63586 21037
rect 64050 20837 64110 21037
rect 71846 21121 72046 21181
rect 71846 20929 72246 20989
rect 71846 20811 72246 20871
rect 71846 20693 72246 20753
rect 71846 20575 72246 20635
rect 71846 20379 72046 20439
rect 40101 18018 40161 18218
rect 40219 18018 40279 18218
rect 40337 18018 40397 18218
rect 43124 18288 43184 18488
rect 41243 18014 41303 18214
rect 41361 18014 41421 18214
rect 41479 18014 41539 18214
rect 43359 18088 43419 18488
rect 43477 18088 43537 18488
rect 46659 18014 46719 18214
rect 46777 18014 46837 18214
rect 46895 18014 46955 18214
rect 49682 18284 49742 18484
rect 47801 18010 47861 18210
rect 47919 18010 47979 18210
rect 48037 18010 48097 18210
rect 49917 18084 49977 18484
rect 50035 18084 50095 18484
rect 53193 18019 53253 18219
rect 53311 18019 53371 18219
rect 53429 18019 53489 18219
rect 56216 18289 56276 18489
rect 54335 18015 54395 18215
rect 54453 18015 54513 18215
rect 54571 18015 54631 18215
rect 56451 18089 56511 18489
rect 56569 18089 56629 18489
rect 59706 18022 59766 18222
rect 59824 18022 59884 18222
rect 59942 18022 60002 18222
rect 62729 18292 62789 18492
rect 60848 18018 60908 18218
rect 60966 18018 61026 18218
rect 61084 18018 61144 18218
rect 62964 18092 63024 18492
rect 63082 18092 63142 18492
rect 71846 17977 72046 18037
rect 71846 17785 72246 17845
rect 71846 17667 72246 17727
rect 71846 17549 72246 17609
rect 71846 17431 72246 17491
rect 5010 15826 5070 16026
rect 5128 15826 5188 16026
rect 5246 15826 5306 16026
rect 6178 15826 6238 16026
rect 6296 15826 6356 16026
rect 6414 15826 6474 16026
rect 7346 15824 7406 16024
rect 7464 15824 7524 16024
rect 7582 15824 7642 16024
rect 8514 15824 8574 16024
rect 8632 15824 8692 16024
rect 8750 15824 8810 16024
rect 9688 15824 9748 16024
rect 9806 15824 9866 16024
rect 9924 15824 9984 16024
rect 10856 15824 10916 16024
rect 10974 15824 11034 16024
rect 11092 15824 11152 16024
rect 12024 15824 12084 16024
rect 12142 15824 12202 16024
rect 12260 15824 12320 16024
rect 13192 15822 13252 16022
rect 13310 15822 13370 16022
rect 13428 15822 13488 16022
rect 14203 15976 14263 16176
rect 14438 15776 14498 16176
rect 14556 15776 14616 16176
rect 15651 15976 15711 16176
rect 15886 15776 15946 16176
rect 16004 15776 16064 16176
rect 43110 16638 43170 16838
rect 17149 15974 17209 16174
rect 17384 15774 17444 16174
rect 17502 15774 17562 16174
rect 18597 15974 18657 16174
rect 18832 15774 18892 16174
rect 18950 15774 19010 16174
rect 20117 15976 20177 16176
rect 20352 15776 20412 16176
rect 20470 15776 20530 16176
rect 21565 15976 21625 16176
rect 21800 15776 21860 16176
rect 21918 15776 21978 16176
rect 23063 15974 23123 16174
rect 23298 15774 23358 16174
rect 23416 15774 23476 16174
rect 24511 15974 24571 16174
rect 24746 15774 24806 16174
rect 24864 15774 24924 16174
rect 43345 16438 43405 16838
rect 43463 16438 43523 16838
rect 49668 16634 49728 16834
rect 38915 15233 38975 15433
rect 39439 15033 39499 15433
rect 39557 15033 39617 15433
rect 39675 15033 39735 15433
rect 39793 15033 39853 15433
rect 40213 15233 40273 15433
rect 40813 15233 40873 15433
rect 41337 15033 41397 15433
rect 41455 15033 41515 15433
rect 41573 15033 41633 15433
rect 41691 15033 41751 15433
rect 42111 15233 42171 15433
rect 49903 16434 49963 16834
rect 50021 16434 50081 16834
rect 56202 16639 56262 16839
rect 43115 15034 43175 15234
rect 1424 13325 1484 13525
rect 1620 13125 1680 13525
rect 1738 13125 1798 13525
rect 1856 13125 1916 13525
rect 1974 13125 2034 13525
rect 2166 13325 2226 13525
rect 4568 13325 4628 13525
rect 4764 13125 4824 13525
rect 4882 13125 4942 13525
rect 5000 13125 5060 13525
rect 5118 13125 5178 13525
rect 5310 13325 5370 13525
rect 43350 14834 43410 15234
rect 43468 14834 43528 15234
rect 45473 15229 45533 15429
rect 45997 15029 46057 15429
rect 46115 15029 46175 15429
rect 46233 15029 46293 15429
rect 46351 15029 46411 15429
rect 46771 15229 46831 15429
rect 47371 15229 47431 15429
rect 47895 15029 47955 15429
rect 48013 15029 48073 15429
rect 48131 15029 48191 15429
rect 48249 15029 48309 15429
rect 48669 15229 48729 15429
rect 56437 16439 56497 16839
rect 56555 16439 56615 16839
rect 71846 17235 72046 17295
rect 62715 16642 62775 16842
rect 52007 15234 52067 15434
rect 49673 15030 49733 15230
rect 49908 14830 49968 15230
rect 50026 14830 50086 15230
rect 52531 15034 52591 15434
rect 52649 15034 52709 15434
rect 52767 15034 52827 15434
rect 52885 15034 52945 15434
rect 53305 15234 53365 15434
rect 53905 15234 53965 15434
rect 54429 15034 54489 15434
rect 54547 15034 54607 15434
rect 54665 15034 54725 15434
rect 54783 15034 54843 15434
rect 55203 15234 55263 15434
rect 62950 16442 63010 16842
rect 63068 16442 63128 16842
rect 58520 15237 58580 15437
rect 56207 15035 56267 15235
rect 56442 14835 56502 15235
rect 56560 14835 56620 15235
rect 59044 15037 59104 15437
rect 59162 15037 59222 15437
rect 59280 15037 59340 15437
rect 59398 15037 59458 15437
rect 59818 15237 59878 15437
rect 60418 15237 60478 15437
rect 60942 15037 61002 15437
rect 61060 15037 61120 15437
rect 61178 15037 61238 15437
rect 61296 15037 61356 15437
rect 61716 15237 61776 15437
rect 62720 15038 62780 15238
rect 62955 14838 63015 15238
rect 63073 14838 63133 15238
rect 71842 14845 72042 14905
rect 71842 14653 72242 14713
rect 7700 13321 7760 13521
rect 7896 13121 7956 13521
rect 8014 13121 8074 13521
rect 8132 13121 8192 13521
rect 8250 13121 8310 13521
rect 8442 13321 8502 13521
rect 10844 13321 10904 13521
rect 11040 13121 11100 13521
rect 11158 13121 11218 13521
rect 11276 13121 11336 13521
rect 11394 13121 11454 13521
rect 11586 13321 11646 13521
rect 14046 13325 14106 13525
rect 14242 13125 14302 13525
rect 14360 13125 14420 13525
rect 14478 13125 14538 13525
rect 14596 13125 14656 13525
rect 14788 13325 14848 13525
rect 17190 13325 17250 13525
rect 17386 13125 17446 13525
rect 17504 13125 17564 13525
rect 17622 13125 17682 13525
rect 17740 13125 17800 13525
rect 17932 13325 17992 13525
rect 71842 14535 72242 14595
rect 71842 14417 72242 14477
rect 71842 14299 72242 14359
rect 71842 14103 72042 14163
rect 20322 13321 20382 13521
rect 20518 13121 20578 13521
rect 20636 13121 20696 13521
rect 20754 13121 20814 13521
rect 20872 13121 20932 13521
rect 21064 13321 21124 13521
rect 23466 13321 23526 13521
rect 23662 13121 23722 13521
rect 23780 13121 23840 13521
rect 23898 13121 23958 13521
rect 24016 13121 24076 13521
rect 24208 13321 24268 13521
rect 31379 12937 31579 12997
rect 31379 12517 31779 12577
rect 31379 12399 31779 12459
rect 1424 10591 1484 10791
rect 1620 10391 1680 10791
rect 1738 10391 1798 10791
rect 1856 10391 1916 10791
rect 1974 10391 2034 10791
rect 2166 10591 2226 10791
rect 4568 10591 4628 10791
rect 4764 10391 4824 10791
rect 4882 10391 4942 10791
rect 5000 10391 5060 10791
rect 5118 10391 5178 10791
rect 5310 10591 5370 10791
rect 31379 12281 31779 12341
rect 31379 12163 31779 12223
rect 7700 10587 7760 10787
rect 7896 10387 7956 10787
rect 8014 10387 8074 10787
rect 8132 10387 8192 10787
rect 8250 10387 8310 10787
rect 8442 10587 8502 10787
rect 10844 10587 10904 10787
rect 11040 10387 11100 10787
rect 11158 10387 11218 10787
rect 11276 10387 11336 10787
rect 11394 10387 11454 10787
rect 11586 10587 11646 10787
rect 14046 10591 14106 10791
rect 14242 10391 14302 10791
rect 14360 10391 14420 10791
rect 14478 10391 14538 10791
rect 14596 10391 14656 10791
rect 14788 10591 14848 10791
rect 17190 10591 17250 10791
rect 17386 10391 17446 10791
rect 17504 10391 17564 10791
rect 17622 10391 17682 10791
rect 17740 10391 17800 10791
rect 17932 10591 17992 10791
rect 31379 11639 31579 11699
rect 41853 11312 41913 11712
rect 41971 11312 42031 11712
rect 42206 11512 42266 11712
rect 48402 11311 48462 11711
rect 48520 11311 48580 11711
rect 48755 11511 48815 11711
rect 55056 11332 55116 11732
rect 55174 11332 55234 11732
rect 55409 11532 55469 11732
rect 63709 11165 63769 11565
rect 63827 11165 63887 11565
rect 64062 11365 64122 11565
rect 71842 11701 72042 11761
rect 71842 11509 72242 11569
rect 31377 10869 31577 10929
rect 20322 10587 20382 10787
rect 20518 10387 20578 10787
rect 20636 10387 20696 10787
rect 20754 10387 20814 10787
rect 20872 10387 20932 10787
rect 21064 10587 21124 10787
rect 23466 10587 23526 10787
rect 23662 10387 23722 10787
rect 23780 10387 23840 10787
rect 23898 10387 23958 10787
rect 24016 10387 24076 10787
rect 24208 10587 24268 10787
rect 31377 10449 31777 10509
rect 31377 10331 31777 10391
rect 31377 10213 31777 10273
rect 31377 10095 31777 10155
rect 71842 11391 72242 11451
rect 71842 11273 72242 11333
rect 67310 10757 67370 11157
rect 67428 10757 67488 11157
rect 67663 10957 67723 11157
rect 71842 11155 72242 11215
rect 71842 10959 72042 11019
rect 31377 9571 31577 9631
rect 35189 9412 35249 9812
rect 35307 9412 35367 9812
rect 35542 9612 35602 9812
rect 1434 7859 1494 8059
rect 1630 7659 1690 8059
rect 1748 7659 1808 8059
rect 1866 7659 1926 8059
rect 1984 7659 2044 8059
rect 2176 7859 2236 8059
rect 4578 7859 4638 8059
rect 4774 7659 4834 8059
rect 4892 7659 4952 8059
rect 5010 7659 5070 8059
rect 5128 7659 5188 8059
rect 5320 7859 5380 8059
rect 38079 9145 38139 9545
rect 38197 9145 38257 9545
rect 38432 9345 38492 9545
rect 65405 10172 65465 10372
rect 40077 9071 40137 9271
rect 40195 9071 40255 9271
rect 40313 9071 40373 9271
rect 41219 9075 41279 9275
rect 41337 9075 41397 9275
rect 41455 9075 41515 9275
rect 44628 9233 44688 9633
rect 44746 9233 44806 9633
rect 44981 9433 45041 9633
rect 46626 9159 46686 9359
rect 46744 9159 46804 9359
rect 46862 9159 46922 9359
rect 47768 9163 47828 9363
rect 47886 9163 47946 9363
rect 48004 9163 48064 9363
rect 51282 9165 51342 9565
rect 51400 9165 51460 9565
rect 51635 9365 51695 9565
rect 65825 9972 65885 10372
rect 65943 9972 66003 10372
rect 66061 9972 66121 10372
rect 66179 9972 66239 10372
rect 66703 10172 66763 10372
rect 53280 9091 53340 9291
rect 53398 9091 53458 9291
rect 53516 9091 53576 9291
rect 54422 9095 54482 9295
rect 54540 9095 54600 9295
rect 54658 9095 54718 9295
rect 57907 9233 57967 9633
rect 58025 9233 58085 9633
rect 58260 9433 58320 9633
rect 59905 9159 59965 9359
rect 60023 9159 60083 9359
rect 60141 9159 60201 9359
rect 61047 9163 61107 9363
rect 61165 9163 61225 9363
rect 61283 9163 61343 9363
rect 7710 7855 7770 8055
rect 7906 7655 7966 8055
rect 8024 7655 8084 8055
rect 8142 7655 8202 8055
rect 8260 7655 8320 8055
rect 8452 7855 8512 8055
rect 10854 7855 10914 8055
rect 11050 7655 11110 8055
rect 11168 7655 11228 8055
rect 11286 7655 11346 8055
rect 11404 7655 11464 8055
rect 11596 7855 11656 8055
rect 14056 7859 14116 8059
rect 14252 7659 14312 8059
rect 14370 7659 14430 8059
rect 14488 7659 14548 8059
rect 14606 7659 14666 8059
rect 14798 7859 14858 8059
rect 17200 7859 17260 8059
rect 17396 7659 17456 8059
rect 17514 7659 17574 8059
rect 17632 7659 17692 8059
rect 17750 7659 17810 8059
rect 17942 7859 18002 8059
rect 31379 8800 31579 8860
rect 63704 8594 63764 8994
rect 63822 8594 63882 8994
rect 64057 8794 64117 8994
rect 31379 8380 31779 8440
rect 31379 8262 31779 8322
rect 20332 7855 20392 8055
rect 20528 7655 20588 8055
rect 20646 7655 20706 8055
rect 20764 7655 20824 8055
rect 20882 7655 20942 8055
rect 21074 7855 21134 8055
rect 23476 7855 23536 8055
rect 23672 7655 23732 8055
rect 23790 7655 23850 8055
rect 23908 7655 23968 8055
rect 24026 7655 24086 8055
rect 24218 7855 24278 8055
rect 31379 8144 31779 8204
rect 31379 8026 31779 8086
rect 71846 8499 72046 8559
rect 71846 8307 72246 8367
rect 31379 7502 31579 7562
rect 38093 7495 38153 7895
rect 38211 7495 38271 7895
rect 38446 7695 38506 7895
rect 44642 7583 44702 7983
rect 44760 7583 44820 7983
rect 44995 7783 45055 7983
rect 35181 6827 35241 7227
rect 35299 6827 35359 7227
rect 35534 7027 35594 7227
rect 31377 6732 31577 6792
rect 3293 5975 3353 6175
rect 4031 5975 4091 6175
rect 4769 5971 4829 6171
rect 5507 5971 5567 6171
rect 6247 5971 6307 6171
rect 6989 5971 7049 6171
rect 7727 5975 7787 6175
rect 8465 5973 8525 6173
rect 9413 4822 9473 5022
rect 9937 4622 9997 5022
rect 10055 4622 10115 5022
rect 10173 4622 10233 5022
rect 10291 4622 10351 5022
rect 10711 4822 10771 5022
rect 11481 4820 11541 5020
rect 12005 4620 12065 5020
rect 12123 4620 12183 5020
rect 12241 4620 12301 5020
rect 12359 4620 12419 5020
rect 12779 4820 12839 5020
rect 13550 4822 13610 5022
rect 14074 4622 14134 5022
rect 14192 4622 14252 5022
rect 14310 4622 14370 5022
rect 14428 4622 14488 5022
rect 14848 4822 14908 5022
rect 31377 6312 31777 6372
rect 71846 8189 72246 8249
rect 71846 8071 72246 8131
rect 31377 6194 31777 6254
rect 15618 4820 15678 5020
rect 16142 4620 16202 5020
rect 16260 4620 16320 5020
rect 16378 4620 16438 5020
rect 16496 4620 16556 5020
rect 16916 4820 16976 5020
rect 17687 4820 17747 5020
rect 18211 4620 18271 5020
rect 18329 4620 18389 5020
rect 18447 4620 18507 5020
rect 18565 4620 18625 5020
rect 18985 4820 19045 5020
rect 31377 6076 31777 6136
rect 31377 5958 31777 6018
rect 38088 5891 38148 6291
rect 38206 5891 38266 6291
rect 38441 6091 38501 6291
rect 39445 6290 39505 6490
rect 39865 6090 39925 6490
rect 39983 6090 40043 6490
rect 40101 6090 40161 6490
rect 40219 6090 40279 6490
rect 40743 6290 40803 6490
rect 41343 6290 41403 6490
rect 41763 6090 41823 6490
rect 41881 6090 41941 6490
rect 41999 6090 42059 6490
rect 42117 6090 42177 6490
rect 42641 6290 42701 6490
rect 51296 7515 51356 7915
rect 51414 7515 51474 7915
rect 51649 7715 51709 7915
rect 57921 7583 57981 7983
rect 58039 7583 58099 7983
rect 58274 7783 58334 7983
rect 44637 5979 44697 6379
rect 44755 5979 44815 6379
rect 44990 6179 45050 6379
rect 45994 6378 46054 6578
rect 46414 6178 46474 6578
rect 46532 6178 46592 6578
rect 46650 6178 46710 6578
rect 46768 6178 46828 6578
rect 47292 6378 47352 6578
rect 47892 6378 47952 6578
rect 48312 6178 48372 6578
rect 48430 6178 48490 6578
rect 48548 6178 48608 6578
rect 48666 6178 48726 6578
rect 49190 6378 49250 6578
rect 71846 7953 72246 8013
rect 19755 4818 19815 5018
rect 20279 4618 20339 5018
rect 20397 4618 20457 5018
rect 20515 4618 20575 5018
rect 20633 4618 20693 5018
rect 21053 4818 21113 5018
rect 21824 4820 21884 5020
rect 22348 4620 22408 5020
rect 22466 4620 22526 5020
rect 22584 4620 22644 5020
rect 22702 4620 22762 5020
rect 23122 4820 23182 5020
rect 51291 5911 51351 6311
rect 51409 5911 51469 6311
rect 51644 6111 51704 6311
rect 52648 6310 52708 6510
rect 53068 6110 53128 6510
rect 53186 6110 53246 6510
rect 53304 6110 53364 6510
rect 53422 6110 53482 6510
rect 53946 6310 54006 6510
rect 54546 6310 54606 6510
rect 54966 6110 55026 6510
rect 55084 6110 55144 6510
rect 55202 6110 55262 6510
rect 55320 6110 55380 6510
rect 55844 6310 55904 6510
rect 71846 7757 72046 7817
rect 57916 5979 57976 6379
rect 58034 5979 58094 6379
rect 58269 6179 58329 6379
rect 59273 6378 59333 6578
rect 59693 6178 59753 6578
rect 59811 6178 59871 6578
rect 59929 6178 59989 6578
rect 60047 6178 60107 6578
rect 60571 6378 60631 6578
rect 61171 6378 61231 6578
rect 61591 6178 61651 6578
rect 61709 6178 61769 6578
rect 61827 6178 61887 6578
rect 61945 6178 62005 6578
rect 62469 6378 62529 6578
rect 67312 6666 67372 7066
rect 67430 6666 67490 7066
rect 67665 6866 67725 7066
rect 65407 6081 65467 6281
rect 63704 5561 63764 5961
rect 63822 5561 63882 5961
rect 64057 5761 64117 5961
rect 65827 5881 65887 6281
rect 65945 5881 66005 6281
rect 66063 5881 66123 6281
rect 66181 5881 66241 6281
rect 66705 6081 66765 6281
rect 31377 5434 31577 5494
rect 71846 5355 72046 5415
rect 71846 5163 72246 5223
rect 23892 4818 23952 5018
rect 24416 4618 24476 5018
rect 24534 4618 24594 5018
rect 24652 4618 24712 5018
rect 24770 4618 24830 5018
rect 25190 4818 25250 5018
rect 71846 5045 72246 5105
rect 71846 4927 72246 4987
rect 71846 4809 72246 4869
rect 31377 4663 31577 4723
rect 31377 4243 31777 4303
rect 31377 4125 31777 4185
rect 31377 4007 31777 4067
rect 31377 3889 31777 3949
rect 35162 3549 35222 3949
rect 35280 3549 35340 3949
rect 35515 3749 35575 3949
rect 31377 3365 31577 3425
rect 38071 3365 38131 3765
rect 38189 3365 38249 3765
rect 38424 3565 38484 3765
rect 40069 3291 40129 3491
rect 40187 3291 40247 3491
rect 40305 3291 40365 3491
rect 41211 3295 41271 3495
rect 41329 3295 41389 3495
rect 41447 3295 41507 3495
rect 44622 3363 44682 3763
rect 44740 3363 44800 3763
rect 44975 3563 45035 3763
rect 71846 4613 72046 4673
rect 46620 3289 46680 3489
rect 46738 3289 46798 3489
rect 46856 3289 46916 3489
rect 47762 3293 47822 3493
rect 47880 3293 47940 3493
rect 47998 3293 48058 3493
rect 51277 3364 51337 3764
rect 51395 3364 51455 3764
rect 51630 3564 51690 3764
rect 53275 3290 53335 3490
rect 53393 3290 53453 3490
rect 53511 3290 53571 3490
rect 54417 3294 54477 3494
rect 54535 3294 54595 3494
rect 54653 3294 54713 3494
rect 57899 3365 57959 3765
rect 58017 3365 58077 3765
rect 58252 3565 58312 3765
rect 63775 3641 63835 4041
rect 63893 3641 63953 4041
rect 64128 3841 64188 4041
rect 59897 3291 59957 3491
rect 60015 3291 60075 3491
rect 60133 3291 60193 3491
rect 61039 3295 61099 3495
rect 61157 3295 61217 3495
rect 61275 3295 61335 3495
rect 67312 3171 67372 3571
rect 67430 3171 67490 3571
rect 67665 3371 67725 3571
rect 31375 2595 31575 2655
rect 31375 2175 31775 2235
rect 31375 2057 31775 2117
rect 65407 2586 65467 2786
rect 65827 2386 65887 2786
rect 65945 2386 66005 2786
rect 66063 2386 66123 2786
rect 66181 2386 66241 2786
rect 66705 2586 66765 2786
rect 1140 607 1200 807
rect 1332 407 1392 807
rect 1450 407 1510 807
rect 1568 407 1628 807
rect 1686 407 1746 807
rect 1882 607 1942 807
rect 4284 607 4344 807
rect 4476 407 4536 807
rect 4594 407 4654 807
rect 4712 407 4772 807
rect 4830 407 4890 807
rect 5026 607 5086 807
rect 7416 611 7476 811
rect 7608 411 7668 811
rect 7726 411 7786 811
rect 7844 411 7904 811
rect 7962 411 8022 811
rect 8158 611 8218 811
rect 10560 611 10620 811
rect 10752 411 10812 811
rect 10870 411 10930 811
rect 10988 411 11048 811
rect 11106 411 11166 811
rect 11302 611 11362 811
rect 31375 1939 31775 1999
rect 31375 1821 31775 1881
rect 38085 1715 38145 2115
rect 38203 1715 38263 2115
rect 38438 1915 38498 2115
rect 31375 1297 31575 1357
rect 13762 607 13822 807
rect 13954 407 14014 807
rect 14072 407 14132 807
rect 14190 407 14250 807
rect 14308 407 14368 807
rect 14504 607 14564 807
rect 16906 607 16966 807
rect 17098 407 17158 807
rect 17216 407 17276 807
rect 17334 407 17394 807
rect 17452 407 17512 807
rect 17648 607 17708 807
rect 20038 611 20098 811
rect 20230 411 20290 811
rect 20348 411 20408 811
rect 20466 411 20526 811
rect 20584 411 20644 811
rect 20780 611 20840 811
rect 23182 611 23242 811
rect 23374 411 23434 811
rect 23492 411 23552 811
rect 23610 411 23670 811
rect 23728 411 23788 811
rect 23924 611 23984 811
rect 35178 789 35238 1189
rect 35296 789 35356 1189
rect 35531 989 35591 1189
rect 31377 526 31577 586
rect 44636 1713 44696 2113
rect 44754 1713 44814 2113
rect 44989 1913 45049 2113
rect 31377 106 31777 166
rect 38080 111 38140 511
rect 38198 111 38258 511
rect 38433 311 38493 511
rect 39437 510 39497 710
rect 39857 310 39917 710
rect 39975 310 40035 710
rect 40093 310 40153 710
rect 40211 310 40271 710
rect 40735 510 40795 710
rect 41335 510 41395 710
rect 41755 310 41815 710
rect 41873 310 41933 710
rect 41991 310 42051 710
rect 42109 310 42169 710
rect 42633 510 42693 710
rect 51291 1714 51351 2114
rect 51409 1714 51469 2114
rect 51644 1914 51704 2114
rect 31377 -12 31777 48
rect 44631 109 44691 509
rect 44749 109 44809 509
rect 44984 309 45044 509
rect 45988 508 46048 708
rect 46408 308 46468 708
rect 46526 308 46586 708
rect 46644 308 46704 708
rect 46762 308 46822 708
rect 47286 508 47346 708
rect 47886 508 47946 708
rect 48306 308 48366 708
rect 48424 308 48484 708
rect 48542 308 48602 708
rect 48660 308 48720 708
rect 49184 508 49244 708
rect 57913 1715 57973 2115
rect 58031 1715 58091 2115
rect 58266 1915 58326 2115
rect 71842 2223 72042 2283
rect 71842 2031 72242 2091
rect 71842 1913 72242 1973
rect 31377 -130 31777 -70
rect 51286 110 51346 510
rect 51404 110 51464 510
rect 51639 310 51699 510
rect 52643 509 52703 709
rect 53063 309 53123 709
rect 53181 309 53241 709
rect 53299 309 53359 709
rect 53417 309 53477 709
rect 53941 509 54001 709
rect 54541 509 54601 709
rect 54961 309 55021 709
rect 55079 309 55139 709
rect 55197 309 55257 709
rect 55315 309 55375 709
rect 55839 509 55899 709
rect 71842 1795 72242 1855
rect 71842 1677 72242 1737
rect 71842 1481 72042 1541
rect 57908 111 57968 511
rect 58026 111 58086 511
rect 58261 311 58321 511
rect 59265 510 59325 710
rect 59685 310 59745 710
rect 59803 310 59863 710
rect 59921 310 59981 710
rect 60039 310 60099 710
rect 60563 510 60623 710
rect 61163 510 61223 710
rect 61583 310 61643 710
rect 61701 310 61761 710
rect 61819 310 61879 710
rect 61937 310 61997 710
rect 62461 510 62521 710
rect 63772 571 63832 971
rect 63890 571 63950 971
rect 64125 771 64185 971
rect 31377 -248 31777 -188
rect 31377 -772 31577 -712
rect 41888 -1318 41948 -918
rect 42006 -1318 42066 -918
rect 42241 -1318 42301 -1118
rect 48442 -1313 48502 -913
rect 48560 -1313 48620 -913
rect 48795 -1313 48855 -1113
rect 31375 -1542 31575 -1482
rect 55091 -1325 55151 -925
rect 55209 -1325 55269 -925
rect 55444 -1325 55504 -1125
rect 67312 -1177 67372 -777
rect 67430 -1177 67490 -777
rect 67665 -977 67725 -777
rect 71842 -921 72042 -861
rect 71842 -1113 72242 -1053
rect 71842 -1231 72242 -1171
rect 71842 -1349 72242 -1289
rect 71842 -1467 72242 -1407
rect 65407 -1762 65467 -1562
rect 1172 -3285 1232 -3085
rect 1364 -3485 1424 -3085
rect 1482 -3485 1542 -3085
rect 1600 -3485 1660 -3085
rect 1718 -3485 1778 -3085
rect 1914 -3285 1974 -3085
rect 4316 -3285 4376 -3085
rect 4508 -3485 4568 -3085
rect 4626 -3485 4686 -3085
rect 4744 -3485 4804 -3085
rect 4862 -3485 4922 -3085
rect 5058 -3285 5118 -3085
rect 7448 -3281 7508 -3081
rect 7640 -3481 7700 -3081
rect 7758 -3481 7818 -3081
rect 7876 -3481 7936 -3081
rect 7994 -3481 8054 -3081
rect 8190 -3281 8250 -3081
rect 10592 -3281 10652 -3081
rect 10784 -3481 10844 -3081
rect 10902 -3481 10962 -3081
rect 11020 -3481 11080 -3081
rect 11138 -3481 11198 -3081
rect 11334 -3281 11394 -3081
rect 31375 -1962 31775 -1902
rect 31375 -2080 31775 -2020
rect 31375 -2198 31775 -2138
rect 31375 -2316 31775 -2256
rect 63779 -2274 63839 -1874
rect 63897 -2274 63957 -1874
rect 64132 -2074 64192 -1874
rect 65827 -1962 65887 -1562
rect 65945 -1962 66005 -1562
rect 66063 -1962 66123 -1562
rect 66181 -1962 66241 -1562
rect 66705 -1762 66765 -1562
rect 71842 -1663 72042 -1603
rect 31375 -2840 31575 -2780
rect 13794 -3285 13854 -3085
rect 13986 -3485 14046 -3085
rect 14104 -3485 14164 -3085
rect 14222 -3485 14282 -3085
rect 14340 -3485 14400 -3085
rect 14536 -3285 14596 -3085
rect 16938 -3285 16998 -3085
rect 17130 -3485 17190 -3085
rect 17248 -3485 17308 -3085
rect 17366 -3485 17426 -3085
rect 17484 -3485 17544 -3085
rect 17680 -3285 17740 -3085
rect 20070 -3281 20130 -3081
rect 20262 -3481 20322 -3081
rect 20380 -3481 20440 -3081
rect 20498 -3481 20558 -3081
rect 20616 -3481 20676 -3081
rect 20812 -3281 20872 -3081
rect 23214 -3281 23274 -3081
rect 23406 -3481 23466 -3081
rect 23524 -3481 23584 -3081
rect 23642 -3481 23702 -3081
rect 23760 -3481 23820 -3081
rect 23956 -3281 24016 -3081
<< pmos >>
rect 39646 24333 39706 24533
rect 39764 24333 39824 24533
rect 39882 24333 39942 24533
rect 40000 24333 40060 24533
rect 40118 24333 40178 24533
rect 40236 24333 40296 24533
rect 40354 24333 40414 24533
rect 40472 24333 40532 24533
rect 40590 24333 40650 24533
rect 41971 24205 42031 24605
rect 42089 24205 42149 24605
rect 42207 24205 42267 24605
rect 42325 24205 42385 24605
rect 42443 24205 42503 24605
rect 42561 24205 42621 24605
rect 43113 24209 43173 24609
rect 43231 24209 43291 24609
rect 43349 24209 43409 24609
rect 43467 24209 43527 24609
rect 43585 24209 43645 24609
rect 43703 24209 43763 24609
rect 46159 24330 46219 24530
rect 46277 24330 46337 24530
rect 46395 24330 46455 24530
rect 46513 24330 46573 24530
rect 46631 24330 46691 24530
rect 46749 24330 46809 24530
rect 46867 24330 46927 24530
rect 46985 24330 47045 24530
rect 47103 24330 47163 24530
rect 48484 24202 48544 24602
rect 48602 24202 48662 24602
rect 48720 24202 48780 24602
rect 48838 24202 48898 24602
rect 48956 24202 49016 24602
rect 49074 24202 49134 24602
rect 49626 24206 49686 24606
rect 49744 24206 49804 24606
rect 49862 24206 49922 24606
rect 49980 24206 50040 24606
rect 50098 24206 50158 24606
rect 50216 24206 50276 24606
rect 52693 24325 52753 24525
rect 52811 24325 52871 24525
rect 52929 24325 52989 24525
rect 53047 24325 53107 24525
rect 53165 24325 53225 24525
rect 53283 24325 53343 24525
rect 53401 24325 53461 24525
rect 53519 24325 53579 24525
rect 53637 24325 53697 24525
rect 42400 23622 42460 23822
rect 42518 23622 42578 23822
rect 42636 23622 42696 23822
rect 43542 23626 43602 23826
rect 43660 23626 43720 23826
rect 43778 23626 43838 23826
rect 55018 24197 55078 24597
rect 55136 24197 55196 24597
rect 55254 24197 55314 24597
rect 55372 24197 55432 24597
rect 55490 24197 55550 24597
rect 55608 24197 55668 24597
rect 56160 24201 56220 24601
rect 56278 24201 56338 24601
rect 56396 24201 56456 24601
rect 56514 24201 56574 24601
rect 56632 24201 56692 24601
rect 56750 24201 56810 24601
rect 59251 24329 59311 24529
rect 59369 24329 59429 24529
rect 59487 24329 59547 24529
rect 59605 24329 59665 24529
rect 59723 24329 59783 24529
rect 59841 24329 59901 24529
rect 59959 24329 60019 24529
rect 60077 24329 60137 24529
rect 60195 24329 60255 24529
rect 48913 23619 48973 23819
rect 49031 23619 49091 23819
rect 49149 23619 49209 23819
rect 50055 23623 50115 23823
rect 50173 23623 50233 23823
rect 50291 23623 50351 23823
rect 61576 24201 61636 24601
rect 61694 24201 61754 24601
rect 61812 24201 61872 24601
rect 61930 24201 61990 24601
rect 62048 24201 62108 24601
rect 62166 24201 62226 24601
rect 62718 24205 62778 24605
rect 62836 24205 62896 24605
rect 62954 24205 63014 24605
rect 63072 24205 63132 24605
rect 63190 24205 63250 24605
rect 63308 24205 63368 24605
rect 55447 23614 55507 23814
rect 55565 23614 55625 23814
rect 55683 23614 55743 23814
rect 56589 23618 56649 23818
rect 56707 23618 56767 23818
rect 56825 23618 56885 23818
rect 62005 23618 62065 23818
rect 62123 23618 62183 23818
rect 62241 23618 62301 23818
rect 63147 23622 63207 23822
rect 63265 23622 63325 23822
rect 63383 23622 63443 23822
rect 39660 22683 39720 22883
rect 39778 22683 39838 22883
rect 39896 22683 39956 22883
rect 40014 22683 40074 22883
rect 40132 22683 40192 22883
rect 40250 22683 40310 22883
rect 40368 22683 40428 22883
rect 40486 22683 40546 22883
rect 40604 22683 40664 22883
rect 46173 22680 46233 22880
rect 46291 22680 46351 22880
rect 46409 22680 46469 22880
rect 46527 22680 46587 22880
rect 46645 22680 46705 22880
rect 46763 22680 46823 22880
rect 46881 22680 46941 22880
rect 46999 22680 47059 22880
rect 47117 22680 47177 22880
rect 3058 21596 3118 21796
rect 3176 21596 3236 21796
rect 3294 21596 3354 21796
rect 3531 21596 3591 21996
rect 3649 21596 3709 21996
rect 3767 21596 3827 21996
rect 4004 21596 4064 21996
rect 4122 21596 4182 21996
rect 4240 21596 4300 21996
rect 4358 21596 4418 21996
rect 4476 21596 4536 21996
rect 4594 21596 4654 21996
rect 4825 21596 4885 21996
rect 4943 21596 5003 21996
rect 5061 21596 5121 21996
rect 5266 21596 5326 21796
rect 5384 21596 5444 21796
rect 5502 21596 5562 21796
rect 6202 21596 6262 21796
rect 6320 21596 6380 21796
rect 6438 21596 6498 21796
rect 6675 21596 6735 21996
rect 6793 21596 6853 21996
rect 6911 21596 6971 21996
rect 7148 21596 7208 21996
rect 7266 21596 7326 21996
rect 7384 21596 7444 21996
rect 7502 21596 7562 21996
rect 7620 21596 7680 21996
rect 7738 21596 7798 21996
rect 7969 21596 8029 21996
rect 8087 21596 8147 21996
rect 8205 21596 8265 21996
rect 8410 21596 8470 21796
rect 8528 21596 8588 21796
rect 8646 21596 8706 21796
rect 9334 21592 9394 21792
rect 9452 21592 9512 21792
rect 9570 21592 9630 21792
rect 9807 21592 9867 21992
rect 9925 21592 9985 21992
rect 10043 21592 10103 21992
rect 10280 21592 10340 21992
rect 10398 21592 10458 21992
rect 10516 21592 10576 21992
rect 10634 21592 10694 21992
rect 10752 21592 10812 21992
rect 10870 21592 10930 21992
rect 11101 21592 11161 21992
rect 11219 21592 11279 21992
rect 11337 21592 11397 21992
rect 11542 21592 11602 21792
rect 11660 21592 11720 21792
rect 11778 21592 11838 21792
rect 12478 21592 12538 21792
rect 12596 21592 12656 21792
rect 12714 21592 12774 21792
rect 12951 21592 13011 21992
rect 13069 21592 13129 21992
rect 13187 21592 13247 21992
rect 13424 21592 13484 21992
rect 13542 21592 13602 21992
rect 13660 21592 13720 21992
rect 13778 21592 13838 21992
rect 13896 21592 13956 21992
rect 14014 21592 14074 21992
rect 14245 21592 14305 21992
rect 14363 21592 14423 21992
rect 14481 21592 14541 21992
rect 14686 21592 14746 21792
rect 14804 21592 14864 21792
rect 14922 21592 14982 21792
rect 15680 21596 15740 21796
rect 15798 21596 15858 21796
rect 15916 21596 15976 21796
rect 16153 21596 16213 21996
rect 16271 21596 16331 21996
rect 16389 21596 16449 21996
rect 16626 21596 16686 21996
rect 16744 21596 16804 21996
rect 16862 21596 16922 21996
rect 16980 21596 17040 21996
rect 17098 21596 17158 21996
rect 17216 21596 17276 21996
rect 17447 21596 17507 21996
rect 17565 21596 17625 21996
rect 17683 21596 17743 21996
rect 17888 21596 17948 21796
rect 18006 21596 18066 21796
rect 18124 21596 18184 21796
rect 18824 21596 18884 21796
rect 18942 21596 19002 21796
rect 19060 21596 19120 21796
rect 19297 21596 19357 21996
rect 19415 21596 19475 21996
rect 19533 21596 19593 21996
rect 19770 21596 19830 21996
rect 19888 21596 19948 21996
rect 20006 21596 20066 21996
rect 20124 21596 20184 21996
rect 20242 21596 20302 21996
rect 20360 21596 20420 21996
rect 20591 21596 20651 21996
rect 20709 21596 20769 21996
rect 20827 21596 20887 21996
rect 21032 21596 21092 21796
rect 21150 21596 21210 21796
rect 21268 21596 21328 21796
rect 21956 21592 22016 21792
rect 22074 21592 22134 21792
rect 22192 21592 22252 21792
rect 22429 21592 22489 21992
rect 22547 21592 22607 21992
rect 22665 21592 22725 21992
rect 22902 21592 22962 21992
rect 23020 21592 23080 21992
rect 23138 21592 23198 21992
rect 23256 21592 23316 21992
rect 23374 21592 23434 21992
rect 23492 21592 23552 21992
rect 23723 21592 23783 21992
rect 23841 21592 23901 21992
rect 23959 21592 24019 21992
rect 24164 21592 24224 21792
rect 24282 21592 24342 21792
rect 24400 21592 24460 21792
rect 25100 21592 25160 21792
rect 25218 21592 25278 21792
rect 25336 21592 25396 21792
rect 25573 21592 25633 21992
rect 25691 21592 25751 21992
rect 25809 21592 25869 21992
rect 26046 21592 26106 21992
rect 26164 21592 26224 21992
rect 26282 21592 26342 21992
rect 26400 21592 26460 21992
rect 26518 21592 26578 21992
rect 26636 21592 26696 21992
rect 26867 21592 26927 21992
rect 26985 21592 27045 21992
rect 27103 21592 27163 21992
rect 41124 22066 41184 22266
rect 41242 22066 41302 22266
rect 41360 22066 41420 22266
rect 41608 22066 41668 22466
rect 41726 22066 41786 22466
rect 41844 22066 41904 22466
rect 41962 22066 42022 22466
rect 42080 22066 42140 22466
rect 42198 22066 42258 22466
rect 42445 22066 42505 22266
rect 42563 22066 42623 22266
rect 42681 22066 42741 22266
rect 43022 22066 43082 22266
rect 43140 22066 43200 22266
rect 43258 22066 43318 22266
rect 43506 22066 43566 22466
rect 43624 22066 43684 22466
rect 43742 22066 43802 22466
rect 43860 22066 43920 22466
rect 43978 22066 44038 22466
rect 44096 22066 44156 22466
rect 52707 22675 52767 22875
rect 52825 22675 52885 22875
rect 52943 22675 53003 22875
rect 53061 22675 53121 22875
rect 53179 22675 53239 22875
rect 53297 22675 53357 22875
rect 53415 22675 53475 22875
rect 53533 22675 53593 22875
rect 53651 22675 53711 22875
rect 59265 22679 59325 22879
rect 59383 22679 59443 22879
rect 59501 22679 59561 22879
rect 59619 22679 59679 22879
rect 59737 22679 59797 22879
rect 59855 22679 59915 22879
rect 59973 22679 60033 22879
rect 60091 22679 60151 22879
rect 60209 22679 60269 22879
rect 44343 22066 44403 22266
rect 44461 22066 44521 22266
rect 44579 22066 44639 22266
rect 27308 21592 27368 21792
rect 27426 21592 27486 21792
rect 27544 21592 27604 21792
rect 39655 21079 39715 21279
rect 39773 21079 39833 21279
rect 39891 21079 39951 21279
rect 40009 21079 40069 21279
rect 40127 21079 40187 21279
rect 40245 21079 40305 21279
rect 40363 21079 40423 21279
rect 40481 21079 40541 21279
rect 40599 21079 40659 21279
rect 41551 21373 41611 21773
rect 41669 21373 41729 21773
rect 41787 21373 41847 21773
rect 41905 21373 41965 21773
rect 42023 21373 42083 21773
rect 42141 21373 42201 21773
rect 47637 22063 47697 22263
rect 47755 22063 47815 22263
rect 47873 22063 47933 22263
rect 48121 22063 48181 22463
rect 48239 22063 48299 22463
rect 48357 22063 48417 22463
rect 48475 22063 48535 22463
rect 48593 22063 48653 22463
rect 48711 22063 48771 22463
rect 48958 22063 49018 22263
rect 49076 22063 49136 22263
rect 49194 22063 49254 22263
rect 49535 22063 49595 22263
rect 49653 22063 49713 22263
rect 49771 22063 49831 22263
rect 50019 22063 50079 22463
rect 50137 22063 50197 22463
rect 50255 22063 50315 22463
rect 50373 22063 50433 22463
rect 50491 22063 50551 22463
rect 50609 22063 50669 22463
rect 50856 22063 50916 22263
rect 50974 22063 51034 22263
rect 51092 22063 51152 22263
rect 43449 21373 43509 21773
rect 43567 21373 43627 21773
rect 43685 21373 43745 21773
rect 43803 21373 43863 21773
rect 43921 21373 43981 21773
rect 44039 21373 44099 21773
rect 46168 21076 46228 21276
rect 46286 21076 46346 21276
rect 46404 21076 46464 21276
rect 46522 21076 46582 21276
rect 46640 21076 46700 21276
rect 46758 21076 46818 21276
rect 46876 21076 46936 21276
rect 46994 21076 47054 21276
rect 47112 21076 47172 21276
rect 48064 21370 48124 21770
rect 48182 21370 48242 21770
rect 48300 21370 48360 21770
rect 48418 21370 48478 21770
rect 48536 21370 48596 21770
rect 48654 21370 48714 21770
rect 54171 22058 54231 22258
rect 54289 22058 54349 22258
rect 54407 22058 54467 22258
rect 54655 22058 54715 22458
rect 54773 22058 54833 22458
rect 54891 22058 54951 22458
rect 55009 22058 55069 22458
rect 55127 22058 55187 22458
rect 55245 22058 55305 22458
rect 55492 22058 55552 22258
rect 55610 22058 55670 22258
rect 55728 22058 55788 22258
rect 56069 22058 56129 22258
rect 56187 22058 56247 22258
rect 56305 22058 56365 22258
rect 56553 22058 56613 22458
rect 56671 22058 56731 22458
rect 56789 22058 56849 22458
rect 56907 22058 56967 22458
rect 57025 22058 57085 22458
rect 57143 22058 57203 22458
rect 57390 22058 57450 22258
rect 57508 22058 57568 22258
rect 57626 22058 57686 22258
rect 49962 21370 50022 21770
rect 50080 21370 50140 21770
rect 50198 21370 50258 21770
rect 50316 21370 50376 21770
rect 50434 21370 50494 21770
rect 50552 21370 50612 21770
rect 52702 21071 52762 21271
rect 52820 21071 52880 21271
rect 52938 21071 52998 21271
rect 53056 21071 53116 21271
rect 53174 21071 53234 21271
rect 53292 21071 53352 21271
rect 53410 21071 53470 21271
rect 53528 21071 53588 21271
rect 53646 21071 53706 21271
rect 54598 21365 54658 21765
rect 54716 21365 54776 21765
rect 54834 21365 54894 21765
rect 54952 21365 55012 21765
rect 55070 21365 55130 21765
rect 55188 21365 55248 21765
rect 60729 22062 60789 22262
rect 60847 22062 60907 22262
rect 60965 22062 61025 22262
rect 61213 22062 61273 22462
rect 61331 22062 61391 22462
rect 61449 22062 61509 22462
rect 61567 22062 61627 22462
rect 61685 22062 61745 22462
rect 61803 22062 61863 22462
rect 62050 22062 62110 22262
rect 62168 22062 62228 22262
rect 62286 22062 62346 22262
rect 62627 22062 62687 22262
rect 62745 22062 62805 22262
rect 62863 22062 62923 22262
rect 63111 22062 63171 22462
rect 63229 22062 63289 22462
rect 63347 22062 63407 22462
rect 63465 22062 63525 22462
rect 63583 22062 63643 22462
rect 63701 22062 63761 22462
rect 63948 22062 64008 22262
rect 64066 22062 64126 22262
rect 64184 22062 64244 22262
rect 56496 21365 56556 21765
rect 56614 21365 56674 21765
rect 56732 21365 56792 21765
rect 56850 21365 56910 21765
rect 56968 21365 57028 21765
rect 57086 21365 57146 21765
rect 59260 21075 59320 21275
rect 59378 21075 59438 21275
rect 59496 21075 59556 21275
rect 59614 21075 59674 21275
rect 59732 21075 59792 21275
rect 59850 21075 59910 21275
rect 59968 21075 60028 21275
rect 60086 21075 60146 21275
rect 60204 21075 60264 21275
rect 61156 21369 61216 21769
rect 61274 21369 61334 21769
rect 61392 21369 61452 21769
rect 61510 21369 61570 21769
rect 61628 21369 61688 21769
rect 61746 21369 61806 21769
rect 70713 21955 70913 22015
rect 63054 21369 63114 21769
rect 63172 21369 63232 21769
rect 63290 21369 63350 21769
rect 63408 21369 63468 21769
rect 63526 21369 63586 21769
rect 63644 21369 63704 21769
rect 70713 21837 70913 21897
rect 70713 21719 70913 21779
rect 70513 21514 70913 21574
rect 70513 21396 70913 21456
rect 70513 21278 70913 21338
rect 70513 21047 70913 21107
rect 70513 20929 70913 20989
rect 70513 20811 70913 20871
rect 70513 20693 70913 20753
rect 70513 20575 70913 20635
rect 70513 20457 70913 20517
rect 70513 20220 70913 20280
rect 70513 20102 70913 20162
rect 70513 19984 70913 20044
rect 70713 19747 70913 19807
rect 70713 19629 70913 19689
rect 70713 19511 70913 19571
rect 39657 18601 39717 19001
rect 39775 18601 39835 19001
rect 39893 18601 39953 19001
rect 40011 18601 40071 19001
rect 40129 18601 40189 19001
rect 40247 18601 40307 19001
rect 40799 18597 40859 18997
rect 40917 18597 40977 18997
rect 41035 18597 41095 18997
rect 41153 18597 41213 18997
rect 41271 18597 41331 18997
rect 41389 18597 41449 18997
rect 42770 18725 42830 18925
rect 42888 18725 42948 18925
rect 43006 18725 43066 18925
rect 43124 18725 43184 18925
rect 43242 18725 43302 18925
rect 43360 18725 43420 18925
rect 43478 18725 43538 18925
rect 43596 18725 43656 18925
rect 43714 18725 43774 18925
rect 46215 18597 46275 18997
rect 46333 18597 46393 18997
rect 46451 18597 46511 18997
rect 46569 18597 46629 18997
rect 46687 18597 46747 18997
rect 46805 18597 46865 18997
rect 39582 18018 39642 18218
rect 39700 18018 39760 18218
rect 39818 18018 39878 18218
rect 40724 18014 40784 18214
rect 40842 18014 40902 18214
rect 40960 18014 41020 18214
rect 47357 18593 47417 18993
rect 47475 18593 47535 18993
rect 47593 18593 47653 18993
rect 47711 18593 47771 18993
rect 47829 18593 47889 18993
rect 47947 18593 48007 18993
rect 49328 18721 49388 18921
rect 49446 18721 49506 18921
rect 49564 18721 49624 18921
rect 49682 18721 49742 18921
rect 49800 18721 49860 18921
rect 49918 18721 49978 18921
rect 50036 18721 50096 18921
rect 50154 18721 50214 18921
rect 50272 18721 50332 18921
rect 52749 18602 52809 19002
rect 52867 18602 52927 19002
rect 52985 18602 53045 19002
rect 53103 18602 53163 19002
rect 53221 18602 53281 19002
rect 53339 18602 53399 19002
rect 46140 18014 46200 18214
rect 46258 18014 46318 18214
rect 46376 18014 46436 18214
rect 47282 18010 47342 18210
rect 47400 18010 47460 18210
rect 47518 18010 47578 18210
rect 53891 18598 53951 18998
rect 54009 18598 54069 18998
rect 54127 18598 54187 18998
rect 54245 18598 54305 18998
rect 54363 18598 54423 18998
rect 54481 18598 54541 18998
rect 55862 18726 55922 18926
rect 55980 18726 56040 18926
rect 56098 18726 56158 18926
rect 56216 18726 56276 18926
rect 56334 18726 56394 18926
rect 56452 18726 56512 18926
rect 56570 18726 56630 18926
rect 56688 18726 56748 18926
rect 56806 18726 56866 18926
rect 59262 18605 59322 19005
rect 59380 18605 59440 19005
rect 59498 18605 59558 19005
rect 59616 18605 59676 19005
rect 59734 18605 59794 19005
rect 59852 18605 59912 19005
rect 52674 18019 52734 18219
rect 52792 18019 52852 18219
rect 52910 18019 52970 18219
rect 53816 18015 53876 18215
rect 53934 18015 53994 18215
rect 54052 18015 54112 18215
rect 60404 18601 60464 19001
rect 60522 18601 60582 19001
rect 60640 18601 60700 19001
rect 60758 18601 60818 19001
rect 60876 18601 60936 19001
rect 60994 18601 61054 19001
rect 62375 18729 62435 18929
rect 62493 18729 62553 18929
rect 62611 18729 62671 18929
rect 62729 18729 62789 18929
rect 62847 18729 62907 18929
rect 62965 18729 63025 18929
rect 63083 18729 63143 18929
rect 63201 18729 63261 18929
rect 63319 18729 63379 18929
rect 70713 18811 70913 18871
rect 70713 18693 70913 18753
rect 70713 18575 70913 18635
rect 59187 18022 59247 18222
rect 59305 18022 59365 18222
rect 59423 18022 59483 18222
rect 60329 18018 60389 18218
rect 60447 18018 60507 18218
rect 60565 18018 60625 18218
rect 70513 18370 70913 18430
rect 70513 18252 70913 18312
rect 70513 18134 70913 18194
rect 70513 17903 70913 17963
rect 70513 17785 70913 17845
rect 70513 17667 70913 17727
rect 70513 17549 70913 17609
rect 70513 17431 70913 17491
rect 4566 16408 4626 16808
rect 4684 16408 4744 16808
rect 4802 16408 4862 16808
rect 4920 16408 4980 16808
rect 5038 16408 5098 16808
rect 5156 16408 5216 16808
rect 5734 16410 5794 16810
rect 5852 16410 5912 16810
rect 5970 16410 6030 16810
rect 6088 16410 6148 16810
rect 6206 16410 6266 16810
rect 6324 16410 6384 16810
rect 42756 17075 42816 17275
rect 42874 17075 42934 17275
rect 42992 17075 43052 17275
rect 43110 17075 43170 17275
rect 43228 17075 43288 17275
rect 43346 17075 43406 17275
rect 43464 17075 43524 17275
rect 43582 17075 43642 17275
rect 43700 17075 43760 17275
rect 49314 17071 49374 17271
rect 49432 17071 49492 17271
rect 49550 17071 49610 17271
rect 49668 17071 49728 17271
rect 49786 17071 49846 17271
rect 49904 17071 49964 17271
rect 50022 17071 50082 17271
rect 50140 17071 50200 17271
rect 50258 17071 50318 17271
rect 55848 17076 55908 17276
rect 55966 17076 56026 17276
rect 56084 17076 56144 17276
rect 56202 17076 56262 17276
rect 56320 17076 56380 17276
rect 56438 17076 56498 17276
rect 56556 17076 56616 17276
rect 56674 17076 56734 17276
rect 56792 17076 56852 17276
rect 70513 17313 70913 17373
rect 62361 17079 62421 17279
rect 62479 17079 62539 17279
rect 62597 17079 62657 17279
rect 62715 17079 62775 17279
rect 62833 17079 62893 17279
rect 62951 17079 63011 17279
rect 63069 17079 63129 17279
rect 63187 17079 63247 17279
rect 63305 17079 63365 17279
rect 6902 16408 6962 16808
rect 7020 16408 7080 16808
rect 7138 16408 7198 16808
rect 7256 16408 7316 16808
rect 7374 16408 7434 16808
rect 7492 16408 7552 16808
rect 8070 16410 8130 16810
rect 8188 16410 8248 16810
rect 8306 16410 8366 16810
rect 8424 16410 8484 16810
rect 8542 16410 8602 16810
rect 8660 16410 8720 16810
rect 4491 15820 4551 16020
rect 4609 15820 4669 16020
rect 4727 15820 4787 16020
rect 5659 15819 5719 16019
rect 5777 15819 5837 16019
rect 5895 15819 5955 16019
rect 9244 16408 9304 16808
rect 9362 16408 9422 16808
rect 9480 16408 9540 16808
rect 9598 16408 9658 16808
rect 9716 16408 9776 16808
rect 9834 16408 9894 16808
rect 6827 15819 6887 16019
rect 6945 15819 7005 16019
rect 7063 15819 7123 16019
rect 10412 16406 10472 16806
rect 10530 16406 10590 16806
rect 10648 16406 10708 16806
rect 10766 16406 10826 16806
rect 10884 16406 10944 16806
rect 11002 16406 11062 16806
rect 11580 16408 11640 16808
rect 11698 16408 11758 16808
rect 11816 16408 11876 16808
rect 11934 16408 11994 16808
rect 12052 16408 12112 16808
rect 12170 16408 12230 16808
rect 12748 16408 12808 16808
rect 12866 16408 12926 16808
rect 12984 16408 13044 16808
rect 13102 16408 13162 16808
rect 13220 16408 13280 16808
rect 13338 16408 13398 16808
rect 13849 16413 13909 16613
rect 13967 16413 14027 16613
rect 14085 16413 14145 16613
rect 14203 16413 14263 16613
rect 14321 16413 14381 16613
rect 14439 16413 14499 16613
rect 14557 16413 14617 16613
rect 14675 16413 14735 16613
rect 14793 16413 14853 16613
rect 15297 16413 15357 16613
rect 15415 16413 15475 16613
rect 15533 16413 15593 16613
rect 15651 16413 15711 16613
rect 15769 16413 15829 16613
rect 15887 16413 15947 16613
rect 16005 16413 16065 16613
rect 16123 16413 16183 16613
rect 16241 16413 16301 16613
rect 7996 15820 8056 16020
rect 8114 15820 8174 16020
rect 8232 15820 8292 16020
rect 9168 15824 9228 16024
rect 9286 15824 9346 16024
rect 9404 15824 9464 16024
rect 10337 15824 10397 16024
rect 10455 15824 10515 16024
rect 10573 15824 10633 16024
rect 11505 15824 11565 16024
rect 11623 15824 11683 16024
rect 11741 15824 11801 16024
rect 16795 16411 16855 16611
rect 16913 16411 16973 16611
rect 17031 16411 17091 16611
rect 17149 16411 17209 16611
rect 17267 16411 17327 16611
rect 17385 16411 17445 16611
rect 17503 16411 17563 16611
rect 17621 16411 17681 16611
rect 17739 16411 17799 16611
rect 18243 16411 18303 16611
rect 18361 16411 18421 16611
rect 18479 16411 18539 16611
rect 18597 16411 18657 16611
rect 18715 16411 18775 16611
rect 18833 16411 18893 16611
rect 18951 16411 19011 16611
rect 19069 16411 19129 16611
rect 19187 16411 19247 16611
rect 19763 16413 19823 16613
rect 19881 16413 19941 16613
rect 19999 16413 20059 16613
rect 20117 16413 20177 16613
rect 20235 16413 20295 16613
rect 20353 16413 20413 16613
rect 20471 16413 20531 16613
rect 20589 16413 20649 16613
rect 20707 16413 20767 16613
rect 21211 16413 21271 16613
rect 21329 16413 21389 16613
rect 21447 16413 21507 16613
rect 21565 16413 21625 16613
rect 21683 16413 21743 16613
rect 21801 16413 21861 16613
rect 21919 16413 21979 16613
rect 22037 16413 22097 16613
rect 22155 16413 22215 16613
rect 12672 15818 12732 16018
rect 12790 15818 12850 16018
rect 12908 15818 12968 16018
rect 22709 16411 22769 16611
rect 22827 16411 22887 16611
rect 22945 16411 23005 16611
rect 23063 16411 23123 16611
rect 23181 16411 23241 16611
rect 23299 16411 23359 16611
rect 23417 16411 23477 16611
rect 23535 16411 23595 16611
rect 23653 16411 23713 16611
rect 24157 16411 24217 16611
rect 24275 16411 24335 16611
rect 24393 16411 24453 16611
rect 24511 16411 24571 16611
rect 24629 16411 24689 16611
rect 24747 16411 24807 16611
rect 24865 16411 24925 16611
rect 24983 16411 25043 16611
rect 25101 16411 25161 16611
rect 38781 16458 38841 16658
rect 38899 16458 38959 16658
rect 39017 16458 39077 16658
rect 39264 16458 39324 16858
rect 39382 16458 39442 16858
rect 39500 16458 39560 16858
rect 39618 16458 39678 16858
rect 39736 16458 39796 16858
rect 39854 16458 39914 16858
rect 40102 16458 40162 16658
rect 40220 16458 40280 16658
rect 40338 16458 40398 16658
rect 40679 16458 40739 16658
rect 40797 16458 40857 16658
rect 40915 16458 40975 16658
rect 41162 16458 41222 16858
rect 41280 16458 41340 16858
rect 41398 16458 41458 16858
rect 41516 16458 41576 16858
rect 41634 16458 41694 16858
rect 41752 16458 41812 16858
rect 42000 16458 42060 16658
rect 42118 16458 42178 16658
rect 42236 16458 42296 16658
rect 39321 15765 39381 16165
rect 39439 15765 39499 16165
rect 39557 15765 39617 16165
rect 39675 15765 39735 16165
rect 39793 15765 39853 16165
rect 39911 15765 39971 16165
rect 45339 16454 45399 16654
rect 45457 16454 45517 16654
rect 45575 16454 45635 16654
rect 45822 16454 45882 16854
rect 45940 16454 46000 16854
rect 46058 16454 46118 16854
rect 46176 16454 46236 16854
rect 46294 16454 46354 16854
rect 46412 16454 46472 16854
rect 46660 16454 46720 16654
rect 46778 16454 46838 16654
rect 46896 16454 46956 16654
rect 47237 16454 47297 16654
rect 47355 16454 47415 16654
rect 47473 16454 47533 16654
rect 47720 16454 47780 16854
rect 47838 16454 47898 16854
rect 47956 16454 48016 16854
rect 48074 16454 48134 16854
rect 48192 16454 48252 16854
rect 48310 16454 48370 16854
rect 48558 16454 48618 16654
rect 48676 16454 48736 16654
rect 48794 16454 48854 16654
rect 41219 15765 41279 16165
rect 41337 15765 41397 16165
rect 41455 15765 41515 16165
rect 41573 15765 41633 16165
rect 41691 15765 41751 16165
rect 41809 15765 41869 16165
rect 42761 15471 42821 15671
rect 42879 15471 42939 15671
rect 42997 15471 43057 15671
rect 43115 15471 43175 15671
rect 43233 15471 43293 15671
rect 43351 15471 43411 15671
rect 43469 15471 43529 15671
rect 43587 15471 43647 15671
rect 43705 15471 43765 15671
rect 45879 15761 45939 16161
rect 45997 15761 46057 16161
rect 46115 15761 46175 16161
rect 46233 15761 46293 16161
rect 46351 15761 46411 16161
rect 46469 15761 46529 16161
rect 51873 16459 51933 16659
rect 51991 16459 52051 16659
rect 52109 16459 52169 16659
rect 52356 16459 52416 16859
rect 52474 16459 52534 16859
rect 52592 16459 52652 16859
rect 52710 16459 52770 16859
rect 52828 16459 52888 16859
rect 52946 16459 53006 16859
rect 53194 16459 53254 16659
rect 53312 16459 53372 16659
rect 53430 16459 53490 16659
rect 53771 16459 53831 16659
rect 53889 16459 53949 16659
rect 54007 16459 54067 16659
rect 54254 16459 54314 16859
rect 54372 16459 54432 16859
rect 54490 16459 54550 16859
rect 54608 16459 54668 16859
rect 54726 16459 54786 16859
rect 54844 16459 54904 16859
rect 70513 17076 70913 17136
rect 55092 16459 55152 16659
rect 55210 16459 55270 16659
rect 55328 16459 55388 16659
rect 47777 15761 47837 16161
rect 47895 15761 47955 16161
rect 48013 15761 48073 16161
rect 48131 15761 48191 16161
rect 48249 15761 48309 16161
rect 48367 15761 48427 16161
rect 49319 15467 49379 15667
rect 49437 15467 49497 15667
rect 49555 15467 49615 15667
rect 49673 15467 49733 15667
rect 49791 15467 49851 15667
rect 49909 15467 49969 15667
rect 50027 15467 50087 15667
rect 50145 15467 50205 15667
rect 50263 15467 50323 15667
rect 52413 15766 52473 16166
rect 52531 15766 52591 16166
rect 52649 15766 52709 16166
rect 52767 15766 52827 16166
rect 52885 15766 52945 16166
rect 53003 15766 53063 16166
rect 556 14458 616 14658
rect 674 14458 734 14658
rect 792 14458 852 14658
rect 1029 14458 1089 14858
rect 1147 14458 1207 14858
rect 1265 14458 1325 14858
rect 1502 14458 1562 14858
rect 1620 14458 1680 14858
rect 1738 14458 1798 14858
rect 1856 14458 1916 14858
rect 1974 14458 2034 14858
rect 2092 14458 2152 14858
rect 2323 14458 2383 14858
rect 2441 14458 2501 14858
rect 2559 14458 2619 14858
rect 2764 14458 2824 14658
rect 2882 14458 2942 14658
rect 3000 14458 3060 14658
rect 3700 14458 3760 14658
rect 3818 14458 3878 14658
rect 3936 14458 3996 14658
rect 4173 14458 4233 14858
rect 4291 14458 4351 14858
rect 4409 14458 4469 14858
rect 4646 14458 4706 14858
rect 4764 14458 4824 14858
rect 4882 14458 4942 14858
rect 5000 14458 5060 14858
rect 5118 14458 5178 14858
rect 5236 14458 5296 14858
rect 5467 14458 5527 14858
rect 5585 14458 5645 14858
rect 5703 14458 5763 14858
rect 5908 14458 5968 14658
rect 6026 14458 6086 14658
rect 6144 14458 6204 14658
rect 6832 14454 6892 14654
rect 6950 14454 7010 14654
rect 7068 14454 7128 14654
rect 7305 14454 7365 14854
rect 7423 14454 7483 14854
rect 7541 14454 7601 14854
rect 7778 14454 7838 14854
rect 7896 14454 7956 14854
rect 8014 14454 8074 14854
rect 8132 14454 8192 14854
rect 8250 14454 8310 14854
rect 8368 14454 8428 14854
rect 8599 14454 8659 14854
rect 8717 14454 8777 14854
rect 8835 14454 8895 14854
rect 9040 14454 9100 14654
rect 9158 14454 9218 14654
rect 9276 14454 9336 14654
rect 9976 14454 10036 14654
rect 10094 14454 10154 14654
rect 10212 14454 10272 14654
rect 10449 14454 10509 14854
rect 10567 14454 10627 14854
rect 10685 14454 10745 14854
rect 10922 14454 10982 14854
rect 11040 14454 11100 14854
rect 11158 14454 11218 14854
rect 11276 14454 11336 14854
rect 11394 14454 11454 14854
rect 11512 14454 11572 14854
rect 11743 14454 11803 14854
rect 11861 14454 11921 14854
rect 11979 14454 12039 14854
rect 12184 14454 12244 14654
rect 12302 14454 12362 14654
rect 12420 14454 12480 14654
rect 13178 14458 13238 14658
rect 13296 14458 13356 14658
rect 13414 14458 13474 14658
rect 13651 14458 13711 14858
rect 13769 14458 13829 14858
rect 13887 14458 13947 14858
rect 14124 14458 14184 14858
rect 14242 14458 14302 14858
rect 14360 14458 14420 14858
rect 14478 14458 14538 14858
rect 14596 14458 14656 14858
rect 14714 14458 14774 14858
rect 14945 14458 15005 14858
rect 15063 14458 15123 14858
rect 15181 14458 15241 14858
rect 15386 14458 15446 14658
rect 15504 14458 15564 14658
rect 15622 14458 15682 14658
rect 16322 14458 16382 14658
rect 16440 14458 16500 14658
rect 16558 14458 16618 14658
rect 16795 14458 16855 14858
rect 16913 14458 16973 14858
rect 17031 14458 17091 14858
rect 17268 14458 17328 14858
rect 17386 14458 17446 14858
rect 17504 14458 17564 14858
rect 17622 14458 17682 14858
rect 17740 14458 17800 14858
rect 17858 14458 17918 14858
rect 18089 14458 18149 14858
rect 18207 14458 18267 14858
rect 18325 14458 18385 14858
rect 18530 14458 18590 14658
rect 18648 14458 18708 14658
rect 18766 14458 18826 14658
rect 19454 14454 19514 14654
rect 19572 14454 19632 14654
rect 19690 14454 19750 14654
rect 19927 14454 19987 14854
rect 20045 14454 20105 14854
rect 20163 14454 20223 14854
rect 20400 14454 20460 14854
rect 20518 14454 20578 14854
rect 20636 14454 20696 14854
rect 20754 14454 20814 14854
rect 20872 14454 20932 14854
rect 20990 14454 21050 14854
rect 21221 14454 21281 14854
rect 21339 14454 21399 14854
rect 21457 14454 21517 14854
rect 21662 14454 21722 14654
rect 21780 14454 21840 14654
rect 21898 14454 21958 14654
rect 22598 14454 22658 14654
rect 22716 14454 22776 14654
rect 22834 14454 22894 14654
rect 23071 14454 23131 14854
rect 23189 14454 23249 14854
rect 23307 14454 23367 14854
rect 23544 14454 23604 14854
rect 23662 14454 23722 14854
rect 23780 14454 23840 14854
rect 23898 14454 23958 14854
rect 24016 14454 24076 14854
rect 24134 14454 24194 14854
rect 24365 14454 24425 14854
rect 24483 14454 24543 14854
rect 24601 14454 24661 14854
rect 58386 16462 58446 16662
rect 58504 16462 58564 16662
rect 58622 16462 58682 16662
rect 58869 16462 58929 16862
rect 58987 16462 59047 16862
rect 59105 16462 59165 16862
rect 59223 16462 59283 16862
rect 59341 16462 59401 16862
rect 59459 16462 59519 16862
rect 59707 16462 59767 16662
rect 59825 16462 59885 16662
rect 59943 16462 60003 16662
rect 60284 16462 60344 16662
rect 60402 16462 60462 16662
rect 60520 16462 60580 16662
rect 60767 16462 60827 16862
rect 60885 16462 60945 16862
rect 61003 16462 61063 16862
rect 61121 16462 61181 16862
rect 61239 16462 61299 16862
rect 61357 16462 61417 16862
rect 70513 16958 70913 17018
rect 61605 16462 61665 16662
rect 61723 16462 61783 16662
rect 61841 16462 61901 16662
rect 54311 15766 54371 16166
rect 54429 15766 54489 16166
rect 54547 15766 54607 16166
rect 54665 15766 54725 16166
rect 54783 15766 54843 16166
rect 54901 15766 54961 16166
rect 55853 15472 55913 15672
rect 55971 15472 56031 15672
rect 56089 15472 56149 15672
rect 56207 15472 56267 15672
rect 56325 15472 56385 15672
rect 56443 15472 56503 15672
rect 56561 15472 56621 15672
rect 56679 15472 56739 15672
rect 56797 15472 56857 15672
rect 58926 15769 58986 16169
rect 59044 15769 59104 16169
rect 59162 15769 59222 16169
rect 59280 15769 59340 16169
rect 59398 15769 59458 16169
rect 59516 15769 59576 16169
rect 70513 16840 70913 16900
rect 70713 16603 70913 16663
rect 70713 16485 70913 16545
rect 70713 16367 70913 16427
rect 60824 15769 60884 16169
rect 60942 15769 61002 16169
rect 61060 15769 61120 16169
rect 61178 15769 61238 16169
rect 61296 15769 61356 16169
rect 61414 15769 61474 16169
rect 70709 15679 70909 15739
rect 62366 15475 62426 15675
rect 62484 15475 62544 15675
rect 62602 15475 62662 15675
rect 62720 15475 62780 15675
rect 62838 15475 62898 15675
rect 62956 15475 63016 15675
rect 63074 15475 63134 15675
rect 63192 15475 63252 15675
rect 63310 15475 63370 15675
rect 70709 15561 70909 15621
rect 24806 14454 24866 14654
rect 24924 14454 24984 14654
rect 25042 14454 25102 14654
rect 70709 15443 70909 15503
rect 70509 15238 70909 15298
rect 70509 15120 70909 15180
rect 70509 15002 70909 15062
rect 70509 14771 70909 14831
rect 70509 14653 70909 14713
rect 70509 14535 70909 14595
rect 70509 14417 70909 14477
rect 70509 14299 70909 14359
rect 70509 14181 70909 14241
rect 70509 13944 70909 14004
rect 70509 13826 70909 13886
rect 70509 13708 70909 13768
rect 70709 13471 70909 13531
rect 70709 13353 70909 13413
rect 70709 13235 70909 13295
rect 30154 13062 30354 13122
rect 30154 12944 30354 13004
rect 30154 12826 30354 12886
rect 29954 12578 30354 12638
rect 30647 12635 31047 12695
rect 29954 12460 30354 12520
rect 30647 12517 31047 12577
rect 70709 12535 70909 12595
rect 29954 12342 30354 12402
rect 30647 12399 31047 12459
rect 556 11724 616 11924
rect 674 11724 734 11924
rect 792 11724 852 11924
rect 1029 11724 1089 12124
rect 1147 11724 1207 12124
rect 1265 11724 1325 12124
rect 1502 11724 1562 12124
rect 1620 11724 1680 12124
rect 1738 11724 1798 12124
rect 1856 11724 1916 12124
rect 1974 11724 2034 12124
rect 2092 11724 2152 12124
rect 2323 11724 2383 12124
rect 2441 11724 2501 12124
rect 2559 11724 2619 12124
rect 2764 11724 2824 11924
rect 2882 11724 2942 11924
rect 3000 11724 3060 11924
rect 3700 11724 3760 11924
rect 3818 11724 3878 11924
rect 3936 11724 3996 11924
rect 4173 11724 4233 12124
rect 4291 11724 4351 12124
rect 4409 11724 4469 12124
rect 4646 11724 4706 12124
rect 4764 11724 4824 12124
rect 4882 11724 4942 12124
rect 5000 11724 5060 12124
rect 5118 11724 5178 12124
rect 5236 11724 5296 12124
rect 5467 11724 5527 12124
rect 5585 11724 5645 12124
rect 5703 11724 5763 12124
rect 5908 11724 5968 11924
rect 6026 11724 6086 11924
rect 6144 11724 6204 11924
rect 6832 11720 6892 11920
rect 6950 11720 7010 11920
rect 7068 11720 7128 11920
rect 7305 11720 7365 12120
rect 7423 11720 7483 12120
rect 7541 11720 7601 12120
rect 7778 11720 7838 12120
rect 7896 11720 7956 12120
rect 8014 11720 8074 12120
rect 8132 11720 8192 12120
rect 8250 11720 8310 12120
rect 8368 11720 8428 12120
rect 8599 11720 8659 12120
rect 8717 11720 8777 12120
rect 8835 11720 8895 12120
rect 9040 11720 9100 11920
rect 9158 11720 9218 11920
rect 9276 11720 9336 11920
rect 9976 11720 10036 11920
rect 10094 11720 10154 11920
rect 10212 11720 10272 11920
rect 10449 11720 10509 12120
rect 10567 11720 10627 12120
rect 10685 11720 10745 12120
rect 10922 11720 10982 12120
rect 11040 11720 11100 12120
rect 11158 11720 11218 12120
rect 11276 11720 11336 12120
rect 11394 11720 11454 12120
rect 11512 11720 11572 12120
rect 11743 11720 11803 12120
rect 11861 11720 11921 12120
rect 11979 11720 12039 12120
rect 12184 11720 12244 11920
rect 12302 11720 12362 11920
rect 12420 11720 12480 11920
rect 13178 11724 13238 11924
rect 13296 11724 13356 11924
rect 13414 11724 13474 11924
rect 13651 11724 13711 12124
rect 13769 11724 13829 12124
rect 13887 11724 13947 12124
rect 14124 11724 14184 12124
rect 14242 11724 14302 12124
rect 14360 11724 14420 12124
rect 14478 11724 14538 12124
rect 14596 11724 14656 12124
rect 14714 11724 14774 12124
rect 14945 11724 15005 12124
rect 15063 11724 15123 12124
rect 15181 11724 15241 12124
rect 15386 11724 15446 11924
rect 15504 11724 15564 11924
rect 15622 11724 15682 11924
rect 16322 11724 16382 11924
rect 16440 11724 16500 11924
rect 16558 11724 16618 11924
rect 16795 11724 16855 12124
rect 16913 11724 16973 12124
rect 17031 11724 17091 12124
rect 17268 11724 17328 12124
rect 17386 11724 17446 12124
rect 17504 11724 17564 12124
rect 17622 11724 17682 12124
rect 17740 11724 17800 12124
rect 17858 11724 17918 12124
rect 18089 11724 18149 12124
rect 18207 11724 18267 12124
rect 18325 11724 18385 12124
rect 18530 11724 18590 11924
rect 18648 11724 18708 11924
rect 18766 11724 18826 11924
rect 19454 11720 19514 11920
rect 19572 11720 19632 11920
rect 19690 11720 19750 11920
rect 19927 11720 19987 12120
rect 20045 11720 20105 12120
rect 20163 11720 20223 12120
rect 20400 11720 20460 12120
rect 20518 11720 20578 12120
rect 20636 11720 20696 12120
rect 20754 11720 20814 12120
rect 20872 11720 20932 12120
rect 20990 11720 21050 12120
rect 21221 11720 21281 12120
rect 21339 11720 21399 12120
rect 21457 11720 21517 12120
rect 21662 11720 21722 11920
rect 21780 11720 21840 11920
rect 21898 11720 21958 11920
rect 22598 11720 22658 11920
rect 22716 11720 22776 11920
rect 22834 11720 22894 11920
rect 23071 11720 23131 12120
rect 23189 11720 23249 12120
rect 23307 11720 23367 12120
rect 23544 11720 23604 12120
rect 23662 11720 23722 12120
rect 23780 11720 23840 12120
rect 23898 11720 23958 12120
rect 24016 11720 24076 12120
rect 24134 11720 24194 12120
rect 24365 11720 24425 12120
rect 24483 11720 24543 12120
rect 24601 11720 24661 12120
rect 29954 12224 30354 12284
rect 29954 12106 30354 12166
rect 29954 11988 30354 12048
rect 30647 12281 31047 12341
rect 70709 12417 70909 12477
rect 70709 12299 70909 12359
rect 30647 12163 31047 12223
rect 30647 12045 31047 12105
rect 24806 11720 24866 11920
rect 24924 11720 24984 11920
rect 25042 11720 25102 11920
rect 41616 11949 41676 12149
rect 41734 11949 41794 12149
rect 41852 11949 41912 12149
rect 41970 11949 42030 12149
rect 42088 11949 42148 12149
rect 42206 11949 42266 12149
rect 42324 11949 42384 12149
rect 42442 11949 42502 12149
rect 42560 11949 42620 12149
rect 30154 11741 30354 11801
rect 48165 11948 48225 12148
rect 48283 11948 48343 12148
rect 48401 11948 48461 12148
rect 48519 11948 48579 12148
rect 48637 11948 48697 12148
rect 48755 11948 48815 12148
rect 48873 11948 48933 12148
rect 48991 11948 49051 12148
rect 49109 11948 49169 12148
rect 54819 11969 54879 12169
rect 54937 11969 54997 12169
rect 55055 11969 55115 12169
rect 55173 11969 55233 12169
rect 55291 11969 55351 12169
rect 55409 11969 55469 12169
rect 55527 11969 55587 12169
rect 55645 11969 55705 12169
rect 55763 11969 55823 12169
rect 70509 12094 70909 12154
rect 30154 11623 30354 11683
rect 30154 11505 30354 11565
rect 63472 11802 63532 12002
rect 63590 11802 63650 12002
rect 63708 11802 63768 12002
rect 63826 11802 63886 12002
rect 63944 11802 64004 12002
rect 64062 11802 64122 12002
rect 64180 11802 64240 12002
rect 64298 11802 64358 12002
rect 64416 11802 64476 12002
rect 70509 11976 70909 12036
rect 70509 11858 70909 11918
rect 65280 11397 65340 11597
rect 65398 11397 65458 11597
rect 65516 11397 65576 11597
rect 65764 11397 65824 11797
rect 65882 11397 65942 11797
rect 66000 11397 66060 11797
rect 66118 11397 66178 11797
rect 66236 11397 66296 11797
rect 66354 11397 66414 11797
rect 66601 11397 66661 11597
rect 66719 11397 66779 11597
rect 66837 11397 66897 11597
rect 70509 11627 70909 11687
rect 67073 11394 67133 11594
rect 67191 11394 67251 11594
rect 67309 11394 67369 11594
rect 67427 11394 67487 11594
rect 67545 11394 67605 11594
rect 67663 11394 67723 11594
rect 67781 11394 67841 11594
rect 67899 11394 67959 11594
rect 68017 11394 68077 11594
rect 70509 11509 70909 11569
rect 30152 10994 30352 11054
rect 30152 10876 30352 10936
rect 30152 10758 30352 10818
rect 29952 10510 30352 10570
rect 30645 10567 31045 10627
rect 29952 10392 30352 10452
rect 30645 10449 31045 10509
rect 29952 10274 30352 10334
rect 30645 10331 31045 10391
rect 29952 10156 30352 10216
rect 29952 10038 30352 10098
rect 29952 9920 30352 9980
rect 30645 10213 31045 10273
rect 30645 10095 31045 10155
rect 30645 9977 31045 10037
rect 34952 10049 35012 10249
rect 35070 10049 35130 10249
rect 35188 10049 35248 10249
rect 35306 10049 35366 10249
rect 35424 10049 35484 10249
rect 35542 10049 35602 10249
rect 35660 10049 35720 10249
rect 35778 10049 35838 10249
rect 35896 10049 35956 10249
rect 65707 10704 65767 11104
rect 65825 10704 65885 11104
rect 65943 10704 66003 11104
rect 66061 10704 66121 11104
rect 66179 10704 66239 11104
rect 66297 10704 66357 11104
rect 70509 11391 70909 11451
rect 70509 11273 70909 11333
rect 70509 11155 70909 11215
rect 70509 11037 70909 11097
rect 70509 10800 70909 10860
rect 70509 10682 70909 10742
rect 70509 10564 70909 10624
rect 30152 9673 30352 9733
rect 30152 9555 30352 9615
rect 566 8992 626 9192
rect 684 8992 744 9192
rect 802 8992 862 9192
rect 1039 8992 1099 9392
rect 1157 8992 1217 9392
rect 1275 8992 1335 9392
rect 1512 8992 1572 9392
rect 1630 8992 1690 9392
rect 1748 8992 1808 9392
rect 1866 8992 1926 9392
rect 1984 8992 2044 9392
rect 2102 8992 2162 9392
rect 2333 8992 2393 9392
rect 2451 8992 2511 9392
rect 2569 8992 2629 9392
rect 2774 8992 2834 9192
rect 2892 8992 2952 9192
rect 3010 8992 3070 9192
rect 3710 8992 3770 9192
rect 3828 8992 3888 9192
rect 3946 8992 4006 9192
rect 4183 8992 4243 9392
rect 4301 8992 4361 9392
rect 4419 8992 4479 9392
rect 4656 8992 4716 9392
rect 4774 8992 4834 9392
rect 4892 8992 4952 9392
rect 5010 8992 5070 9392
rect 5128 8992 5188 9392
rect 5246 8992 5306 9392
rect 5477 8992 5537 9392
rect 5595 8992 5655 9392
rect 5713 8992 5773 9392
rect 5918 8992 5978 9192
rect 6036 8992 6096 9192
rect 6154 8992 6214 9192
rect 6842 8988 6902 9188
rect 6960 8988 7020 9188
rect 7078 8988 7138 9188
rect 7315 8988 7375 9388
rect 7433 8988 7493 9388
rect 7551 8988 7611 9388
rect 7788 8988 7848 9388
rect 7906 8988 7966 9388
rect 8024 8988 8084 9388
rect 8142 8988 8202 9388
rect 8260 8988 8320 9388
rect 8378 8988 8438 9388
rect 8609 8988 8669 9388
rect 8727 8988 8787 9388
rect 8845 8988 8905 9388
rect 9050 8988 9110 9188
rect 9168 8988 9228 9188
rect 9286 8988 9346 9188
rect 9986 8988 10046 9188
rect 10104 8988 10164 9188
rect 10222 8988 10282 9188
rect 10459 8988 10519 9388
rect 10577 8988 10637 9388
rect 10695 8988 10755 9388
rect 10932 8988 10992 9388
rect 11050 8988 11110 9388
rect 11168 8988 11228 9388
rect 11286 8988 11346 9388
rect 11404 8988 11464 9388
rect 11522 8988 11582 9388
rect 11753 8988 11813 9388
rect 11871 8988 11931 9388
rect 11989 8988 12049 9388
rect 12194 8988 12254 9188
rect 12312 8988 12372 9188
rect 12430 8988 12490 9188
rect 13188 8992 13248 9192
rect 13306 8992 13366 9192
rect 13424 8992 13484 9192
rect 13661 8992 13721 9392
rect 13779 8992 13839 9392
rect 13897 8992 13957 9392
rect 14134 8992 14194 9392
rect 14252 8992 14312 9392
rect 14370 8992 14430 9392
rect 14488 8992 14548 9392
rect 14606 8992 14666 9392
rect 14724 8992 14784 9392
rect 14955 8992 15015 9392
rect 15073 8992 15133 9392
rect 15191 8992 15251 9392
rect 15396 8992 15456 9192
rect 15514 8992 15574 9192
rect 15632 8992 15692 9192
rect 16332 8992 16392 9192
rect 16450 8992 16510 9192
rect 16568 8992 16628 9192
rect 16805 8992 16865 9392
rect 16923 8992 16983 9392
rect 17041 8992 17101 9392
rect 17278 8992 17338 9392
rect 17396 8992 17456 9392
rect 17514 8992 17574 9392
rect 17632 8992 17692 9392
rect 17750 8992 17810 9392
rect 17868 8992 17928 9392
rect 18099 8992 18159 9392
rect 18217 8992 18277 9392
rect 18335 8992 18395 9392
rect 30152 9437 30352 9497
rect 37842 9782 37902 9982
rect 37960 9782 38020 9982
rect 38078 9782 38138 9982
rect 38196 9782 38256 9982
rect 38314 9782 38374 9982
rect 38432 9782 38492 9982
rect 38550 9782 38610 9982
rect 38668 9782 38728 9982
rect 38786 9782 38846 9982
rect 40167 9654 40227 10054
rect 40285 9654 40345 10054
rect 40403 9654 40463 10054
rect 40521 9654 40581 10054
rect 40639 9654 40699 10054
rect 40757 9654 40817 10054
rect 41309 9658 41369 10058
rect 41427 9658 41487 10058
rect 41545 9658 41605 10058
rect 41663 9658 41723 10058
rect 41781 9658 41841 10058
rect 41899 9658 41959 10058
rect 44391 9870 44451 10070
rect 44509 9870 44569 10070
rect 44627 9870 44687 10070
rect 44745 9870 44805 10070
rect 44863 9870 44923 10070
rect 44981 9870 45041 10070
rect 45099 9870 45159 10070
rect 45217 9870 45277 10070
rect 45335 9870 45395 10070
rect 18540 8992 18600 9192
rect 18658 8992 18718 9192
rect 18776 8992 18836 9192
rect 19464 8988 19524 9188
rect 19582 8988 19642 9188
rect 19700 8988 19760 9188
rect 19937 8988 19997 9388
rect 20055 8988 20115 9388
rect 20173 8988 20233 9388
rect 20410 8988 20470 9388
rect 20528 8988 20588 9388
rect 20646 8988 20706 9388
rect 20764 8988 20824 9388
rect 20882 8988 20942 9388
rect 21000 8988 21060 9388
rect 21231 8988 21291 9388
rect 21349 8988 21409 9388
rect 21467 8988 21527 9388
rect 21672 8988 21732 9188
rect 21790 8988 21850 9188
rect 21908 8988 21968 9188
rect 22608 8988 22668 9188
rect 22726 8988 22786 9188
rect 22844 8988 22904 9188
rect 23081 8988 23141 9388
rect 23199 8988 23259 9388
rect 23317 8988 23377 9388
rect 23554 8988 23614 9388
rect 23672 8988 23732 9388
rect 23790 8988 23850 9388
rect 23908 8988 23968 9388
rect 24026 8988 24086 9388
rect 24144 8988 24204 9388
rect 24375 8988 24435 9388
rect 24493 8988 24553 9388
rect 24611 8988 24671 9388
rect 24816 8988 24876 9188
rect 24934 8988 24994 9188
rect 25052 8988 25112 9188
rect 46716 9742 46776 10142
rect 46834 9742 46894 10142
rect 46952 9742 47012 10142
rect 47070 9742 47130 10142
rect 47188 9742 47248 10142
rect 47306 9742 47366 10142
rect 47858 9746 47918 10146
rect 47976 9746 48036 10146
rect 48094 9746 48154 10146
rect 48212 9746 48272 10146
rect 48330 9746 48390 10146
rect 48448 9746 48508 10146
rect 51045 9802 51105 10002
rect 51163 9802 51223 10002
rect 51281 9802 51341 10002
rect 51399 9802 51459 10002
rect 51517 9802 51577 10002
rect 51635 9802 51695 10002
rect 51753 9802 51813 10002
rect 51871 9802 51931 10002
rect 51989 9802 52049 10002
rect 40596 9071 40656 9271
rect 40714 9071 40774 9271
rect 40832 9071 40892 9271
rect 41738 9075 41798 9275
rect 41856 9075 41916 9275
rect 41974 9075 42034 9275
rect 53370 9674 53430 10074
rect 53488 9674 53548 10074
rect 53606 9674 53666 10074
rect 53724 9674 53784 10074
rect 53842 9674 53902 10074
rect 53960 9674 54020 10074
rect 54512 9678 54572 10078
rect 54630 9678 54690 10078
rect 54748 9678 54808 10078
rect 54866 9678 54926 10078
rect 54984 9678 55044 10078
rect 55102 9678 55162 10078
rect 57670 9870 57730 10070
rect 57788 9870 57848 10070
rect 57906 9870 57966 10070
rect 58024 9870 58084 10070
rect 58142 9870 58202 10070
rect 58260 9870 58320 10070
rect 58378 9870 58438 10070
rect 58496 9870 58556 10070
rect 58614 9870 58674 10070
rect 47145 9159 47205 9359
rect 47263 9159 47323 9359
rect 47381 9159 47441 9359
rect 48287 9163 48347 9363
rect 48405 9163 48465 9363
rect 48523 9163 48583 9363
rect 59995 9742 60055 10142
rect 60113 9742 60173 10142
rect 60231 9742 60291 10142
rect 60349 9742 60409 10142
rect 60467 9742 60527 10142
rect 60585 9742 60645 10142
rect 61137 9746 61197 10146
rect 61255 9746 61315 10146
rect 61373 9746 61433 10146
rect 61491 9746 61551 10146
rect 61609 9746 61669 10146
rect 61727 9746 61787 10146
rect 70709 10327 70909 10387
rect 70709 10209 70909 10269
rect 70709 10091 70909 10151
rect 53799 9091 53859 9291
rect 53917 9091 53977 9291
rect 54035 9091 54095 9291
rect 54941 9095 55001 9295
rect 55059 9095 55119 9295
rect 55177 9095 55237 9295
rect 60424 9159 60484 9359
rect 60542 9159 60602 9359
rect 60660 9159 60720 9359
rect 61566 9163 61626 9363
rect 61684 9163 61744 9363
rect 61802 9163 61862 9363
rect 63467 9231 63527 9431
rect 63585 9231 63645 9431
rect 63703 9231 63763 9431
rect 63821 9231 63881 9431
rect 63939 9231 63999 9431
rect 64057 9231 64117 9431
rect 64175 9231 64235 9431
rect 64293 9231 64353 9431
rect 64411 9231 64471 9431
rect 70713 9333 70913 9393
rect 30154 8925 30354 8985
rect 30154 8807 30354 8867
rect 70713 9215 70913 9275
rect 70713 9097 70913 9157
rect 30154 8689 30354 8749
rect 29954 8441 30354 8501
rect 30647 8498 31047 8558
rect 70513 8892 70913 8952
rect 70513 8774 70913 8834
rect 70513 8656 70913 8716
rect 29954 8323 30354 8383
rect 30647 8380 31047 8440
rect 29954 8205 30354 8265
rect 30647 8262 31047 8322
rect 29954 8087 30354 8147
rect 29954 7969 30354 8029
rect 29954 7851 30354 7911
rect 30647 8144 31047 8204
rect 37856 8132 37916 8332
rect 37974 8132 38034 8332
rect 38092 8132 38152 8332
rect 38210 8132 38270 8332
rect 38328 8132 38388 8332
rect 38446 8132 38506 8332
rect 38564 8132 38624 8332
rect 38682 8132 38742 8332
rect 38800 8132 38860 8332
rect 44405 8220 44465 8420
rect 44523 8220 44583 8420
rect 44641 8220 44701 8420
rect 44759 8220 44819 8420
rect 44877 8220 44937 8420
rect 44995 8220 45055 8420
rect 45113 8220 45173 8420
rect 45231 8220 45291 8420
rect 45349 8220 45409 8420
rect 30647 8026 31047 8086
rect 30647 7908 31047 7968
rect 51059 8152 51119 8352
rect 51177 8152 51237 8352
rect 51295 8152 51355 8352
rect 51413 8152 51473 8352
rect 51531 8152 51591 8352
rect 51649 8152 51709 8352
rect 51767 8152 51827 8352
rect 51885 8152 51945 8352
rect 52003 8152 52063 8352
rect 57684 8220 57744 8420
rect 57802 8220 57862 8420
rect 57920 8220 57980 8420
rect 58038 8220 58098 8420
rect 58156 8220 58216 8420
rect 58274 8220 58334 8420
rect 58392 8220 58452 8420
rect 58510 8220 58570 8420
rect 58628 8220 58688 8420
rect 70513 8425 70913 8485
rect 70513 8307 70913 8367
rect 30154 7604 30354 7664
rect 30154 7486 30354 7546
rect 34944 7464 35004 7664
rect 35062 7464 35122 7664
rect 35180 7464 35240 7664
rect 35298 7464 35358 7664
rect 35416 7464 35476 7664
rect 35534 7464 35594 7664
rect 35652 7464 35712 7664
rect 35770 7464 35830 7664
rect 35888 7464 35948 7664
rect 30154 7368 30354 7428
rect 39320 7515 39380 7715
rect 39438 7515 39498 7715
rect 39556 7515 39616 7715
rect 39804 7515 39864 7915
rect 39922 7515 39982 7915
rect 40040 7515 40100 7915
rect 40158 7515 40218 7915
rect 40276 7515 40336 7915
rect 40394 7515 40454 7915
rect 40641 7515 40701 7715
rect 40759 7515 40819 7715
rect 40877 7515 40937 7715
rect 41218 7515 41278 7715
rect 41336 7515 41396 7715
rect 41454 7515 41514 7715
rect 41702 7515 41762 7915
rect 41820 7515 41880 7915
rect 41938 7515 41998 7915
rect 42056 7515 42116 7915
rect 42174 7515 42234 7915
rect 42292 7515 42352 7915
rect 42539 7515 42599 7715
rect 42657 7515 42717 7715
rect 42775 7515 42835 7715
rect 30152 6857 30352 6917
rect 30152 6739 30352 6799
rect 30152 6621 30352 6681
rect 3175 6357 3235 6557
rect 3293 6357 3353 6557
rect 3411 6357 3471 6557
rect 3913 6357 3973 6557
rect 4031 6357 4091 6557
rect 4149 6357 4209 6557
rect 4651 6357 4711 6557
rect 4769 6357 4829 6557
rect 4887 6357 4947 6557
rect 5389 6357 5449 6557
rect 5507 6357 5567 6557
rect 5625 6357 5685 6557
rect 6129 6357 6189 6557
rect 6247 6357 6307 6557
rect 6365 6357 6425 6557
rect 6871 6359 6931 6559
rect 6989 6359 7049 6559
rect 7107 6359 7167 6559
rect 7609 6363 7669 6563
rect 7727 6363 7787 6563
rect 7845 6363 7905 6563
rect 8347 6359 8407 6559
rect 8465 6359 8525 6559
rect 8583 6359 8643 6559
rect 9279 6047 9339 6247
rect 9397 6047 9457 6247
rect 9515 6047 9575 6247
rect 9762 6047 9822 6447
rect 9880 6047 9940 6447
rect 9998 6047 10058 6447
rect 10116 6047 10176 6447
rect 10234 6047 10294 6447
rect 10352 6047 10412 6447
rect 10600 6047 10660 6247
rect 10718 6047 10778 6247
rect 10836 6047 10896 6247
rect 11347 6045 11407 6245
rect 11465 6045 11525 6245
rect 11583 6045 11643 6245
rect 11830 6045 11890 6445
rect 11948 6045 12008 6445
rect 12066 6045 12126 6445
rect 12184 6045 12244 6445
rect 12302 6045 12362 6445
rect 12420 6045 12480 6445
rect 12668 6045 12728 6245
rect 12786 6045 12846 6245
rect 12904 6045 12964 6245
rect 13416 6047 13476 6247
rect 13534 6047 13594 6247
rect 13652 6047 13712 6247
rect 13899 6047 13959 6447
rect 14017 6047 14077 6447
rect 14135 6047 14195 6447
rect 14253 6047 14313 6447
rect 14371 6047 14431 6447
rect 14489 6047 14549 6447
rect 14737 6047 14797 6247
rect 14855 6047 14915 6247
rect 14973 6047 15033 6247
rect 9819 5354 9879 5754
rect 9937 5354 9997 5754
rect 10055 5354 10115 5754
rect 10173 5354 10233 5754
rect 10291 5354 10351 5754
rect 10409 5354 10469 5754
rect 15484 6045 15544 6245
rect 15602 6045 15662 6245
rect 15720 6045 15780 6245
rect 15967 6045 16027 6445
rect 16085 6045 16145 6445
rect 16203 6045 16263 6445
rect 16321 6045 16381 6445
rect 16439 6045 16499 6445
rect 16557 6045 16617 6445
rect 16805 6045 16865 6245
rect 16923 6045 16983 6245
rect 17041 6045 17101 6245
rect 17553 6045 17613 6245
rect 17671 6045 17731 6245
rect 17789 6045 17849 6245
rect 18036 6045 18096 6445
rect 18154 6045 18214 6445
rect 18272 6045 18332 6445
rect 18390 6045 18450 6445
rect 18508 6045 18568 6445
rect 18626 6045 18686 6445
rect 18874 6045 18934 6245
rect 18992 6045 19052 6245
rect 19110 6045 19170 6245
rect 11887 5352 11947 5752
rect 12005 5352 12065 5752
rect 12123 5352 12183 5752
rect 12241 5352 12301 5752
rect 12359 5352 12419 5752
rect 12477 5352 12537 5752
rect 13956 5354 14016 5754
rect 14074 5354 14134 5754
rect 14192 5354 14252 5754
rect 14310 5354 14370 5754
rect 14428 5354 14488 5754
rect 14546 5354 14606 5754
rect 16024 5352 16084 5752
rect 16142 5352 16202 5752
rect 16260 5352 16320 5752
rect 16378 5352 16438 5752
rect 16496 5352 16556 5752
rect 16614 5352 16674 5752
rect 19621 6043 19681 6243
rect 19739 6043 19799 6243
rect 19857 6043 19917 6243
rect 20104 6043 20164 6443
rect 20222 6043 20282 6443
rect 20340 6043 20400 6443
rect 20458 6043 20518 6443
rect 20576 6043 20636 6443
rect 20694 6043 20754 6443
rect 20942 6043 21002 6243
rect 21060 6043 21120 6243
rect 21178 6043 21238 6243
rect 21690 6045 21750 6245
rect 21808 6045 21868 6245
rect 21926 6045 21986 6245
rect 22173 6045 22233 6445
rect 22291 6045 22351 6445
rect 22409 6045 22469 6445
rect 22527 6045 22587 6445
rect 22645 6045 22705 6445
rect 22763 6045 22823 6445
rect 23011 6045 23071 6245
rect 23129 6045 23189 6245
rect 23247 6045 23307 6245
rect 18093 5352 18153 5752
rect 18211 5352 18271 5752
rect 18329 5352 18389 5752
rect 18447 5352 18507 5752
rect 18565 5352 18625 5752
rect 18683 5352 18743 5752
rect 23758 6043 23818 6243
rect 23876 6043 23936 6243
rect 23994 6043 24054 6243
rect 24241 6043 24301 6443
rect 24359 6043 24419 6443
rect 24477 6043 24537 6443
rect 24595 6043 24655 6443
rect 24713 6043 24773 6443
rect 24831 6043 24891 6443
rect 37851 6528 37911 6728
rect 37969 6528 38029 6728
rect 38087 6528 38147 6728
rect 38205 6528 38265 6728
rect 38323 6528 38383 6728
rect 38441 6528 38501 6728
rect 38559 6528 38619 6728
rect 38677 6528 38737 6728
rect 38795 6528 38855 6728
rect 39747 6822 39807 7222
rect 39865 6822 39925 7222
rect 39983 6822 40043 7222
rect 40101 6822 40161 7222
rect 40219 6822 40279 7222
rect 40337 6822 40397 7222
rect 29952 6373 30352 6433
rect 30645 6430 31045 6490
rect 25079 6043 25139 6243
rect 25197 6043 25257 6243
rect 25315 6043 25375 6243
rect 29952 6255 30352 6315
rect 30645 6312 31045 6372
rect 45869 7603 45929 7803
rect 45987 7603 46047 7803
rect 46105 7603 46165 7803
rect 46353 7603 46413 8003
rect 46471 7603 46531 8003
rect 46589 7603 46649 8003
rect 46707 7603 46767 8003
rect 46825 7603 46885 8003
rect 46943 7603 47003 8003
rect 47190 7603 47250 7803
rect 47308 7603 47368 7803
rect 47426 7603 47486 7803
rect 47767 7603 47827 7803
rect 47885 7603 47945 7803
rect 48003 7603 48063 7803
rect 48251 7603 48311 8003
rect 48369 7603 48429 8003
rect 48487 7603 48547 8003
rect 48605 7603 48665 8003
rect 48723 7603 48783 8003
rect 48841 7603 48901 8003
rect 70513 8189 70913 8249
rect 70513 8071 70913 8131
rect 49088 7603 49148 7803
rect 49206 7603 49266 7803
rect 49324 7603 49384 7803
rect 41645 6822 41705 7222
rect 41763 6822 41823 7222
rect 41881 6822 41941 7222
rect 41999 6822 42059 7222
rect 42117 6822 42177 7222
rect 42235 6822 42295 7222
rect 44400 6616 44460 6816
rect 44518 6616 44578 6816
rect 44636 6616 44696 6816
rect 44754 6616 44814 6816
rect 44872 6616 44932 6816
rect 44990 6616 45050 6816
rect 45108 6616 45168 6816
rect 45226 6616 45286 6816
rect 45344 6616 45404 6816
rect 46296 6910 46356 7310
rect 46414 6910 46474 7310
rect 46532 6910 46592 7310
rect 46650 6910 46710 7310
rect 46768 6910 46828 7310
rect 46886 6910 46946 7310
rect 29952 6137 30352 6197
rect 30645 6194 31045 6254
rect 20161 5350 20221 5750
rect 20279 5350 20339 5750
rect 20397 5350 20457 5750
rect 20515 5350 20575 5750
rect 20633 5350 20693 5750
rect 20751 5350 20811 5750
rect 22230 5352 22290 5752
rect 22348 5352 22408 5752
rect 22466 5352 22526 5752
rect 22584 5352 22644 5752
rect 22702 5352 22762 5752
rect 22820 5352 22880 5752
rect 24298 5350 24358 5750
rect 24416 5350 24476 5750
rect 24534 5350 24594 5750
rect 24652 5350 24712 5750
rect 24770 5350 24830 5750
rect 24888 5350 24948 5750
rect 29952 6019 30352 6079
rect 29952 5901 30352 5961
rect 29952 5783 30352 5843
rect 30645 6076 31045 6136
rect 30645 5958 31045 6018
rect 30645 5840 31045 5900
rect 52523 7535 52583 7735
rect 52641 7535 52701 7735
rect 52759 7535 52819 7735
rect 53007 7535 53067 7935
rect 53125 7535 53185 7935
rect 53243 7535 53303 7935
rect 53361 7535 53421 7935
rect 53479 7535 53539 7935
rect 53597 7535 53657 7935
rect 53844 7535 53904 7735
rect 53962 7535 54022 7735
rect 54080 7535 54140 7735
rect 54421 7535 54481 7735
rect 54539 7535 54599 7735
rect 54657 7535 54717 7735
rect 54905 7535 54965 7935
rect 55023 7535 55083 7935
rect 55141 7535 55201 7935
rect 55259 7535 55319 7935
rect 55377 7535 55437 7935
rect 55495 7535 55555 7935
rect 55742 7535 55802 7735
rect 55860 7535 55920 7735
rect 55978 7535 56038 7735
rect 48194 6910 48254 7310
rect 48312 6910 48372 7310
rect 48430 6910 48490 7310
rect 48548 6910 48608 7310
rect 48666 6910 48726 7310
rect 48784 6910 48844 7310
rect 51054 6548 51114 6748
rect 51172 6548 51232 6748
rect 51290 6548 51350 6748
rect 51408 6548 51468 6748
rect 51526 6548 51586 6748
rect 51644 6548 51704 6748
rect 51762 6548 51822 6748
rect 51880 6548 51940 6748
rect 51998 6548 52058 6748
rect 52950 6842 53010 7242
rect 53068 6842 53128 7242
rect 53186 6842 53246 7242
rect 53304 6842 53364 7242
rect 53422 6842 53482 7242
rect 53540 6842 53600 7242
rect 59148 7603 59208 7803
rect 59266 7603 59326 7803
rect 59384 7603 59444 7803
rect 59632 7603 59692 8003
rect 59750 7603 59810 8003
rect 59868 7603 59928 8003
rect 59986 7603 60046 8003
rect 60104 7603 60164 8003
rect 60222 7603 60282 8003
rect 60469 7603 60529 7803
rect 60587 7603 60647 7803
rect 60705 7603 60765 7803
rect 61046 7603 61106 7803
rect 61164 7603 61224 7803
rect 61282 7603 61342 7803
rect 61530 7603 61590 8003
rect 61648 7603 61708 8003
rect 61766 7603 61826 8003
rect 61884 7603 61944 8003
rect 62002 7603 62062 8003
rect 62120 7603 62180 8003
rect 70513 7953 70913 8013
rect 70513 7835 70913 7895
rect 62367 7603 62427 7803
rect 62485 7603 62545 7803
rect 62603 7603 62663 7803
rect 54848 6842 54908 7242
rect 54966 6842 55026 7242
rect 55084 6842 55144 7242
rect 55202 6842 55262 7242
rect 55320 6842 55380 7242
rect 55438 6842 55498 7242
rect 57679 6616 57739 6816
rect 57797 6616 57857 6816
rect 57915 6616 57975 6816
rect 58033 6616 58093 6816
rect 58151 6616 58211 6816
rect 58269 6616 58329 6816
rect 58387 6616 58447 6816
rect 58505 6616 58565 6816
rect 58623 6616 58683 6816
rect 59575 6910 59635 7310
rect 59693 6910 59753 7310
rect 59811 6910 59871 7310
rect 59929 6910 59989 7310
rect 60047 6910 60107 7310
rect 60165 6910 60225 7310
rect 61473 6910 61533 7310
rect 61591 6910 61651 7310
rect 61709 6910 61769 7310
rect 61827 6910 61887 7310
rect 61945 6910 62005 7310
rect 62063 6910 62123 7310
rect 65282 7306 65342 7506
rect 65400 7306 65460 7506
rect 65518 7306 65578 7506
rect 65766 7306 65826 7706
rect 65884 7306 65944 7706
rect 66002 7306 66062 7706
rect 66120 7306 66180 7706
rect 66238 7306 66298 7706
rect 66356 7306 66416 7706
rect 70513 7598 70913 7658
rect 66603 7306 66663 7506
rect 66721 7306 66781 7506
rect 66839 7306 66899 7506
rect 67075 7303 67135 7503
rect 67193 7303 67253 7503
rect 67311 7303 67371 7503
rect 67429 7303 67489 7503
rect 67547 7303 67607 7503
rect 67665 7303 67725 7503
rect 67783 7303 67843 7503
rect 67901 7303 67961 7503
rect 68019 7303 68079 7503
rect 70513 7480 70913 7540
rect 70513 7362 70913 7422
rect 63467 6198 63527 6398
rect 63585 6198 63645 6398
rect 63703 6198 63763 6398
rect 63821 6198 63881 6398
rect 63939 6198 63999 6398
rect 64057 6198 64117 6398
rect 64175 6198 64235 6398
rect 64293 6198 64353 6398
rect 64411 6198 64471 6398
rect 65709 6613 65769 7013
rect 65827 6613 65887 7013
rect 65945 6613 66005 7013
rect 66063 6613 66123 7013
rect 66181 6613 66241 7013
rect 66299 6613 66359 7013
rect 70713 7125 70913 7185
rect 70713 7007 70913 7067
rect 70713 6889 70913 6949
rect 30152 5536 30352 5596
rect 70713 6189 70913 6249
rect 70713 6071 70913 6131
rect 70713 5953 70913 6013
rect 70513 5748 70913 5808
rect 70513 5630 70913 5690
rect 30152 5418 30352 5478
rect 70513 5512 70913 5572
rect 30152 5300 30352 5360
rect 70513 5281 70913 5341
rect 70513 5163 70913 5223
rect 70513 5045 70913 5105
rect 30152 4788 30352 4848
rect 30152 4670 30352 4730
rect 70513 4927 70913 4987
rect 70513 4809 70913 4869
rect 30152 4552 30352 4612
rect 29952 4304 30352 4364
rect 30645 4361 31045 4421
rect 29952 4186 30352 4246
rect 30645 4243 31045 4303
rect 29952 4068 30352 4128
rect 30645 4125 31045 4185
rect 34925 4186 34985 4386
rect 35043 4186 35103 4386
rect 35161 4186 35221 4386
rect 35279 4186 35339 4386
rect 35397 4186 35457 4386
rect 35515 4186 35575 4386
rect 35633 4186 35693 4386
rect 35751 4186 35811 4386
rect 35869 4186 35929 4386
rect 29952 3950 30352 4010
rect 29952 3832 30352 3892
rect 29952 3714 30352 3774
rect 30645 4007 31045 4067
rect 37834 4002 37894 4202
rect 37952 4002 38012 4202
rect 38070 4002 38130 4202
rect 38188 4002 38248 4202
rect 38306 4002 38366 4202
rect 38424 4002 38484 4202
rect 38542 4002 38602 4202
rect 38660 4002 38720 4202
rect 38778 4002 38838 4202
rect 30645 3889 31045 3949
rect 30645 3771 31045 3831
rect 40159 3874 40219 4274
rect 40277 3874 40337 4274
rect 40395 3874 40455 4274
rect 40513 3874 40573 4274
rect 40631 3874 40691 4274
rect 40749 3874 40809 4274
rect 41301 3878 41361 4278
rect 41419 3878 41479 4278
rect 41537 3878 41597 4278
rect 41655 3878 41715 4278
rect 41773 3878 41833 4278
rect 41891 3878 41951 4278
rect 70513 4691 70913 4751
rect 44385 4000 44445 4200
rect 44503 4000 44563 4200
rect 44621 4000 44681 4200
rect 44739 4000 44799 4200
rect 44857 4000 44917 4200
rect 44975 4000 45035 4200
rect 45093 4000 45153 4200
rect 45211 4000 45271 4200
rect 45329 4000 45389 4200
rect 30152 3467 30352 3527
rect 30152 3349 30352 3409
rect 46710 3872 46770 4272
rect 46828 3872 46888 4272
rect 46946 3872 47006 4272
rect 47064 3872 47124 4272
rect 47182 3872 47242 4272
rect 47300 3872 47360 4272
rect 47852 3876 47912 4276
rect 47970 3876 48030 4276
rect 48088 3876 48148 4276
rect 48206 3876 48266 4276
rect 48324 3876 48384 4276
rect 48442 3876 48502 4276
rect 51040 4001 51100 4201
rect 51158 4001 51218 4201
rect 51276 4001 51336 4201
rect 51394 4001 51454 4201
rect 51512 4001 51572 4201
rect 51630 4001 51690 4201
rect 51748 4001 51808 4201
rect 51866 4001 51926 4201
rect 51984 4001 52044 4201
rect 30152 3231 30352 3291
rect 40588 3291 40648 3491
rect 40706 3291 40766 3491
rect 40824 3291 40884 3491
rect 41730 3295 41790 3495
rect 41848 3295 41908 3495
rect 41966 3295 42026 3495
rect 53365 3873 53425 4273
rect 53483 3873 53543 4273
rect 53601 3873 53661 4273
rect 53719 3873 53779 4273
rect 53837 3873 53897 4273
rect 53955 3873 54015 4273
rect 54507 3877 54567 4277
rect 54625 3877 54685 4277
rect 54743 3877 54803 4277
rect 54861 3877 54921 4277
rect 54979 3877 55039 4277
rect 55097 3877 55157 4277
rect 63538 4278 63598 4478
rect 63656 4278 63716 4478
rect 63774 4278 63834 4478
rect 63892 4278 63952 4478
rect 64010 4278 64070 4478
rect 64128 4278 64188 4478
rect 64246 4278 64306 4478
rect 64364 4278 64424 4478
rect 64482 4278 64542 4478
rect 70513 4454 70913 4514
rect 70513 4336 70913 4396
rect 57662 4002 57722 4202
rect 57780 4002 57840 4202
rect 57898 4002 57958 4202
rect 58016 4002 58076 4202
rect 58134 4002 58194 4202
rect 58252 4002 58312 4202
rect 58370 4002 58430 4202
rect 58488 4002 58548 4202
rect 58606 4002 58666 4202
rect 47139 3289 47199 3489
rect 47257 3289 47317 3489
rect 47375 3289 47435 3489
rect 48281 3293 48341 3493
rect 48399 3293 48459 3493
rect 48517 3293 48577 3493
rect 59987 3874 60047 4274
rect 60105 3874 60165 4274
rect 60223 3874 60283 4274
rect 60341 3874 60401 4274
rect 60459 3874 60519 4274
rect 60577 3874 60637 4274
rect 61129 3878 61189 4278
rect 61247 3878 61307 4278
rect 61365 3878 61425 4278
rect 61483 3878 61543 4278
rect 61601 3878 61661 4278
rect 61719 3878 61779 4278
rect 53794 3290 53854 3490
rect 53912 3290 53972 3490
rect 54030 3290 54090 3490
rect 54936 3294 54996 3494
rect 55054 3294 55114 3494
rect 55172 3294 55232 3494
rect 65282 3811 65342 4011
rect 65400 3811 65460 4011
rect 65518 3811 65578 4011
rect 65766 3811 65826 4211
rect 65884 3811 65944 4211
rect 66002 3811 66062 4211
rect 66120 3811 66180 4211
rect 66238 3811 66298 4211
rect 66356 3811 66416 4211
rect 70513 4218 70913 4278
rect 66603 3811 66663 4011
rect 66721 3811 66781 4011
rect 66839 3811 66899 4011
rect 67075 3808 67135 4008
rect 67193 3808 67253 4008
rect 67311 3808 67371 4008
rect 67429 3808 67489 4008
rect 67547 3808 67607 4008
rect 67665 3808 67725 4008
rect 67783 3808 67843 4008
rect 67901 3808 67961 4008
rect 68019 3808 68079 4008
rect 70713 3981 70913 4041
rect 70713 3863 70913 3923
rect 60416 3291 60476 3491
rect 60534 3291 60594 3491
rect 60652 3291 60712 3491
rect 61558 3295 61618 3495
rect 61676 3295 61736 3495
rect 61794 3295 61854 3495
rect 30150 2720 30350 2780
rect 30150 2602 30350 2662
rect 65709 3118 65769 3518
rect 65827 3118 65887 3518
rect 65945 3118 66005 3518
rect 66063 3118 66123 3518
rect 66181 3118 66241 3518
rect 66299 3118 66359 3518
rect 70713 3745 70913 3805
rect 70709 3057 70909 3117
rect 70709 2939 70909 2999
rect 70709 2821 70909 2881
rect 30150 2484 30350 2544
rect 29950 2236 30350 2296
rect 30643 2293 31043 2353
rect 37848 2352 37908 2552
rect 37966 2352 38026 2552
rect 38084 2352 38144 2552
rect 38202 2352 38262 2552
rect 38320 2352 38380 2552
rect 38438 2352 38498 2552
rect 38556 2352 38616 2552
rect 38674 2352 38734 2552
rect 38792 2352 38852 2552
rect 306 1740 366 1940
rect 424 1740 484 1940
rect 542 1740 602 1940
rect 747 1740 807 2140
rect 865 1740 925 2140
rect 983 1740 1043 2140
rect 1214 1740 1274 2140
rect 1332 1740 1392 2140
rect 1450 1740 1510 2140
rect 1568 1740 1628 2140
rect 1686 1740 1746 2140
rect 1804 1740 1864 2140
rect 2041 1740 2101 2140
rect 2159 1740 2219 2140
rect 2277 1740 2337 2140
rect 2514 1740 2574 1940
rect 2632 1740 2692 1940
rect 2750 1740 2810 1940
rect 3450 1740 3510 1940
rect 3568 1740 3628 1940
rect 3686 1740 3746 1940
rect 3891 1740 3951 2140
rect 4009 1740 4069 2140
rect 4127 1740 4187 2140
rect 4358 1740 4418 2140
rect 4476 1740 4536 2140
rect 4594 1740 4654 2140
rect 4712 1740 4772 2140
rect 4830 1740 4890 2140
rect 4948 1740 5008 2140
rect 5185 1740 5245 2140
rect 5303 1740 5363 2140
rect 5421 1740 5481 2140
rect 5658 1740 5718 1940
rect 5776 1740 5836 1940
rect 5894 1740 5954 1940
rect 6582 1744 6642 1944
rect 6700 1744 6760 1944
rect 6818 1744 6878 1944
rect 7023 1744 7083 2144
rect 7141 1744 7201 2144
rect 7259 1744 7319 2144
rect 7490 1744 7550 2144
rect 7608 1744 7668 2144
rect 7726 1744 7786 2144
rect 7844 1744 7904 2144
rect 7962 1744 8022 2144
rect 8080 1744 8140 2144
rect 8317 1744 8377 2144
rect 8435 1744 8495 2144
rect 8553 1744 8613 2144
rect 8790 1744 8850 1944
rect 8908 1744 8968 1944
rect 9026 1744 9086 1944
rect 9726 1744 9786 1944
rect 9844 1744 9904 1944
rect 9962 1744 10022 1944
rect 10167 1744 10227 2144
rect 10285 1744 10345 2144
rect 10403 1744 10463 2144
rect 10634 1744 10694 2144
rect 10752 1744 10812 2144
rect 10870 1744 10930 2144
rect 10988 1744 11048 2144
rect 11106 1744 11166 2144
rect 11224 1744 11284 2144
rect 11461 1744 11521 2144
rect 11579 1744 11639 2144
rect 11697 1744 11757 2144
rect 11934 1744 11994 1944
rect 12052 1744 12112 1944
rect 12170 1744 12230 1944
rect 12928 1740 12988 1940
rect 13046 1740 13106 1940
rect 13164 1740 13224 1940
rect 13369 1740 13429 2140
rect 13487 1740 13547 2140
rect 13605 1740 13665 2140
rect 13836 1740 13896 2140
rect 13954 1740 14014 2140
rect 14072 1740 14132 2140
rect 14190 1740 14250 2140
rect 14308 1740 14368 2140
rect 14426 1740 14486 2140
rect 14663 1740 14723 2140
rect 14781 1740 14841 2140
rect 14899 1740 14959 2140
rect 15136 1740 15196 1940
rect 15254 1740 15314 1940
rect 15372 1740 15432 1940
rect 16072 1740 16132 1940
rect 16190 1740 16250 1940
rect 16308 1740 16368 1940
rect 16513 1740 16573 2140
rect 16631 1740 16691 2140
rect 16749 1740 16809 2140
rect 16980 1740 17040 2140
rect 17098 1740 17158 2140
rect 17216 1740 17276 2140
rect 17334 1740 17394 2140
rect 17452 1740 17512 2140
rect 17570 1740 17630 2140
rect 17807 1740 17867 2140
rect 17925 1740 17985 2140
rect 18043 1740 18103 2140
rect 18280 1740 18340 1940
rect 18398 1740 18458 1940
rect 18516 1740 18576 1940
rect 19204 1744 19264 1944
rect 19322 1744 19382 1944
rect 19440 1744 19500 1944
rect 19645 1744 19705 2144
rect 19763 1744 19823 2144
rect 19881 1744 19941 2144
rect 20112 1744 20172 2144
rect 20230 1744 20290 2144
rect 20348 1744 20408 2144
rect 20466 1744 20526 2144
rect 20584 1744 20644 2144
rect 20702 1744 20762 2144
rect 20939 1744 20999 2144
rect 21057 1744 21117 2144
rect 21175 1744 21235 2144
rect 21412 1744 21472 1944
rect 21530 1744 21590 1944
rect 21648 1744 21708 1944
rect 22348 1744 22408 1944
rect 22466 1744 22526 1944
rect 22584 1744 22644 1944
rect 22789 1744 22849 2144
rect 22907 1744 22967 2144
rect 23025 1744 23085 2144
rect 23256 1744 23316 2144
rect 23374 1744 23434 2144
rect 23492 1744 23552 2144
rect 23610 1744 23670 2144
rect 23728 1744 23788 2144
rect 23846 1744 23906 2144
rect 24083 1744 24143 2144
rect 24201 1744 24261 2144
rect 24319 1744 24379 2144
rect 24556 1744 24616 1944
rect 24674 1744 24734 1944
rect 24792 1744 24852 1944
rect 29950 2118 30350 2178
rect 30643 2175 31043 2235
rect 29950 2000 30350 2060
rect 30643 2057 31043 2117
rect 44399 2350 44459 2550
rect 44517 2350 44577 2550
rect 44635 2350 44695 2550
rect 44753 2350 44813 2550
rect 44871 2350 44931 2550
rect 44989 2350 45049 2550
rect 45107 2350 45167 2550
rect 45225 2350 45285 2550
rect 45343 2350 45403 2550
rect 51054 2351 51114 2551
rect 51172 2351 51232 2551
rect 51290 2351 51350 2551
rect 51408 2351 51468 2551
rect 51526 2351 51586 2551
rect 51644 2351 51704 2551
rect 51762 2351 51822 2551
rect 51880 2351 51940 2551
rect 51998 2351 52058 2551
rect 57676 2352 57736 2552
rect 57794 2352 57854 2552
rect 57912 2352 57972 2552
rect 58030 2352 58090 2552
rect 58148 2352 58208 2552
rect 58266 2352 58326 2552
rect 58384 2352 58444 2552
rect 58502 2352 58562 2552
rect 58620 2352 58680 2552
rect 70509 2616 70909 2676
rect 70509 2498 70909 2558
rect 70509 2380 70909 2440
rect 29950 1882 30350 1942
rect 29950 1764 30350 1824
rect 29950 1646 30350 1706
rect 30643 1939 31043 1999
rect 30643 1821 31043 1881
rect 30643 1703 31043 1763
rect 39312 1735 39372 1935
rect 39430 1735 39490 1935
rect 39548 1735 39608 1935
rect 39796 1735 39856 2135
rect 39914 1735 39974 2135
rect 40032 1735 40092 2135
rect 40150 1735 40210 2135
rect 40268 1735 40328 2135
rect 40386 1735 40446 2135
rect 40633 1735 40693 1935
rect 40751 1735 40811 1935
rect 40869 1735 40929 1935
rect 41210 1735 41270 1935
rect 41328 1735 41388 1935
rect 41446 1735 41506 1935
rect 41694 1735 41754 2135
rect 41812 1735 41872 2135
rect 41930 1735 41990 2135
rect 42048 1735 42108 2135
rect 42166 1735 42226 2135
rect 42284 1735 42344 2135
rect 42531 1735 42591 1935
rect 42649 1735 42709 1935
rect 42767 1735 42827 1935
rect 30150 1399 30350 1459
rect 34941 1426 35001 1626
rect 35059 1426 35119 1626
rect 35177 1426 35237 1626
rect 35295 1426 35355 1626
rect 35413 1426 35473 1626
rect 35531 1426 35591 1626
rect 35649 1426 35709 1626
rect 35767 1426 35827 1626
rect 35885 1426 35945 1626
rect 30150 1281 30350 1341
rect 30150 1163 30350 1223
rect 30152 651 30352 711
rect 30152 533 30352 593
rect 37843 748 37903 948
rect 37961 748 38021 948
rect 38079 748 38139 948
rect 38197 748 38257 948
rect 38315 748 38375 948
rect 38433 748 38493 948
rect 38551 748 38611 948
rect 38669 748 38729 948
rect 38787 748 38847 948
rect 39739 1042 39799 1442
rect 39857 1042 39917 1442
rect 39975 1042 40035 1442
rect 40093 1042 40153 1442
rect 40211 1042 40271 1442
rect 40329 1042 40389 1442
rect 30152 415 30352 475
rect 45863 1733 45923 1933
rect 45981 1733 46041 1933
rect 46099 1733 46159 1933
rect 46347 1733 46407 2133
rect 46465 1733 46525 2133
rect 46583 1733 46643 2133
rect 46701 1733 46761 2133
rect 46819 1733 46879 2133
rect 46937 1733 46997 2133
rect 47184 1733 47244 1933
rect 47302 1733 47362 1933
rect 47420 1733 47480 1933
rect 47761 1733 47821 1933
rect 47879 1733 47939 1933
rect 47997 1733 48057 1933
rect 48245 1733 48305 2133
rect 48363 1733 48423 2133
rect 48481 1733 48541 2133
rect 48599 1733 48659 2133
rect 48717 1733 48777 2133
rect 48835 1733 48895 2133
rect 49082 1733 49142 1933
rect 49200 1733 49260 1933
rect 49318 1733 49378 1933
rect 41637 1042 41697 1442
rect 41755 1042 41815 1442
rect 41873 1042 41933 1442
rect 41991 1042 42051 1442
rect 42109 1042 42169 1442
rect 42227 1042 42287 1442
rect 44394 746 44454 946
rect 44512 746 44572 946
rect 44630 746 44690 946
rect 44748 746 44808 946
rect 44866 746 44926 946
rect 44984 746 45044 946
rect 45102 746 45162 946
rect 45220 746 45280 946
rect 45338 746 45398 946
rect 46290 1040 46350 1440
rect 46408 1040 46468 1440
rect 46526 1040 46586 1440
rect 46644 1040 46704 1440
rect 46762 1040 46822 1440
rect 46880 1040 46940 1440
rect 29952 167 30352 227
rect 30645 224 31045 284
rect 29952 49 30352 109
rect 30645 106 31045 166
rect 52518 1734 52578 1934
rect 52636 1734 52696 1934
rect 52754 1734 52814 1934
rect 53002 1734 53062 2134
rect 53120 1734 53180 2134
rect 53238 1734 53298 2134
rect 53356 1734 53416 2134
rect 53474 1734 53534 2134
rect 53592 1734 53652 2134
rect 53839 1734 53899 1934
rect 53957 1734 54017 1934
rect 54075 1734 54135 1934
rect 54416 1734 54476 1934
rect 54534 1734 54594 1934
rect 54652 1734 54712 1934
rect 54900 1734 54960 2134
rect 55018 1734 55078 2134
rect 55136 1734 55196 2134
rect 55254 1734 55314 2134
rect 55372 1734 55432 2134
rect 55490 1734 55550 2134
rect 55737 1734 55797 1934
rect 55855 1734 55915 1934
rect 55973 1734 56033 1934
rect 48188 1040 48248 1440
rect 48306 1040 48366 1440
rect 48424 1040 48484 1440
rect 48542 1040 48602 1440
rect 48660 1040 48720 1440
rect 48778 1040 48838 1440
rect 51049 747 51109 947
rect 51167 747 51227 947
rect 51285 747 51345 947
rect 51403 747 51463 947
rect 51521 747 51581 947
rect 51639 747 51699 947
rect 51757 747 51817 947
rect 51875 747 51935 947
rect 51993 747 52053 947
rect 52945 1041 53005 1441
rect 53063 1041 53123 1441
rect 53181 1041 53241 1441
rect 53299 1041 53359 1441
rect 53417 1041 53477 1441
rect 53535 1041 53595 1441
rect 29952 -69 30352 -9
rect 30645 -12 31045 48
rect 59140 1735 59200 1935
rect 59258 1735 59318 1935
rect 59376 1735 59436 1935
rect 59624 1735 59684 2135
rect 59742 1735 59802 2135
rect 59860 1735 59920 2135
rect 59978 1735 60038 2135
rect 60096 1735 60156 2135
rect 60214 1735 60274 2135
rect 60461 1735 60521 1935
rect 60579 1735 60639 1935
rect 60697 1735 60757 1935
rect 61038 1735 61098 1935
rect 61156 1735 61216 1935
rect 61274 1735 61334 1935
rect 61522 1735 61582 2135
rect 61640 1735 61700 2135
rect 61758 1735 61818 2135
rect 61876 1735 61936 2135
rect 61994 1735 62054 2135
rect 62112 1735 62172 2135
rect 70509 2149 70909 2209
rect 70509 2031 70909 2091
rect 62359 1735 62419 1935
rect 62477 1735 62537 1935
rect 62595 1735 62655 1935
rect 70509 1913 70909 1973
rect 54843 1041 54903 1441
rect 54961 1041 55021 1441
rect 55079 1041 55139 1441
rect 55197 1041 55257 1441
rect 55315 1041 55375 1441
rect 55433 1041 55493 1441
rect 57671 748 57731 948
rect 57789 748 57849 948
rect 57907 748 57967 948
rect 58025 748 58085 948
rect 58143 748 58203 948
rect 58261 748 58321 948
rect 58379 748 58439 948
rect 58497 748 58557 948
rect 58615 748 58675 948
rect 59567 1042 59627 1442
rect 59685 1042 59745 1442
rect 59803 1042 59863 1442
rect 59921 1042 59981 1442
rect 60039 1042 60099 1442
rect 60157 1042 60217 1442
rect 29952 -187 30352 -127
rect 29952 -305 30352 -245
rect 29952 -423 30352 -363
rect 30645 -130 31045 -70
rect 70509 1795 70909 1855
rect 70509 1677 70909 1737
rect 70509 1559 70909 1619
rect 61465 1042 61525 1442
rect 61583 1042 61643 1442
rect 61701 1042 61761 1442
rect 61819 1042 61879 1442
rect 61937 1042 61997 1442
rect 62055 1042 62115 1442
rect 63535 1208 63595 1408
rect 63653 1208 63713 1408
rect 63771 1208 63831 1408
rect 63889 1208 63949 1408
rect 64007 1208 64067 1408
rect 64125 1208 64185 1408
rect 64243 1208 64303 1408
rect 64361 1208 64421 1408
rect 64479 1208 64539 1408
rect 70509 1322 70909 1382
rect 70509 1204 70909 1264
rect 70509 1086 70909 1146
rect 70709 849 70909 909
rect 70709 731 70909 791
rect 70709 613 70909 673
rect 30645 -248 31045 -188
rect 30645 -366 31045 -306
rect 65282 -537 65342 -337
rect 65400 -537 65460 -337
rect 65518 -537 65578 -337
rect 65766 -537 65826 -137
rect 65884 -537 65944 -137
rect 66002 -537 66062 -137
rect 66120 -537 66180 -137
rect 66238 -537 66298 -137
rect 66356 -537 66416 -137
rect 70709 -87 70909 -27
rect 70709 -205 70909 -145
rect 66603 -537 66663 -337
rect 66721 -537 66781 -337
rect 66839 -537 66899 -337
rect 70709 -323 70909 -263
rect 30152 -670 30352 -610
rect 30152 -788 30352 -728
rect 67075 -540 67135 -340
rect 67193 -540 67253 -340
rect 67311 -540 67371 -340
rect 67429 -540 67489 -340
rect 67547 -540 67607 -340
rect 67665 -540 67725 -340
rect 67783 -540 67843 -340
rect 67901 -540 67961 -340
rect 68019 -540 68079 -340
rect 70509 -528 70909 -468
rect 30152 -906 30352 -846
rect 30150 -1417 30350 -1357
rect 30150 -1535 30350 -1475
rect 30150 -1653 30350 -1593
rect 338 -2152 398 -1952
rect 456 -2152 516 -1952
rect 574 -2152 634 -1952
rect 779 -2152 839 -1752
rect 897 -2152 957 -1752
rect 1015 -2152 1075 -1752
rect 1246 -2152 1306 -1752
rect 1364 -2152 1424 -1752
rect 1482 -2152 1542 -1752
rect 1600 -2152 1660 -1752
rect 1718 -2152 1778 -1752
rect 1836 -2152 1896 -1752
rect 2073 -2152 2133 -1752
rect 2191 -2152 2251 -1752
rect 2309 -2152 2369 -1752
rect 2546 -2152 2606 -1952
rect 2664 -2152 2724 -1952
rect 2782 -2152 2842 -1952
rect 3482 -2152 3542 -1952
rect 3600 -2152 3660 -1952
rect 3718 -2152 3778 -1952
rect 3923 -2152 3983 -1752
rect 4041 -2152 4101 -1752
rect 4159 -2152 4219 -1752
rect 4390 -2152 4450 -1752
rect 4508 -2152 4568 -1752
rect 4626 -2152 4686 -1752
rect 4744 -2152 4804 -1752
rect 4862 -2152 4922 -1752
rect 4980 -2152 5040 -1752
rect 5217 -2152 5277 -1752
rect 5335 -2152 5395 -1752
rect 5453 -2152 5513 -1752
rect 5690 -2152 5750 -1952
rect 5808 -2152 5868 -1952
rect 5926 -2152 5986 -1952
rect 6614 -2148 6674 -1948
rect 6732 -2148 6792 -1948
rect 6850 -2148 6910 -1948
rect 7055 -2148 7115 -1748
rect 7173 -2148 7233 -1748
rect 7291 -2148 7351 -1748
rect 7522 -2148 7582 -1748
rect 7640 -2148 7700 -1748
rect 7758 -2148 7818 -1748
rect 7876 -2148 7936 -1748
rect 7994 -2148 8054 -1748
rect 8112 -2148 8172 -1748
rect 8349 -2148 8409 -1748
rect 8467 -2148 8527 -1748
rect 8585 -2148 8645 -1748
rect 8822 -2148 8882 -1948
rect 8940 -2148 9000 -1948
rect 9058 -2148 9118 -1948
rect 9758 -2148 9818 -1948
rect 9876 -2148 9936 -1948
rect 9994 -2148 10054 -1948
rect 10199 -2148 10259 -1748
rect 10317 -2148 10377 -1748
rect 10435 -2148 10495 -1748
rect 10666 -2148 10726 -1748
rect 10784 -2148 10844 -1748
rect 10902 -2148 10962 -1748
rect 11020 -2148 11080 -1748
rect 11138 -2148 11198 -1748
rect 11256 -2148 11316 -1748
rect 11493 -2148 11553 -1748
rect 11611 -2148 11671 -1748
rect 11729 -2148 11789 -1748
rect 11966 -2148 12026 -1948
rect 12084 -2148 12144 -1948
rect 12202 -2148 12262 -1948
rect 12960 -2152 13020 -1952
rect 13078 -2152 13138 -1952
rect 13196 -2152 13256 -1952
rect 13401 -2152 13461 -1752
rect 13519 -2152 13579 -1752
rect 13637 -2152 13697 -1752
rect 13868 -2152 13928 -1752
rect 13986 -2152 14046 -1752
rect 14104 -2152 14164 -1752
rect 14222 -2152 14282 -1752
rect 14340 -2152 14400 -1752
rect 14458 -2152 14518 -1752
rect 14695 -2152 14755 -1752
rect 14813 -2152 14873 -1752
rect 14931 -2152 14991 -1752
rect 15168 -2152 15228 -1952
rect 15286 -2152 15346 -1952
rect 15404 -2152 15464 -1952
rect 16104 -2152 16164 -1952
rect 16222 -2152 16282 -1952
rect 16340 -2152 16400 -1952
rect 16545 -2152 16605 -1752
rect 16663 -2152 16723 -1752
rect 16781 -2152 16841 -1752
rect 17012 -2152 17072 -1752
rect 17130 -2152 17190 -1752
rect 17248 -2152 17308 -1752
rect 17366 -2152 17426 -1752
rect 17484 -2152 17544 -1752
rect 17602 -2152 17662 -1752
rect 17839 -2152 17899 -1752
rect 17957 -2152 18017 -1752
rect 18075 -2152 18135 -1752
rect 18312 -2152 18372 -1952
rect 18430 -2152 18490 -1952
rect 18548 -2152 18608 -1952
rect 19236 -2148 19296 -1948
rect 19354 -2148 19414 -1948
rect 19472 -2148 19532 -1948
rect 19677 -2148 19737 -1748
rect 19795 -2148 19855 -1748
rect 19913 -2148 19973 -1748
rect 20144 -2148 20204 -1748
rect 20262 -2148 20322 -1748
rect 20380 -2148 20440 -1748
rect 20498 -2148 20558 -1748
rect 20616 -2148 20676 -1748
rect 20734 -2148 20794 -1748
rect 20971 -2148 21031 -1748
rect 21089 -2148 21149 -1748
rect 21207 -2148 21267 -1748
rect 21444 -2148 21504 -1948
rect 21562 -2148 21622 -1948
rect 21680 -2148 21740 -1948
rect 22380 -2148 22440 -1948
rect 22498 -2148 22558 -1948
rect 22616 -2148 22676 -1948
rect 22821 -2148 22881 -1748
rect 22939 -2148 22999 -1748
rect 23057 -2148 23117 -1748
rect 23288 -2148 23348 -1748
rect 23406 -2148 23466 -1748
rect 23524 -2148 23584 -1748
rect 23642 -2148 23702 -1748
rect 23760 -2148 23820 -1748
rect 23878 -2148 23938 -1748
rect 24115 -2148 24175 -1748
rect 24233 -2148 24293 -1748
rect 24351 -2148 24411 -1748
rect 41651 -1755 41711 -1555
rect 41769 -1755 41829 -1555
rect 41887 -1755 41947 -1555
rect 42005 -1755 42065 -1555
rect 42123 -1755 42183 -1555
rect 42241 -1755 42301 -1555
rect 42359 -1755 42419 -1555
rect 42477 -1755 42537 -1555
rect 42595 -1755 42655 -1555
rect 48205 -1750 48265 -1550
rect 48323 -1750 48383 -1550
rect 48441 -1750 48501 -1550
rect 48559 -1750 48619 -1550
rect 48677 -1750 48737 -1550
rect 48795 -1750 48855 -1550
rect 48913 -1750 48973 -1550
rect 49031 -1750 49091 -1550
rect 49149 -1750 49209 -1550
rect 29950 -1901 30350 -1841
rect 30643 -1844 31043 -1784
rect 54854 -1762 54914 -1562
rect 54972 -1762 55032 -1562
rect 55090 -1762 55150 -1562
rect 55208 -1762 55268 -1562
rect 55326 -1762 55386 -1562
rect 55444 -1762 55504 -1562
rect 55562 -1762 55622 -1562
rect 55680 -1762 55740 -1562
rect 55798 -1762 55858 -1562
rect 63542 -1637 63602 -1437
rect 63660 -1637 63720 -1437
rect 63778 -1637 63838 -1437
rect 63896 -1637 63956 -1437
rect 64014 -1637 64074 -1437
rect 64132 -1637 64192 -1437
rect 64250 -1637 64310 -1437
rect 64368 -1637 64428 -1437
rect 64486 -1637 64546 -1437
rect 65709 -1230 65769 -830
rect 65827 -1230 65887 -830
rect 65945 -1230 66005 -830
rect 66063 -1230 66123 -830
rect 66181 -1230 66241 -830
rect 66299 -1230 66359 -830
rect 70509 -646 70909 -586
rect 70509 -764 70909 -704
rect 70509 -995 70909 -935
rect 70509 -1113 70909 -1053
rect 70509 -1231 70909 -1171
rect 70509 -1349 70909 -1289
rect 70509 -1467 70909 -1407
rect 24588 -2148 24648 -1948
rect 24706 -2148 24766 -1948
rect 24824 -2148 24884 -1948
rect 29950 -2019 30350 -1959
rect 30643 -1962 31043 -1902
rect 29950 -2137 30350 -2077
rect 30643 -2080 31043 -2020
rect 29950 -2255 30350 -2195
rect 29950 -2373 30350 -2313
rect 29950 -2491 30350 -2431
rect 30643 -2198 31043 -2138
rect 30643 -2316 31043 -2256
rect 70509 -1585 70909 -1525
rect 70509 -1822 70909 -1762
rect 70509 -1940 70909 -1880
rect 70509 -2058 70909 -1998
rect 70709 -2295 70909 -2235
rect 30643 -2434 31043 -2374
rect 70709 -2413 70909 -2353
rect 70709 -2531 70909 -2471
rect 30150 -2738 30350 -2678
rect 30150 -2856 30350 -2796
rect 30150 -2974 30350 -2914
<< ndiff >>
rect 39825 24084 39883 24096
rect 39825 23708 39837 24084
rect 39871 23708 39883 24084
rect 39825 23696 39883 23708
rect 39943 24084 40001 24096
rect 39943 23708 39955 24084
rect 39989 23708 40001 24084
rect 39943 23696 40001 23708
rect 40061 24084 40119 24096
rect 40061 23708 40073 24084
rect 40107 23708 40119 24084
rect 40178 24084 40236 24096
rect 40178 23908 40190 24084
rect 40224 23908 40236 24084
rect 40178 23896 40236 23908
rect 40296 24084 40354 24096
rect 40296 23908 40308 24084
rect 40342 23908 40354 24084
rect 40296 23896 40354 23908
rect 46338 24081 46396 24093
rect 41823 23810 41881 23822
rect 40061 23696 40119 23708
rect 41823 23634 41835 23810
rect 41869 23634 41881 23810
rect 41823 23622 41881 23634
rect 41941 23810 41999 23822
rect 41941 23634 41953 23810
rect 41987 23634 41999 23810
rect 41941 23622 41999 23634
rect 42059 23810 42117 23822
rect 42059 23634 42071 23810
rect 42105 23634 42117 23810
rect 42059 23622 42117 23634
rect 42177 23810 42235 23822
rect 42177 23634 42189 23810
rect 42223 23634 42235 23810
rect 42177 23622 42235 23634
rect 42965 23814 43023 23826
rect 42965 23638 42977 23814
rect 43011 23638 43023 23814
rect 42965 23626 43023 23638
rect 43083 23814 43141 23826
rect 43083 23638 43095 23814
rect 43129 23638 43141 23814
rect 43083 23626 43141 23638
rect 43201 23814 43259 23826
rect 43201 23638 43213 23814
rect 43247 23638 43259 23814
rect 43201 23626 43259 23638
rect 43319 23814 43377 23826
rect 43319 23638 43331 23814
rect 43365 23638 43377 23814
rect 43319 23626 43377 23638
rect 46338 23705 46350 24081
rect 46384 23705 46396 24081
rect 46338 23693 46396 23705
rect 46456 24081 46514 24093
rect 46456 23705 46468 24081
rect 46502 23705 46514 24081
rect 46456 23693 46514 23705
rect 46574 24081 46632 24093
rect 46574 23705 46586 24081
rect 46620 23705 46632 24081
rect 46691 24081 46749 24093
rect 46691 23905 46703 24081
rect 46737 23905 46749 24081
rect 46691 23893 46749 23905
rect 46809 24081 46867 24093
rect 46809 23905 46821 24081
rect 46855 23905 46867 24081
rect 46809 23893 46867 23905
rect 52872 24076 52930 24088
rect 48336 23807 48394 23819
rect 46574 23693 46632 23705
rect 48336 23631 48348 23807
rect 48382 23631 48394 23807
rect 48336 23619 48394 23631
rect 48454 23807 48512 23819
rect 48454 23631 48466 23807
rect 48500 23631 48512 23807
rect 48454 23619 48512 23631
rect 48572 23807 48630 23819
rect 48572 23631 48584 23807
rect 48618 23631 48630 23807
rect 48572 23619 48630 23631
rect 48690 23807 48748 23819
rect 48690 23631 48702 23807
rect 48736 23631 48748 23807
rect 48690 23619 48748 23631
rect 49478 23811 49536 23823
rect 49478 23635 49490 23811
rect 49524 23635 49536 23811
rect 49478 23623 49536 23635
rect 49596 23811 49654 23823
rect 49596 23635 49608 23811
rect 49642 23635 49654 23811
rect 49596 23623 49654 23635
rect 49714 23811 49772 23823
rect 49714 23635 49726 23811
rect 49760 23635 49772 23811
rect 49714 23623 49772 23635
rect 49832 23811 49890 23823
rect 49832 23635 49844 23811
rect 49878 23635 49890 23811
rect 49832 23623 49890 23635
rect 52872 23700 52884 24076
rect 52918 23700 52930 24076
rect 52872 23688 52930 23700
rect 52990 24076 53048 24088
rect 52990 23700 53002 24076
rect 53036 23700 53048 24076
rect 52990 23688 53048 23700
rect 53108 24076 53166 24088
rect 53108 23700 53120 24076
rect 53154 23700 53166 24076
rect 53225 24076 53283 24088
rect 53225 23900 53237 24076
rect 53271 23900 53283 24076
rect 53225 23888 53283 23900
rect 53343 24076 53401 24088
rect 53343 23900 53355 24076
rect 53389 23900 53401 24076
rect 53343 23888 53401 23900
rect 59430 24080 59488 24092
rect 54870 23802 54928 23814
rect 53108 23688 53166 23700
rect 54870 23626 54882 23802
rect 54916 23626 54928 23802
rect 54870 23614 54928 23626
rect 54988 23802 55046 23814
rect 54988 23626 55000 23802
rect 55034 23626 55046 23802
rect 54988 23614 55046 23626
rect 55106 23802 55164 23814
rect 55106 23626 55118 23802
rect 55152 23626 55164 23802
rect 55106 23614 55164 23626
rect 55224 23802 55282 23814
rect 55224 23626 55236 23802
rect 55270 23626 55282 23802
rect 55224 23614 55282 23626
rect 56012 23806 56070 23818
rect 56012 23630 56024 23806
rect 56058 23630 56070 23806
rect 56012 23618 56070 23630
rect 56130 23806 56188 23818
rect 56130 23630 56142 23806
rect 56176 23630 56188 23806
rect 56130 23618 56188 23630
rect 56248 23806 56306 23818
rect 56248 23630 56260 23806
rect 56294 23630 56306 23806
rect 56248 23618 56306 23630
rect 56366 23806 56424 23818
rect 56366 23630 56378 23806
rect 56412 23630 56424 23806
rect 56366 23618 56424 23630
rect 59430 23704 59442 24080
rect 59476 23704 59488 24080
rect 59430 23692 59488 23704
rect 59548 24080 59606 24092
rect 59548 23704 59560 24080
rect 59594 23704 59606 24080
rect 59548 23692 59606 23704
rect 59666 24080 59724 24092
rect 59666 23704 59678 24080
rect 59712 23704 59724 24080
rect 59783 24080 59841 24092
rect 59783 23904 59795 24080
rect 59829 23904 59841 24080
rect 59783 23892 59841 23904
rect 59901 24080 59959 24092
rect 59901 23904 59913 24080
rect 59947 23904 59959 24080
rect 59901 23892 59959 23904
rect 61428 23806 61486 23818
rect 59666 23692 59724 23704
rect 61428 23630 61440 23806
rect 61474 23630 61486 23806
rect 61428 23618 61486 23630
rect 61546 23806 61604 23818
rect 61546 23630 61558 23806
rect 61592 23630 61604 23806
rect 61546 23618 61604 23630
rect 61664 23806 61722 23818
rect 61664 23630 61676 23806
rect 61710 23630 61722 23806
rect 61664 23618 61722 23630
rect 61782 23806 61840 23818
rect 61782 23630 61794 23806
rect 61828 23630 61840 23806
rect 61782 23618 61840 23630
rect 62570 23810 62628 23822
rect 62570 23634 62582 23810
rect 62616 23634 62628 23810
rect 62570 23622 62628 23634
rect 62688 23810 62746 23822
rect 62688 23634 62700 23810
rect 62734 23634 62746 23810
rect 62688 23622 62746 23634
rect 62806 23810 62864 23822
rect 62806 23634 62818 23810
rect 62852 23634 62864 23810
rect 62806 23622 62864 23634
rect 62924 23810 62982 23822
rect 62924 23634 62936 23810
rect 62970 23634 62982 23810
rect 62924 23622 62982 23634
rect 39839 22434 39897 22446
rect 39839 22058 39851 22434
rect 39885 22058 39897 22434
rect 39839 22046 39897 22058
rect 39957 22434 40015 22446
rect 39957 22058 39969 22434
rect 40003 22058 40015 22434
rect 39957 22046 40015 22058
rect 40075 22434 40133 22446
rect 40075 22058 40087 22434
rect 40121 22058 40133 22434
rect 40192 22434 40250 22446
rect 40192 22258 40204 22434
rect 40238 22258 40250 22434
rect 40192 22246 40250 22258
rect 40310 22434 40368 22446
rect 40310 22258 40322 22434
rect 40356 22258 40368 22434
rect 40310 22246 40368 22258
rect 40075 22046 40133 22058
rect 3868 20651 3926 20663
rect 3868 20475 3880 20651
rect 3914 20475 3926 20651
rect 3868 20463 3926 20475
rect 3986 20651 4122 20663
rect 3986 20475 3998 20651
rect 4032 20475 4076 20651
rect 3986 20463 4076 20475
rect 4064 20275 4076 20463
rect 4110 20275 4122 20651
rect 4064 20263 4122 20275
rect 4182 20651 4240 20663
rect 4182 20275 4194 20651
rect 4228 20275 4240 20651
rect 4182 20263 4240 20275
rect 4300 20651 4358 20663
rect 4300 20275 4312 20651
rect 4346 20275 4358 20651
rect 4300 20263 4358 20275
rect 4418 20651 4476 20663
rect 4418 20275 4430 20651
rect 4464 20275 4476 20651
rect 4418 20263 4476 20275
rect 4536 20651 4668 20663
rect 4536 20275 4548 20651
rect 4582 20475 4622 20651
rect 4656 20475 4668 20651
rect 4582 20463 4668 20475
rect 4728 20651 4786 20663
rect 4728 20475 4740 20651
rect 4774 20475 4786 20651
rect 4728 20463 4786 20475
rect 7012 20651 7070 20663
rect 7012 20475 7024 20651
rect 7058 20475 7070 20651
rect 7012 20463 7070 20475
rect 7130 20651 7266 20663
rect 7130 20475 7142 20651
rect 7176 20475 7220 20651
rect 7130 20463 7220 20475
rect 4582 20275 4594 20463
rect 4536 20263 4594 20275
rect 7208 20275 7220 20463
rect 7254 20275 7266 20651
rect 7208 20263 7266 20275
rect 7326 20651 7384 20663
rect 7326 20275 7338 20651
rect 7372 20275 7384 20651
rect 7326 20263 7384 20275
rect 7444 20651 7502 20663
rect 7444 20275 7456 20651
rect 7490 20275 7502 20651
rect 7444 20263 7502 20275
rect 7562 20651 7620 20663
rect 7562 20275 7574 20651
rect 7608 20275 7620 20651
rect 7562 20263 7620 20275
rect 7680 20651 7812 20663
rect 7680 20275 7692 20651
rect 7726 20475 7766 20651
rect 7800 20475 7812 20651
rect 7726 20463 7812 20475
rect 7872 20651 7930 20663
rect 46352 22431 46410 22443
rect 7872 20475 7884 20651
rect 7918 20475 7930 20651
rect 7872 20463 7930 20475
rect 10144 20647 10202 20659
rect 10144 20471 10156 20647
rect 10190 20471 10202 20647
rect 7726 20275 7738 20463
rect 10144 20459 10202 20471
rect 10262 20647 10398 20659
rect 10262 20471 10274 20647
rect 10308 20471 10352 20647
rect 10262 20459 10352 20471
rect 7680 20263 7738 20275
rect 10340 20271 10352 20459
rect 10386 20271 10398 20647
rect 10340 20259 10398 20271
rect 10458 20647 10516 20659
rect 10458 20271 10470 20647
rect 10504 20271 10516 20647
rect 10458 20259 10516 20271
rect 10576 20647 10634 20659
rect 10576 20271 10588 20647
rect 10622 20271 10634 20647
rect 10576 20259 10634 20271
rect 10694 20647 10752 20659
rect 10694 20271 10706 20647
rect 10740 20271 10752 20647
rect 10694 20259 10752 20271
rect 10812 20647 10944 20659
rect 10812 20271 10824 20647
rect 10858 20471 10898 20647
rect 10932 20471 10944 20647
rect 10858 20459 10944 20471
rect 11004 20647 11062 20659
rect 11004 20471 11016 20647
rect 11050 20471 11062 20647
rect 11004 20459 11062 20471
rect 13288 20647 13346 20659
rect 13288 20471 13300 20647
rect 13334 20471 13346 20647
rect 13288 20459 13346 20471
rect 13406 20647 13542 20659
rect 13406 20471 13418 20647
rect 13452 20471 13496 20647
rect 13406 20459 13496 20471
rect 10858 20271 10870 20459
rect 10812 20259 10870 20271
rect 13484 20271 13496 20459
rect 13530 20271 13542 20647
rect 13484 20259 13542 20271
rect 13602 20647 13660 20659
rect 13602 20271 13614 20647
rect 13648 20271 13660 20647
rect 13602 20259 13660 20271
rect 13720 20647 13778 20659
rect 13720 20271 13732 20647
rect 13766 20271 13778 20647
rect 13720 20259 13778 20271
rect 13838 20647 13896 20659
rect 13838 20271 13850 20647
rect 13884 20271 13896 20647
rect 13838 20259 13896 20271
rect 13956 20647 14088 20659
rect 13956 20271 13968 20647
rect 14002 20471 14042 20647
rect 14076 20471 14088 20647
rect 14002 20459 14088 20471
rect 14148 20647 14206 20659
rect 14148 20471 14160 20647
rect 14194 20471 14206 20647
rect 14148 20459 14206 20471
rect 16490 20651 16548 20663
rect 16490 20475 16502 20651
rect 16536 20475 16548 20651
rect 16490 20463 16548 20475
rect 16608 20651 16744 20663
rect 16608 20475 16620 20651
rect 16654 20475 16698 20651
rect 16608 20463 16698 20475
rect 14002 20271 14014 20459
rect 13956 20259 14014 20271
rect 16686 20275 16698 20463
rect 16732 20275 16744 20651
rect 16686 20263 16744 20275
rect 16804 20651 16862 20663
rect 16804 20275 16816 20651
rect 16850 20275 16862 20651
rect 16804 20263 16862 20275
rect 16922 20651 16980 20663
rect 16922 20275 16934 20651
rect 16968 20275 16980 20651
rect 16922 20263 16980 20275
rect 17040 20651 17098 20663
rect 17040 20275 17052 20651
rect 17086 20275 17098 20651
rect 17040 20263 17098 20275
rect 17158 20651 17290 20663
rect 17158 20275 17170 20651
rect 17204 20475 17244 20651
rect 17278 20475 17290 20651
rect 17204 20463 17290 20475
rect 17350 20651 17408 20663
rect 17350 20475 17362 20651
rect 17396 20475 17408 20651
rect 17350 20463 17408 20475
rect 19634 20651 19692 20663
rect 19634 20475 19646 20651
rect 19680 20475 19692 20651
rect 19634 20463 19692 20475
rect 19752 20651 19888 20663
rect 19752 20475 19764 20651
rect 19798 20475 19842 20651
rect 19752 20463 19842 20475
rect 17204 20275 17216 20463
rect 17158 20263 17216 20275
rect 19830 20275 19842 20463
rect 19876 20275 19888 20651
rect 19830 20263 19888 20275
rect 19948 20651 20006 20663
rect 19948 20275 19960 20651
rect 19994 20275 20006 20651
rect 19948 20263 20006 20275
rect 20066 20651 20124 20663
rect 20066 20275 20078 20651
rect 20112 20275 20124 20651
rect 20066 20263 20124 20275
rect 20184 20651 20242 20663
rect 20184 20275 20196 20651
rect 20230 20275 20242 20651
rect 20184 20263 20242 20275
rect 20302 20651 20434 20663
rect 20302 20275 20314 20651
rect 20348 20475 20388 20651
rect 20422 20475 20434 20651
rect 20348 20463 20434 20475
rect 20494 20651 20552 20663
rect 46352 22055 46364 22431
rect 46398 22055 46410 22431
rect 46352 22043 46410 22055
rect 46470 22431 46528 22443
rect 46470 22055 46482 22431
rect 46516 22055 46528 22431
rect 46470 22043 46528 22055
rect 46588 22431 46646 22443
rect 46588 22055 46600 22431
rect 46634 22055 46646 22431
rect 46705 22431 46763 22443
rect 46705 22255 46717 22431
rect 46751 22255 46763 22431
rect 46705 22243 46763 22255
rect 46823 22431 46881 22443
rect 46823 22255 46835 22431
rect 46869 22255 46881 22431
rect 46823 22243 46881 22255
rect 46588 22043 46646 22055
rect 52886 22426 52944 22438
rect 41191 21029 41249 21041
rect 41191 20853 41203 21029
rect 41237 20853 41249 21029
rect 39834 20830 39892 20842
rect 20494 20475 20506 20651
rect 20540 20475 20552 20651
rect 20494 20463 20552 20475
rect 22766 20647 22824 20659
rect 22766 20471 22778 20647
rect 22812 20471 22824 20647
rect 20348 20275 20360 20463
rect 22766 20459 22824 20471
rect 22884 20647 23020 20659
rect 22884 20471 22896 20647
rect 22930 20471 22974 20647
rect 22884 20459 22974 20471
rect 20302 20263 20360 20275
rect 22962 20271 22974 20459
rect 23008 20271 23020 20647
rect 22962 20259 23020 20271
rect 23080 20647 23138 20659
rect 23080 20271 23092 20647
rect 23126 20271 23138 20647
rect 23080 20259 23138 20271
rect 23198 20647 23256 20659
rect 23198 20271 23210 20647
rect 23244 20271 23256 20647
rect 23198 20259 23256 20271
rect 23316 20647 23374 20659
rect 23316 20271 23328 20647
rect 23362 20271 23374 20647
rect 23316 20259 23374 20271
rect 23434 20647 23566 20659
rect 23434 20271 23446 20647
rect 23480 20471 23520 20647
rect 23554 20471 23566 20647
rect 23480 20459 23566 20471
rect 23626 20647 23684 20659
rect 23626 20471 23638 20647
rect 23672 20471 23684 20647
rect 23626 20459 23684 20471
rect 25910 20647 25968 20659
rect 25910 20471 25922 20647
rect 25956 20471 25968 20647
rect 25910 20459 25968 20471
rect 26028 20647 26164 20659
rect 26028 20471 26040 20647
rect 26074 20471 26118 20647
rect 26028 20459 26118 20471
rect 23480 20271 23492 20459
rect 23434 20259 23492 20271
rect 26106 20271 26118 20459
rect 26152 20271 26164 20647
rect 26106 20259 26164 20271
rect 26224 20647 26282 20659
rect 26224 20271 26236 20647
rect 26270 20271 26282 20647
rect 26224 20259 26282 20271
rect 26342 20647 26400 20659
rect 26342 20271 26354 20647
rect 26388 20271 26400 20647
rect 26342 20259 26400 20271
rect 26460 20647 26518 20659
rect 26460 20271 26472 20647
rect 26506 20271 26518 20647
rect 26460 20259 26518 20271
rect 26578 20647 26710 20659
rect 26578 20271 26590 20647
rect 26624 20471 26664 20647
rect 26698 20471 26710 20647
rect 26624 20459 26710 20471
rect 26770 20647 26828 20659
rect 26770 20471 26782 20647
rect 26816 20471 26828 20647
rect 26770 20459 26828 20471
rect 26624 20271 26636 20459
rect 39834 20454 39846 20830
rect 39880 20454 39892 20830
rect 39834 20442 39892 20454
rect 39952 20830 40010 20842
rect 39952 20454 39964 20830
rect 39998 20454 40010 20830
rect 39952 20442 40010 20454
rect 40070 20830 40128 20842
rect 40070 20454 40082 20830
rect 40116 20454 40128 20830
rect 40187 20830 40245 20842
rect 40187 20654 40199 20830
rect 40233 20654 40245 20830
rect 40187 20642 40245 20654
rect 40305 20830 40363 20842
rect 41191 20841 41249 20853
rect 41309 21029 41367 21041
rect 41309 20853 41321 21029
rect 41355 20853 41367 21029
rect 41309 20841 41367 20853
rect 41611 21029 41669 21041
rect 40305 20654 40317 20830
rect 40351 20654 40363 20830
rect 40305 20642 40363 20654
rect 41611 20653 41623 21029
rect 41657 20653 41669 21029
rect 41611 20641 41669 20653
rect 41729 21029 41787 21041
rect 41729 20653 41741 21029
rect 41775 20653 41787 21029
rect 41729 20641 41787 20653
rect 41847 21029 41905 21041
rect 41847 20653 41859 21029
rect 41893 20653 41905 21029
rect 41847 20641 41905 20653
rect 41965 21029 42023 21041
rect 41965 20653 41977 21029
rect 42011 20653 42023 21029
rect 41965 20641 42023 20653
rect 42083 21029 42141 21041
rect 42083 20653 42095 21029
rect 42129 20653 42141 21029
rect 42489 21029 42547 21041
rect 42489 20853 42501 21029
rect 42535 20853 42547 21029
rect 42489 20841 42547 20853
rect 42607 21029 42665 21041
rect 42607 20853 42619 21029
rect 42653 20853 42665 21029
rect 42607 20841 42665 20853
rect 43089 21029 43147 21041
rect 43089 20853 43101 21029
rect 43135 20853 43147 21029
rect 43089 20841 43147 20853
rect 43207 21029 43265 21041
rect 43207 20853 43219 21029
rect 43253 20853 43265 21029
rect 43207 20841 43265 20853
rect 43509 21029 43567 21041
rect 42083 20641 42141 20653
rect 43509 20653 43521 21029
rect 43555 20653 43567 21029
rect 43509 20641 43567 20653
rect 43627 21029 43685 21041
rect 43627 20653 43639 21029
rect 43673 20653 43685 21029
rect 43627 20641 43685 20653
rect 43745 21029 43803 21041
rect 43745 20653 43757 21029
rect 43791 20653 43803 21029
rect 43745 20641 43803 20653
rect 43863 21029 43921 21041
rect 43863 20653 43875 21029
rect 43909 20653 43921 21029
rect 43863 20641 43921 20653
rect 43981 21029 44039 21041
rect 43981 20653 43993 21029
rect 44027 20653 44039 21029
rect 44387 21029 44445 21041
rect 44387 20853 44399 21029
rect 44433 20853 44445 21029
rect 44387 20841 44445 20853
rect 44505 21029 44563 21041
rect 44505 20853 44517 21029
rect 44551 20853 44563 21029
rect 44505 20841 44563 20853
rect 52886 22050 52898 22426
rect 52932 22050 52944 22426
rect 52886 22038 52944 22050
rect 53004 22426 53062 22438
rect 53004 22050 53016 22426
rect 53050 22050 53062 22426
rect 53004 22038 53062 22050
rect 53122 22426 53180 22438
rect 53122 22050 53134 22426
rect 53168 22050 53180 22426
rect 53239 22426 53297 22438
rect 53239 22250 53251 22426
rect 53285 22250 53297 22426
rect 53239 22238 53297 22250
rect 53357 22426 53415 22438
rect 53357 22250 53369 22426
rect 53403 22250 53415 22426
rect 53357 22238 53415 22250
rect 53122 22038 53180 22050
rect 59444 22430 59502 22442
rect 47704 21026 47762 21038
rect 47704 20850 47716 21026
rect 47750 20850 47762 21026
rect 46347 20827 46405 20839
rect 43981 20641 44039 20653
rect 40070 20442 40128 20454
rect 46347 20451 46359 20827
rect 46393 20451 46405 20827
rect 46347 20439 46405 20451
rect 46465 20827 46523 20839
rect 46465 20451 46477 20827
rect 46511 20451 46523 20827
rect 46465 20439 46523 20451
rect 46583 20827 46641 20839
rect 46583 20451 46595 20827
rect 46629 20451 46641 20827
rect 46700 20827 46758 20839
rect 46700 20651 46712 20827
rect 46746 20651 46758 20827
rect 46700 20639 46758 20651
rect 46818 20827 46876 20839
rect 47704 20838 47762 20850
rect 47822 21026 47880 21038
rect 47822 20850 47834 21026
rect 47868 20850 47880 21026
rect 47822 20838 47880 20850
rect 48124 21026 48182 21038
rect 46818 20651 46830 20827
rect 46864 20651 46876 20827
rect 46818 20639 46876 20651
rect 48124 20650 48136 21026
rect 48170 20650 48182 21026
rect 48124 20638 48182 20650
rect 48242 21026 48300 21038
rect 48242 20650 48254 21026
rect 48288 20650 48300 21026
rect 48242 20638 48300 20650
rect 48360 21026 48418 21038
rect 48360 20650 48372 21026
rect 48406 20650 48418 21026
rect 48360 20638 48418 20650
rect 48478 21026 48536 21038
rect 48478 20650 48490 21026
rect 48524 20650 48536 21026
rect 48478 20638 48536 20650
rect 48596 21026 48654 21038
rect 48596 20650 48608 21026
rect 48642 20650 48654 21026
rect 49002 21026 49060 21038
rect 49002 20850 49014 21026
rect 49048 20850 49060 21026
rect 49002 20838 49060 20850
rect 49120 21026 49178 21038
rect 49120 20850 49132 21026
rect 49166 20850 49178 21026
rect 49120 20838 49178 20850
rect 49602 21026 49660 21038
rect 49602 20850 49614 21026
rect 49648 20850 49660 21026
rect 49602 20838 49660 20850
rect 49720 21026 49778 21038
rect 49720 20850 49732 21026
rect 49766 20850 49778 21026
rect 49720 20838 49778 20850
rect 50022 21026 50080 21038
rect 48596 20638 48654 20650
rect 50022 20650 50034 21026
rect 50068 20650 50080 21026
rect 50022 20638 50080 20650
rect 50140 21026 50198 21038
rect 50140 20650 50152 21026
rect 50186 20650 50198 21026
rect 50140 20638 50198 20650
rect 50258 21026 50316 21038
rect 50258 20650 50270 21026
rect 50304 20650 50316 21026
rect 50258 20638 50316 20650
rect 50376 21026 50434 21038
rect 50376 20650 50388 21026
rect 50422 20650 50434 21026
rect 50376 20638 50434 20650
rect 50494 21026 50552 21038
rect 50494 20650 50506 21026
rect 50540 20650 50552 21026
rect 50900 21026 50958 21038
rect 50900 20850 50912 21026
rect 50946 20850 50958 21026
rect 50900 20838 50958 20850
rect 51018 21026 51076 21038
rect 51018 20850 51030 21026
rect 51064 20850 51076 21026
rect 51018 20838 51076 20850
rect 59444 22054 59456 22430
rect 59490 22054 59502 22430
rect 59444 22042 59502 22054
rect 59562 22430 59620 22442
rect 59562 22054 59574 22430
rect 59608 22054 59620 22430
rect 59562 22042 59620 22054
rect 59680 22430 59738 22442
rect 59680 22054 59692 22430
rect 59726 22054 59738 22430
rect 59797 22430 59855 22442
rect 59797 22254 59809 22430
rect 59843 22254 59855 22430
rect 59797 22242 59855 22254
rect 59915 22430 59973 22442
rect 59915 22254 59927 22430
rect 59961 22254 59973 22430
rect 59915 22242 59973 22254
rect 59680 22042 59738 22054
rect 54238 21021 54296 21033
rect 54238 20845 54250 21021
rect 54284 20845 54296 21021
rect 52881 20822 52939 20834
rect 50494 20638 50552 20650
rect 46583 20439 46641 20451
rect 26578 20259 26636 20271
rect 52881 20446 52893 20822
rect 52927 20446 52939 20822
rect 52881 20434 52939 20446
rect 52999 20822 53057 20834
rect 52999 20446 53011 20822
rect 53045 20446 53057 20822
rect 52999 20434 53057 20446
rect 53117 20822 53175 20834
rect 53117 20446 53129 20822
rect 53163 20446 53175 20822
rect 53234 20822 53292 20834
rect 53234 20646 53246 20822
rect 53280 20646 53292 20822
rect 53234 20634 53292 20646
rect 53352 20822 53410 20834
rect 54238 20833 54296 20845
rect 54356 21021 54414 21033
rect 54356 20845 54368 21021
rect 54402 20845 54414 21021
rect 54356 20833 54414 20845
rect 54658 21021 54716 21033
rect 53352 20646 53364 20822
rect 53398 20646 53410 20822
rect 53352 20634 53410 20646
rect 54658 20645 54670 21021
rect 54704 20645 54716 21021
rect 54658 20633 54716 20645
rect 54776 21021 54834 21033
rect 54776 20645 54788 21021
rect 54822 20645 54834 21021
rect 54776 20633 54834 20645
rect 54894 21021 54952 21033
rect 54894 20645 54906 21021
rect 54940 20645 54952 21021
rect 54894 20633 54952 20645
rect 55012 21021 55070 21033
rect 55012 20645 55024 21021
rect 55058 20645 55070 21021
rect 55012 20633 55070 20645
rect 55130 21021 55188 21033
rect 55130 20645 55142 21021
rect 55176 20645 55188 21021
rect 55536 21021 55594 21033
rect 55536 20845 55548 21021
rect 55582 20845 55594 21021
rect 55536 20833 55594 20845
rect 55654 21021 55712 21033
rect 55654 20845 55666 21021
rect 55700 20845 55712 21021
rect 55654 20833 55712 20845
rect 56136 21021 56194 21033
rect 56136 20845 56148 21021
rect 56182 20845 56194 21021
rect 56136 20833 56194 20845
rect 56254 21021 56312 21033
rect 56254 20845 56266 21021
rect 56300 20845 56312 21021
rect 56254 20833 56312 20845
rect 56556 21021 56614 21033
rect 55130 20633 55188 20645
rect 56556 20645 56568 21021
rect 56602 20645 56614 21021
rect 56556 20633 56614 20645
rect 56674 21021 56732 21033
rect 56674 20645 56686 21021
rect 56720 20645 56732 21021
rect 56674 20633 56732 20645
rect 56792 21021 56850 21033
rect 56792 20645 56804 21021
rect 56838 20645 56850 21021
rect 56792 20633 56850 20645
rect 56910 21021 56968 21033
rect 56910 20645 56922 21021
rect 56956 20645 56968 21021
rect 56910 20633 56968 20645
rect 57028 21021 57086 21033
rect 57028 20645 57040 21021
rect 57074 20645 57086 21021
rect 57434 21021 57492 21033
rect 57434 20845 57446 21021
rect 57480 20845 57492 21021
rect 57434 20833 57492 20845
rect 57552 21021 57610 21033
rect 57552 20845 57564 21021
rect 57598 20845 57610 21021
rect 57552 20833 57610 20845
rect 60796 21025 60854 21037
rect 60796 20849 60808 21025
rect 60842 20849 60854 21025
rect 59439 20826 59497 20838
rect 57028 20633 57086 20645
rect 53117 20434 53175 20446
rect 59439 20450 59451 20826
rect 59485 20450 59497 20826
rect 59439 20438 59497 20450
rect 59557 20826 59615 20838
rect 59557 20450 59569 20826
rect 59603 20450 59615 20826
rect 59557 20438 59615 20450
rect 59675 20826 59733 20838
rect 59675 20450 59687 20826
rect 59721 20450 59733 20826
rect 59792 20826 59850 20838
rect 59792 20650 59804 20826
rect 59838 20650 59850 20826
rect 59792 20638 59850 20650
rect 59910 20826 59968 20838
rect 60796 20837 60854 20849
rect 60914 21025 60972 21037
rect 60914 20849 60926 21025
rect 60960 20849 60972 21025
rect 60914 20837 60972 20849
rect 61216 21025 61274 21037
rect 59910 20650 59922 20826
rect 59956 20650 59968 20826
rect 59910 20638 59968 20650
rect 61216 20649 61228 21025
rect 61262 20649 61274 21025
rect 61216 20637 61274 20649
rect 61334 21025 61392 21037
rect 61334 20649 61346 21025
rect 61380 20649 61392 21025
rect 61334 20637 61392 20649
rect 61452 21025 61510 21037
rect 61452 20649 61464 21025
rect 61498 20649 61510 21025
rect 61452 20637 61510 20649
rect 61570 21025 61628 21037
rect 61570 20649 61582 21025
rect 61616 20649 61628 21025
rect 61570 20637 61628 20649
rect 61688 21025 61746 21037
rect 61688 20649 61700 21025
rect 61734 20649 61746 21025
rect 62094 21025 62152 21037
rect 62094 20849 62106 21025
rect 62140 20849 62152 21025
rect 62094 20837 62152 20849
rect 62212 21025 62270 21037
rect 62212 20849 62224 21025
rect 62258 20849 62270 21025
rect 62212 20837 62270 20849
rect 62694 21025 62752 21037
rect 62694 20849 62706 21025
rect 62740 20849 62752 21025
rect 62694 20837 62752 20849
rect 62812 21025 62870 21037
rect 62812 20849 62824 21025
rect 62858 20849 62870 21025
rect 62812 20837 62870 20849
rect 63114 21025 63172 21037
rect 61688 20637 61746 20649
rect 63114 20649 63126 21025
rect 63160 20649 63172 21025
rect 63114 20637 63172 20649
rect 63232 21025 63290 21037
rect 63232 20649 63244 21025
rect 63278 20649 63290 21025
rect 63232 20637 63290 20649
rect 63350 21025 63408 21037
rect 63350 20649 63362 21025
rect 63396 20649 63408 21025
rect 63350 20637 63408 20649
rect 63468 21025 63526 21037
rect 63468 20649 63480 21025
rect 63514 20649 63526 21025
rect 63468 20637 63526 20649
rect 63586 21025 63644 21037
rect 63586 20649 63598 21025
rect 63632 20649 63644 21025
rect 63992 21025 64050 21037
rect 63992 20849 64004 21025
rect 64038 20849 64050 21025
rect 63992 20837 64050 20849
rect 64110 21025 64168 21037
rect 64110 20849 64122 21025
rect 64156 20849 64168 21025
rect 71846 21227 72046 21239
rect 71846 21193 71858 21227
rect 72034 21193 72046 21227
rect 71846 21181 72046 21193
rect 71846 21109 72046 21121
rect 71846 21075 71858 21109
rect 72034 21075 72046 21109
rect 71846 21047 72046 21075
rect 71846 21035 72246 21047
rect 71846 21001 71858 21035
rect 72234 21001 72246 21035
rect 71846 20989 72246 21001
rect 64110 20837 64168 20849
rect 63586 20637 63644 20649
rect 71846 20917 72246 20929
rect 71846 20883 71858 20917
rect 72234 20883 72246 20917
rect 71846 20871 72246 20883
rect 71846 20799 72246 20811
rect 71846 20765 71858 20799
rect 72234 20765 72246 20799
rect 71846 20753 72246 20765
rect 71846 20681 72246 20693
rect 71846 20647 71858 20681
rect 72234 20647 72246 20681
rect 71846 20635 72246 20647
rect 59675 20438 59733 20450
rect 71846 20563 72246 20575
rect 71846 20529 71858 20563
rect 72234 20529 72246 20563
rect 71846 20517 72246 20529
rect 71846 20485 72046 20517
rect 71846 20451 71858 20485
rect 72034 20451 72046 20485
rect 71846 20439 72046 20451
rect 71846 20367 72046 20379
rect 71846 20333 71858 20367
rect 72034 20333 72046 20367
rect 71846 20321 72046 20333
rect 40043 18206 40101 18218
rect 40043 18030 40055 18206
rect 40089 18030 40101 18206
rect 40043 18018 40101 18030
rect 40161 18206 40219 18218
rect 40161 18030 40173 18206
rect 40207 18030 40219 18206
rect 40161 18018 40219 18030
rect 40279 18206 40337 18218
rect 40279 18030 40291 18206
rect 40325 18030 40337 18206
rect 40279 18018 40337 18030
rect 40397 18206 40455 18218
rect 43066 18476 43124 18488
rect 43066 18300 43078 18476
rect 43112 18300 43124 18476
rect 43066 18288 43124 18300
rect 43184 18476 43242 18488
rect 43184 18300 43196 18476
rect 43230 18300 43242 18476
rect 43184 18288 43242 18300
rect 43301 18476 43359 18488
rect 40397 18030 40409 18206
rect 40443 18030 40455 18206
rect 40397 18018 40455 18030
rect 41185 18202 41243 18214
rect 41185 18026 41197 18202
rect 41231 18026 41243 18202
rect 41185 18014 41243 18026
rect 41303 18202 41361 18214
rect 41303 18026 41315 18202
rect 41349 18026 41361 18202
rect 41303 18014 41361 18026
rect 41421 18202 41479 18214
rect 41421 18026 41433 18202
rect 41467 18026 41479 18202
rect 41421 18014 41479 18026
rect 41539 18202 41597 18214
rect 41539 18026 41551 18202
rect 41585 18026 41597 18202
rect 43301 18100 43313 18476
rect 43347 18100 43359 18476
rect 43301 18088 43359 18100
rect 43419 18476 43477 18488
rect 43419 18100 43431 18476
rect 43465 18100 43477 18476
rect 43419 18088 43477 18100
rect 43537 18476 43595 18488
rect 43537 18100 43549 18476
rect 43583 18100 43595 18476
rect 43537 18088 43595 18100
rect 41539 18014 41597 18026
rect 46601 18202 46659 18214
rect 46601 18026 46613 18202
rect 46647 18026 46659 18202
rect 46601 18014 46659 18026
rect 46719 18202 46777 18214
rect 46719 18026 46731 18202
rect 46765 18026 46777 18202
rect 46719 18014 46777 18026
rect 46837 18202 46895 18214
rect 46837 18026 46849 18202
rect 46883 18026 46895 18202
rect 46837 18014 46895 18026
rect 46955 18202 47013 18214
rect 49624 18472 49682 18484
rect 49624 18296 49636 18472
rect 49670 18296 49682 18472
rect 49624 18284 49682 18296
rect 49742 18472 49800 18484
rect 49742 18296 49754 18472
rect 49788 18296 49800 18472
rect 49742 18284 49800 18296
rect 49859 18472 49917 18484
rect 46955 18026 46967 18202
rect 47001 18026 47013 18202
rect 46955 18014 47013 18026
rect 47743 18198 47801 18210
rect 47743 18022 47755 18198
rect 47789 18022 47801 18198
rect 47743 18010 47801 18022
rect 47861 18198 47919 18210
rect 47861 18022 47873 18198
rect 47907 18022 47919 18198
rect 47861 18010 47919 18022
rect 47979 18198 48037 18210
rect 47979 18022 47991 18198
rect 48025 18022 48037 18198
rect 47979 18010 48037 18022
rect 48097 18198 48155 18210
rect 48097 18022 48109 18198
rect 48143 18022 48155 18198
rect 49859 18096 49871 18472
rect 49905 18096 49917 18472
rect 49859 18084 49917 18096
rect 49977 18472 50035 18484
rect 49977 18096 49989 18472
rect 50023 18096 50035 18472
rect 49977 18084 50035 18096
rect 50095 18472 50153 18484
rect 50095 18096 50107 18472
rect 50141 18096 50153 18472
rect 50095 18084 50153 18096
rect 48097 18010 48155 18022
rect 53135 18207 53193 18219
rect 53135 18031 53147 18207
rect 53181 18031 53193 18207
rect 53135 18019 53193 18031
rect 53253 18207 53311 18219
rect 53253 18031 53265 18207
rect 53299 18031 53311 18207
rect 53253 18019 53311 18031
rect 53371 18207 53429 18219
rect 53371 18031 53383 18207
rect 53417 18031 53429 18207
rect 53371 18019 53429 18031
rect 53489 18207 53547 18219
rect 56158 18477 56216 18489
rect 56158 18301 56170 18477
rect 56204 18301 56216 18477
rect 56158 18289 56216 18301
rect 56276 18477 56334 18489
rect 56276 18301 56288 18477
rect 56322 18301 56334 18477
rect 56276 18289 56334 18301
rect 56393 18477 56451 18489
rect 53489 18031 53501 18207
rect 53535 18031 53547 18207
rect 53489 18019 53547 18031
rect 54277 18203 54335 18215
rect 54277 18027 54289 18203
rect 54323 18027 54335 18203
rect 54277 18015 54335 18027
rect 54395 18203 54453 18215
rect 54395 18027 54407 18203
rect 54441 18027 54453 18203
rect 54395 18015 54453 18027
rect 54513 18203 54571 18215
rect 54513 18027 54525 18203
rect 54559 18027 54571 18203
rect 54513 18015 54571 18027
rect 54631 18203 54689 18215
rect 54631 18027 54643 18203
rect 54677 18027 54689 18203
rect 56393 18101 56405 18477
rect 56439 18101 56451 18477
rect 56393 18089 56451 18101
rect 56511 18477 56569 18489
rect 56511 18101 56523 18477
rect 56557 18101 56569 18477
rect 56511 18089 56569 18101
rect 56629 18477 56687 18489
rect 56629 18101 56641 18477
rect 56675 18101 56687 18477
rect 56629 18089 56687 18101
rect 54631 18015 54689 18027
rect 59648 18210 59706 18222
rect 59648 18034 59660 18210
rect 59694 18034 59706 18210
rect 59648 18022 59706 18034
rect 59766 18210 59824 18222
rect 59766 18034 59778 18210
rect 59812 18034 59824 18210
rect 59766 18022 59824 18034
rect 59884 18210 59942 18222
rect 59884 18034 59896 18210
rect 59930 18034 59942 18210
rect 59884 18022 59942 18034
rect 60002 18210 60060 18222
rect 62671 18480 62729 18492
rect 62671 18304 62683 18480
rect 62717 18304 62729 18480
rect 62671 18292 62729 18304
rect 62789 18480 62847 18492
rect 62789 18304 62801 18480
rect 62835 18304 62847 18480
rect 62789 18292 62847 18304
rect 62906 18480 62964 18492
rect 60002 18034 60014 18210
rect 60048 18034 60060 18210
rect 60002 18022 60060 18034
rect 60790 18206 60848 18218
rect 60790 18030 60802 18206
rect 60836 18030 60848 18206
rect 60790 18018 60848 18030
rect 60908 18206 60966 18218
rect 60908 18030 60920 18206
rect 60954 18030 60966 18206
rect 60908 18018 60966 18030
rect 61026 18206 61084 18218
rect 61026 18030 61038 18206
rect 61072 18030 61084 18206
rect 61026 18018 61084 18030
rect 61144 18206 61202 18218
rect 61144 18030 61156 18206
rect 61190 18030 61202 18206
rect 62906 18104 62918 18480
rect 62952 18104 62964 18480
rect 62906 18092 62964 18104
rect 63024 18480 63082 18492
rect 63024 18104 63036 18480
rect 63070 18104 63082 18480
rect 63024 18092 63082 18104
rect 63142 18480 63200 18492
rect 63142 18104 63154 18480
rect 63188 18104 63200 18480
rect 63142 18092 63200 18104
rect 61144 18018 61202 18030
rect 71846 18083 72046 18095
rect 71846 18049 71858 18083
rect 72034 18049 72046 18083
rect 71846 18037 72046 18049
rect 71846 17965 72046 17977
rect 71846 17931 71858 17965
rect 72034 17931 72046 17965
rect 71846 17903 72046 17931
rect 71846 17891 72246 17903
rect 71846 17857 71858 17891
rect 72234 17857 72246 17891
rect 71846 17845 72246 17857
rect 71846 17773 72246 17785
rect 71846 17739 71858 17773
rect 72234 17739 72246 17773
rect 71846 17727 72246 17739
rect 71846 17655 72246 17667
rect 71846 17621 71858 17655
rect 72234 17621 72246 17655
rect 71846 17609 72246 17621
rect 71846 17537 72246 17549
rect 71846 17503 71858 17537
rect 72234 17503 72246 17537
rect 71846 17491 72246 17503
rect 4952 16014 5010 16026
rect 4952 15838 4964 16014
rect 4998 15838 5010 16014
rect 4952 15826 5010 15838
rect 5070 16014 5128 16026
rect 5070 15838 5082 16014
rect 5116 15838 5128 16014
rect 5070 15826 5128 15838
rect 5188 16014 5246 16026
rect 5188 15838 5200 16014
rect 5234 15838 5246 16014
rect 5188 15826 5246 15838
rect 5306 16014 5364 16026
rect 5306 15838 5318 16014
rect 5352 15838 5364 16014
rect 5306 15826 5364 15838
rect 6120 16014 6178 16026
rect 6120 15838 6132 16014
rect 6166 15838 6178 16014
rect 6120 15826 6178 15838
rect 6238 16014 6296 16026
rect 6238 15838 6250 16014
rect 6284 15838 6296 16014
rect 6238 15826 6296 15838
rect 6356 16014 6414 16026
rect 6356 15838 6368 16014
rect 6402 15838 6414 16014
rect 6356 15826 6414 15838
rect 6474 16014 6532 16026
rect 6474 15838 6486 16014
rect 6520 15838 6532 16014
rect 6474 15826 6532 15838
rect 7288 16012 7346 16024
rect 7288 15836 7300 16012
rect 7334 15836 7346 16012
rect 7288 15824 7346 15836
rect 7406 16012 7464 16024
rect 7406 15836 7418 16012
rect 7452 15836 7464 16012
rect 7406 15824 7464 15836
rect 7524 16012 7582 16024
rect 7524 15836 7536 16012
rect 7570 15836 7582 16012
rect 7524 15824 7582 15836
rect 7642 16012 7700 16024
rect 7642 15836 7654 16012
rect 7688 15836 7700 16012
rect 7642 15824 7700 15836
rect 8456 16012 8514 16024
rect 8456 15836 8468 16012
rect 8502 15836 8514 16012
rect 8456 15824 8514 15836
rect 8574 16012 8632 16024
rect 8574 15836 8586 16012
rect 8620 15836 8632 16012
rect 8574 15824 8632 15836
rect 8692 16012 8750 16024
rect 8692 15836 8704 16012
rect 8738 15836 8750 16012
rect 8692 15824 8750 15836
rect 8810 16012 8868 16024
rect 8810 15836 8822 16012
rect 8856 15836 8868 16012
rect 8810 15824 8868 15836
rect 9630 16012 9688 16024
rect 9630 15836 9642 16012
rect 9676 15836 9688 16012
rect 9630 15824 9688 15836
rect 9748 16012 9806 16024
rect 9748 15836 9760 16012
rect 9794 15836 9806 16012
rect 9748 15824 9806 15836
rect 9866 16012 9924 16024
rect 9866 15836 9878 16012
rect 9912 15836 9924 16012
rect 9866 15824 9924 15836
rect 9984 16012 10042 16024
rect 9984 15836 9996 16012
rect 10030 15836 10042 16012
rect 9984 15824 10042 15836
rect 10798 16012 10856 16024
rect 10798 15836 10810 16012
rect 10844 15836 10856 16012
rect 10798 15824 10856 15836
rect 10916 16012 10974 16024
rect 10916 15836 10928 16012
rect 10962 15836 10974 16012
rect 10916 15824 10974 15836
rect 11034 16012 11092 16024
rect 11034 15836 11046 16012
rect 11080 15836 11092 16012
rect 11034 15824 11092 15836
rect 11152 16012 11210 16024
rect 11152 15836 11164 16012
rect 11198 15836 11210 16012
rect 11152 15824 11210 15836
rect 11966 16012 12024 16024
rect 11966 15836 11978 16012
rect 12012 15836 12024 16012
rect 11966 15824 12024 15836
rect 12084 16012 12142 16024
rect 12084 15836 12096 16012
rect 12130 15836 12142 16012
rect 12084 15824 12142 15836
rect 12202 16012 12260 16024
rect 12202 15836 12214 16012
rect 12248 15836 12260 16012
rect 12202 15824 12260 15836
rect 12320 16012 12378 16024
rect 14145 16164 14203 16176
rect 12320 15836 12332 16012
rect 12366 15836 12378 16012
rect 12320 15824 12378 15836
rect 13134 16010 13192 16022
rect 13134 15834 13146 16010
rect 13180 15834 13192 16010
rect 13134 15822 13192 15834
rect 13252 16010 13310 16022
rect 13252 15834 13264 16010
rect 13298 15834 13310 16010
rect 13252 15822 13310 15834
rect 13370 16010 13428 16022
rect 13370 15834 13382 16010
rect 13416 15834 13428 16010
rect 13370 15822 13428 15834
rect 13488 16010 13546 16022
rect 13488 15834 13500 16010
rect 13534 15834 13546 16010
rect 14145 15988 14157 16164
rect 14191 15988 14203 16164
rect 14145 15976 14203 15988
rect 14263 16164 14321 16176
rect 14263 15988 14275 16164
rect 14309 15988 14321 16164
rect 14263 15976 14321 15988
rect 14380 16164 14438 16176
rect 13488 15822 13546 15834
rect 14380 15788 14392 16164
rect 14426 15788 14438 16164
rect 14380 15776 14438 15788
rect 14498 16164 14556 16176
rect 14498 15788 14510 16164
rect 14544 15788 14556 16164
rect 14498 15776 14556 15788
rect 14616 16164 14674 16176
rect 14616 15788 14628 16164
rect 14662 15788 14674 16164
rect 15593 16164 15651 16176
rect 15593 15988 15605 16164
rect 15639 15988 15651 16164
rect 15593 15976 15651 15988
rect 15711 16164 15769 16176
rect 15711 15988 15723 16164
rect 15757 15988 15769 16164
rect 15711 15976 15769 15988
rect 15828 16164 15886 16176
rect 14616 15776 14674 15788
rect 15828 15788 15840 16164
rect 15874 15788 15886 16164
rect 15828 15776 15886 15788
rect 15946 16164 16004 16176
rect 15946 15788 15958 16164
rect 15992 15788 16004 16164
rect 15946 15776 16004 15788
rect 16064 16164 16122 16176
rect 43052 16826 43110 16838
rect 43052 16650 43064 16826
rect 43098 16650 43110 16826
rect 43052 16638 43110 16650
rect 43170 16826 43228 16838
rect 43170 16650 43182 16826
rect 43216 16650 43228 16826
rect 43170 16638 43228 16650
rect 43287 16826 43345 16838
rect 16064 15788 16076 16164
rect 16110 15788 16122 16164
rect 17091 16162 17149 16174
rect 17091 15986 17103 16162
rect 17137 15986 17149 16162
rect 17091 15974 17149 15986
rect 17209 16162 17267 16174
rect 17209 15986 17221 16162
rect 17255 15986 17267 16162
rect 17209 15974 17267 15986
rect 17326 16162 17384 16174
rect 16064 15776 16122 15788
rect 17326 15786 17338 16162
rect 17372 15786 17384 16162
rect 17326 15774 17384 15786
rect 17444 16162 17502 16174
rect 17444 15786 17456 16162
rect 17490 15786 17502 16162
rect 17444 15774 17502 15786
rect 17562 16162 17620 16174
rect 17562 15786 17574 16162
rect 17608 15786 17620 16162
rect 18539 16162 18597 16174
rect 18539 15986 18551 16162
rect 18585 15986 18597 16162
rect 18539 15974 18597 15986
rect 18657 16162 18715 16174
rect 18657 15986 18669 16162
rect 18703 15986 18715 16162
rect 18657 15974 18715 15986
rect 18774 16162 18832 16174
rect 17562 15774 17620 15786
rect 18774 15786 18786 16162
rect 18820 15786 18832 16162
rect 18774 15774 18832 15786
rect 18892 16162 18950 16174
rect 18892 15786 18904 16162
rect 18938 15786 18950 16162
rect 18892 15774 18950 15786
rect 19010 16162 19068 16174
rect 19010 15786 19022 16162
rect 19056 15786 19068 16162
rect 20059 16164 20117 16176
rect 20059 15988 20071 16164
rect 20105 15988 20117 16164
rect 20059 15976 20117 15988
rect 20177 16164 20235 16176
rect 20177 15988 20189 16164
rect 20223 15988 20235 16164
rect 20177 15976 20235 15988
rect 20294 16164 20352 16176
rect 19010 15774 19068 15786
rect 20294 15788 20306 16164
rect 20340 15788 20352 16164
rect 20294 15776 20352 15788
rect 20412 16164 20470 16176
rect 20412 15788 20424 16164
rect 20458 15788 20470 16164
rect 20412 15776 20470 15788
rect 20530 16164 20588 16176
rect 20530 15788 20542 16164
rect 20576 15788 20588 16164
rect 21507 16164 21565 16176
rect 21507 15988 21519 16164
rect 21553 15988 21565 16164
rect 21507 15976 21565 15988
rect 21625 16164 21683 16176
rect 21625 15988 21637 16164
rect 21671 15988 21683 16164
rect 21625 15976 21683 15988
rect 21742 16164 21800 16176
rect 20530 15776 20588 15788
rect 21742 15788 21754 16164
rect 21788 15788 21800 16164
rect 21742 15776 21800 15788
rect 21860 16164 21918 16176
rect 21860 15788 21872 16164
rect 21906 15788 21918 16164
rect 21860 15776 21918 15788
rect 21978 16164 22036 16176
rect 21978 15788 21990 16164
rect 22024 15788 22036 16164
rect 23005 16162 23063 16174
rect 23005 15986 23017 16162
rect 23051 15986 23063 16162
rect 23005 15974 23063 15986
rect 23123 16162 23181 16174
rect 23123 15986 23135 16162
rect 23169 15986 23181 16162
rect 23123 15974 23181 15986
rect 23240 16162 23298 16174
rect 21978 15776 22036 15788
rect 23240 15786 23252 16162
rect 23286 15786 23298 16162
rect 23240 15774 23298 15786
rect 23358 16162 23416 16174
rect 23358 15786 23370 16162
rect 23404 15786 23416 16162
rect 23358 15774 23416 15786
rect 23476 16162 23534 16174
rect 23476 15786 23488 16162
rect 23522 15786 23534 16162
rect 24453 16162 24511 16174
rect 24453 15986 24465 16162
rect 24499 15986 24511 16162
rect 24453 15974 24511 15986
rect 24571 16162 24629 16174
rect 24571 15986 24583 16162
rect 24617 15986 24629 16162
rect 24571 15974 24629 15986
rect 24688 16162 24746 16174
rect 23476 15774 23534 15786
rect 24688 15786 24700 16162
rect 24734 15786 24746 16162
rect 24688 15774 24746 15786
rect 24806 16162 24864 16174
rect 24806 15786 24818 16162
rect 24852 15786 24864 16162
rect 24806 15774 24864 15786
rect 24924 16162 24982 16174
rect 24924 15786 24936 16162
rect 24970 15786 24982 16162
rect 24924 15774 24982 15786
rect 43287 16450 43299 16826
rect 43333 16450 43345 16826
rect 43287 16438 43345 16450
rect 43405 16826 43463 16838
rect 43405 16450 43417 16826
rect 43451 16450 43463 16826
rect 43405 16438 43463 16450
rect 43523 16826 43581 16838
rect 43523 16450 43535 16826
rect 43569 16450 43581 16826
rect 49610 16822 49668 16834
rect 49610 16646 49622 16822
rect 49656 16646 49668 16822
rect 49610 16634 49668 16646
rect 49728 16822 49786 16834
rect 49728 16646 49740 16822
rect 49774 16646 49786 16822
rect 49728 16634 49786 16646
rect 49845 16822 49903 16834
rect 43523 16438 43581 16450
rect 38857 15421 38915 15433
rect 38857 15245 38869 15421
rect 38903 15245 38915 15421
rect 38857 15233 38915 15245
rect 38975 15421 39033 15433
rect 38975 15245 38987 15421
rect 39021 15245 39033 15421
rect 38975 15233 39033 15245
rect 39381 15421 39439 15433
rect 39381 15045 39393 15421
rect 39427 15045 39439 15421
rect 39381 15033 39439 15045
rect 39499 15421 39557 15433
rect 39499 15045 39511 15421
rect 39545 15045 39557 15421
rect 39499 15033 39557 15045
rect 39617 15421 39675 15433
rect 39617 15045 39629 15421
rect 39663 15045 39675 15421
rect 39617 15033 39675 15045
rect 39735 15421 39793 15433
rect 39735 15045 39747 15421
rect 39781 15045 39793 15421
rect 39735 15033 39793 15045
rect 39853 15421 39911 15433
rect 39853 15045 39865 15421
rect 39899 15045 39911 15421
rect 40155 15421 40213 15433
rect 40155 15245 40167 15421
rect 40201 15245 40213 15421
rect 40155 15233 40213 15245
rect 40273 15421 40331 15433
rect 40273 15245 40285 15421
rect 40319 15245 40331 15421
rect 40273 15233 40331 15245
rect 40755 15421 40813 15433
rect 40755 15245 40767 15421
rect 40801 15245 40813 15421
rect 40755 15233 40813 15245
rect 40873 15421 40931 15433
rect 40873 15245 40885 15421
rect 40919 15245 40931 15421
rect 40873 15233 40931 15245
rect 41279 15421 41337 15433
rect 39853 15033 39911 15045
rect 41279 15045 41291 15421
rect 41325 15045 41337 15421
rect 41279 15033 41337 15045
rect 41397 15421 41455 15433
rect 41397 15045 41409 15421
rect 41443 15045 41455 15421
rect 41397 15033 41455 15045
rect 41515 15421 41573 15433
rect 41515 15045 41527 15421
rect 41561 15045 41573 15421
rect 41515 15033 41573 15045
rect 41633 15421 41691 15433
rect 41633 15045 41645 15421
rect 41679 15045 41691 15421
rect 41633 15033 41691 15045
rect 41751 15421 41809 15433
rect 41751 15045 41763 15421
rect 41797 15045 41809 15421
rect 42053 15421 42111 15433
rect 42053 15245 42065 15421
rect 42099 15245 42111 15421
rect 42053 15233 42111 15245
rect 42171 15421 42229 15433
rect 42171 15245 42183 15421
rect 42217 15245 42229 15421
rect 42171 15233 42229 15245
rect 49845 16446 49857 16822
rect 49891 16446 49903 16822
rect 49845 16434 49903 16446
rect 49963 16822 50021 16834
rect 49963 16446 49975 16822
rect 50009 16446 50021 16822
rect 49963 16434 50021 16446
rect 50081 16822 50139 16834
rect 50081 16446 50093 16822
rect 50127 16446 50139 16822
rect 56144 16827 56202 16839
rect 56144 16651 56156 16827
rect 56190 16651 56202 16827
rect 56144 16639 56202 16651
rect 56262 16827 56320 16839
rect 56262 16651 56274 16827
rect 56308 16651 56320 16827
rect 56262 16639 56320 16651
rect 56379 16827 56437 16839
rect 50081 16434 50139 16446
rect 45415 15417 45473 15429
rect 45415 15241 45427 15417
rect 45461 15241 45473 15417
rect 43057 15222 43115 15234
rect 41751 15033 41809 15045
rect 43057 15046 43069 15222
rect 43103 15046 43115 15222
rect 43057 15034 43115 15046
rect 43175 15222 43233 15234
rect 43175 15046 43187 15222
rect 43221 15046 43233 15222
rect 43175 15034 43233 15046
rect 43292 15222 43350 15234
rect 1366 13513 1424 13525
rect 1366 13337 1378 13513
rect 1412 13337 1424 13513
rect 1366 13325 1424 13337
rect 1484 13513 1620 13525
rect 1484 13337 1496 13513
rect 1530 13337 1574 13513
rect 1484 13325 1574 13337
rect 1562 13137 1574 13325
rect 1608 13137 1620 13513
rect 1562 13125 1620 13137
rect 1680 13513 1738 13525
rect 1680 13137 1692 13513
rect 1726 13137 1738 13513
rect 1680 13125 1738 13137
rect 1798 13513 1856 13525
rect 1798 13137 1810 13513
rect 1844 13137 1856 13513
rect 1798 13125 1856 13137
rect 1916 13513 1974 13525
rect 1916 13137 1928 13513
rect 1962 13137 1974 13513
rect 1916 13125 1974 13137
rect 2034 13513 2166 13525
rect 2034 13137 2046 13513
rect 2080 13337 2120 13513
rect 2154 13337 2166 13513
rect 2080 13325 2166 13337
rect 2226 13513 2284 13525
rect 2226 13337 2238 13513
rect 2272 13337 2284 13513
rect 2226 13325 2284 13337
rect 4510 13513 4568 13525
rect 4510 13337 4522 13513
rect 4556 13337 4568 13513
rect 4510 13325 4568 13337
rect 4628 13513 4764 13525
rect 4628 13337 4640 13513
rect 4674 13337 4718 13513
rect 4628 13325 4718 13337
rect 2080 13137 2092 13325
rect 2034 13125 2092 13137
rect 4706 13137 4718 13325
rect 4752 13137 4764 13513
rect 4706 13125 4764 13137
rect 4824 13513 4882 13525
rect 4824 13137 4836 13513
rect 4870 13137 4882 13513
rect 4824 13125 4882 13137
rect 4942 13513 5000 13525
rect 4942 13137 4954 13513
rect 4988 13137 5000 13513
rect 4942 13125 5000 13137
rect 5060 13513 5118 13525
rect 5060 13137 5072 13513
rect 5106 13137 5118 13513
rect 5060 13125 5118 13137
rect 5178 13513 5310 13525
rect 5178 13137 5190 13513
rect 5224 13337 5264 13513
rect 5298 13337 5310 13513
rect 5224 13325 5310 13337
rect 5370 13513 5428 13525
rect 43292 14846 43304 15222
rect 43338 14846 43350 15222
rect 43292 14834 43350 14846
rect 43410 15222 43468 15234
rect 43410 14846 43422 15222
rect 43456 14846 43468 15222
rect 43410 14834 43468 14846
rect 43528 15222 43586 15234
rect 45415 15229 45473 15241
rect 45533 15417 45591 15429
rect 45533 15241 45545 15417
rect 45579 15241 45591 15417
rect 45533 15229 45591 15241
rect 45939 15417 45997 15429
rect 43528 14846 43540 15222
rect 43574 14846 43586 15222
rect 45939 15041 45951 15417
rect 45985 15041 45997 15417
rect 45939 15029 45997 15041
rect 46057 15417 46115 15429
rect 46057 15041 46069 15417
rect 46103 15041 46115 15417
rect 46057 15029 46115 15041
rect 46175 15417 46233 15429
rect 46175 15041 46187 15417
rect 46221 15041 46233 15417
rect 46175 15029 46233 15041
rect 46293 15417 46351 15429
rect 46293 15041 46305 15417
rect 46339 15041 46351 15417
rect 46293 15029 46351 15041
rect 46411 15417 46469 15429
rect 46411 15041 46423 15417
rect 46457 15041 46469 15417
rect 46713 15417 46771 15429
rect 46713 15241 46725 15417
rect 46759 15241 46771 15417
rect 46713 15229 46771 15241
rect 46831 15417 46889 15429
rect 46831 15241 46843 15417
rect 46877 15241 46889 15417
rect 46831 15229 46889 15241
rect 47313 15417 47371 15429
rect 47313 15241 47325 15417
rect 47359 15241 47371 15417
rect 47313 15229 47371 15241
rect 47431 15417 47489 15429
rect 47431 15241 47443 15417
rect 47477 15241 47489 15417
rect 47431 15229 47489 15241
rect 47837 15417 47895 15429
rect 46411 15029 46469 15041
rect 47837 15041 47849 15417
rect 47883 15041 47895 15417
rect 47837 15029 47895 15041
rect 47955 15417 48013 15429
rect 47955 15041 47967 15417
rect 48001 15041 48013 15417
rect 47955 15029 48013 15041
rect 48073 15417 48131 15429
rect 48073 15041 48085 15417
rect 48119 15041 48131 15417
rect 48073 15029 48131 15041
rect 48191 15417 48249 15429
rect 48191 15041 48203 15417
rect 48237 15041 48249 15417
rect 48191 15029 48249 15041
rect 48309 15417 48367 15429
rect 48309 15041 48321 15417
rect 48355 15041 48367 15417
rect 48611 15417 48669 15429
rect 48611 15241 48623 15417
rect 48657 15241 48669 15417
rect 48611 15229 48669 15241
rect 48729 15417 48787 15429
rect 48729 15241 48741 15417
rect 48775 15241 48787 15417
rect 48729 15229 48787 15241
rect 56379 16451 56391 16827
rect 56425 16451 56437 16827
rect 56379 16439 56437 16451
rect 56497 16827 56555 16839
rect 56497 16451 56509 16827
rect 56543 16451 56555 16827
rect 56497 16439 56555 16451
rect 56615 16827 56673 16839
rect 56615 16451 56627 16827
rect 56661 16451 56673 16827
rect 71846 17419 72246 17431
rect 71846 17385 71858 17419
rect 72234 17385 72246 17419
rect 71846 17373 72246 17385
rect 71846 17341 72046 17373
rect 71846 17307 71858 17341
rect 72034 17307 72046 17341
rect 71846 17295 72046 17307
rect 62657 16830 62715 16842
rect 62657 16654 62669 16830
rect 62703 16654 62715 16830
rect 62657 16642 62715 16654
rect 62775 16830 62833 16842
rect 62775 16654 62787 16830
rect 62821 16654 62833 16830
rect 62775 16642 62833 16654
rect 62892 16830 62950 16842
rect 56615 16439 56673 16451
rect 51949 15422 52007 15434
rect 51949 15246 51961 15422
rect 51995 15246 52007 15422
rect 51949 15234 52007 15246
rect 52067 15422 52125 15434
rect 52067 15246 52079 15422
rect 52113 15246 52125 15422
rect 52067 15234 52125 15246
rect 52473 15422 52531 15434
rect 49615 15218 49673 15230
rect 48309 15029 48367 15041
rect 49615 15042 49627 15218
rect 49661 15042 49673 15218
rect 49615 15030 49673 15042
rect 49733 15218 49791 15230
rect 49733 15042 49745 15218
rect 49779 15042 49791 15218
rect 49733 15030 49791 15042
rect 49850 15218 49908 15230
rect 43528 14834 43586 14846
rect 49850 14842 49862 15218
rect 49896 14842 49908 15218
rect 49850 14830 49908 14842
rect 49968 15218 50026 15230
rect 49968 14842 49980 15218
rect 50014 14842 50026 15218
rect 49968 14830 50026 14842
rect 50086 15218 50144 15230
rect 50086 14842 50098 15218
rect 50132 14842 50144 15218
rect 52473 15046 52485 15422
rect 52519 15046 52531 15422
rect 52473 15034 52531 15046
rect 52591 15422 52649 15434
rect 52591 15046 52603 15422
rect 52637 15046 52649 15422
rect 52591 15034 52649 15046
rect 52709 15422 52767 15434
rect 52709 15046 52721 15422
rect 52755 15046 52767 15422
rect 52709 15034 52767 15046
rect 52827 15422 52885 15434
rect 52827 15046 52839 15422
rect 52873 15046 52885 15422
rect 52827 15034 52885 15046
rect 52945 15422 53003 15434
rect 52945 15046 52957 15422
rect 52991 15046 53003 15422
rect 53247 15422 53305 15434
rect 53247 15246 53259 15422
rect 53293 15246 53305 15422
rect 53247 15234 53305 15246
rect 53365 15422 53423 15434
rect 53365 15246 53377 15422
rect 53411 15246 53423 15422
rect 53365 15234 53423 15246
rect 53847 15422 53905 15434
rect 53847 15246 53859 15422
rect 53893 15246 53905 15422
rect 53847 15234 53905 15246
rect 53965 15422 54023 15434
rect 53965 15246 53977 15422
rect 54011 15246 54023 15422
rect 53965 15234 54023 15246
rect 54371 15422 54429 15434
rect 52945 15034 53003 15046
rect 54371 15046 54383 15422
rect 54417 15046 54429 15422
rect 54371 15034 54429 15046
rect 54489 15422 54547 15434
rect 54489 15046 54501 15422
rect 54535 15046 54547 15422
rect 54489 15034 54547 15046
rect 54607 15422 54665 15434
rect 54607 15046 54619 15422
rect 54653 15046 54665 15422
rect 54607 15034 54665 15046
rect 54725 15422 54783 15434
rect 54725 15046 54737 15422
rect 54771 15046 54783 15422
rect 54725 15034 54783 15046
rect 54843 15422 54901 15434
rect 54843 15046 54855 15422
rect 54889 15046 54901 15422
rect 55145 15422 55203 15434
rect 55145 15246 55157 15422
rect 55191 15246 55203 15422
rect 55145 15234 55203 15246
rect 55263 15422 55321 15434
rect 55263 15246 55275 15422
rect 55309 15246 55321 15422
rect 55263 15234 55321 15246
rect 62892 16454 62904 16830
rect 62938 16454 62950 16830
rect 62892 16442 62950 16454
rect 63010 16830 63068 16842
rect 63010 16454 63022 16830
rect 63056 16454 63068 16830
rect 63010 16442 63068 16454
rect 63128 16830 63186 16842
rect 63128 16454 63140 16830
rect 63174 16454 63186 16830
rect 63128 16442 63186 16454
rect 71846 17223 72046 17235
rect 71846 17189 71858 17223
rect 72034 17189 72046 17223
rect 71846 17177 72046 17189
rect 58462 15425 58520 15437
rect 58462 15249 58474 15425
rect 58508 15249 58520 15425
rect 58462 15237 58520 15249
rect 58580 15425 58638 15437
rect 58580 15249 58592 15425
rect 58626 15249 58638 15425
rect 58580 15237 58638 15249
rect 58986 15425 59044 15437
rect 56149 15223 56207 15235
rect 54843 15034 54901 15046
rect 56149 15047 56161 15223
rect 56195 15047 56207 15223
rect 56149 15035 56207 15047
rect 56267 15223 56325 15235
rect 56267 15047 56279 15223
rect 56313 15047 56325 15223
rect 56267 15035 56325 15047
rect 56384 15223 56442 15235
rect 50086 14830 50144 14842
rect 56384 14847 56396 15223
rect 56430 14847 56442 15223
rect 56384 14835 56442 14847
rect 56502 15223 56560 15235
rect 56502 14847 56514 15223
rect 56548 14847 56560 15223
rect 56502 14835 56560 14847
rect 56620 15223 56678 15235
rect 56620 14847 56632 15223
rect 56666 14847 56678 15223
rect 58986 15049 58998 15425
rect 59032 15049 59044 15425
rect 58986 15037 59044 15049
rect 59104 15425 59162 15437
rect 59104 15049 59116 15425
rect 59150 15049 59162 15425
rect 59104 15037 59162 15049
rect 59222 15425 59280 15437
rect 59222 15049 59234 15425
rect 59268 15049 59280 15425
rect 59222 15037 59280 15049
rect 59340 15425 59398 15437
rect 59340 15049 59352 15425
rect 59386 15049 59398 15425
rect 59340 15037 59398 15049
rect 59458 15425 59516 15437
rect 59458 15049 59470 15425
rect 59504 15049 59516 15425
rect 59760 15425 59818 15437
rect 59760 15249 59772 15425
rect 59806 15249 59818 15425
rect 59760 15237 59818 15249
rect 59878 15425 59936 15437
rect 59878 15249 59890 15425
rect 59924 15249 59936 15425
rect 59878 15237 59936 15249
rect 60360 15425 60418 15437
rect 60360 15249 60372 15425
rect 60406 15249 60418 15425
rect 60360 15237 60418 15249
rect 60478 15425 60536 15437
rect 60478 15249 60490 15425
rect 60524 15249 60536 15425
rect 60478 15237 60536 15249
rect 60884 15425 60942 15437
rect 59458 15037 59516 15049
rect 60884 15049 60896 15425
rect 60930 15049 60942 15425
rect 60884 15037 60942 15049
rect 61002 15425 61060 15437
rect 61002 15049 61014 15425
rect 61048 15049 61060 15425
rect 61002 15037 61060 15049
rect 61120 15425 61178 15437
rect 61120 15049 61132 15425
rect 61166 15049 61178 15425
rect 61120 15037 61178 15049
rect 61238 15425 61296 15437
rect 61238 15049 61250 15425
rect 61284 15049 61296 15425
rect 61238 15037 61296 15049
rect 61356 15425 61414 15437
rect 61356 15049 61368 15425
rect 61402 15049 61414 15425
rect 61658 15425 61716 15437
rect 61658 15249 61670 15425
rect 61704 15249 61716 15425
rect 61658 15237 61716 15249
rect 61776 15425 61834 15437
rect 61776 15249 61788 15425
rect 61822 15249 61834 15425
rect 61776 15237 61834 15249
rect 62662 15226 62720 15238
rect 61356 15037 61414 15049
rect 62662 15050 62674 15226
rect 62708 15050 62720 15226
rect 62662 15038 62720 15050
rect 62780 15226 62838 15238
rect 62780 15050 62792 15226
rect 62826 15050 62838 15226
rect 62780 15038 62838 15050
rect 62897 15226 62955 15238
rect 56620 14835 56678 14847
rect 62897 14850 62909 15226
rect 62943 14850 62955 15226
rect 62897 14838 62955 14850
rect 63015 15226 63073 15238
rect 63015 14850 63027 15226
rect 63061 14850 63073 15226
rect 63015 14838 63073 14850
rect 63133 15226 63191 15238
rect 63133 14850 63145 15226
rect 63179 14850 63191 15226
rect 63133 14838 63191 14850
rect 71842 14951 72042 14963
rect 71842 14917 71854 14951
rect 72030 14917 72042 14951
rect 71842 14905 72042 14917
rect 71842 14833 72042 14845
rect 71842 14799 71854 14833
rect 72030 14799 72042 14833
rect 71842 14771 72042 14799
rect 71842 14759 72242 14771
rect 71842 14725 71854 14759
rect 72230 14725 72242 14759
rect 71842 14713 72242 14725
rect 5370 13337 5382 13513
rect 5416 13337 5428 13513
rect 5370 13325 5428 13337
rect 7642 13509 7700 13521
rect 7642 13333 7654 13509
rect 7688 13333 7700 13509
rect 5224 13137 5236 13325
rect 7642 13321 7700 13333
rect 7760 13509 7896 13521
rect 7760 13333 7772 13509
rect 7806 13333 7850 13509
rect 7760 13321 7850 13333
rect 5178 13125 5236 13137
rect 7838 13133 7850 13321
rect 7884 13133 7896 13509
rect 7838 13121 7896 13133
rect 7956 13509 8014 13521
rect 7956 13133 7968 13509
rect 8002 13133 8014 13509
rect 7956 13121 8014 13133
rect 8074 13509 8132 13521
rect 8074 13133 8086 13509
rect 8120 13133 8132 13509
rect 8074 13121 8132 13133
rect 8192 13509 8250 13521
rect 8192 13133 8204 13509
rect 8238 13133 8250 13509
rect 8192 13121 8250 13133
rect 8310 13509 8442 13521
rect 8310 13133 8322 13509
rect 8356 13333 8396 13509
rect 8430 13333 8442 13509
rect 8356 13321 8442 13333
rect 8502 13509 8560 13521
rect 8502 13333 8514 13509
rect 8548 13333 8560 13509
rect 8502 13321 8560 13333
rect 10786 13509 10844 13521
rect 10786 13333 10798 13509
rect 10832 13333 10844 13509
rect 10786 13321 10844 13333
rect 10904 13509 11040 13521
rect 10904 13333 10916 13509
rect 10950 13333 10994 13509
rect 10904 13321 10994 13333
rect 8356 13133 8368 13321
rect 8310 13121 8368 13133
rect 10982 13133 10994 13321
rect 11028 13133 11040 13509
rect 10982 13121 11040 13133
rect 11100 13509 11158 13521
rect 11100 13133 11112 13509
rect 11146 13133 11158 13509
rect 11100 13121 11158 13133
rect 11218 13509 11276 13521
rect 11218 13133 11230 13509
rect 11264 13133 11276 13509
rect 11218 13121 11276 13133
rect 11336 13509 11394 13521
rect 11336 13133 11348 13509
rect 11382 13133 11394 13509
rect 11336 13121 11394 13133
rect 11454 13509 11586 13521
rect 11454 13133 11466 13509
rect 11500 13333 11540 13509
rect 11574 13333 11586 13509
rect 11500 13321 11586 13333
rect 11646 13509 11704 13521
rect 11646 13333 11658 13509
rect 11692 13333 11704 13509
rect 11646 13321 11704 13333
rect 13988 13513 14046 13525
rect 13988 13337 14000 13513
rect 14034 13337 14046 13513
rect 13988 13325 14046 13337
rect 14106 13513 14242 13525
rect 14106 13337 14118 13513
rect 14152 13337 14196 13513
rect 14106 13325 14196 13337
rect 11500 13133 11512 13321
rect 11454 13121 11512 13133
rect 14184 13137 14196 13325
rect 14230 13137 14242 13513
rect 14184 13125 14242 13137
rect 14302 13513 14360 13525
rect 14302 13137 14314 13513
rect 14348 13137 14360 13513
rect 14302 13125 14360 13137
rect 14420 13513 14478 13525
rect 14420 13137 14432 13513
rect 14466 13137 14478 13513
rect 14420 13125 14478 13137
rect 14538 13513 14596 13525
rect 14538 13137 14550 13513
rect 14584 13137 14596 13513
rect 14538 13125 14596 13137
rect 14656 13513 14788 13525
rect 14656 13137 14668 13513
rect 14702 13337 14742 13513
rect 14776 13337 14788 13513
rect 14702 13325 14788 13337
rect 14848 13513 14906 13525
rect 14848 13337 14860 13513
rect 14894 13337 14906 13513
rect 14848 13325 14906 13337
rect 17132 13513 17190 13525
rect 17132 13337 17144 13513
rect 17178 13337 17190 13513
rect 17132 13325 17190 13337
rect 17250 13513 17386 13525
rect 17250 13337 17262 13513
rect 17296 13337 17340 13513
rect 17250 13325 17340 13337
rect 14702 13137 14714 13325
rect 14656 13125 14714 13137
rect 17328 13137 17340 13325
rect 17374 13137 17386 13513
rect 17328 13125 17386 13137
rect 17446 13513 17504 13525
rect 17446 13137 17458 13513
rect 17492 13137 17504 13513
rect 17446 13125 17504 13137
rect 17564 13513 17622 13525
rect 17564 13137 17576 13513
rect 17610 13137 17622 13513
rect 17564 13125 17622 13137
rect 17682 13513 17740 13525
rect 17682 13137 17694 13513
rect 17728 13137 17740 13513
rect 17682 13125 17740 13137
rect 17800 13513 17932 13525
rect 17800 13137 17812 13513
rect 17846 13337 17886 13513
rect 17920 13337 17932 13513
rect 17846 13325 17932 13337
rect 17992 13513 18050 13525
rect 71842 14641 72242 14653
rect 71842 14607 71854 14641
rect 72230 14607 72242 14641
rect 71842 14595 72242 14607
rect 71842 14523 72242 14535
rect 71842 14489 71854 14523
rect 72230 14489 72242 14523
rect 71842 14477 72242 14489
rect 71842 14405 72242 14417
rect 71842 14371 71854 14405
rect 72230 14371 72242 14405
rect 71842 14359 72242 14371
rect 71842 14287 72242 14299
rect 71842 14253 71854 14287
rect 72230 14253 72242 14287
rect 71842 14241 72242 14253
rect 71842 14209 72042 14241
rect 71842 14175 71854 14209
rect 72030 14175 72042 14209
rect 71842 14163 72042 14175
rect 17992 13337 18004 13513
rect 18038 13337 18050 13513
rect 17992 13325 18050 13337
rect 20264 13509 20322 13521
rect 20264 13333 20276 13509
rect 20310 13333 20322 13509
rect 17846 13137 17858 13325
rect 20264 13321 20322 13333
rect 20382 13509 20518 13521
rect 20382 13333 20394 13509
rect 20428 13333 20472 13509
rect 20382 13321 20472 13333
rect 17800 13125 17858 13137
rect 20460 13133 20472 13321
rect 20506 13133 20518 13509
rect 20460 13121 20518 13133
rect 20578 13509 20636 13521
rect 20578 13133 20590 13509
rect 20624 13133 20636 13509
rect 20578 13121 20636 13133
rect 20696 13509 20754 13521
rect 20696 13133 20708 13509
rect 20742 13133 20754 13509
rect 20696 13121 20754 13133
rect 20814 13509 20872 13521
rect 20814 13133 20826 13509
rect 20860 13133 20872 13509
rect 20814 13121 20872 13133
rect 20932 13509 21064 13521
rect 20932 13133 20944 13509
rect 20978 13333 21018 13509
rect 21052 13333 21064 13509
rect 20978 13321 21064 13333
rect 21124 13509 21182 13521
rect 21124 13333 21136 13509
rect 21170 13333 21182 13509
rect 21124 13321 21182 13333
rect 23408 13509 23466 13521
rect 23408 13333 23420 13509
rect 23454 13333 23466 13509
rect 23408 13321 23466 13333
rect 23526 13509 23662 13521
rect 23526 13333 23538 13509
rect 23572 13333 23616 13509
rect 23526 13321 23616 13333
rect 20978 13133 20990 13321
rect 20932 13121 20990 13133
rect 23604 13133 23616 13321
rect 23650 13133 23662 13509
rect 23604 13121 23662 13133
rect 23722 13509 23780 13521
rect 23722 13133 23734 13509
rect 23768 13133 23780 13509
rect 23722 13121 23780 13133
rect 23840 13509 23898 13521
rect 23840 13133 23852 13509
rect 23886 13133 23898 13509
rect 23840 13121 23898 13133
rect 23958 13509 24016 13521
rect 23958 13133 23970 13509
rect 24004 13133 24016 13509
rect 23958 13121 24016 13133
rect 24076 13509 24208 13521
rect 24076 13133 24088 13509
rect 24122 13333 24162 13509
rect 24196 13333 24208 13509
rect 24122 13321 24208 13333
rect 24268 13509 24326 13521
rect 24268 13333 24280 13509
rect 24314 13333 24326 13509
rect 24268 13321 24326 13333
rect 24122 13133 24134 13321
rect 71842 14091 72042 14103
rect 71842 14057 71854 14091
rect 72030 14057 72042 14091
rect 71842 14045 72042 14057
rect 24076 13121 24134 13133
rect 31379 13043 31579 13055
rect 31379 13009 31391 13043
rect 31567 13009 31579 13043
rect 31379 12997 31579 13009
rect 31379 12925 31579 12937
rect 31379 12891 31391 12925
rect 31567 12891 31579 12925
rect 31379 12879 31579 12891
rect 31379 12623 31779 12635
rect 31379 12589 31391 12623
rect 31767 12589 31779 12623
rect 31379 12577 31779 12589
rect 31379 12505 31779 12517
rect 31379 12471 31391 12505
rect 31767 12471 31779 12505
rect 31379 12459 31779 12471
rect 31379 12387 31779 12399
rect 31379 12353 31391 12387
rect 31767 12353 31779 12387
rect 31379 12341 31779 12353
rect 1366 10779 1424 10791
rect 1366 10603 1378 10779
rect 1412 10603 1424 10779
rect 1366 10591 1424 10603
rect 1484 10779 1620 10791
rect 1484 10603 1496 10779
rect 1530 10603 1574 10779
rect 1484 10591 1574 10603
rect 1562 10403 1574 10591
rect 1608 10403 1620 10779
rect 1562 10391 1620 10403
rect 1680 10779 1738 10791
rect 1680 10403 1692 10779
rect 1726 10403 1738 10779
rect 1680 10391 1738 10403
rect 1798 10779 1856 10791
rect 1798 10403 1810 10779
rect 1844 10403 1856 10779
rect 1798 10391 1856 10403
rect 1916 10779 1974 10791
rect 1916 10403 1928 10779
rect 1962 10403 1974 10779
rect 1916 10391 1974 10403
rect 2034 10779 2166 10791
rect 2034 10403 2046 10779
rect 2080 10603 2120 10779
rect 2154 10603 2166 10779
rect 2080 10591 2166 10603
rect 2226 10779 2284 10791
rect 2226 10603 2238 10779
rect 2272 10603 2284 10779
rect 2226 10591 2284 10603
rect 4510 10779 4568 10791
rect 4510 10603 4522 10779
rect 4556 10603 4568 10779
rect 4510 10591 4568 10603
rect 4628 10779 4764 10791
rect 4628 10603 4640 10779
rect 4674 10603 4718 10779
rect 4628 10591 4718 10603
rect 2080 10403 2092 10591
rect 2034 10391 2092 10403
rect 4706 10403 4718 10591
rect 4752 10403 4764 10779
rect 4706 10391 4764 10403
rect 4824 10779 4882 10791
rect 4824 10403 4836 10779
rect 4870 10403 4882 10779
rect 4824 10391 4882 10403
rect 4942 10779 5000 10791
rect 4942 10403 4954 10779
rect 4988 10403 5000 10779
rect 4942 10391 5000 10403
rect 5060 10779 5118 10791
rect 5060 10403 5072 10779
rect 5106 10403 5118 10779
rect 5060 10391 5118 10403
rect 5178 10779 5310 10791
rect 5178 10403 5190 10779
rect 5224 10603 5264 10779
rect 5298 10603 5310 10779
rect 5224 10591 5310 10603
rect 5370 10779 5428 10791
rect 31379 12269 31779 12281
rect 31379 12235 31391 12269
rect 31767 12235 31779 12269
rect 31379 12223 31779 12235
rect 31379 12151 31779 12163
rect 31379 12117 31391 12151
rect 31767 12117 31779 12151
rect 31379 12105 31779 12117
rect 5370 10603 5382 10779
rect 5416 10603 5428 10779
rect 5370 10591 5428 10603
rect 7642 10775 7700 10787
rect 7642 10599 7654 10775
rect 7688 10599 7700 10775
rect 5224 10403 5236 10591
rect 7642 10587 7700 10599
rect 7760 10775 7896 10787
rect 7760 10599 7772 10775
rect 7806 10599 7850 10775
rect 7760 10587 7850 10599
rect 5178 10391 5236 10403
rect 7838 10399 7850 10587
rect 7884 10399 7896 10775
rect 7838 10387 7896 10399
rect 7956 10775 8014 10787
rect 7956 10399 7968 10775
rect 8002 10399 8014 10775
rect 7956 10387 8014 10399
rect 8074 10775 8132 10787
rect 8074 10399 8086 10775
rect 8120 10399 8132 10775
rect 8074 10387 8132 10399
rect 8192 10775 8250 10787
rect 8192 10399 8204 10775
rect 8238 10399 8250 10775
rect 8192 10387 8250 10399
rect 8310 10775 8442 10787
rect 8310 10399 8322 10775
rect 8356 10599 8396 10775
rect 8430 10599 8442 10775
rect 8356 10587 8442 10599
rect 8502 10775 8560 10787
rect 8502 10599 8514 10775
rect 8548 10599 8560 10775
rect 8502 10587 8560 10599
rect 10786 10775 10844 10787
rect 10786 10599 10798 10775
rect 10832 10599 10844 10775
rect 10786 10587 10844 10599
rect 10904 10775 11040 10787
rect 10904 10599 10916 10775
rect 10950 10599 10994 10775
rect 10904 10587 10994 10599
rect 8356 10399 8368 10587
rect 8310 10387 8368 10399
rect 10982 10399 10994 10587
rect 11028 10399 11040 10775
rect 10982 10387 11040 10399
rect 11100 10775 11158 10787
rect 11100 10399 11112 10775
rect 11146 10399 11158 10775
rect 11100 10387 11158 10399
rect 11218 10775 11276 10787
rect 11218 10399 11230 10775
rect 11264 10399 11276 10775
rect 11218 10387 11276 10399
rect 11336 10775 11394 10787
rect 11336 10399 11348 10775
rect 11382 10399 11394 10775
rect 11336 10387 11394 10399
rect 11454 10775 11586 10787
rect 11454 10399 11466 10775
rect 11500 10599 11540 10775
rect 11574 10599 11586 10775
rect 11500 10587 11586 10599
rect 11646 10775 11704 10787
rect 11646 10599 11658 10775
rect 11692 10599 11704 10775
rect 11646 10587 11704 10599
rect 13988 10779 14046 10791
rect 13988 10603 14000 10779
rect 14034 10603 14046 10779
rect 13988 10591 14046 10603
rect 14106 10779 14242 10791
rect 14106 10603 14118 10779
rect 14152 10603 14196 10779
rect 14106 10591 14196 10603
rect 11500 10399 11512 10587
rect 11454 10387 11512 10399
rect 14184 10403 14196 10591
rect 14230 10403 14242 10779
rect 14184 10391 14242 10403
rect 14302 10779 14360 10791
rect 14302 10403 14314 10779
rect 14348 10403 14360 10779
rect 14302 10391 14360 10403
rect 14420 10779 14478 10791
rect 14420 10403 14432 10779
rect 14466 10403 14478 10779
rect 14420 10391 14478 10403
rect 14538 10779 14596 10791
rect 14538 10403 14550 10779
rect 14584 10403 14596 10779
rect 14538 10391 14596 10403
rect 14656 10779 14788 10791
rect 14656 10403 14668 10779
rect 14702 10603 14742 10779
rect 14776 10603 14788 10779
rect 14702 10591 14788 10603
rect 14848 10779 14906 10791
rect 14848 10603 14860 10779
rect 14894 10603 14906 10779
rect 14848 10591 14906 10603
rect 17132 10779 17190 10791
rect 17132 10603 17144 10779
rect 17178 10603 17190 10779
rect 17132 10591 17190 10603
rect 17250 10779 17386 10791
rect 17250 10603 17262 10779
rect 17296 10603 17340 10779
rect 17250 10591 17340 10603
rect 14702 10403 14714 10591
rect 14656 10391 14714 10403
rect 17328 10403 17340 10591
rect 17374 10403 17386 10779
rect 17328 10391 17386 10403
rect 17446 10779 17504 10791
rect 17446 10403 17458 10779
rect 17492 10403 17504 10779
rect 17446 10391 17504 10403
rect 17564 10779 17622 10791
rect 17564 10403 17576 10779
rect 17610 10403 17622 10779
rect 17564 10391 17622 10403
rect 17682 10779 17740 10791
rect 17682 10403 17694 10779
rect 17728 10403 17740 10779
rect 17682 10391 17740 10403
rect 17800 10779 17932 10791
rect 17800 10403 17812 10779
rect 17846 10603 17886 10779
rect 17920 10603 17932 10779
rect 17846 10591 17932 10603
rect 17992 10779 18050 10791
rect 31379 11745 31579 11757
rect 31379 11711 31391 11745
rect 31567 11711 31579 11745
rect 31379 11699 31579 11711
rect 41795 11700 41853 11712
rect 31379 11627 31579 11639
rect 31379 11593 31391 11627
rect 31567 11593 31579 11627
rect 31379 11581 31579 11593
rect 41795 11324 41807 11700
rect 41841 11324 41853 11700
rect 41795 11312 41853 11324
rect 41913 11700 41971 11712
rect 41913 11324 41925 11700
rect 41959 11324 41971 11700
rect 41913 11312 41971 11324
rect 42031 11700 42089 11712
rect 42031 11324 42043 11700
rect 42077 11324 42089 11700
rect 42148 11700 42206 11712
rect 42148 11524 42160 11700
rect 42194 11524 42206 11700
rect 42148 11512 42206 11524
rect 42266 11700 42324 11712
rect 54998 11720 55056 11732
rect 42266 11524 42278 11700
rect 42312 11524 42324 11700
rect 42266 11512 42324 11524
rect 48344 11699 48402 11711
rect 42031 11312 42089 11324
rect 48344 11323 48356 11699
rect 48390 11323 48402 11699
rect 48344 11311 48402 11323
rect 48462 11699 48520 11711
rect 48462 11323 48474 11699
rect 48508 11323 48520 11699
rect 48462 11311 48520 11323
rect 48580 11699 48638 11711
rect 48580 11323 48592 11699
rect 48626 11323 48638 11699
rect 48697 11699 48755 11711
rect 48697 11523 48709 11699
rect 48743 11523 48755 11699
rect 48697 11511 48755 11523
rect 48815 11699 48873 11711
rect 48815 11523 48827 11699
rect 48861 11523 48873 11699
rect 48815 11511 48873 11523
rect 54998 11344 55010 11720
rect 55044 11344 55056 11720
rect 54998 11332 55056 11344
rect 55116 11720 55174 11732
rect 55116 11344 55128 11720
rect 55162 11344 55174 11720
rect 55116 11332 55174 11344
rect 55234 11720 55292 11732
rect 55234 11344 55246 11720
rect 55280 11344 55292 11720
rect 55351 11720 55409 11732
rect 55351 11544 55363 11720
rect 55397 11544 55409 11720
rect 55351 11532 55409 11544
rect 55469 11720 55527 11732
rect 55469 11544 55481 11720
rect 55515 11544 55527 11720
rect 55469 11532 55527 11544
rect 63651 11553 63709 11565
rect 55234 11332 55292 11344
rect 48580 11311 48638 11323
rect 63651 11177 63663 11553
rect 63697 11177 63709 11553
rect 63651 11165 63709 11177
rect 63769 11553 63827 11565
rect 63769 11177 63781 11553
rect 63815 11177 63827 11553
rect 63769 11165 63827 11177
rect 63887 11553 63945 11565
rect 63887 11177 63899 11553
rect 63933 11177 63945 11553
rect 64004 11553 64062 11565
rect 64004 11377 64016 11553
rect 64050 11377 64062 11553
rect 64004 11365 64062 11377
rect 64122 11553 64180 11565
rect 64122 11377 64134 11553
rect 64168 11377 64180 11553
rect 64122 11365 64180 11377
rect 63887 11165 63945 11177
rect 71842 11807 72042 11819
rect 71842 11773 71854 11807
rect 72030 11773 72042 11807
rect 71842 11761 72042 11773
rect 71842 11689 72042 11701
rect 71842 11655 71854 11689
rect 72030 11655 72042 11689
rect 71842 11627 72042 11655
rect 71842 11615 72242 11627
rect 71842 11581 71854 11615
rect 72230 11581 72242 11615
rect 71842 11569 72242 11581
rect 31377 10975 31577 10987
rect 31377 10941 31389 10975
rect 31565 10941 31577 10975
rect 31377 10929 31577 10941
rect 17992 10603 18004 10779
rect 18038 10603 18050 10779
rect 17992 10591 18050 10603
rect 20264 10775 20322 10787
rect 20264 10599 20276 10775
rect 20310 10599 20322 10775
rect 17846 10403 17858 10591
rect 20264 10587 20322 10599
rect 20382 10775 20518 10787
rect 20382 10599 20394 10775
rect 20428 10599 20472 10775
rect 20382 10587 20472 10599
rect 17800 10391 17858 10403
rect 20460 10399 20472 10587
rect 20506 10399 20518 10775
rect 20460 10387 20518 10399
rect 20578 10775 20636 10787
rect 20578 10399 20590 10775
rect 20624 10399 20636 10775
rect 20578 10387 20636 10399
rect 20696 10775 20754 10787
rect 20696 10399 20708 10775
rect 20742 10399 20754 10775
rect 20696 10387 20754 10399
rect 20814 10775 20872 10787
rect 20814 10399 20826 10775
rect 20860 10399 20872 10775
rect 20814 10387 20872 10399
rect 20932 10775 21064 10787
rect 20932 10399 20944 10775
rect 20978 10599 21018 10775
rect 21052 10599 21064 10775
rect 20978 10587 21064 10599
rect 21124 10775 21182 10787
rect 21124 10599 21136 10775
rect 21170 10599 21182 10775
rect 21124 10587 21182 10599
rect 23408 10775 23466 10787
rect 23408 10599 23420 10775
rect 23454 10599 23466 10775
rect 23408 10587 23466 10599
rect 23526 10775 23662 10787
rect 23526 10599 23538 10775
rect 23572 10599 23616 10775
rect 23526 10587 23616 10599
rect 20978 10399 20990 10587
rect 20932 10387 20990 10399
rect 23604 10399 23616 10587
rect 23650 10399 23662 10775
rect 23604 10387 23662 10399
rect 23722 10775 23780 10787
rect 23722 10399 23734 10775
rect 23768 10399 23780 10775
rect 23722 10387 23780 10399
rect 23840 10775 23898 10787
rect 23840 10399 23852 10775
rect 23886 10399 23898 10775
rect 23840 10387 23898 10399
rect 23958 10775 24016 10787
rect 23958 10399 23970 10775
rect 24004 10399 24016 10775
rect 23958 10387 24016 10399
rect 24076 10775 24208 10787
rect 24076 10399 24088 10775
rect 24122 10599 24162 10775
rect 24196 10599 24208 10775
rect 24122 10587 24208 10599
rect 24268 10775 24326 10787
rect 24268 10599 24280 10775
rect 24314 10599 24326 10775
rect 31377 10857 31577 10869
rect 31377 10823 31389 10857
rect 31565 10823 31577 10857
rect 31377 10811 31577 10823
rect 24268 10587 24326 10599
rect 24122 10399 24134 10587
rect 31377 10555 31777 10567
rect 31377 10521 31389 10555
rect 31765 10521 31777 10555
rect 31377 10509 31777 10521
rect 24076 10387 24134 10399
rect 31377 10437 31777 10449
rect 31377 10403 31389 10437
rect 31765 10403 31777 10437
rect 31377 10391 31777 10403
rect 31377 10319 31777 10331
rect 31377 10285 31389 10319
rect 31765 10285 31777 10319
rect 31377 10273 31777 10285
rect 31377 10201 31777 10213
rect 31377 10167 31389 10201
rect 31765 10167 31777 10201
rect 31377 10155 31777 10167
rect 31377 10083 31777 10095
rect 31377 10049 31389 10083
rect 31765 10049 31777 10083
rect 71842 11497 72242 11509
rect 71842 11463 71854 11497
rect 72230 11463 72242 11497
rect 71842 11451 72242 11463
rect 71842 11379 72242 11391
rect 71842 11345 71854 11379
rect 72230 11345 72242 11379
rect 71842 11333 72242 11345
rect 71842 11261 72242 11273
rect 71842 11227 71854 11261
rect 72230 11227 72242 11261
rect 67252 11145 67310 11157
rect 67252 10769 67264 11145
rect 67298 10769 67310 11145
rect 67252 10757 67310 10769
rect 67370 11145 67428 11157
rect 67370 10769 67382 11145
rect 67416 10769 67428 11145
rect 67370 10757 67428 10769
rect 67488 11145 67546 11157
rect 67488 10769 67500 11145
rect 67534 10769 67546 11145
rect 67605 11145 67663 11157
rect 67605 10969 67617 11145
rect 67651 10969 67663 11145
rect 67605 10957 67663 10969
rect 67723 11145 67781 11157
rect 67723 10969 67735 11145
rect 67769 10969 67781 11145
rect 71842 11215 72242 11227
rect 67723 10957 67781 10969
rect 67488 10757 67546 10769
rect 71842 11143 72242 11155
rect 71842 11109 71854 11143
rect 72230 11109 72242 11143
rect 71842 11097 72242 11109
rect 71842 11065 72042 11097
rect 71842 11031 71854 11065
rect 72030 11031 72042 11065
rect 71842 11019 72042 11031
rect 65347 10360 65405 10372
rect 31377 10037 31777 10049
rect 35131 9800 35189 9812
rect 31377 9677 31577 9689
rect 31377 9643 31389 9677
rect 31565 9643 31577 9677
rect 31377 9631 31577 9643
rect 31377 9559 31577 9571
rect 31377 9525 31389 9559
rect 31565 9525 31577 9559
rect 31377 9513 31577 9525
rect 35131 9424 35143 9800
rect 35177 9424 35189 9800
rect 35131 9412 35189 9424
rect 35249 9800 35307 9812
rect 35249 9424 35261 9800
rect 35295 9424 35307 9800
rect 35249 9412 35307 9424
rect 35367 9800 35425 9812
rect 35367 9424 35379 9800
rect 35413 9424 35425 9800
rect 35484 9800 35542 9812
rect 35484 9624 35496 9800
rect 35530 9624 35542 9800
rect 35484 9612 35542 9624
rect 35602 9800 35660 9812
rect 35602 9624 35614 9800
rect 35648 9624 35660 9800
rect 35602 9612 35660 9624
rect 35367 9412 35425 9424
rect 38021 9533 38079 9545
rect 1376 8047 1434 8059
rect 1376 7871 1388 8047
rect 1422 7871 1434 8047
rect 1376 7859 1434 7871
rect 1494 8047 1630 8059
rect 1494 7871 1506 8047
rect 1540 7871 1584 8047
rect 1494 7859 1584 7871
rect 1572 7671 1584 7859
rect 1618 7671 1630 8047
rect 1572 7659 1630 7671
rect 1690 8047 1748 8059
rect 1690 7671 1702 8047
rect 1736 7671 1748 8047
rect 1690 7659 1748 7671
rect 1808 8047 1866 8059
rect 1808 7671 1820 8047
rect 1854 7671 1866 8047
rect 1808 7659 1866 7671
rect 1926 8047 1984 8059
rect 1926 7671 1938 8047
rect 1972 7671 1984 8047
rect 1926 7659 1984 7671
rect 2044 8047 2176 8059
rect 2044 7671 2056 8047
rect 2090 7871 2130 8047
rect 2164 7871 2176 8047
rect 2090 7859 2176 7871
rect 2236 8047 2294 8059
rect 2236 7871 2248 8047
rect 2282 7871 2294 8047
rect 2236 7859 2294 7871
rect 4520 8047 4578 8059
rect 4520 7871 4532 8047
rect 4566 7871 4578 8047
rect 4520 7859 4578 7871
rect 4638 8047 4774 8059
rect 4638 7871 4650 8047
rect 4684 7871 4728 8047
rect 4638 7859 4728 7871
rect 2090 7671 2102 7859
rect 2044 7659 2102 7671
rect 4716 7671 4728 7859
rect 4762 7671 4774 8047
rect 4716 7659 4774 7671
rect 4834 8047 4892 8059
rect 4834 7671 4846 8047
rect 4880 7671 4892 8047
rect 4834 7659 4892 7671
rect 4952 8047 5010 8059
rect 4952 7671 4964 8047
rect 4998 7671 5010 8047
rect 4952 7659 5010 7671
rect 5070 8047 5128 8059
rect 5070 7671 5082 8047
rect 5116 7671 5128 8047
rect 5070 7659 5128 7671
rect 5188 8047 5320 8059
rect 5188 7671 5200 8047
rect 5234 7871 5274 8047
rect 5308 7871 5320 8047
rect 5234 7859 5320 7871
rect 5380 8047 5438 8059
rect 38021 9157 38033 9533
rect 38067 9157 38079 9533
rect 38021 9145 38079 9157
rect 38139 9533 38197 9545
rect 38139 9157 38151 9533
rect 38185 9157 38197 9533
rect 38139 9145 38197 9157
rect 38257 9533 38315 9545
rect 38257 9157 38269 9533
rect 38303 9157 38315 9533
rect 38374 9533 38432 9545
rect 38374 9357 38386 9533
rect 38420 9357 38432 9533
rect 38374 9345 38432 9357
rect 38492 9533 38550 9545
rect 38492 9357 38504 9533
rect 38538 9357 38550 9533
rect 38492 9345 38550 9357
rect 65347 10184 65359 10360
rect 65393 10184 65405 10360
rect 65347 10172 65405 10184
rect 65465 10360 65523 10372
rect 65465 10184 65477 10360
rect 65511 10184 65523 10360
rect 65465 10172 65523 10184
rect 65767 10360 65825 10372
rect 44570 9621 44628 9633
rect 40019 9259 40077 9271
rect 38257 9145 38315 9157
rect 40019 9083 40031 9259
rect 40065 9083 40077 9259
rect 40019 9071 40077 9083
rect 40137 9259 40195 9271
rect 40137 9083 40149 9259
rect 40183 9083 40195 9259
rect 40137 9071 40195 9083
rect 40255 9259 40313 9271
rect 40255 9083 40267 9259
rect 40301 9083 40313 9259
rect 40255 9071 40313 9083
rect 40373 9259 40431 9271
rect 40373 9083 40385 9259
rect 40419 9083 40431 9259
rect 40373 9071 40431 9083
rect 41161 9263 41219 9275
rect 41161 9087 41173 9263
rect 41207 9087 41219 9263
rect 41161 9075 41219 9087
rect 41279 9263 41337 9275
rect 41279 9087 41291 9263
rect 41325 9087 41337 9263
rect 41279 9075 41337 9087
rect 41397 9263 41455 9275
rect 41397 9087 41409 9263
rect 41443 9087 41455 9263
rect 41397 9075 41455 9087
rect 41515 9263 41573 9275
rect 41515 9087 41527 9263
rect 41561 9087 41573 9263
rect 41515 9075 41573 9087
rect 44570 9245 44582 9621
rect 44616 9245 44628 9621
rect 44570 9233 44628 9245
rect 44688 9621 44746 9633
rect 44688 9245 44700 9621
rect 44734 9245 44746 9621
rect 44688 9233 44746 9245
rect 44806 9621 44864 9633
rect 44806 9245 44818 9621
rect 44852 9245 44864 9621
rect 44923 9621 44981 9633
rect 44923 9445 44935 9621
rect 44969 9445 44981 9621
rect 44923 9433 44981 9445
rect 45041 9621 45099 9633
rect 45041 9445 45053 9621
rect 45087 9445 45099 9621
rect 45041 9433 45099 9445
rect 51224 9553 51282 9565
rect 46568 9347 46626 9359
rect 44806 9233 44864 9245
rect 46568 9171 46580 9347
rect 46614 9171 46626 9347
rect 46568 9159 46626 9171
rect 46686 9347 46744 9359
rect 46686 9171 46698 9347
rect 46732 9171 46744 9347
rect 46686 9159 46744 9171
rect 46804 9347 46862 9359
rect 46804 9171 46816 9347
rect 46850 9171 46862 9347
rect 46804 9159 46862 9171
rect 46922 9347 46980 9359
rect 46922 9171 46934 9347
rect 46968 9171 46980 9347
rect 46922 9159 46980 9171
rect 47710 9351 47768 9363
rect 47710 9175 47722 9351
rect 47756 9175 47768 9351
rect 47710 9163 47768 9175
rect 47828 9351 47886 9363
rect 47828 9175 47840 9351
rect 47874 9175 47886 9351
rect 47828 9163 47886 9175
rect 47946 9351 48004 9363
rect 47946 9175 47958 9351
rect 47992 9175 48004 9351
rect 47946 9163 48004 9175
rect 48064 9351 48122 9363
rect 48064 9175 48076 9351
rect 48110 9175 48122 9351
rect 48064 9163 48122 9175
rect 51224 9177 51236 9553
rect 51270 9177 51282 9553
rect 51224 9165 51282 9177
rect 51342 9553 51400 9565
rect 51342 9177 51354 9553
rect 51388 9177 51400 9553
rect 51342 9165 51400 9177
rect 51460 9553 51518 9565
rect 51460 9177 51472 9553
rect 51506 9177 51518 9553
rect 51577 9553 51635 9565
rect 51577 9377 51589 9553
rect 51623 9377 51635 9553
rect 51577 9365 51635 9377
rect 51695 9553 51753 9565
rect 51695 9377 51707 9553
rect 51741 9377 51753 9553
rect 51695 9365 51753 9377
rect 65767 9984 65779 10360
rect 65813 9984 65825 10360
rect 65767 9972 65825 9984
rect 65885 10360 65943 10372
rect 65885 9984 65897 10360
rect 65931 9984 65943 10360
rect 65885 9972 65943 9984
rect 66003 10360 66061 10372
rect 66003 9984 66015 10360
rect 66049 9984 66061 10360
rect 66003 9972 66061 9984
rect 66121 10360 66179 10372
rect 66121 9984 66133 10360
rect 66167 9984 66179 10360
rect 66121 9972 66179 9984
rect 66239 10360 66297 10372
rect 66239 9984 66251 10360
rect 66285 9984 66297 10360
rect 66645 10360 66703 10372
rect 66645 10184 66657 10360
rect 66691 10184 66703 10360
rect 66645 10172 66703 10184
rect 66763 10360 66821 10372
rect 66763 10184 66775 10360
rect 66809 10184 66821 10360
rect 66763 10172 66821 10184
rect 71842 10947 72042 10959
rect 71842 10913 71854 10947
rect 72030 10913 72042 10947
rect 71842 10901 72042 10913
rect 66239 9972 66297 9984
rect 57849 9621 57907 9633
rect 53222 9279 53280 9291
rect 51460 9165 51518 9177
rect 53222 9103 53234 9279
rect 53268 9103 53280 9279
rect 53222 9091 53280 9103
rect 53340 9279 53398 9291
rect 53340 9103 53352 9279
rect 53386 9103 53398 9279
rect 53340 9091 53398 9103
rect 53458 9279 53516 9291
rect 53458 9103 53470 9279
rect 53504 9103 53516 9279
rect 53458 9091 53516 9103
rect 53576 9279 53634 9291
rect 53576 9103 53588 9279
rect 53622 9103 53634 9279
rect 53576 9091 53634 9103
rect 54364 9283 54422 9295
rect 54364 9107 54376 9283
rect 54410 9107 54422 9283
rect 54364 9095 54422 9107
rect 54482 9283 54540 9295
rect 54482 9107 54494 9283
rect 54528 9107 54540 9283
rect 54482 9095 54540 9107
rect 54600 9283 54658 9295
rect 54600 9107 54612 9283
rect 54646 9107 54658 9283
rect 54600 9095 54658 9107
rect 54718 9283 54776 9295
rect 54718 9107 54730 9283
rect 54764 9107 54776 9283
rect 54718 9095 54776 9107
rect 57849 9245 57861 9621
rect 57895 9245 57907 9621
rect 57849 9233 57907 9245
rect 57967 9621 58025 9633
rect 57967 9245 57979 9621
rect 58013 9245 58025 9621
rect 57967 9233 58025 9245
rect 58085 9621 58143 9633
rect 58085 9245 58097 9621
rect 58131 9245 58143 9621
rect 58202 9621 58260 9633
rect 58202 9445 58214 9621
rect 58248 9445 58260 9621
rect 58202 9433 58260 9445
rect 58320 9621 58378 9633
rect 58320 9445 58332 9621
rect 58366 9445 58378 9621
rect 58320 9433 58378 9445
rect 59847 9347 59905 9359
rect 58085 9233 58143 9245
rect 59847 9171 59859 9347
rect 59893 9171 59905 9347
rect 59847 9159 59905 9171
rect 59965 9347 60023 9359
rect 59965 9171 59977 9347
rect 60011 9171 60023 9347
rect 59965 9159 60023 9171
rect 60083 9347 60141 9359
rect 60083 9171 60095 9347
rect 60129 9171 60141 9347
rect 60083 9159 60141 9171
rect 60201 9347 60259 9359
rect 60201 9171 60213 9347
rect 60247 9171 60259 9347
rect 60201 9159 60259 9171
rect 60989 9351 61047 9363
rect 60989 9175 61001 9351
rect 61035 9175 61047 9351
rect 60989 9163 61047 9175
rect 61107 9351 61165 9363
rect 61107 9175 61119 9351
rect 61153 9175 61165 9351
rect 61107 9163 61165 9175
rect 61225 9351 61283 9363
rect 61225 9175 61237 9351
rect 61271 9175 61283 9351
rect 61225 9163 61283 9175
rect 61343 9351 61401 9363
rect 61343 9175 61355 9351
rect 61389 9175 61401 9351
rect 61343 9163 61401 9175
rect 5380 7871 5392 8047
rect 5426 7871 5438 8047
rect 5380 7859 5438 7871
rect 7652 8043 7710 8055
rect 7652 7867 7664 8043
rect 7698 7867 7710 8043
rect 5234 7671 5246 7859
rect 7652 7855 7710 7867
rect 7770 8043 7906 8055
rect 7770 7867 7782 8043
rect 7816 7867 7860 8043
rect 7770 7855 7860 7867
rect 5188 7659 5246 7671
rect 7848 7667 7860 7855
rect 7894 7667 7906 8043
rect 7848 7655 7906 7667
rect 7966 8043 8024 8055
rect 7966 7667 7978 8043
rect 8012 7667 8024 8043
rect 7966 7655 8024 7667
rect 8084 8043 8142 8055
rect 8084 7667 8096 8043
rect 8130 7667 8142 8043
rect 8084 7655 8142 7667
rect 8202 8043 8260 8055
rect 8202 7667 8214 8043
rect 8248 7667 8260 8043
rect 8202 7655 8260 7667
rect 8320 8043 8452 8055
rect 8320 7667 8332 8043
rect 8366 7867 8406 8043
rect 8440 7867 8452 8043
rect 8366 7855 8452 7867
rect 8512 8043 8570 8055
rect 8512 7867 8524 8043
rect 8558 7867 8570 8043
rect 8512 7855 8570 7867
rect 10796 8043 10854 8055
rect 10796 7867 10808 8043
rect 10842 7867 10854 8043
rect 10796 7855 10854 7867
rect 10914 8043 11050 8055
rect 10914 7867 10926 8043
rect 10960 7867 11004 8043
rect 10914 7855 11004 7867
rect 8366 7667 8378 7855
rect 8320 7655 8378 7667
rect 10992 7667 11004 7855
rect 11038 7667 11050 8043
rect 10992 7655 11050 7667
rect 11110 8043 11168 8055
rect 11110 7667 11122 8043
rect 11156 7667 11168 8043
rect 11110 7655 11168 7667
rect 11228 8043 11286 8055
rect 11228 7667 11240 8043
rect 11274 7667 11286 8043
rect 11228 7655 11286 7667
rect 11346 8043 11404 8055
rect 11346 7667 11358 8043
rect 11392 7667 11404 8043
rect 11346 7655 11404 7667
rect 11464 8043 11596 8055
rect 11464 7667 11476 8043
rect 11510 7867 11550 8043
rect 11584 7867 11596 8043
rect 11510 7855 11596 7867
rect 11656 8043 11714 8055
rect 11656 7867 11668 8043
rect 11702 7867 11714 8043
rect 11656 7855 11714 7867
rect 13998 8047 14056 8059
rect 13998 7871 14010 8047
rect 14044 7871 14056 8047
rect 13998 7859 14056 7871
rect 14116 8047 14252 8059
rect 14116 7871 14128 8047
rect 14162 7871 14206 8047
rect 14116 7859 14206 7871
rect 11510 7667 11522 7855
rect 11464 7655 11522 7667
rect 14194 7671 14206 7859
rect 14240 7671 14252 8047
rect 14194 7659 14252 7671
rect 14312 8047 14370 8059
rect 14312 7671 14324 8047
rect 14358 7671 14370 8047
rect 14312 7659 14370 7671
rect 14430 8047 14488 8059
rect 14430 7671 14442 8047
rect 14476 7671 14488 8047
rect 14430 7659 14488 7671
rect 14548 8047 14606 8059
rect 14548 7671 14560 8047
rect 14594 7671 14606 8047
rect 14548 7659 14606 7671
rect 14666 8047 14798 8059
rect 14666 7671 14678 8047
rect 14712 7871 14752 8047
rect 14786 7871 14798 8047
rect 14712 7859 14798 7871
rect 14858 8047 14916 8059
rect 14858 7871 14870 8047
rect 14904 7871 14916 8047
rect 14858 7859 14916 7871
rect 17142 8047 17200 8059
rect 17142 7871 17154 8047
rect 17188 7871 17200 8047
rect 17142 7859 17200 7871
rect 17260 8047 17396 8059
rect 17260 7871 17272 8047
rect 17306 7871 17350 8047
rect 17260 7859 17350 7871
rect 14712 7671 14724 7859
rect 14666 7659 14724 7671
rect 17338 7671 17350 7859
rect 17384 7671 17396 8047
rect 17338 7659 17396 7671
rect 17456 8047 17514 8059
rect 17456 7671 17468 8047
rect 17502 7671 17514 8047
rect 17456 7659 17514 7671
rect 17574 8047 17632 8059
rect 17574 7671 17586 8047
rect 17620 7671 17632 8047
rect 17574 7659 17632 7671
rect 17692 8047 17750 8059
rect 17692 7671 17704 8047
rect 17738 7671 17750 8047
rect 17692 7659 17750 7671
rect 17810 8047 17942 8059
rect 17810 7671 17822 8047
rect 17856 7871 17896 8047
rect 17930 7871 17942 8047
rect 17856 7859 17942 7871
rect 18002 8047 18060 8059
rect 63646 8982 63704 8994
rect 31379 8906 31579 8918
rect 31379 8872 31391 8906
rect 31567 8872 31579 8906
rect 31379 8860 31579 8872
rect 31379 8788 31579 8800
rect 31379 8754 31391 8788
rect 31567 8754 31579 8788
rect 31379 8742 31579 8754
rect 63646 8606 63658 8982
rect 63692 8606 63704 8982
rect 63646 8594 63704 8606
rect 63764 8982 63822 8994
rect 63764 8606 63776 8982
rect 63810 8606 63822 8982
rect 63764 8594 63822 8606
rect 63882 8982 63940 8994
rect 63882 8606 63894 8982
rect 63928 8606 63940 8982
rect 63999 8982 64057 8994
rect 63999 8806 64011 8982
rect 64045 8806 64057 8982
rect 63999 8794 64057 8806
rect 64117 8982 64175 8994
rect 64117 8806 64129 8982
rect 64163 8806 64175 8982
rect 64117 8794 64175 8806
rect 63882 8594 63940 8606
rect 31379 8486 31779 8498
rect 31379 8452 31391 8486
rect 31767 8452 31779 8486
rect 31379 8440 31779 8452
rect 31379 8368 31779 8380
rect 31379 8334 31391 8368
rect 31767 8334 31779 8368
rect 31379 8322 31779 8334
rect 31379 8250 31779 8262
rect 31379 8216 31391 8250
rect 31767 8216 31779 8250
rect 31379 8204 31779 8216
rect 18002 7871 18014 8047
rect 18048 7871 18060 8047
rect 18002 7859 18060 7871
rect 20274 8043 20332 8055
rect 20274 7867 20286 8043
rect 20320 7867 20332 8043
rect 17856 7671 17868 7859
rect 20274 7855 20332 7867
rect 20392 8043 20528 8055
rect 20392 7867 20404 8043
rect 20438 7867 20482 8043
rect 20392 7855 20482 7867
rect 17810 7659 17868 7671
rect 20470 7667 20482 7855
rect 20516 7667 20528 8043
rect 20470 7655 20528 7667
rect 20588 8043 20646 8055
rect 20588 7667 20600 8043
rect 20634 7667 20646 8043
rect 20588 7655 20646 7667
rect 20706 8043 20764 8055
rect 20706 7667 20718 8043
rect 20752 7667 20764 8043
rect 20706 7655 20764 7667
rect 20824 8043 20882 8055
rect 20824 7667 20836 8043
rect 20870 7667 20882 8043
rect 20824 7655 20882 7667
rect 20942 8043 21074 8055
rect 20942 7667 20954 8043
rect 20988 7867 21028 8043
rect 21062 7867 21074 8043
rect 20988 7855 21074 7867
rect 21134 8043 21192 8055
rect 21134 7867 21146 8043
rect 21180 7867 21192 8043
rect 21134 7855 21192 7867
rect 23418 8043 23476 8055
rect 23418 7867 23430 8043
rect 23464 7867 23476 8043
rect 23418 7855 23476 7867
rect 23536 8043 23672 8055
rect 23536 7867 23548 8043
rect 23582 7867 23626 8043
rect 23536 7855 23626 7867
rect 20988 7667 21000 7855
rect 20942 7655 21000 7667
rect 23614 7667 23626 7855
rect 23660 7667 23672 8043
rect 23614 7655 23672 7667
rect 23732 8043 23790 8055
rect 23732 7667 23744 8043
rect 23778 7667 23790 8043
rect 23732 7655 23790 7667
rect 23850 8043 23908 8055
rect 23850 7667 23862 8043
rect 23896 7667 23908 8043
rect 23850 7655 23908 7667
rect 23968 8043 24026 8055
rect 23968 7667 23980 8043
rect 24014 7667 24026 8043
rect 23968 7655 24026 7667
rect 24086 8043 24218 8055
rect 24086 7667 24098 8043
rect 24132 7867 24172 8043
rect 24206 7867 24218 8043
rect 24132 7855 24218 7867
rect 24278 8043 24336 8055
rect 24278 7867 24290 8043
rect 24324 7867 24336 8043
rect 24278 7855 24336 7867
rect 24132 7667 24144 7855
rect 31379 8132 31779 8144
rect 31379 8098 31391 8132
rect 31767 8098 31779 8132
rect 31379 8086 31779 8098
rect 31379 8014 31779 8026
rect 31379 7980 31391 8014
rect 31767 7980 31779 8014
rect 31379 7968 31779 7980
rect 24086 7655 24144 7667
rect 71846 8605 72046 8617
rect 71846 8571 71858 8605
rect 72034 8571 72046 8605
rect 71846 8559 72046 8571
rect 71846 8487 72046 8499
rect 71846 8453 71858 8487
rect 72034 8453 72046 8487
rect 71846 8425 72046 8453
rect 71846 8413 72246 8425
rect 71846 8379 71858 8413
rect 72234 8379 72246 8413
rect 71846 8367 72246 8379
rect 44584 7971 44642 7983
rect 38035 7883 38093 7895
rect 31379 7608 31579 7620
rect 31379 7574 31391 7608
rect 31567 7574 31579 7608
rect 31379 7562 31579 7574
rect 31379 7490 31579 7502
rect 31379 7456 31391 7490
rect 31567 7456 31579 7490
rect 38035 7507 38047 7883
rect 38081 7507 38093 7883
rect 38035 7495 38093 7507
rect 38153 7883 38211 7895
rect 38153 7507 38165 7883
rect 38199 7507 38211 7883
rect 38153 7495 38211 7507
rect 38271 7883 38329 7895
rect 38271 7507 38283 7883
rect 38317 7507 38329 7883
rect 38388 7883 38446 7895
rect 38388 7707 38400 7883
rect 38434 7707 38446 7883
rect 38388 7695 38446 7707
rect 38506 7883 38564 7895
rect 38506 7707 38518 7883
rect 38552 7707 38564 7883
rect 38506 7695 38564 7707
rect 38271 7495 38329 7507
rect 31379 7444 31579 7456
rect 44584 7595 44596 7971
rect 44630 7595 44642 7971
rect 44584 7583 44642 7595
rect 44702 7971 44760 7983
rect 44702 7595 44714 7971
rect 44748 7595 44760 7971
rect 44702 7583 44760 7595
rect 44820 7971 44878 7983
rect 44820 7595 44832 7971
rect 44866 7595 44878 7971
rect 44937 7971 44995 7983
rect 44937 7795 44949 7971
rect 44983 7795 44995 7971
rect 44937 7783 44995 7795
rect 45055 7971 45113 7983
rect 45055 7795 45067 7971
rect 45101 7795 45113 7971
rect 45055 7783 45113 7795
rect 44820 7583 44878 7595
rect 35123 7215 35181 7227
rect 31377 6838 31577 6850
rect 31377 6804 31389 6838
rect 31565 6804 31577 6838
rect 35123 6839 35135 7215
rect 35169 6839 35181 7215
rect 35123 6827 35181 6839
rect 35241 7215 35299 7227
rect 35241 6839 35253 7215
rect 35287 6839 35299 7215
rect 35241 6827 35299 6839
rect 35359 7215 35417 7227
rect 35359 6839 35371 7215
rect 35405 6839 35417 7215
rect 35476 7215 35534 7227
rect 35476 7039 35488 7215
rect 35522 7039 35534 7215
rect 35476 7027 35534 7039
rect 35594 7215 35652 7227
rect 35594 7039 35606 7215
rect 35640 7039 35652 7215
rect 35594 7027 35652 7039
rect 35359 6827 35417 6839
rect 31377 6792 31577 6804
rect 31377 6720 31577 6732
rect 31377 6686 31389 6720
rect 31565 6686 31577 6720
rect 31377 6674 31577 6686
rect 3235 6163 3293 6175
rect 3235 5987 3247 6163
rect 3281 5987 3293 6163
rect 3235 5975 3293 5987
rect 3353 6163 3411 6175
rect 3353 5987 3365 6163
rect 3399 5987 3411 6163
rect 3353 5975 3411 5987
rect 3973 6163 4031 6175
rect 3973 5987 3985 6163
rect 4019 5987 4031 6163
rect 3973 5975 4031 5987
rect 4091 6163 4149 6175
rect 4091 5987 4103 6163
rect 4137 5987 4149 6163
rect 4091 5975 4149 5987
rect 4711 6159 4769 6171
rect 4711 5983 4723 6159
rect 4757 5983 4769 6159
rect 4711 5971 4769 5983
rect 4829 6159 4887 6171
rect 4829 5983 4841 6159
rect 4875 5983 4887 6159
rect 4829 5971 4887 5983
rect 5449 6159 5507 6171
rect 5449 5983 5461 6159
rect 5495 5983 5507 6159
rect 5449 5971 5507 5983
rect 5567 6159 5625 6171
rect 5567 5983 5579 6159
rect 5613 5983 5625 6159
rect 5567 5971 5625 5983
rect 6189 6159 6247 6171
rect 6189 5983 6201 6159
rect 6235 5983 6247 6159
rect 6189 5971 6247 5983
rect 6307 6159 6365 6171
rect 6307 5983 6319 6159
rect 6353 5983 6365 6159
rect 6307 5971 6365 5983
rect 6931 6159 6989 6171
rect 6931 5983 6943 6159
rect 6977 5983 6989 6159
rect 6931 5971 6989 5983
rect 7049 6159 7107 6171
rect 7049 5983 7061 6159
rect 7095 5983 7107 6159
rect 7049 5971 7107 5983
rect 7669 6163 7727 6175
rect 7669 5987 7681 6163
rect 7715 5987 7727 6163
rect 7669 5975 7727 5987
rect 7787 6163 7845 6175
rect 7787 5987 7799 6163
rect 7833 5987 7845 6163
rect 7787 5975 7845 5987
rect 8407 6161 8465 6173
rect 8407 5985 8419 6161
rect 8453 5985 8465 6161
rect 8407 5973 8465 5985
rect 8525 6161 8583 6173
rect 8525 5985 8537 6161
rect 8571 5985 8583 6161
rect 8525 5973 8583 5985
rect 9355 5010 9413 5022
rect 9355 4834 9367 5010
rect 9401 4834 9413 5010
rect 9355 4822 9413 4834
rect 9473 5010 9531 5022
rect 9473 4834 9485 5010
rect 9519 4834 9531 5010
rect 9473 4822 9531 4834
rect 9879 5010 9937 5022
rect 9879 4634 9891 5010
rect 9925 4634 9937 5010
rect 9879 4622 9937 4634
rect 9997 5010 10055 5022
rect 9997 4634 10009 5010
rect 10043 4634 10055 5010
rect 9997 4622 10055 4634
rect 10115 5010 10173 5022
rect 10115 4634 10127 5010
rect 10161 4634 10173 5010
rect 10115 4622 10173 4634
rect 10233 5010 10291 5022
rect 10233 4634 10245 5010
rect 10279 4634 10291 5010
rect 10233 4622 10291 4634
rect 10351 5010 10409 5022
rect 10351 4634 10363 5010
rect 10397 4634 10409 5010
rect 10653 5010 10711 5022
rect 10653 4834 10665 5010
rect 10699 4834 10711 5010
rect 10653 4822 10711 4834
rect 10771 5010 10829 5022
rect 10771 4834 10783 5010
rect 10817 4834 10829 5010
rect 10771 4822 10829 4834
rect 11423 5008 11481 5020
rect 11423 4832 11435 5008
rect 11469 4832 11481 5008
rect 11423 4820 11481 4832
rect 11541 5008 11599 5020
rect 11541 4832 11553 5008
rect 11587 4832 11599 5008
rect 11541 4820 11599 4832
rect 11947 5008 12005 5020
rect 10351 4622 10409 4634
rect 11947 4632 11959 5008
rect 11993 4632 12005 5008
rect 11947 4620 12005 4632
rect 12065 5008 12123 5020
rect 12065 4632 12077 5008
rect 12111 4632 12123 5008
rect 12065 4620 12123 4632
rect 12183 5008 12241 5020
rect 12183 4632 12195 5008
rect 12229 4632 12241 5008
rect 12183 4620 12241 4632
rect 12301 5008 12359 5020
rect 12301 4632 12313 5008
rect 12347 4632 12359 5008
rect 12301 4620 12359 4632
rect 12419 5008 12477 5020
rect 12419 4632 12431 5008
rect 12465 4632 12477 5008
rect 12721 5008 12779 5020
rect 12721 4832 12733 5008
rect 12767 4832 12779 5008
rect 12721 4820 12779 4832
rect 12839 5008 12897 5020
rect 12839 4832 12851 5008
rect 12885 4832 12897 5008
rect 12839 4820 12897 4832
rect 13492 5010 13550 5022
rect 13492 4834 13504 5010
rect 13538 4834 13550 5010
rect 13492 4822 13550 4834
rect 13610 5010 13668 5022
rect 13610 4834 13622 5010
rect 13656 4834 13668 5010
rect 13610 4822 13668 4834
rect 14016 5010 14074 5022
rect 12419 4620 12477 4632
rect 14016 4634 14028 5010
rect 14062 4634 14074 5010
rect 14016 4622 14074 4634
rect 14134 5010 14192 5022
rect 14134 4634 14146 5010
rect 14180 4634 14192 5010
rect 14134 4622 14192 4634
rect 14252 5010 14310 5022
rect 14252 4634 14264 5010
rect 14298 4634 14310 5010
rect 14252 4622 14310 4634
rect 14370 5010 14428 5022
rect 14370 4634 14382 5010
rect 14416 4634 14428 5010
rect 14370 4622 14428 4634
rect 14488 5010 14546 5022
rect 14488 4634 14500 5010
rect 14534 4634 14546 5010
rect 14790 5010 14848 5022
rect 14790 4834 14802 5010
rect 14836 4834 14848 5010
rect 14790 4822 14848 4834
rect 14908 5010 14966 5022
rect 31377 6418 31777 6430
rect 31377 6384 31389 6418
rect 31765 6384 31777 6418
rect 31377 6372 31777 6384
rect 31377 6300 31777 6312
rect 31377 6266 31389 6300
rect 31765 6266 31777 6300
rect 71846 8295 72246 8307
rect 71846 8261 71858 8295
rect 72234 8261 72246 8295
rect 71846 8249 72246 8261
rect 71846 8177 72246 8189
rect 71846 8143 71858 8177
rect 72234 8143 72246 8177
rect 71846 8131 72246 8143
rect 71846 8059 72246 8071
rect 71846 8025 71858 8059
rect 72234 8025 72246 8059
rect 57863 7971 57921 7983
rect 51238 7903 51296 7915
rect 39387 6478 39445 6490
rect 39387 6302 39399 6478
rect 39433 6302 39445 6478
rect 31377 6254 31777 6266
rect 31377 6182 31777 6194
rect 31377 6148 31389 6182
rect 31765 6148 31777 6182
rect 31377 6136 31777 6148
rect 14908 4834 14920 5010
rect 14954 4834 14966 5010
rect 14908 4822 14966 4834
rect 15560 5008 15618 5020
rect 15560 4832 15572 5008
rect 15606 4832 15618 5008
rect 15560 4820 15618 4832
rect 15678 5008 15736 5020
rect 15678 4832 15690 5008
rect 15724 4832 15736 5008
rect 15678 4820 15736 4832
rect 16084 5008 16142 5020
rect 14488 4622 14546 4634
rect 16084 4632 16096 5008
rect 16130 4632 16142 5008
rect 16084 4620 16142 4632
rect 16202 5008 16260 5020
rect 16202 4632 16214 5008
rect 16248 4632 16260 5008
rect 16202 4620 16260 4632
rect 16320 5008 16378 5020
rect 16320 4632 16332 5008
rect 16366 4632 16378 5008
rect 16320 4620 16378 4632
rect 16438 5008 16496 5020
rect 16438 4632 16450 5008
rect 16484 4632 16496 5008
rect 16438 4620 16496 4632
rect 16556 5008 16614 5020
rect 16556 4632 16568 5008
rect 16602 4632 16614 5008
rect 16858 5008 16916 5020
rect 16858 4832 16870 5008
rect 16904 4832 16916 5008
rect 16858 4820 16916 4832
rect 16976 5008 17034 5020
rect 16976 4832 16988 5008
rect 17022 4832 17034 5008
rect 16976 4820 17034 4832
rect 17629 5008 17687 5020
rect 17629 4832 17641 5008
rect 17675 4832 17687 5008
rect 17629 4820 17687 4832
rect 17747 5008 17805 5020
rect 17747 4832 17759 5008
rect 17793 4832 17805 5008
rect 17747 4820 17805 4832
rect 18153 5008 18211 5020
rect 16556 4620 16614 4632
rect 18153 4632 18165 5008
rect 18199 4632 18211 5008
rect 18153 4620 18211 4632
rect 18271 5008 18329 5020
rect 18271 4632 18283 5008
rect 18317 4632 18329 5008
rect 18271 4620 18329 4632
rect 18389 5008 18447 5020
rect 18389 4632 18401 5008
rect 18435 4632 18447 5008
rect 18389 4620 18447 4632
rect 18507 5008 18565 5020
rect 18507 4632 18519 5008
rect 18553 4632 18565 5008
rect 18507 4620 18565 4632
rect 18625 5008 18683 5020
rect 18625 4632 18637 5008
rect 18671 4632 18683 5008
rect 18927 5008 18985 5020
rect 18927 4832 18939 5008
rect 18973 4832 18985 5008
rect 18927 4820 18985 4832
rect 19045 5008 19103 5020
rect 31377 6064 31777 6076
rect 31377 6030 31389 6064
rect 31765 6030 31777 6064
rect 38030 6279 38088 6291
rect 31377 6018 31777 6030
rect 31377 5946 31777 5958
rect 31377 5912 31389 5946
rect 31765 5912 31777 5946
rect 31377 5900 31777 5912
rect 38030 5903 38042 6279
rect 38076 5903 38088 6279
rect 38030 5891 38088 5903
rect 38148 6279 38206 6291
rect 38148 5903 38160 6279
rect 38194 5903 38206 6279
rect 38148 5891 38206 5903
rect 38266 6279 38324 6291
rect 38266 5903 38278 6279
rect 38312 5903 38324 6279
rect 38383 6279 38441 6291
rect 38383 6103 38395 6279
rect 38429 6103 38441 6279
rect 38383 6091 38441 6103
rect 38501 6279 38559 6291
rect 39387 6290 39445 6302
rect 39505 6478 39563 6490
rect 39505 6302 39517 6478
rect 39551 6302 39563 6478
rect 39505 6290 39563 6302
rect 39807 6478 39865 6490
rect 38501 6103 38513 6279
rect 38547 6103 38559 6279
rect 38501 6091 38559 6103
rect 39807 6102 39819 6478
rect 39853 6102 39865 6478
rect 39807 6090 39865 6102
rect 39925 6478 39983 6490
rect 39925 6102 39937 6478
rect 39971 6102 39983 6478
rect 39925 6090 39983 6102
rect 40043 6478 40101 6490
rect 40043 6102 40055 6478
rect 40089 6102 40101 6478
rect 40043 6090 40101 6102
rect 40161 6478 40219 6490
rect 40161 6102 40173 6478
rect 40207 6102 40219 6478
rect 40161 6090 40219 6102
rect 40279 6478 40337 6490
rect 40279 6102 40291 6478
rect 40325 6102 40337 6478
rect 40685 6478 40743 6490
rect 40685 6302 40697 6478
rect 40731 6302 40743 6478
rect 40685 6290 40743 6302
rect 40803 6478 40861 6490
rect 40803 6302 40815 6478
rect 40849 6302 40861 6478
rect 40803 6290 40861 6302
rect 41285 6478 41343 6490
rect 41285 6302 41297 6478
rect 41331 6302 41343 6478
rect 41285 6290 41343 6302
rect 41403 6478 41461 6490
rect 41403 6302 41415 6478
rect 41449 6302 41461 6478
rect 41403 6290 41461 6302
rect 41705 6478 41763 6490
rect 40279 6090 40337 6102
rect 41705 6102 41717 6478
rect 41751 6102 41763 6478
rect 41705 6090 41763 6102
rect 41823 6478 41881 6490
rect 41823 6102 41835 6478
rect 41869 6102 41881 6478
rect 41823 6090 41881 6102
rect 41941 6478 41999 6490
rect 41941 6102 41953 6478
rect 41987 6102 41999 6478
rect 41941 6090 41999 6102
rect 42059 6478 42117 6490
rect 42059 6102 42071 6478
rect 42105 6102 42117 6478
rect 42059 6090 42117 6102
rect 42177 6478 42235 6490
rect 42177 6102 42189 6478
rect 42223 6102 42235 6478
rect 42583 6478 42641 6490
rect 42583 6302 42595 6478
rect 42629 6302 42641 6478
rect 42583 6290 42641 6302
rect 42701 6478 42759 6490
rect 42701 6302 42713 6478
rect 42747 6302 42759 6478
rect 51238 7527 51250 7903
rect 51284 7527 51296 7903
rect 51238 7515 51296 7527
rect 51356 7903 51414 7915
rect 51356 7527 51368 7903
rect 51402 7527 51414 7903
rect 51356 7515 51414 7527
rect 51474 7903 51532 7915
rect 51474 7527 51486 7903
rect 51520 7527 51532 7903
rect 51591 7903 51649 7915
rect 51591 7727 51603 7903
rect 51637 7727 51649 7903
rect 51591 7715 51649 7727
rect 51709 7903 51767 7915
rect 51709 7727 51721 7903
rect 51755 7727 51767 7903
rect 51709 7715 51767 7727
rect 51474 7515 51532 7527
rect 57863 7595 57875 7971
rect 57909 7595 57921 7971
rect 57863 7583 57921 7595
rect 57981 7971 58039 7983
rect 57981 7595 57993 7971
rect 58027 7595 58039 7971
rect 57981 7583 58039 7595
rect 58099 7971 58157 7983
rect 58099 7595 58111 7971
rect 58145 7595 58157 7971
rect 58216 7971 58274 7983
rect 58216 7795 58228 7971
rect 58262 7795 58274 7971
rect 58216 7783 58274 7795
rect 58334 7971 58392 7983
rect 58334 7795 58346 7971
rect 58380 7795 58392 7971
rect 58334 7783 58392 7795
rect 58099 7583 58157 7595
rect 45936 6566 45994 6578
rect 45936 6390 45948 6566
rect 45982 6390 45994 6566
rect 42701 6290 42759 6302
rect 44579 6367 44637 6379
rect 42177 6090 42235 6102
rect 44579 5991 44591 6367
rect 44625 5991 44637 6367
rect 38266 5891 38324 5903
rect 44579 5979 44637 5991
rect 44697 6367 44755 6379
rect 44697 5991 44709 6367
rect 44743 5991 44755 6367
rect 44697 5979 44755 5991
rect 44815 6367 44873 6379
rect 44815 5991 44827 6367
rect 44861 5991 44873 6367
rect 44932 6367 44990 6379
rect 44932 6191 44944 6367
rect 44978 6191 44990 6367
rect 44932 6179 44990 6191
rect 45050 6367 45108 6379
rect 45936 6378 45994 6390
rect 46054 6566 46112 6578
rect 46054 6390 46066 6566
rect 46100 6390 46112 6566
rect 46054 6378 46112 6390
rect 46356 6566 46414 6578
rect 45050 6191 45062 6367
rect 45096 6191 45108 6367
rect 45050 6179 45108 6191
rect 46356 6190 46368 6566
rect 46402 6190 46414 6566
rect 46356 6178 46414 6190
rect 46474 6566 46532 6578
rect 46474 6190 46486 6566
rect 46520 6190 46532 6566
rect 46474 6178 46532 6190
rect 46592 6566 46650 6578
rect 46592 6190 46604 6566
rect 46638 6190 46650 6566
rect 46592 6178 46650 6190
rect 46710 6566 46768 6578
rect 46710 6190 46722 6566
rect 46756 6190 46768 6566
rect 46710 6178 46768 6190
rect 46828 6566 46886 6578
rect 46828 6190 46840 6566
rect 46874 6190 46886 6566
rect 47234 6566 47292 6578
rect 47234 6390 47246 6566
rect 47280 6390 47292 6566
rect 47234 6378 47292 6390
rect 47352 6566 47410 6578
rect 47352 6390 47364 6566
rect 47398 6390 47410 6566
rect 47352 6378 47410 6390
rect 47834 6566 47892 6578
rect 47834 6390 47846 6566
rect 47880 6390 47892 6566
rect 47834 6378 47892 6390
rect 47952 6566 48010 6578
rect 47952 6390 47964 6566
rect 47998 6390 48010 6566
rect 47952 6378 48010 6390
rect 48254 6566 48312 6578
rect 46828 6178 46886 6190
rect 48254 6190 48266 6566
rect 48300 6190 48312 6566
rect 48254 6178 48312 6190
rect 48372 6566 48430 6578
rect 48372 6190 48384 6566
rect 48418 6190 48430 6566
rect 48372 6178 48430 6190
rect 48490 6566 48548 6578
rect 48490 6190 48502 6566
rect 48536 6190 48548 6566
rect 48490 6178 48548 6190
rect 48608 6566 48666 6578
rect 48608 6190 48620 6566
rect 48654 6190 48666 6566
rect 48608 6178 48666 6190
rect 48726 6566 48784 6578
rect 48726 6190 48738 6566
rect 48772 6190 48784 6566
rect 49132 6566 49190 6578
rect 49132 6390 49144 6566
rect 49178 6390 49190 6566
rect 49132 6378 49190 6390
rect 49250 6566 49308 6578
rect 49250 6390 49262 6566
rect 49296 6390 49308 6566
rect 49250 6378 49308 6390
rect 71846 8013 72246 8025
rect 52590 6498 52648 6510
rect 52590 6322 52602 6498
rect 52636 6322 52648 6498
rect 48726 6178 48784 6190
rect 51233 6299 51291 6311
rect 44815 5979 44873 5991
rect 19045 4832 19057 5008
rect 19091 4832 19103 5008
rect 19045 4820 19103 4832
rect 19697 5006 19755 5018
rect 19697 4830 19709 5006
rect 19743 4830 19755 5006
rect 19697 4818 19755 4830
rect 19815 5006 19873 5018
rect 19815 4830 19827 5006
rect 19861 4830 19873 5006
rect 19815 4818 19873 4830
rect 20221 5006 20279 5018
rect 18625 4620 18683 4632
rect 20221 4630 20233 5006
rect 20267 4630 20279 5006
rect 20221 4618 20279 4630
rect 20339 5006 20397 5018
rect 20339 4630 20351 5006
rect 20385 4630 20397 5006
rect 20339 4618 20397 4630
rect 20457 5006 20515 5018
rect 20457 4630 20469 5006
rect 20503 4630 20515 5006
rect 20457 4618 20515 4630
rect 20575 5006 20633 5018
rect 20575 4630 20587 5006
rect 20621 4630 20633 5006
rect 20575 4618 20633 4630
rect 20693 5006 20751 5018
rect 20693 4630 20705 5006
rect 20739 4630 20751 5006
rect 20995 5006 21053 5018
rect 20995 4830 21007 5006
rect 21041 4830 21053 5006
rect 20995 4818 21053 4830
rect 21113 5006 21171 5018
rect 21113 4830 21125 5006
rect 21159 4830 21171 5006
rect 21113 4818 21171 4830
rect 21766 5008 21824 5020
rect 21766 4832 21778 5008
rect 21812 4832 21824 5008
rect 21766 4820 21824 4832
rect 21884 5008 21942 5020
rect 21884 4832 21896 5008
rect 21930 4832 21942 5008
rect 21884 4820 21942 4832
rect 22290 5008 22348 5020
rect 20693 4618 20751 4630
rect 22290 4632 22302 5008
rect 22336 4632 22348 5008
rect 22290 4620 22348 4632
rect 22408 5008 22466 5020
rect 22408 4632 22420 5008
rect 22454 4632 22466 5008
rect 22408 4620 22466 4632
rect 22526 5008 22584 5020
rect 22526 4632 22538 5008
rect 22572 4632 22584 5008
rect 22526 4620 22584 4632
rect 22644 5008 22702 5020
rect 22644 4632 22656 5008
rect 22690 4632 22702 5008
rect 22644 4620 22702 4632
rect 22762 5008 22820 5020
rect 22762 4632 22774 5008
rect 22808 4632 22820 5008
rect 23064 5008 23122 5020
rect 23064 4832 23076 5008
rect 23110 4832 23122 5008
rect 23064 4820 23122 4832
rect 23182 5008 23240 5020
rect 51233 5923 51245 6299
rect 51279 5923 51291 6299
rect 51233 5911 51291 5923
rect 51351 6299 51409 6311
rect 51351 5923 51363 6299
rect 51397 5923 51409 6299
rect 51351 5911 51409 5923
rect 51469 6299 51527 6311
rect 51469 5923 51481 6299
rect 51515 5923 51527 6299
rect 51586 6299 51644 6311
rect 51586 6123 51598 6299
rect 51632 6123 51644 6299
rect 51586 6111 51644 6123
rect 51704 6299 51762 6311
rect 52590 6310 52648 6322
rect 52708 6498 52766 6510
rect 52708 6322 52720 6498
rect 52754 6322 52766 6498
rect 52708 6310 52766 6322
rect 53010 6498 53068 6510
rect 51704 6123 51716 6299
rect 51750 6123 51762 6299
rect 51704 6111 51762 6123
rect 53010 6122 53022 6498
rect 53056 6122 53068 6498
rect 53010 6110 53068 6122
rect 53128 6498 53186 6510
rect 53128 6122 53140 6498
rect 53174 6122 53186 6498
rect 53128 6110 53186 6122
rect 53246 6498 53304 6510
rect 53246 6122 53258 6498
rect 53292 6122 53304 6498
rect 53246 6110 53304 6122
rect 53364 6498 53422 6510
rect 53364 6122 53376 6498
rect 53410 6122 53422 6498
rect 53364 6110 53422 6122
rect 53482 6498 53540 6510
rect 53482 6122 53494 6498
rect 53528 6122 53540 6498
rect 53888 6498 53946 6510
rect 53888 6322 53900 6498
rect 53934 6322 53946 6498
rect 53888 6310 53946 6322
rect 54006 6498 54064 6510
rect 54006 6322 54018 6498
rect 54052 6322 54064 6498
rect 54006 6310 54064 6322
rect 54488 6498 54546 6510
rect 54488 6322 54500 6498
rect 54534 6322 54546 6498
rect 54488 6310 54546 6322
rect 54606 6498 54664 6510
rect 54606 6322 54618 6498
rect 54652 6322 54664 6498
rect 54606 6310 54664 6322
rect 54908 6498 54966 6510
rect 53482 6110 53540 6122
rect 54908 6122 54920 6498
rect 54954 6122 54966 6498
rect 54908 6110 54966 6122
rect 55026 6498 55084 6510
rect 55026 6122 55038 6498
rect 55072 6122 55084 6498
rect 55026 6110 55084 6122
rect 55144 6498 55202 6510
rect 55144 6122 55156 6498
rect 55190 6122 55202 6498
rect 55144 6110 55202 6122
rect 55262 6498 55320 6510
rect 55262 6122 55274 6498
rect 55308 6122 55320 6498
rect 55262 6110 55320 6122
rect 55380 6498 55438 6510
rect 55380 6122 55392 6498
rect 55426 6122 55438 6498
rect 55786 6498 55844 6510
rect 55786 6322 55798 6498
rect 55832 6322 55844 6498
rect 55786 6310 55844 6322
rect 55904 6498 55962 6510
rect 55904 6322 55916 6498
rect 55950 6322 55962 6498
rect 71846 7941 72246 7953
rect 71846 7907 71858 7941
rect 72234 7907 72246 7941
rect 71846 7895 72246 7907
rect 71846 7863 72046 7895
rect 71846 7829 71858 7863
rect 72034 7829 72046 7863
rect 71846 7817 72046 7829
rect 59215 6566 59273 6578
rect 59215 6390 59227 6566
rect 59261 6390 59273 6566
rect 55904 6310 55962 6322
rect 57858 6367 57916 6379
rect 55380 6110 55438 6122
rect 51469 5911 51527 5923
rect 57858 5991 57870 6367
rect 57904 5991 57916 6367
rect 57858 5979 57916 5991
rect 57976 6367 58034 6379
rect 57976 5991 57988 6367
rect 58022 5991 58034 6367
rect 57976 5979 58034 5991
rect 58094 6367 58152 6379
rect 58094 5991 58106 6367
rect 58140 5991 58152 6367
rect 58211 6367 58269 6379
rect 58211 6191 58223 6367
rect 58257 6191 58269 6367
rect 58211 6179 58269 6191
rect 58329 6367 58387 6379
rect 59215 6378 59273 6390
rect 59333 6566 59391 6578
rect 59333 6390 59345 6566
rect 59379 6390 59391 6566
rect 59333 6378 59391 6390
rect 59635 6566 59693 6578
rect 58329 6191 58341 6367
rect 58375 6191 58387 6367
rect 58329 6179 58387 6191
rect 59635 6190 59647 6566
rect 59681 6190 59693 6566
rect 59635 6178 59693 6190
rect 59753 6566 59811 6578
rect 59753 6190 59765 6566
rect 59799 6190 59811 6566
rect 59753 6178 59811 6190
rect 59871 6566 59929 6578
rect 59871 6190 59883 6566
rect 59917 6190 59929 6566
rect 59871 6178 59929 6190
rect 59989 6566 60047 6578
rect 59989 6190 60001 6566
rect 60035 6190 60047 6566
rect 59989 6178 60047 6190
rect 60107 6566 60165 6578
rect 60107 6190 60119 6566
rect 60153 6190 60165 6566
rect 60513 6566 60571 6578
rect 60513 6390 60525 6566
rect 60559 6390 60571 6566
rect 60513 6378 60571 6390
rect 60631 6566 60689 6578
rect 60631 6390 60643 6566
rect 60677 6390 60689 6566
rect 60631 6378 60689 6390
rect 61113 6566 61171 6578
rect 61113 6390 61125 6566
rect 61159 6390 61171 6566
rect 61113 6378 61171 6390
rect 61231 6566 61289 6578
rect 61231 6390 61243 6566
rect 61277 6390 61289 6566
rect 61231 6378 61289 6390
rect 61533 6566 61591 6578
rect 60107 6178 60165 6190
rect 61533 6190 61545 6566
rect 61579 6190 61591 6566
rect 61533 6178 61591 6190
rect 61651 6566 61709 6578
rect 61651 6190 61663 6566
rect 61697 6190 61709 6566
rect 61651 6178 61709 6190
rect 61769 6566 61827 6578
rect 61769 6190 61781 6566
rect 61815 6190 61827 6566
rect 61769 6178 61827 6190
rect 61887 6566 61945 6578
rect 61887 6190 61899 6566
rect 61933 6190 61945 6566
rect 61887 6178 61945 6190
rect 62005 6566 62063 6578
rect 62005 6190 62017 6566
rect 62051 6190 62063 6566
rect 62411 6566 62469 6578
rect 62411 6390 62423 6566
rect 62457 6390 62469 6566
rect 62411 6378 62469 6390
rect 62529 6566 62587 6578
rect 62529 6390 62541 6566
rect 62575 6390 62587 6566
rect 62529 6378 62587 6390
rect 67254 7054 67312 7066
rect 67254 6678 67266 7054
rect 67300 6678 67312 7054
rect 67254 6666 67312 6678
rect 67372 7054 67430 7066
rect 67372 6678 67384 7054
rect 67418 6678 67430 7054
rect 67372 6666 67430 6678
rect 67490 7054 67548 7066
rect 67490 6678 67502 7054
rect 67536 6678 67548 7054
rect 67607 7054 67665 7066
rect 67607 6878 67619 7054
rect 67653 6878 67665 7054
rect 67607 6866 67665 6878
rect 67725 7054 67783 7066
rect 67725 6878 67737 7054
rect 67771 6878 67783 7054
rect 71846 7745 72046 7757
rect 71846 7711 71858 7745
rect 72034 7711 72046 7745
rect 71846 7699 72046 7711
rect 67725 6866 67783 6878
rect 67490 6666 67548 6678
rect 65349 6269 65407 6281
rect 62005 6178 62063 6190
rect 58094 5979 58152 5991
rect 65349 6093 65361 6269
rect 65395 6093 65407 6269
rect 65349 6081 65407 6093
rect 65467 6269 65525 6281
rect 65467 6093 65479 6269
rect 65513 6093 65525 6269
rect 65467 6081 65525 6093
rect 65769 6269 65827 6281
rect 63646 5949 63704 5961
rect 63646 5573 63658 5949
rect 63692 5573 63704 5949
rect 63646 5561 63704 5573
rect 63764 5949 63822 5961
rect 63764 5573 63776 5949
rect 63810 5573 63822 5949
rect 63764 5561 63822 5573
rect 63882 5949 63940 5961
rect 63882 5573 63894 5949
rect 63928 5573 63940 5949
rect 63999 5949 64057 5961
rect 63999 5773 64011 5949
rect 64045 5773 64057 5949
rect 63999 5761 64057 5773
rect 64117 5949 64175 5961
rect 64117 5773 64129 5949
rect 64163 5773 64175 5949
rect 65769 5893 65781 6269
rect 65815 5893 65827 6269
rect 65769 5881 65827 5893
rect 65887 6269 65945 6281
rect 65887 5893 65899 6269
rect 65933 5893 65945 6269
rect 65887 5881 65945 5893
rect 66005 6269 66063 6281
rect 66005 5893 66017 6269
rect 66051 5893 66063 6269
rect 66005 5881 66063 5893
rect 66123 6269 66181 6281
rect 66123 5893 66135 6269
rect 66169 5893 66181 6269
rect 66123 5881 66181 5893
rect 66241 6269 66299 6281
rect 66241 5893 66253 6269
rect 66287 5893 66299 6269
rect 66647 6269 66705 6281
rect 66647 6093 66659 6269
rect 66693 6093 66705 6269
rect 66647 6081 66705 6093
rect 66765 6269 66823 6281
rect 66765 6093 66777 6269
rect 66811 6093 66823 6269
rect 66765 6081 66823 6093
rect 66241 5881 66299 5893
rect 64117 5761 64175 5773
rect 63882 5561 63940 5573
rect 31377 5540 31577 5552
rect 31377 5506 31389 5540
rect 31565 5506 31577 5540
rect 31377 5494 31577 5506
rect 31377 5422 31577 5434
rect 31377 5388 31389 5422
rect 31565 5388 31577 5422
rect 31377 5376 31577 5388
rect 71846 5461 72046 5473
rect 71846 5427 71858 5461
rect 72034 5427 72046 5461
rect 71846 5415 72046 5427
rect 71846 5343 72046 5355
rect 71846 5309 71858 5343
rect 72034 5309 72046 5343
rect 71846 5281 72046 5309
rect 71846 5269 72246 5281
rect 71846 5235 71858 5269
rect 72234 5235 72246 5269
rect 71846 5223 72246 5235
rect 23182 4832 23194 5008
rect 23228 4832 23240 5008
rect 23182 4820 23240 4832
rect 23834 5006 23892 5018
rect 23834 4830 23846 5006
rect 23880 4830 23892 5006
rect 23834 4818 23892 4830
rect 23952 5006 24010 5018
rect 23952 4830 23964 5006
rect 23998 4830 24010 5006
rect 23952 4818 24010 4830
rect 24358 5006 24416 5018
rect 22762 4620 22820 4632
rect 24358 4630 24370 5006
rect 24404 4630 24416 5006
rect 24358 4618 24416 4630
rect 24476 5006 24534 5018
rect 24476 4630 24488 5006
rect 24522 4630 24534 5006
rect 24476 4618 24534 4630
rect 24594 5006 24652 5018
rect 24594 4630 24606 5006
rect 24640 4630 24652 5006
rect 24594 4618 24652 4630
rect 24712 5006 24770 5018
rect 24712 4630 24724 5006
rect 24758 4630 24770 5006
rect 24712 4618 24770 4630
rect 24830 5006 24888 5018
rect 24830 4630 24842 5006
rect 24876 4630 24888 5006
rect 25132 5006 25190 5018
rect 25132 4830 25144 5006
rect 25178 4830 25190 5006
rect 25132 4818 25190 4830
rect 25250 5006 25308 5018
rect 25250 4830 25262 5006
rect 25296 4830 25308 5006
rect 71846 5151 72246 5163
rect 71846 5117 71858 5151
rect 72234 5117 72246 5151
rect 71846 5105 72246 5117
rect 25250 4818 25308 4830
rect 71846 5033 72246 5045
rect 71846 4999 71858 5033
rect 72234 4999 72246 5033
rect 71846 4987 72246 4999
rect 71846 4915 72246 4927
rect 71846 4881 71858 4915
rect 72234 4881 72246 4915
rect 71846 4869 72246 4881
rect 31377 4769 31577 4781
rect 31377 4735 31389 4769
rect 31565 4735 31577 4769
rect 31377 4723 31577 4735
rect 24830 4618 24888 4630
rect 31377 4651 31577 4663
rect 31377 4617 31389 4651
rect 31565 4617 31577 4651
rect 31377 4605 31577 4617
rect 31377 4349 31777 4361
rect 31377 4315 31389 4349
rect 31765 4315 31777 4349
rect 31377 4303 31777 4315
rect 31377 4231 31777 4243
rect 31377 4197 31389 4231
rect 31765 4197 31777 4231
rect 31377 4185 31777 4197
rect 31377 4113 31777 4125
rect 31377 4079 31389 4113
rect 31765 4079 31777 4113
rect 31377 4067 31777 4079
rect 31377 3995 31777 4007
rect 31377 3961 31389 3995
rect 31765 3961 31777 3995
rect 31377 3949 31777 3961
rect 35104 3937 35162 3949
rect 31377 3877 31777 3889
rect 31377 3843 31389 3877
rect 31765 3843 31777 3877
rect 31377 3831 31777 3843
rect 35104 3561 35116 3937
rect 35150 3561 35162 3937
rect 35104 3549 35162 3561
rect 35222 3937 35280 3949
rect 35222 3561 35234 3937
rect 35268 3561 35280 3937
rect 35222 3549 35280 3561
rect 35340 3937 35398 3949
rect 35340 3561 35352 3937
rect 35386 3561 35398 3937
rect 35457 3937 35515 3949
rect 35457 3761 35469 3937
rect 35503 3761 35515 3937
rect 35457 3749 35515 3761
rect 35575 3937 35633 3949
rect 35575 3761 35587 3937
rect 35621 3761 35633 3937
rect 35575 3749 35633 3761
rect 38013 3753 38071 3765
rect 35340 3549 35398 3561
rect 31377 3471 31577 3483
rect 31377 3437 31389 3471
rect 31565 3437 31577 3471
rect 31377 3425 31577 3437
rect 31377 3353 31577 3365
rect 31377 3319 31389 3353
rect 31565 3319 31577 3353
rect 38013 3377 38025 3753
rect 38059 3377 38071 3753
rect 38013 3365 38071 3377
rect 38131 3753 38189 3765
rect 38131 3377 38143 3753
rect 38177 3377 38189 3753
rect 38131 3365 38189 3377
rect 38249 3753 38307 3765
rect 38249 3377 38261 3753
rect 38295 3377 38307 3753
rect 38366 3753 38424 3765
rect 38366 3577 38378 3753
rect 38412 3577 38424 3753
rect 38366 3565 38424 3577
rect 38484 3753 38542 3765
rect 38484 3577 38496 3753
rect 38530 3577 38542 3753
rect 38484 3565 38542 3577
rect 44564 3751 44622 3763
rect 40011 3479 40069 3491
rect 38249 3365 38307 3377
rect 31377 3307 31577 3319
rect 40011 3303 40023 3479
rect 40057 3303 40069 3479
rect 40011 3291 40069 3303
rect 40129 3479 40187 3491
rect 40129 3303 40141 3479
rect 40175 3303 40187 3479
rect 40129 3291 40187 3303
rect 40247 3479 40305 3491
rect 40247 3303 40259 3479
rect 40293 3303 40305 3479
rect 40247 3291 40305 3303
rect 40365 3479 40423 3491
rect 40365 3303 40377 3479
rect 40411 3303 40423 3479
rect 40365 3291 40423 3303
rect 41153 3483 41211 3495
rect 41153 3307 41165 3483
rect 41199 3307 41211 3483
rect 41153 3295 41211 3307
rect 41271 3483 41329 3495
rect 41271 3307 41283 3483
rect 41317 3307 41329 3483
rect 41271 3295 41329 3307
rect 41389 3483 41447 3495
rect 41389 3307 41401 3483
rect 41435 3307 41447 3483
rect 41389 3295 41447 3307
rect 41507 3483 41565 3495
rect 41507 3307 41519 3483
rect 41553 3307 41565 3483
rect 41507 3295 41565 3307
rect 44564 3375 44576 3751
rect 44610 3375 44622 3751
rect 44564 3363 44622 3375
rect 44682 3751 44740 3763
rect 44682 3375 44694 3751
rect 44728 3375 44740 3751
rect 44682 3363 44740 3375
rect 44800 3751 44858 3763
rect 44800 3375 44812 3751
rect 44846 3375 44858 3751
rect 44917 3751 44975 3763
rect 44917 3575 44929 3751
rect 44963 3575 44975 3751
rect 44917 3563 44975 3575
rect 45035 3751 45093 3763
rect 45035 3575 45047 3751
rect 45081 3575 45093 3751
rect 45035 3563 45093 3575
rect 71846 4797 72246 4809
rect 71846 4763 71858 4797
rect 72234 4763 72246 4797
rect 71846 4751 72246 4763
rect 71846 4719 72046 4751
rect 71846 4685 71858 4719
rect 72034 4685 72046 4719
rect 71846 4673 72046 4685
rect 51219 3752 51277 3764
rect 46562 3477 46620 3489
rect 44800 3363 44858 3375
rect 46562 3301 46574 3477
rect 46608 3301 46620 3477
rect 46562 3289 46620 3301
rect 46680 3477 46738 3489
rect 46680 3301 46692 3477
rect 46726 3301 46738 3477
rect 46680 3289 46738 3301
rect 46798 3477 46856 3489
rect 46798 3301 46810 3477
rect 46844 3301 46856 3477
rect 46798 3289 46856 3301
rect 46916 3477 46974 3489
rect 46916 3301 46928 3477
rect 46962 3301 46974 3477
rect 46916 3289 46974 3301
rect 47704 3481 47762 3493
rect 47704 3305 47716 3481
rect 47750 3305 47762 3481
rect 47704 3293 47762 3305
rect 47822 3481 47880 3493
rect 47822 3305 47834 3481
rect 47868 3305 47880 3481
rect 47822 3293 47880 3305
rect 47940 3481 47998 3493
rect 47940 3305 47952 3481
rect 47986 3305 47998 3481
rect 47940 3293 47998 3305
rect 48058 3481 48116 3493
rect 48058 3305 48070 3481
rect 48104 3305 48116 3481
rect 48058 3293 48116 3305
rect 51219 3376 51231 3752
rect 51265 3376 51277 3752
rect 51219 3364 51277 3376
rect 51337 3752 51395 3764
rect 51337 3376 51349 3752
rect 51383 3376 51395 3752
rect 51337 3364 51395 3376
rect 51455 3752 51513 3764
rect 51455 3376 51467 3752
rect 51501 3376 51513 3752
rect 51572 3752 51630 3764
rect 51572 3576 51584 3752
rect 51618 3576 51630 3752
rect 51572 3564 51630 3576
rect 51690 3752 51748 3764
rect 51690 3576 51702 3752
rect 51736 3576 51748 3752
rect 51690 3564 51748 3576
rect 63717 4029 63775 4041
rect 57841 3753 57899 3765
rect 53217 3478 53275 3490
rect 51455 3364 51513 3376
rect 53217 3302 53229 3478
rect 53263 3302 53275 3478
rect 53217 3290 53275 3302
rect 53335 3478 53393 3490
rect 53335 3302 53347 3478
rect 53381 3302 53393 3478
rect 53335 3290 53393 3302
rect 53453 3478 53511 3490
rect 53453 3302 53465 3478
rect 53499 3302 53511 3478
rect 53453 3290 53511 3302
rect 53571 3478 53629 3490
rect 53571 3302 53583 3478
rect 53617 3302 53629 3478
rect 53571 3290 53629 3302
rect 54359 3482 54417 3494
rect 54359 3306 54371 3482
rect 54405 3306 54417 3482
rect 54359 3294 54417 3306
rect 54477 3482 54535 3494
rect 54477 3306 54489 3482
rect 54523 3306 54535 3482
rect 54477 3294 54535 3306
rect 54595 3482 54653 3494
rect 54595 3306 54607 3482
rect 54641 3306 54653 3482
rect 54595 3294 54653 3306
rect 54713 3482 54771 3494
rect 54713 3306 54725 3482
rect 54759 3306 54771 3482
rect 54713 3294 54771 3306
rect 57841 3377 57853 3753
rect 57887 3377 57899 3753
rect 57841 3365 57899 3377
rect 57959 3753 58017 3765
rect 57959 3377 57971 3753
rect 58005 3377 58017 3753
rect 57959 3365 58017 3377
rect 58077 3753 58135 3765
rect 58077 3377 58089 3753
rect 58123 3377 58135 3753
rect 58194 3753 58252 3765
rect 58194 3577 58206 3753
rect 58240 3577 58252 3753
rect 58194 3565 58252 3577
rect 58312 3753 58370 3765
rect 58312 3577 58324 3753
rect 58358 3577 58370 3753
rect 58312 3565 58370 3577
rect 63717 3653 63729 4029
rect 63763 3653 63775 4029
rect 63717 3641 63775 3653
rect 63835 4029 63893 4041
rect 63835 3653 63847 4029
rect 63881 3653 63893 4029
rect 63835 3641 63893 3653
rect 63953 4029 64011 4041
rect 63953 3653 63965 4029
rect 63999 3653 64011 4029
rect 64070 4029 64128 4041
rect 64070 3853 64082 4029
rect 64116 3853 64128 4029
rect 64070 3841 64128 3853
rect 64188 4029 64246 4041
rect 64188 3853 64200 4029
rect 64234 3853 64246 4029
rect 64188 3841 64246 3853
rect 63953 3641 64011 3653
rect 59839 3479 59897 3491
rect 58077 3365 58135 3377
rect 59839 3303 59851 3479
rect 59885 3303 59897 3479
rect 59839 3291 59897 3303
rect 59957 3479 60015 3491
rect 59957 3303 59969 3479
rect 60003 3303 60015 3479
rect 59957 3291 60015 3303
rect 60075 3479 60133 3491
rect 60075 3303 60087 3479
rect 60121 3303 60133 3479
rect 60075 3291 60133 3303
rect 60193 3479 60251 3491
rect 60193 3303 60205 3479
rect 60239 3303 60251 3479
rect 60193 3291 60251 3303
rect 60981 3483 61039 3495
rect 60981 3307 60993 3483
rect 61027 3307 61039 3483
rect 60981 3295 61039 3307
rect 61099 3483 61157 3495
rect 61099 3307 61111 3483
rect 61145 3307 61157 3483
rect 61099 3295 61157 3307
rect 61217 3483 61275 3495
rect 61217 3307 61229 3483
rect 61263 3307 61275 3483
rect 61217 3295 61275 3307
rect 61335 3483 61393 3495
rect 61335 3307 61347 3483
rect 61381 3307 61393 3483
rect 61335 3295 61393 3307
rect 71846 4601 72046 4613
rect 71846 4567 71858 4601
rect 72034 4567 72046 4601
rect 71846 4555 72046 4567
rect 67254 3559 67312 3571
rect 67254 3183 67266 3559
rect 67300 3183 67312 3559
rect 67254 3171 67312 3183
rect 67372 3559 67430 3571
rect 67372 3183 67384 3559
rect 67418 3183 67430 3559
rect 67372 3171 67430 3183
rect 67490 3559 67548 3571
rect 67490 3183 67502 3559
rect 67536 3183 67548 3559
rect 67607 3559 67665 3571
rect 67607 3383 67619 3559
rect 67653 3383 67665 3559
rect 67607 3371 67665 3383
rect 67725 3559 67783 3571
rect 67725 3383 67737 3559
rect 67771 3383 67783 3559
rect 67725 3371 67783 3383
rect 67490 3171 67548 3183
rect 65349 2774 65407 2786
rect 31375 2701 31575 2713
rect 31375 2667 31387 2701
rect 31563 2667 31575 2701
rect 31375 2655 31575 2667
rect 31375 2583 31575 2595
rect 31375 2549 31387 2583
rect 31563 2549 31575 2583
rect 31375 2537 31575 2549
rect 31375 2281 31775 2293
rect 31375 2247 31387 2281
rect 31763 2247 31775 2281
rect 31375 2235 31775 2247
rect 31375 2163 31775 2175
rect 31375 2129 31387 2163
rect 31763 2129 31775 2163
rect 31375 2117 31775 2129
rect 65349 2598 65361 2774
rect 65395 2598 65407 2774
rect 65349 2586 65407 2598
rect 65467 2774 65525 2786
rect 65467 2598 65479 2774
rect 65513 2598 65525 2774
rect 65467 2586 65525 2598
rect 65769 2774 65827 2786
rect 65769 2398 65781 2774
rect 65815 2398 65827 2774
rect 65769 2386 65827 2398
rect 65887 2774 65945 2786
rect 65887 2398 65899 2774
rect 65933 2398 65945 2774
rect 65887 2386 65945 2398
rect 66005 2774 66063 2786
rect 66005 2398 66017 2774
rect 66051 2398 66063 2774
rect 66005 2386 66063 2398
rect 66123 2774 66181 2786
rect 66123 2398 66135 2774
rect 66169 2398 66181 2774
rect 66123 2386 66181 2398
rect 66241 2774 66299 2786
rect 66241 2398 66253 2774
rect 66287 2398 66299 2774
rect 66647 2774 66705 2786
rect 66647 2598 66659 2774
rect 66693 2598 66705 2774
rect 66647 2586 66705 2598
rect 66765 2774 66823 2786
rect 66765 2598 66777 2774
rect 66811 2598 66823 2774
rect 66765 2586 66823 2598
rect 66241 2386 66299 2398
rect 31375 2045 31775 2057
rect 31375 2011 31387 2045
rect 31763 2011 31775 2045
rect 31375 1999 31775 2011
rect 1082 795 1140 807
rect 1082 619 1094 795
rect 1128 619 1140 795
rect 1082 607 1140 619
rect 1200 795 1332 807
rect 1200 619 1212 795
rect 1246 619 1286 795
rect 1200 607 1286 619
rect 1274 419 1286 607
rect 1320 419 1332 795
rect 1274 407 1332 419
rect 1392 795 1450 807
rect 1392 419 1404 795
rect 1438 419 1450 795
rect 1392 407 1450 419
rect 1510 795 1568 807
rect 1510 419 1522 795
rect 1556 419 1568 795
rect 1510 407 1568 419
rect 1628 795 1686 807
rect 1628 419 1640 795
rect 1674 419 1686 795
rect 1628 407 1686 419
rect 1746 795 1882 807
rect 1746 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1882 795
rect 1792 607 1882 619
rect 1942 795 2000 807
rect 1942 619 1954 795
rect 1988 619 2000 795
rect 1942 607 2000 619
rect 4226 795 4284 807
rect 4226 619 4238 795
rect 4272 619 4284 795
rect 4226 607 4284 619
rect 4344 795 4476 807
rect 4344 619 4356 795
rect 4390 619 4430 795
rect 4344 607 4430 619
rect 1792 419 1804 607
rect 1746 407 1804 419
rect 4418 419 4430 607
rect 4464 419 4476 795
rect 4418 407 4476 419
rect 4536 795 4594 807
rect 4536 419 4548 795
rect 4582 419 4594 795
rect 4536 407 4594 419
rect 4654 795 4712 807
rect 4654 419 4666 795
rect 4700 419 4712 795
rect 4654 407 4712 419
rect 4772 795 4830 807
rect 4772 419 4784 795
rect 4818 419 4830 795
rect 4772 407 4830 419
rect 4890 795 5026 807
rect 4890 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5026 795
rect 4936 607 5026 619
rect 5086 795 5144 807
rect 5086 619 5098 795
rect 5132 619 5144 795
rect 5086 607 5144 619
rect 7358 799 7416 811
rect 7358 623 7370 799
rect 7404 623 7416 799
rect 7358 611 7416 623
rect 7476 799 7608 811
rect 7476 623 7488 799
rect 7522 623 7562 799
rect 7476 611 7562 623
rect 4936 419 4948 607
rect 4890 407 4948 419
rect 7550 423 7562 611
rect 7596 423 7608 799
rect 7550 411 7608 423
rect 7668 799 7726 811
rect 7668 423 7680 799
rect 7714 423 7726 799
rect 7668 411 7726 423
rect 7786 799 7844 811
rect 7786 423 7798 799
rect 7832 423 7844 799
rect 7786 411 7844 423
rect 7904 799 7962 811
rect 7904 423 7916 799
rect 7950 423 7962 799
rect 7904 411 7962 423
rect 8022 799 8158 811
rect 8022 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8158 799
rect 8068 611 8158 623
rect 8218 799 8276 811
rect 8218 623 8230 799
rect 8264 623 8276 799
rect 8218 611 8276 623
rect 10502 799 10560 811
rect 10502 623 10514 799
rect 10548 623 10560 799
rect 10502 611 10560 623
rect 10620 799 10752 811
rect 10620 623 10632 799
rect 10666 623 10706 799
rect 10620 611 10706 623
rect 8068 423 8080 611
rect 8022 411 8080 423
rect 10694 423 10706 611
rect 10740 423 10752 799
rect 10694 411 10752 423
rect 10812 799 10870 811
rect 10812 423 10824 799
rect 10858 423 10870 799
rect 10812 411 10870 423
rect 10930 799 10988 811
rect 10930 423 10942 799
rect 10976 423 10988 799
rect 10930 411 10988 423
rect 11048 799 11106 811
rect 11048 423 11060 799
rect 11094 423 11106 799
rect 11048 411 11106 423
rect 11166 799 11302 811
rect 11166 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11302 799
rect 11212 611 11302 623
rect 11362 799 11420 811
rect 31375 1927 31775 1939
rect 31375 1893 31387 1927
rect 31763 1893 31775 1927
rect 38027 2103 38085 2115
rect 31375 1881 31775 1893
rect 31375 1809 31775 1821
rect 31375 1775 31387 1809
rect 31763 1775 31775 1809
rect 31375 1763 31775 1775
rect 38027 1727 38039 2103
rect 38073 1727 38085 2103
rect 38027 1715 38085 1727
rect 38145 2103 38203 2115
rect 38145 1727 38157 2103
rect 38191 1727 38203 2103
rect 38145 1715 38203 1727
rect 38263 2103 38321 2115
rect 38263 1727 38275 2103
rect 38309 1727 38321 2103
rect 38380 2103 38438 2115
rect 38380 1927 38392 2103
rect 38426 1927 38438 2103
rect 38380 1915 38438 1927
rect 38498 2103 38556 2115
rect 38498 1927 38510 2103
rect 38544 1927 38556 2103
rect 38498 1915 38556 1927
rect 38263 1715 38321 1727
rect 44578 2101 44636 2113
rect 31375 1403 31575 1415
rect 31375 1369 31387 1403
rect 31563 1369 31575 1403
rect 31375 1357 31575 1369
rect 31375 1285 31575 1297
rect 31375 1251 31387 1285
rect 31563 1251 31575 1285
rect 31375 1239 31575 1251
rect 35120 1177 35178 1189
rect 11362 623 11374 799
rect 11408 623 11420 799
rect 11362 611 11420 623
rect 13704 795 13762 807
rect 13704 619 13716 795
rect 13750 619 13762 795
rect 11212 423 11224 611
rect 11166 411 11224 423
rect 13704 607 13762 619
rect 13822 795 13954 807
rect 13822 619 13834 795
rect 13868 619 13908 795
rect 13822 607 13908 619
rect 13896 419 13908 607
rect 13942 419 13954 795
rect 13896 407 13954 419
rect 14014 795 14072 807
rect 14014 419 14026 795
rect 14060 419 14072 795
rect 14014 407 14072 419
rect 14132 795 14190 807
rect 14132 419 14144 795
rect 14178 419 14190 795
rect 14132 407 14190 419
rect 14250 795 14308 807
rect 14250 419 14262 795
rect 14296 419 14308 795
rect 14250 407 14308 419
rect 14368 795 14504 807
rect 14368 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14504 795
rect 14414 607 14504 619
rect 14564 795 14622 807
rect 14564 619 14576 795
rect 14610 619 14622 795
rect 14564 607 14622 619
rect 16848 795 16906 807
rect 16848 619 16860 795
rect 16894 619 16906 795
rect 16848 607 16906 619
rect 16966 795 17098 807
rect 16966 619 16978 795
rect 17012 619 17052 795
rect 16966 607 17052 619
rect 14414 419 14426 607
rect 14368 407 14426 419
rect 17040 419 17052 607
rect 17086 419 17098 795
rect 17040 407 17098 419
rect 17158 795 17216 807
rect 17158 419 17170 795
rect 17204 419 17216 795
rect 17158 407 17216 419
rect 17276 795 17334 807
rect 17276 419 17288 795
rect 17322 419 17334 795
rect 17276 407 17334 419
rect 17394 795 17452 807
rect 17394 419 17406 795
rect 17440 419 17452 795
rect 17394 407 17452 419
rect 17512 795 17648 807
rect 17512 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17648 795
rect 17558 607 17648 619
rect 17708 795 17766 807
rect 17708 619 17720 795
rect 17754 619 17766 795
rect 17708 607 17766 619
rect 19980 799 20038 811
rect 19980 623 19992 799
rect 20026 623 20038 799
rect 19980 611 20038 623
rect 20098 799 20230 811
rect 20098 623 20110 799
rect 20144 623 20184 799
rect 20098 611 20184 623
rect 17558 419 17570 607
rect 17512 407 17570 419
rect 20172 423 20184 611
rect 20218 423 20230 799
rect 20172 411 20230 423
rect 20290 799 20348 811
rect 20290 423 20302 799
rect 20336 423 20348 799
rect 20290 411 20348 423
rect 20408 799 20466 811
rect 20408 423 20420 799
rect 20454 423 20466 799
rect 20408 411 20466 423
rect 20526 799 20584 811
rect 20526 423 20538 799
rect 20572 423 20584 799
rect 20526 411 20584 423
rect 20644 799 20780 811
rect 20644 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20780 799
rect 20690 611 20780 623
rect 20840 799 20898 811
rect 20840 623 20852 799
rect 20886 623 20898 799
rect 20840 611 20898 623
rect 23124 799 23182 811
rect 23124 623 23136 799
rect 23170 623 23182 799
rect 23124 611 23182 623
rect 23242 799 23374 811
rect 23242 623 23254 799
rect 23288 623 23328 799
rect 23242 611 23328 623
rect 20690 423 20702 611
rect 20644 411 20702 423
rect 23316 423 23328 611
rect 23362 423 23374 799
rect 23316 411 23374 423
rect 23434 799 23492 811
rect 23434 423 23446 799
rect 23480 423 23492 799
rect 23434 411 23492 423
rect 23552 799 23610 811
rect 23552 423 23564 799
rect 23598 423 23610 799
rect 23552 411 23610 423
rect 23670 799 23728 811
rect 23670 423 23682 799
rect 23716 423 23728 799
rect 23670 411 23728 423
rect 23788 799 23924 811
rect 23788 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23924 799
rect 23834 611 23924 623
rect 23984 799 24042 811
rect 23984 623 23996 799
rect 24030 623 24042 799
rect 35120 801 35132 1177
rect 35166 801 35178 1177
rect 35120 789 35178 801
rect 35238 1177 35296 1189
rect 35238 801 35250 1177
rect 35284 801 35296 1177
rect 35238 789 35296 801
rect 35356 1177 35414 1189
rect 35356 801 35368 1177
rect 35402 801 35414 1177
rect 35473 1177 35531 1189
rect 35473 1001 35485 1177
rect 35519 1001 35531 1177
rect 35473 989 35531 1001
rect 35591 1177 35649 1189
rect 35591 1001 35603 1177
rect 35637 1001 35649 1177
rect 35591 989 35649 1001
rect 35356 789 35414 801
rect 23984 611 24042 623
rect 23834 423 23846 611
rect 23788 411 23846 423
rect 31377 632 31577 644
rect 31377 598 31389 632
rect 31565 598 31577 632
rect 31377 586 31577 598
rect 31377 514 31577 526
rect 31377 480 31389 514
rect 31565 480 31577 514
rect 44578 1725 44590 2101
rect 44624 1725 44636 2101
rect 44578 1713 44636 1725
rect 44696 2101 44754 2113
rect 44696 1725 44708 2101
rect 44742 1725 44754 2101
rect 44696 1713 44754 1725
rect 44814 2101 44872 2113
rect 44814 1725 44826 2101
rect 44860 1725 44872 2101
rect 44931 2101 44989 2113
rect 44931 1925 44943 2101
rect 44977 1925 44989 2101
rect 44931 1913 44989 1925
rect 45049 2101 45107 2113
rect 45049 1925 45061 2101
rect 45095 1925 45107 2101
rect 45049 1913 45107 1925
rect 44814 1713 44872 1725
rect 51233 2102 51291 2114
rect 39379 698 39437 710
rect 39379 522 39391 698
rect 39425 522 39437 698
rect 31377 468 31577 480
rect 38022 499 38080 511
rect 31377 212 31777 224
rect 31377 178 31389 212
rect 31765 178 31777 212
rect 31377 166 31777 178
rect 38022 123 38034 499
rect 38068 123 38080 499
rect 38022 111 38080 123
rect 38140 499 38198 511
rect 38140 123 38152 499
rect 38186 123 38198 499
rect 38140 111 38198 123
rect 38258 499 38316 511
rect 38258 123 38270 499
rect 38304 123 38316 499
rect 38375 499 38433 511
rect 38375 323 38387 499
rect 38421 323 38433 499
rect 38375 311 38433 323
rect 38493 499 38551 511
rect 39379 510 39437 522
rect 39497 698 39555 710
rect 39497 522 39509 698
rect 39543 522 39555 698
rect 39497 510 39555 522
rect 39799 698 39857 710
rect 38493 323 38505 499
rect 38539 323 38551 499
rect 38493 311 38551 323
rect 39799 322 39811 698
rect 39845 322 39857 698
rect 39799 310 39857 322
rect 39917 698 39975 710
rect 39917 322 39929 698
rect 39963 322 39975 698
rect 39917 310 39975 322
rect 40035 698 40093 710
rect 40035 322 40047 698
rect 40081 322 40093 698
rect 40035 310 40093 322
rect 40153 698 40211 710
rect 40153 322 40165 698
rect 40199 322 40211 698
rect 40153 310 40211 322
rect 40271 698 40329 710
rect 40271 322 40283 698
rect 40317 322 40329 698
rect 40677 698 40735 710
rect 40677 522 40689 698
rect 40723 522 40735 698
rect 40677 510 40735 522
rect 40795 698 40853 710
rect 40795 522 40807 698
rect 40841 522 40853 698
rect 40795 510 40853 522
rect 41277 698 41335 710
rect 41277 522 41289 698
rect 41323 522 41335 698
rect 41277 510 41335 522
rect 41395 698 41453 710
rect 41395 522 41407 698
rect 41441 522 41453 698
rect 41395 510 41453 522
rect 41697 698 41755 710
rect 40271 310 40329 322
rect 41697 322 41709 698
rect 41743 322 41755 698
rect 41697 310 41755 322
rect 41815 698 41873 710
rect 41815 322 41827 698
rect 41861 322 41873 698
rect 41815 310 41873 322
rect 41933 698 41991 710
rect 41933 322 41945 698
rect 41979 322 41991 698
rect 41933 310 41991 322
rect 42051 698 42109 710
rect 42051 322 42063 698
rect 42097 322 42109 698
rect 42051 310 42109 322
rect 42169 698 42227 710
rect 42169 322 42181 698
rect 42215 322 42227 698
rect 42575 698 42633 710
rect 42575 522 42587 698
rect 42621 522 42633 698
rect 42575 510 42633 522
rect 42693 698 42751 710
rect 42693 522 42705 698
rect 42739 522 42751 698
rect 42693 510 42751 522
rect 51233 1726 51245 2102
rect 51279 1726 51291 2102
rect 51233 1714 51291 1726
rect 51351 2102 51409 2114
rect 51351 1726 51363 2102
rect 51397 1726 51409 2102
rect 51351 1714 51409 1726
rect 51469 2102 51527 2114
rect 51469 1726 51481 2102
rect 51515 1726 51527 2102
rect 51586 2102 51644 2114
rect 51586 1926 51598 2102
rect 51632 1926 51644 2102
rect 51586 1914 51644 1926
rect 51704 2102 51762 2114
rect 51704 1926 51716 2102
rect 51750 1926 51762 2102
rect 51704 1914 51762 1926
rect 51469 1714 51527 1726
rect 57855 2103 57913 2115
rect 45930 696 45988 708
rect 45930 520 45942 696
rect 45976 520 45988 696
rect 44573 497 44631 509
rect 42169 310 42227 322
rect 38258 111 38316 123
rect 31377 94 31777 106
rect 31377 60 31389 94
rect 31765 60 31777 94
rect 31377 48 31777 60
rect 44573 121 44585 497
rect 44619 121 44631 497
rect 44573 109 44631 121
rect 44691 497 44749 509
rect 44691 121 44703 497
rect 44737 121 44749 497
rect 44691 109 44749 121
rect 44809 497 44867 509
rect 44809 121 44821 497
rect 44855 121 44867 497
rect 44926 497 44984 509
rect 44926 321 44938 497
rect 44972 321 44984 497
rect 44926 309 44984 321
rect 45044 497 45102 509
rect 45930 508 45988 520
rect 46048 696 46106 708
rect 46048 520 46060 696
rect 46094 520 46106 696
rect 46048 508 46106 520
rect 46350 696 46408 708
rect 45044 321 45056 497
rect 45090 321 45102 497
rect 45044 309 45102 321
rect 46350 320 46362 696
rect 46396 320 46408 696
rect 46350 308 46408 320
rect 46468 696 46526 708
rect 46468 320 46480 696
rect 46514 320 46526 696
rect 46468 308 46526 320
rect 46586 696 46644 708
rect 46586 320 46598 696
rect 46632 320 46644 696
rect 46586 308 46644 320
rect 46704 696 46762 708
rect 46704 320 46716 696
rect 46750 320 46762 696
rect 46704 308 46762 320
rect 46822 696 46880 708
rect 46822 320 46834 696
rect 46868 320 46880 696
rect 47228 696 47286 708
rect 47228 520 47240 696
rect 47274 520 47286 696
rect 47228 508 47286 520
rect 47346 696 47404 708
rect 47346 520 47358 696
rect 47392 520 47404 696
rect 47346 508 47404 520
rect 47828 696 47886 708
rect 47828 520 47840 696
rect 47874 520 47886 696
rect 47828 508 47886 520
rect 47946 696 48004 708
rect 47946 520 47958 696
rect 47992 520 48004 696
rect 47946 508 48004 520
rect 48248 696 48306 708
rect 46822 308 46880 320
rect 48248 320 48260 696
rect 48294 320 48306 696
rect 48248 308 48306 320
rect 48366 696 48424 708
rect 48366 320 48378 696
rect 48412 320 48424 696
rect 48366 308 48424 320
rect 48484 696 48542 708
rect 48484 320 48496 696
rect 48530 320 48542 696
rect 48484 308 48542 320
rect 48602 696 48660 708
rect 48602 320 48614 696
rect 48648 320 48660 696
rect 48602 308 48660 320
rect 48720 696 48778 708
rect 48720 320 48732 696
rect 48766 320 48778 696
rect 49126 696 49184 708
rect 49126 520 49138 696
rect 49172 520 49184 696
rect 49126 508 49184 520
rect 49244 696 49302 708
rect 49244 520 49256 696
rect 49290 520 49302 696
rect 49244 508 49302 520
rect 57855 1727 57867 2103
rect 57901 1727 57913 2103
rect 57855 1715 57913 1727
rect 57973 2103 58031 2115
rect 57973 1727 57985 2103
rect 58019 1727 58031 2103
rect 57973 1715 58031 1727
rect 58091 2103 58149 2115
rect 58091 1727 58103 2103
rect 58137 1727 58149 2103
rect 58208 2103 58266 2115
rect 58208 1927 58220 2103
rect 58254 1927 58266 2103
rect 58208 1915 58266 1927
rect 58326 2103 58384 2115
rect 58326 1927 58338 2103
rect 58372 1927 58384 2103
rect 58326 1915 58384 1927
rect 58091 1715 58149 1727
rect 71842 2329 72042 2341
rect 71842 2295 71854 2329
rect 72030 2295 72042 2329
rect 71842 2283 72042 2295
rect 71842 2211 72042 2223
rect 71842 2177 71854 2211
rect 72030 2177 72042 2211
rect 71842 2149 72042 2177
rect 71842 2137 72242 2149
rect 71842 2103 71854 2137
rect 72230 2103 72242 2137
rect 71842 2091 72242 2103
rect 71842 2019 72242 2031
rect 71842 1985 71854 2019
rect 72230 1985 72242 2019
rect 71842 1973 72242 1985
rect 52585 697 52643 709
rect 52585 521 52597 697
rect 52631 521 52643 697
rect 51228 498 51286 510
rect 48720 308 48778 320
rect 44809 109 44867 121
rect 31377 -24 31777 -12
rect 31377 -58 31389 -24
rect 31765 -58 31777 -24
rect 31377 -70 31777 -58
rect 31377 -142 31777 -130
rect 31377 -176 31389 -142
rect 31765 -176 31777 -142
rect 51228 122 51240 498
rect 51274 122 51286 498
rect 51228 110 51286 122
rect 51346 498 51404 510
rect 51346 122 51358 498
rect 51392 122 51404 498
rect 51346 110 51404 122
rect 51464 498 51522 510
rect 51464 122 51476 498
rect 51510 122 51522 498
rect 51581 498 51639 510
rect 51581 322 51593 498
rect 51627 322 51639 498
rect 51581 310 51639 322
rect 51699 498 51757 510
rect 52585 509 52643 521
rect 52703 697 52761 709
rect 52703 521 52715 697
rect 52749 521 52761 697
rect 52703 509 52761 521
rect 53005 697 53063 709
rect 51699 322 51711 498
rect 51745 322 51757 498
rect 51699 310 51757 322
rect 53005 321 53017 697
rect 53051 321 53063 697
rect 53005 309 53063 321
rect 53123 697 53181 709
rect 53123 321 53135 697
rect 53169 321 53181 697
rect 53123 309 53181 321
rect 53241 697 53299 709
rect 53241 321 53253 697
rect 53287 321 53299 697
rect 53241 309 53299 321
rect 53359 697 53417 709
rect 53359 321 53371 697
rect 53405 321 53417 697
rect 53359 309 53417 321
rect 53477 697 53535 709
rect 53477 321 53489 697
rect 53523 321 53535 697
rect 53883 697 53941 709
rect 53883 521 53895 697
rect 53929 521 53941 697
rect 53883 509 53941 521
rect 54001 697 54059 709
rect 54001 521 54013 697
rect 54047 521 54059 697
rect 54001 509 54059 521
rect 54483 697 54541 709
rect 54483 521 54495 697
rect 54529 521 54541 697
rect 54483 509 54541 521
rect 54601 697 54659 709
rect 54601 521 54613 697
rect 54647 521 54659 697
rect 54601 509 54659 521
rect 54903 697 54961 709
rect 53477 309 53535 321
rect 54903 321 54915 697
rect 54949 321 54961 697
rect 54903 309 54961 321
rect 55021 697 55079 709
rect 55021 321 55033 697
rect 55067 321 55079 697
rect 55021 309 55079 321
rect 55139 697 55197 709
rect 55139 321 55151 697
rect 55185 321 55197 697
rect 55139 309 55197 321
rect 55257 697 55315 709
rect 55257 321 55269 697
rect 55303 321 55315 697
rect 55257 309 55315 321
rect 55375 697 55433 709
rect 55375 321 55387 697
rect 55421 321 55433 697
rect 55781 697 55839 709
rect 55781 521 55793 697
rect 55827 521 55839 697
rect 55781 509 55839 521
rect 55899 697 55957 709
rect 55899 521 55911 697
rect 55945 521 55957 697
rect 55899 509 55957 521
rect 71842 1901 72242 1913
rect 71842 1867 71854 1901
rect 72230 1867 72242 1901
rect 71842 1855 72242 1867
rect 71842 1783 72242 1795
rect 71842 1749 71854 1783
rect 72230 1749 72242 1783
rect 71842 1737 72242 1749
rect 71842 1665 72242 1677
rect 71842 1631 71854 1665
rect 72230 1631 72242 1665
rect 71842 1619 72242 1631
rect 71842 1587 72042 1619
rect 71842 1553 71854 1587
rect 72030 1553 72042 1587
rect 71842 1541 72042 1553
rect 63714 959 63772 971
rect 59207 698 59265 710
rect 59207 522 59219 698
rect 59253 522 59265 698
rect 57850 499 57908 511
rect 55375 309 55433 321
rect 51464 110 51522 122
rect 57850 123 57862 499
rect 57896 123 57908 499
rect 57850 111 57908 123
rect 57968 499 58026 511
rect 57968 123 57980 499
rect 58014 123 58026 499
rect 57968 111 58026 123
rect 58086 499 58144 511
rect 58086 123 58098 499
rect 58132 123 58144 499
rect 58203 499 58261 511
rect 58203 323 58215 499
rect 58249 323 58261 499
rect 58203 311 58261 323
rect 58321 499 58379 511
rect 59207 510 59265 522
rect 59325 698 59383 710
rect 59325 522 59337 698
rect 59371 522 59383 698
rect 59325 510 59383 522
rect 59627 698 59685 710
rect 58321 323 58333 499
rect 58367 323 58379 499
rect 58321 311 58379 323
rect 59627 322 59639 698
rect 59673 322 59685 698
rect 59627 310 59685 322
rect 59745 698 59803 710
rect 59745 322 59757 698
rect 59791 322 59803 698
rect 59745 310 59803 322
rect 59863 698 59921 710
rect 59863 322 59875 698
rect 59909 322 59921 698
rect 59863 310 59921 322
rect 59981 698 60039 710
rect 59981 322 59993 698
rect 60027 322 60039 698
rect 59981 310 60039 322
rect 60099 698 60157 710
rect 60099 322 60111 698
rect 60145 322 60157 698
rect 60505 698 60563 710
rect 60505 522 60517 698
rect 60551 522 60563 698
rect 60505 510 60563 522
rect 60623 698 60681 710
rect 60623 522 60635 698
rect 60669 522 60681 698
rect 60623 510 60681 522
rect 61105 698 61163 710
rect 61105 522 61117 698
rect 61151 522 61163 698
rect 61105 510 61163 522
rect 61223 698 61281 710
rect 61223 522 61235 698
rect 61269 522 61281 698
rect 61223 510 61281 522
rect 61525 698 61583 710
rect 60099 310 60157 322
rect 61525 322 61537 698
rect 61571 322 61583 698
rect 61525 310 61583 322
rect 61643 698 61701 710
rect 61643 322 61655 698
rect 61689 322 61701 698
rect 61643 310 61701 322
rect 61761 698 61819 710
rect 61761 322 61773 698
rect 61807 322 61819 698
rect 61761 310 61819 322
rect 61879 698 61937 710
rect 61879 322 61891 698
rect 61925 322 61937 698
rect 61879 310 61937 322
rect 61997 698 62055 710
rect 61997 322 62009 698
rect 62043 322 62055 698
rect 62403 698 62461 710
rect 62403 522 62415 698
rect 62449 522 62461 698
rect 62403 510 62461 522
rect 62521 698 62579 710
rect 62521 522 62533 698
rect 62567 522 62579 698
rect 63714 583 63726 959
rect 63760 583 63772 959
rect 63714 571 63772 583
rect 63832 959 63890 971
rect 63832 583 63844 959
rect 63878 583 63890 959
rect 63832 571 63890 583
rect 63950 959 64008 971
rect 63950 583 63962 959
rect 63996 583 64008 959
rect 64067 959 64125 971
rect 64067 783 64079 959
rect 64113 783 64125 959
rect 64067 771 64125 783
rect 64185 959 64243 971
rect 64185 783 64197 959
rect 64231 783 64243 959
rect 64185 771 64243 783
rect 71842 1469 72042 1481
rect 71842 1435 71854 1469
rect 72030 1435 72042 1469
rect 71842 1423 72042 1435
rect 63950 571 64008 583
rect 62521 510 62579 522
rect 61997 310 62055 322
rect 58086 111 58144 123
rect 31377 -188 31777 -176
rect 31377 -260 31777 -248
rect 31377 -294 31389 -260
rect 31765 -294 31777 -260
rect 31377 -306 31777 -294
rect 31377 -666 31577 -654
rect 31377 -700 31389 -666
rect 31565 -700 31577 -666
rect 31377 -712 31577 -700
rect 31377 -784 31577 -772
rect 31377 -818 31389 -784
rect 31565 -818 31577 -784
rect 31377 -830 31577 -818
rect 41830 -930 41888 -918
rect 41830 -1306 41842 -930
rect 41876 -1306 41888 -930
rect 41830 -1318 41888 -1306
rect 41948 -930 42006 -918
rect 41948 -1306 41960 -930
rect 41994 -1306 42006 -930
rect 41948 -1318 42006 -1306
rect 42066 -930 42124 -918
rect 42066 -1306 42078 -930
rect 42112 -1306 42124 -930
rect 48384 -925 48442 -913
rect 42066 -1318 42124 -1306
rect 42183 -1130 42241 -1118
rect 42183 -1306 42195 -1130
rect 42229 -1306 42241 -1130
rect 42183 -1318 42241 -1306
rect 42301 -1130 42359 -1118
rect 42301 -1306 42313 -1130
rect 42347 -1306 42359 -1130
rect 42301 -1318 42359 -1306
rect 48384 -1301 48396 -925
rect 48430 -1301 48442 -925
rect 48384 -1313 48442 -1301
rect 48502 -925 48560 -913
rect 48502 -1301 48514 -925
rect 48548 -1301 48560 -925
rect 48502 -1313 48560 -1301
rect 48620 -925 48678 -913
rect 48620 -1301 48632 -925
rect 48666 -1301 48678 -925
rect 55033 -937 55091 -925
rect 48620 -1313 48678 -1301
rect 48737 -1125 48795 -1113
rect 48737 -1301 48749 -1125
rect 48783 -1301 48795 -1125
rect 48737 -1313 48795 -1301
rect 48855 -1125 48913 -1113
rect 48855 -1301 48867 -1125
rect 48901 -1301 48913 -1125
rect 48855 -1313 48913 -1301
rect 55033 -1313 55045 -937
rect 55079 -1313 55091 -937
rect 31375 -1436 31575 -1424
rect 31375 -1470 31387 -1436
rect 31563 -1470 31575 -1436
rect 31375 -1482 31575 -1470
rect 31375 -1554 31575 -1542
rect 31375 -1588 31387 -1554
rect 31563 -1588 31575 -1554
rect 55033 -1325 55091 -1313
rect 55151 -937 55209 -925
rect 55151 -1313 55163 -937
rect 55197 -1313 55209 -937
rect 55151 -1325 55209 -1313
rect 55269 -937 55327 -925
rect 55269 -1313 55281 -937
rect 55315 -1313 55327 -937
rect 55269 -1325 55327 -1313
rect 55386 -1137 55444 -1125
rect 55386 -1313 55398 -1137
rect 55432 -1313 55444 -1137
rect 55386 -1325 55444 -1313
rect 55504 -1137 55562 -1125
rect 55504 -1313 55516 -1137
rect 55550 -1313 55562 -1137
rect 55504 -1325 55562 -1313
rect 31375 -1600 31575 -1588
rect 67254 -789 67312 -777
rect 67254 -1165 67266 -789
rect 67300 -1165 67312 -789
rect 67254 -1177 67312 -1165
rect 67372 -789 67430 -777
rect 67372 -1165 67384 -789
rect 67418 -1165 67430 -789
rect 67372 -1177 67430 -1165
rect 67490 -789 67548 -777
rect 67490 -1165 67502 -789
rect 67536 -1165 67548 -789
rect 67607 -789 67665 -777
rect 67607 -965 67619 -789
rect 67653 -965 67665 -789
rect 67607 -977 67665 -965
rect 67725 -789 67783 -777
rect 67725 -965 67737 -789
rect 67771 -965 67783 -789
rect 67725 -977 67783 -965
rect 71842 -815 72042 -803
rect 71842 -849 71854 -815
rect 72030 -849 72042 -815
rect 71842 -861 72042 -849
rect 71842 -933 72042 -921
rect 71842 -967 71854 -933
rect 72030 -967 72042 -933
rect 71842 -995 72042 -967
rect 71842 -1007 72242 -995
rect 71842 -1041 71854 -1007
rect 72230 -1041 72242 -1007
rect 71842 -1053 72242 -1041
rect 67490 -1177 67548 -1165
rect 71842 -1125 72242 -1113
rect 71842 -1159 71854 -1125
rect 72230 -1159 72242 -1125
rect 71842 -1171 72242 -1159
rect 71842 -1243 72242 -1231
rect 71842 -1277 71854 -1243
rect 72230 -1277 72242 -1243
rect 71842 -1289 72242 -1277
rect 71842 -1361 72242 -1349
rect 71842 -1395 71854 -1361
rect 72230 -1395 72242 -1361
rect 71842 -1407 72242 -1395
rect 65349 -1574 65407 -1562
rect 31375 -1856 31775 -1844
rect 31375 -1890 31387 -1856
rect 31763 -1890 31775 -1856
rect 65349 -1750 65361 -1574
rect 65395 -1750 65407 -1574
rect 65349 -1762 65407 -1750
rect 65467 -1574 65525 -1562
rect 65467 -1750 65479 -1574
rect 65513 -1750 65525 -1574
rect 65467 -1762 65525 -1750
rect 65769 -1574 65827 -1562
rect 63721 -1886 63779 -1874
rect 31375 -1902 31775 -1890
rect 1114 -3097 1172 -3085
rect 1114 -3273 1126 -3097
rect 1160 -3273 1172 -3097
rect 1114 -3285 1172 -3273
rect 1232 -3097 1364 -3085
rect 1232 -3273 1244 -3097
rect 1278 -3273 1318 -3097
rect 1232 -3285 1318 -3273
rect 1306 -3473 1318 -3285
rect 1352 -3473 1364 -3097
rect 1306 -3485 1364 -3473
rect 1424 -3097 1482 -3085
rect 1424 -3473 1436 -3097
rect 1470 -3473 1482 -3097
rect 1424 -3485 1482 -3473
rect 1542 -3097 1600 -3085
rect 1542 -3473 1554 -3097
rect 1588 -3473 1600 -3097
rect 1542 -3485 1600 -3473
rect 1660 -3097 1718 -3085
rect 1660 -3473 1672 -3097
rect 1706 -3473 1718 -3097
rect 1660 -3485 1718 -3473
rect 1778 -3097 1914 -3085
rect 1778 -3473 1790 -3097
rect 1824 -3273 1868 -3097
rect 1902 -3273 1914 -3097
rect 1824 -3285 1914 -3273
rect 1974 -3097 2032 -3085
rect 1974 -3273 1986 -3097
rect 2020 -3273 2032 -3097
rect 1974 -3285 2032 -3273
rect 4258 -3097 4316 -3085
rect 4258 -3273 4270 -3097
rect 4304 -3273 4316 -3097
rect 4258 -3285 4316 -3273
rect 4376 -3097 4508 -3085
rect 4376 -3273 4388 -3097
rect 4422 -3273 4462 -3097
rect 4376 -3285 4462 -3273
rect 1824 -3473 1836 -3285
rect 1778 -3485 1836 -3473
rect 4450 -3473 4462 -3285
rect 4496 -3473 4508 -3097
rect 4450 -3485 4508 -3473
rect 4568 -3097 4626 -3085
rect 4568 -3473 4580 -3097
rect 4614 -3473 4626 -3097
rect 4568 -3485 4626 -3473
rect 4686 -3097 4744 -3085
rect 4686 -3473 4698 -3097
rect 4732 -3473 4744 -3097
rect 4686 -3485 4744 -3473
rect 4804 -3097 4862 -3085
rect 4804 -3473 4816 -3097
rect 4850 -3473 4862 -3097
rect 4804 -3485 4862 -3473
rect 4922 -3097 5058 -3085
rect 4922 -3473 4934 -3097
rect 4968 -3273 5012 -3097
rect 5046 -3273 5058 -3097
rect 4968 -3285 5058 -3273
rect 5118 -3097 5176 -3085
rect 5118 -3273 5130 -3097
rect 5164 -3273 5176 -3097
rect 5118 -3285 5176 -3273
rect 7390 -3093 7448 -3081
rect 7390 -3269 7402 -3093
rect 7436 -3269 7448 -3093
rect 7390 -3281 7448 -3269
rect 7508 -3093 7640 -3081
rect 7508 -3269 7520 -3093
rect 7554 -3269 7594 -3093
rect 7508 -3281 7594 -3269
rect 4968 -3473 4980 -3285
rect 4922 -3485 4980 -3473
rect 7582 -3469 7594 -3281
rect 7628 -3469 7640 -3093
rect 7582 -3481 7640 -3469
rect 7700 -3093 7758 -3081
rect 7700 -3469 7712 -3093
rect 7746 -3469 7758 -3093
rect 7700 -3481 7758 -3469
rect 7818 -3093 7876 -3081
rect 7818 -3469 7830 -3093
rect 7864 -3469 7876 -3093
rect 7818 -3481 7876 -3469
rect 7936 -3093 7994 -3081
rect 7936 -3469 7948 -3093
rect 7982 -3469 7994 -3093
rect 7936 -3481 7994 -3469
rect 8054 -3093 8190 -3081
rect 8054 -3469 8066 -3093
rect 8100 -3269 8144 -3093
rect 8178 -3269 8190 -3093
rect 8100 -3281 8190 -3269
rect 8250 -3093 8308 -3081
rect 8250 -3269 8262 -3093
rect 8296 -3269 8308 -3093
rect 8250 -3281 8308 -3269
rect 10534 -3093 10592 -3081
rect 10534 -3269 10546 -3093
rect 10580 -3269 10592 -3093
rect 10534 -3281 10592 -3269
rect 10652 -3093 10784 -3081
rect 10652 -3269 10664 -3093
rect 10698 -3269 10738 -3093
rect 10652 -3281 10738 -3269
rect 8100 -3469 8112 -3281
rect 8054 -3481 8112 -3469
rect 10726 -3469 10738 -3281
rect 10772 -3469 10784 -3093
rect 10726 -3481 10784 -3469
rect 10844 -3093 10902 -3081
rect 10844 -3469 10856 -3093
rect 10890 -3469 10902 -3093
rect 10844 -3481 10902 -3469
rect 10962 -3093 11020 -3081
rect 10962 -3469 10974 -3093
rect 11008 -3469 11020 -3093
rect 10962 -3481 11020 -3469
rect 11080 -3093 11138 -3081
rect 11080 -3469 11092 -3093
rect 11126 -3469 11138 -3093
rect 11080 -3481 11138 -3469
rect 11198 -3093 11334 -3081
rect 11198 -3469 11210 -3093
rect 11244 -3269 11288 -3093
rect 11322 -3269 11334 -3093
rect 11244 -3281 11334 -3269
rect 11394 -3093 11452 -3081
rect 31375 -1974 31775 -1962
rect 31375 -2008 31387 -1974
rect 31763 -2008 31775 -1974
rect 31375 -2020 31775 -2008
rect 31375 -2092 31775 -2080
rect 31375 -2126 31387 -2092
rect 31763 -2126 31775 -2092
rect 31375 -2138 31775 -2126
rect 31375 -2210 31775 -2198
rect 31375 -2244 31387 -2210
rect 31763 -2244 31775 -2210
rect 31375 -2256 31775 -2244
rect 63721 -2262 63733 -1886
rect 63767 -2262 63779 -1886
rect 63721 -2274 63779 -2262
rect 63839 -1886 63897 -1874
rect 63839 -2262 63851 -1886
rect 63885 -2262 63897 -1886
rect 63839 -2274 63897 -2262
rect 63957 -1886 64015 -1874
rect 63957 -2262 63969 -1886
rect 64003 -2262 64015 -1886
rect 64074 -1886 64132 -1874
rect 64074 -2062 64086 -1886
rect 64120 -2062 64132 -1886
rect 64074 -2074 64132 -2062
rect 64192 -1886 64250 -1874
rect 64192 -2062 64204 -1886
rect 64238 -2062 64250 -1886
rect 65769 -1950 65781 -1574
rect 65815 -1950 65827 -1574
rect 65769 -1962 65827 -1950
rect 65887 -1574 65945 -1562
rect 65887 -1950 65899 -1574
rect 65933 -1950 65945 -1574
rect 65887 -1962 65945 -1950
rect 66005 -1574 66063 -1562
rect 66005 -1950 66017 -1574
rect 66051 -1950 66063 -1574
rect 66005 -1962 66063 -1950
rect 66123 -1574 66181 -1562
rect 66123 -1950 66135 -1574
rect 66169 -1950 66181 -1574
rect 66123 -1962 66181 -1950
rect 66241 -1574 66299 -1562
rect 66241 -1950 66253 -1574
rect 66287 -1950 66299 -1574
rect 66647 -1574 66705 -1562
rect 66647 -1750 66659 -1574
rect 66693 -1750 66705 -1574
rect 66647 -1762 66705 -1750
rect 66765 -1574 66823 -1562
rect 66765 -1750 66777 -1574
rect 66811 -1750 66823 -1574
rect 66765 -1762 66823 -1750
rect 66241 -1962 66299 -1950
rect 71842 -1479 72242 -1467
rect 71842 -1513 71854 -1479
rect 72230 -1513 72242 -1479
rect 71842 -1525 72242 -1513
rect 71842 -1557 72042 -1525
rect 71842 -1591 71854 -1557
rect 72030 -1591 72042 -1557
rect 71842 -1603 72042 -1591
rect 64192 -2074 64250 -2062
rect 63957 -2274 64015 -2262
rect 31375 -2328 31775 -2316
rect 31375 -2362 31387 -2328
rect 31763 -2362 31775 -2328
rect 31375 -2374 31775 -2362
rect 71842 -1675 72042 -1663
rect 71842 -1709 71854 -1675
rect 72030 -1709 72042 -1675
rect 71842 -1721 72042 -1709
rect 31375 -2734 31575 -2722
rect 31375 -2768 31387 -2734
rect 31563 -2768 31575 -2734
rect 31375 -2780 31575 -2768
rect 31375 -2852 31575 -2840
rect 31375 -2886 31387 -2852
rect 31563 -2886 31575 -2852
rect 31375 -2898 31575 -2886
rect 11394 -3269 11406 -3093
rect 11440 -3269 11452 -3093
rect 11394 -3281 11452 -3269
rect 13736 -3097 13794 -3085
rect 13736 -3273 13748 -3097
rect 13782 -3273 13794 -3097
rect 11244 -3469 11256 -3281
rect 11198 -3481 11256 -3469
rect 13736 -3285 13794 -3273
rect 13854 -3097 13986 -3085
rect 13854 -3273 13866 -3097
rect 13900 -3273 13940 -3097
rect 13854 -3285 13940 -3273
rect 13928 -3473 13940 -3285
rect 13974 -3473 13986 -3097
rect 13928 -3485 13986 -3473
rect 14046 -3097 14104 -3085
rect 14046 -3473 14058 -3097
rect 14092 -3473 14104 -3097
rect 14046 -3485 14104 -3473
rect 14164 -3097 14222 -3085
rect 14164 -3473 14176 -3097
rect 14210 -3473 14222 -3097
rect 14164 -3485 14222 -3473
rect 14282 -3097 14340 -3085
rect 14282 -3473 14294 -3097
rect 14328 -3473 14340 -3097
rect 14282 -3485 14340 -3473
rect 14400 -3097 14536 -3085
rect 14400 -3473 14412 -3097
rect 14446 -3273 14490 -3097
rect 14524 -3273 14536 -3097
rect 14446 -3285 14536 -3273
rect 14596 -3097 14654 -3085
rect 14596 -3273 14608 -3097
rect 14642 -3273 14654 -3097
rect 14596 -3285 14654 -3273
rect 16880 -3097 16938 -3085
rect 16880 -3273 16892 -3097
rect 16926 -3273 16938 -3097
rect 16880 -3285 16938 -3273
rect 16998 -3097 17130 -3085
rect 16998 -3273 17010 -3097
rect 17044 -3273 17084 -3097
rect 16998 -3285 17084 -3273
rect 14446 -3473 14458 -3285
rect 14400 -3485 14458 -3473
rect 17072 -3473 17084 -3285
rect 17118 -3473 17130 -3097
rect 17072 -3485 17130 -3473
rect 17190 -3097 17248 -3085
rect 17190 -3473 17202 -3097
rect 17236 -3473 17248 -3097
rect 17190 -3485 17248 -3473
rect 17308 -3097 17366 -3085
rect 17308 -3473 17320 -3097
rect 17354 -3473 17366 -3097
rect 17308 -3485 17366 -3473
rect 17426 -3097 17484 -3085
rect 17426 -3473 17438 -3097
rect 17472 -3473 17484 -3097
rect 17426 -3485 17484 -3473
rect 17544 -3097 17680 -3085
rect 17544 -3473 17556 -3097
rect 17590 -3273 17634 -3097
rect 17668 -3273 17680 -3097
rect 17590 -3285 17680 -3273
rect 17740 -3097 17798 -3085
rect 17740 -3273 17752 -3097
rect 17786 -3273 17798 -3097
rect 17740 -3285 17798 -3273
rect 20012 -3093 20070 -3081
rect 20012 -3269 20024 -3093
rect 20058 -3269 20070 -3093
rect 20012 -3281 20070 -3269
rect 20130 -3093 20262 -3081
rect 20130 -3269 20142 -3093
rect 20176 -3269 20216 -3093
rect 20130 -3281 20216 -3269
rect 17590 -3473 17602 -3285
rect 17544 -3485 17602 -3473
rect 20204 -3469 20216 -3281
rect 20250 -3469 20262 -3093
rect 20204 -3481 20262 -3469
rect 20322 -3093 20380 -3081
rect 20322 -3469 20334 -3093
rect 20368 -3469 20380 -3093
rect 20322 -3481 20380 -3469
rect 20440 -3093 20498 -3081
rect 20440 -3469 20452 -3093
rect 20486 -3469 20498 -3093
rect 20440 -3481 20498 -3469
rect 20558 -3093 20616 -3081
rect 20558 -3469 20570 -3093
rect 20604 -3469 20616 -3093
rect 20558 -3481 20616 -3469
rect 20676 -3093 20812 -3081
rect 20676 -3469 20688 -3093
rect 20722 -3269 20766 -3093
rect 20800 -3269 20812 -3093
rect 20722 -3281 20812 -3269
rect 20872 -3093 20930 -3081
rect 20872 -3269 20884 -3093
rect 20918 -3269 20930 -3093
rect 20872 -3281 20930 -3269
rect 23156 -3093 23214 -3081
rect 23156 -3269 23168 -3093
rect 23202 -3269 23214 -3093
rect 23156 -3281 23214 -3269
rect 23274 -3093 23406 -3081
rect 23274 -3269 23286 -3093
rect 23320 -3269 23360 -3093
rect 23274 -3281 23360 -3269
rect 20722 -3469 20734 -3281
rect 20676 -3481 20734 -3469
rect 23348 -3469 23360 -3281
rect 23394 -3469 23406 -3093
rect 23348 -3481 23406 -3469
rect 23466 -3093 23524 -3081
rect 23466 -3469 23478 -3093
rect 23512 -3469 23524 -3093
rect 23466 -3481 23524 -3469
rect 23584 -3093 23642 -3081
rect 23584 -3469 23596 -3093
rect 23630 -3469 23642 -3093
rect 23584 -3481 23642 -3469
rect 23702 -3093 23760 -3081
rect 23702 -3469 23714 -3093
rect 23748 -3469 23760 -3093
rect 23702 -3481 23760 -3469
rect 23820 -3093 23956 -3081
rect 23820 -3469 23832 -3093
rect 23866 -3269 23910 -3093
rect 23944 -3269 23956 -3093
rect 23866 -3281 23956 -3269
rect 24016 -3093 24074 -3081
rect 24016 -3269 24028 -3093
rect 24062 -3269 24074 -3093
rect 24016 -3281 24074 -3269
rect 23866 -3469 23878 -3281
rect 23820 -3481 23878 -3469
<< pdiff >>
rect 41913 24593 41971 24605
rect 39588 24521 39646 24533
rect 39588 24345 39600 24521
rect 39634 24345 39646 24521
rect 39588 24333 39646 24345
rect 39706 24521 39764 24533
rect 39706 24345 39718 24521
rect 39752 24345 39764 24521
rect 39706 24333 39764 24345
rect 39824 24521 39882 24533
rect 39824 24345 39836 24521
rect 39870 24345 39882 24521
rect 39824 24333 39882 24345
rect 39942 24521 40000 24533
rect 39942 24345 39954 24521
rect 39988 24345 40000 24521
rect 39942 24333 40000 24345
rect 40060 24521 40118 24533
rect 40060 24345 40072 24521
rect 40106 24345 40118 24521
rect 40060 24333 40118 24345
rect 40178 24521 40236 24533
rect 40178 24345 40190 24521
rect 40224 24345 40236 24521
rect 40178 24333 40236 24345
rect 40296 24521 40354 24533
rect 40296 24345 40308 24521
rect 40342 24345 40354 24521
rect 40296 24333 40354 24345
rect 40414 24521 40472 24533
rect 40414 24345 40426 24521
rect 40460 24345 40472 24521
rect 40414 24333 40472 24345
rect 40532 24521 40590 24533
rect 40532 24345 40544 24521
rect 40578 24345 40590 24521
rect 40532 24333 40590 24345
rect 40650 24521 40708 24533
rect 40650 24345 40662 24521
rect 40696 24345 40708 24521
rect 40650 24333 40708 24345
rect 41913 24217 41925 24593
rect 41959 24217 41971 24593
rect 41913 24205 41971 24217
rect 42031 24593 42089 24605
rect 42031 24217 42043 24593
rect 42077 24217 42089 24593
rect 42031 24205 42089 24217
rect 42149 24593 42207 24605
rect 42149 24217 42161 24593
rect 42195 24217 42207 24593
rect 42149 24205 42207 24217
rect 42267 24593 42325 24605
rect 42267 24217 42279 24593
rect 42313 24217 42325 24593
rect 42267 24205 42325 24217
rect 42385 24593 42443 24605
rect 42385 24217 42397 24593
rect 42431 24217 42443 24593
rect 42385 24205 42443 24217
rect 42503 24593 42561 24605
rect 42503 24217 42515 24593
rect 42549 24217 42561 24593
rect 42503 24205 42561 24217
rect 42621 24593 42679 24605
rect 42621 24217 42633 24593
rect 42667 24217 42679 24593
rect 42621 24205 42679 24217
rect 43055 24597 43113 24609
rect 43055 24221 43067 24597
rect 43101 24221 43113 24597
rect 43055 24209 43113 24221
rect 43173 24597 43231 24609
rect 43173 24221 43185 24597
rect 43219 24221 43231 24597
rect 43173 24209 43231 24221
rect 43291 24597 43349 24609
rect 43291 24221 43303 24597
rect 43337 24221 43349 24597
rect 43291 24209 43349 24221
rect 43409 24597 43467 24609
rect 43409 24221 43421 24597
rect 43455 24221 43467 24597
rect 43409 24209 43467 24221
rect 43527 24597 43585 24609
rect 43527 24221 43539 24597
rect 43573 24221 43585 24597
rect 43527 24209 43585 24221
rect 43645 24597 43703 24609
rect 43645 24221 43657 24597
rect 43691 24221 43703 24597
rect 43645 24209 43703 24221
rect 43763 24597 43821 24609
rect 43763 24221 43775 24597
rect 43809 24221 43821 24597
rect 48426 24590 48484 24602
rect 46101 24518 46159 24530
rect 46101 24342 46113 24518
rect 46147 24342 46159 24518
rect 46101 24330 46159 24342
rect 46219 24518 46277 24530
rect 46219 24342 46231 24518
rect 46265 24342 46277 24518
rect 46219 24330 46277 24342
rect 46337 24518 46395 24530
rect 46337 24342 46349 24518
rect 46383 24342 46395 24518
rect 46337 24330 46395 24342
rect 46455 24518 46513 24530
rect 46455 24342 46467 24518
rect 46501 24342 46513 24518
rect 46455 24330 46513 24342
rect 46573 24518 46631 24530
rect 46573 24342 46585 24518
rect 46619 24342 46631 24518
rect 46573 24330 46631 24342
rect 46691 24518 46749 24530
rect 46691 24342 46703 24518
rect 46737 24342 46749 24518
rect 46691 24330 46749 24342
rect 46809 24518 46867 24530
rect 46809 24342 46821 24518
rect 46855 24342 46867 24518
rect 46809 24330 46867 24342
rect 46927 24518 46985 24530
rect 46927 24342 46939 24518
rect 46973 24342 46985 24518
rect 46927 24330 46985 24342
rect 47045 24518 47103 24530
rect 47045 24342 47057 24518
rect 47091 24342 47103 24518
rect 47045 24330 47103 24342
rect 47163 24518 47221 24530
rect 47163 24342 47175 24518
rect 47209 24342 47221 24518
rect 47163 24330 47221 24342
rect 43763 24209 43821 24221
rect 48426 24214 48438 24590
rect 48472 24214 48484 24590
rect 48426 24202 48484 24214
rect 48544 24590 48602 24602
rect 48544 24214 48556 24590
rect 48590 24214 48602 24590
rect 48544 24202 48602 24214
rect 48662 24590 48720 24602
rect 48662 24214 48674 24590
rect 48708 24214 48720 24590
rect 48662 24202 48720 24214
rect 48780 24590 48838 24602
rect 48780 24214 48792 24590
rect 48826 24214 48838 24590
rect 48780 24202 48838 24214
rect 48898 24590 48956 24602
rect 48898 24214 48910 24590
rect 48944 24214 48956 24590
rect 48898 24202 48956 24214
rect 49016 24590 49074 24602
rect 49016 24214 49028 24590
rect 49062 24214 49074 24590
rect 49016 24202 49074 24214
rect 49134 24590 49192 24602
rect 49134 24214 49146 24590
rect 49180 24214 49192 24590
rect 49134 24202 49192 24214
rect 49568 24594 49626 24606
rect 49568 24218 49580 24594
rect 49614 24218 49626 24594
rect 49568 24206 49626 24218
rect 49686 24594 49744 24606
rect 49686 24218 49698 24594
rect 49732 24218 49744 24594
rect 49686 24206 49744 24218
rect 49804 24594 49862 24606
rect 49804 24218 49816 24594
rect 49850 24218 49862 24594
rect 49804 24206 49862 24218
rect 49922 24594 49980 24606
rect 49922 24218 49934 24594
rect 49968 24218 49980 24594
rect 49922 24206 49980 24218
rect 50040 24594 50098 24606
rect 50040 24218 50052 24594
rect 50086 24218 50098 24594
rect 50040 24206 50098 24218
rect 50158 24594 50216 24606
rect 50158 24218 50170 24594
rect 50204 24218 50216 24594
rect 50158 24206 50216 24218
rect 50276 24594 50334 24606
rect 50276 24218 50288 24594
rect 50322 24218 50334 24594
rect 54960 24585 55018 24597
rect 52635 24513 52693 24525
rect 52635 24337 52647 24513
rect 52681 24337 52693 24513
rect 52635 24325 52693 24337
rect 52753 24513 52811 24525
rect 52753 24337 52765 24513
rect 52799 24337 52811 24513
rect 52753 24325 52811 24337
rect 52871 24513 52929 24525
rect 52871 24337 52883 24513
rect 52917 24337 52929 24513
rect 52871 24325 52929 24337
rect 52989 24513 53047 24525
rect 52989 24337 53001 24513
rect 53035 24337 53047 24513
rect 52989 24325 53047 24337
rect 53107 24513 53165 24525
rect 53107 24337 53119 24513
rect 53153 24337 53165 24513
rect 53107 24325 53165 24337
rect 53225 24513 53283 24525
rect 53225 24337 53237 24513
rect 53271 24337 53283 24513
rect 53225 24325 53283 24337
rect 53343 24513 53401 24525
rect 53343 24337 53355 24513
rect 53389 24337 53401 24513
rect 53343 24325 53401 24337
rect 53461 24513 53519 24525
rect 53461 24337 53473 24513
rect 53507 24337 53519 24513
rect 53461 24325 53519 24337
rect 53579 24513 53637 24525
rect 53579 24337 53591 24513
rect 53625 24337 53637 24513
rect 53579 24325 53637 24337
rect 53697 24513 53755 24525
rect 53697 24337 53709 24513
rect 53743 24337 53755 24513
rect 53697 24325 53755 24337
rect 50276 24206 50334 24218
rect 42342 23810 42400 23822
rect 42342 23634 42354 23810
rect 42388 23634 42400 23810
rect 42342 23622 42400 23634
rect 42460 23810 42518 23822
rect 42460 23634 42472 23810
rect 42506 23634 42518 23810
rect 42460 23622 42518 23634
rect 42578 23810 42636 23822
rect 42578 23634 42590 23810
rect 42624 23634 42636 23810
rect 42578 23622 42636 23634
rect 42696 23810 42754 23822
rect 42696 23634 42708 23810
rect 42742 23634 42754 23810
rect 42696 23622 42754 23634
rect 43484 23814 43542 23826
rect 43484 23638 43496 23814
rect 43530 23638 43542 23814
rect 43484 23626 43542 23638
rect 43602 23814 43660 23826
rect 43602 23638 43614 23814
rect 43648 23638 43660 23814
rect 43602 23626 43660 23638
rect 43720 23814 43778 23826
rect 43720 23638 43732 23814
rect 43766 23638 43778 23814
rect 43720 23626 43778 23638
rect 43838 23814 43896 23826
rect 43838 23638 43850 23814
rect 43884 23638 43896 23814
rect 54960 24209 54972 24585
rect 55006 24209 55018 24585
rect 54960 24197 55018 24209
rect 55078 24585 55136 24597
rect 55078 24209 55090 24585
rect 55124 24209 55136 24585
rect 55078 24197 55136 24209
rect 55196 24585 55254 24597
rect 55196 24209 55208 24585
rect 55242 24209 55254 24585
rect 55196 24197 55254 24209
rect 55314 24585 55372 24597
rect 55314 24209 55326 24585
rect 55360 24209 55372 24585
rect 55314 24197 55372 24209
rect 55432 24585 55490 24597
rect 55432 24209 55444 24585
rect 55478 24209 55490 24585
rect 55432 24197 55490 24209
rect 55550 24585 55608 24597
rect 55550 24209 55562 24585
rect 55596 24209 55608 24585
rect 55550 24197 55608 24209
rect 55668 24585 55726 24597
rect 55668 24209 55680 24585
rect 55714 24209 55726 24585
rect 55668 24197 55726 24209
rect 56102 24589 56160 24601
rect 56102 24213 56114 24589
rect 56148 24213 56160 24589
rect 56102 24201 56160 24213
rect 56220 24589 56278 24601
rect 56220 24213 56232 24589
rect 56266 24213 56278 24589
rect 56220 24201 56278 24213
rect 56338 24589 56396 24601
rect 56338 24213 56350 24589
rect 56384 24213 56396 24589
rect 56338 24201 56396 24213
rect 56456 24589 56514 24601
rect 56456 24213 56468 24589
rect 56502 24213 56514 24589
rect 56456 24201 56514 24213
rect 56574 24589 56632 24601
rect 56574 24213 56586 24589
rect 56620 24213 56632 24589
rect 56574 24201 56632 24213
rect 56692 24589 56750 24601
rect 56692 24213 56704 24589
rect 56738 24213 56750 24589
rect 56692 24201 56750 24213
rect 56810 24589 56868 24601
rect 56810 24213 56822 24589
rect 56856 24213 56868 24589
rect 61518 24589 61576 24601
rect 59193 24517 59251 24529
rect 59193 24341 59205 24517
rect 59239 24341 59251 24517
rect 59193 24329 59251 24341
rect 59311 24517 59369 24529
rect 59311 24341 59323 24517
rect 59357 24341 59369 24517
rect 59311 24329 59369 24341
rect 59429 24517 59487 24529
rect 59429 24341 59441 24517
rect 59475 24341 59487 24517
rect 59429 24329 59487 24341
rect 59547 24517 59605 24529
rect 59547 24341 59559 24517
rect 59593 24341 59605 24517
rect 59547 24329 59605 24341
rect 59665 24517 59723 24529
rect 59665 24341 59677 24517
rect 59711 24341 59723 24517
rect 59665 24329 59723 24341
rect 59783 24517 59841 24529
rect 59783 24341 59795 24517
rect 59829 24341 59841 24517
rect 59783 24329 59841 24341
rect 59901 24517 59959 24529
rect 59901 24341 59913 24517
rect 59947 24341 59959 24517
rect 59901 24329 59959 24341
rect 60019 24517 60077 24529
rect 60019 24341 60031 24517
rect 60065 24341 60077 24517
rect 60019 24329 60077 24341
rect 60137 24517 60195 24529
rect 60137 24341 60149 24517
rect 60183 24341 60195 24517
rect 60137 24329 60195 24341
rect 60255 24517 60313 24529
rect 60255 24341 60267 24517
rect 60301 24341 60313 24517
rect 60255 24329 60313 24341
rect 56810 24201 56868 24213
rect 43838 23626 43896 23638
rect 48855 23807 48913 23819
rect 48855 23631 48867 23807
rect 48901 23631 48913 23807
rect 48855 23619 48913 23631
rect 48973 23807 49031 23819
rect 48973 23631 48985 23807
rect 49019 23631 49031 23807
rect 48973 23619 49031 23631
rect 49091 23807 49149 23819
rect 49091 23631 49103 23807
rect 49137 23631 49149 23807
rect 49091 23619 49149 23631
rect 49209 23807 49267 23819
rect 49209 23631 49221 23807
rect 49255 23631 49267 23807
rect 49209 23619 49267 23631
rect 49997 23811 50055 23823
rect 49997 23635 50009 23811
rect 50043 23635 50055 23811
rect 49997 23623 50055 23635
rect 50115 23811 50173 23823
rect 50115 23635 50127 23811
rect 50161 23635 50173 23811
rect 50115 23623 50173 23635
rect 50233 23811 50291 23823
rect 50233 23635 50245 23811
rect 50279 23635 50291 23811
rect 50233 23623 50291 23635
rect 50351 23811 50409 23823
rect 50351 23635 50363 23811
rect 50397 23635 50409 23811
rect 61518 24213 61530 24589
rect 61564 24213 61576 24589
rect 61518 24201 61576 24213
rect 61636 24589 61694 24601
rect 61636 24213 61648 24589
rect 61682 24213 61694 24589
rect 61636 24201 61694 24213
rect 61754 24589 61812 24601
rect 61754 24213 61766 24589
rect 61800 24213 61812 24589
rect 61754 24201 61812 24213
rect 61872 24589 61930 24601
rect 61872 24213 61884 24589
rect 61918 24213 61930 24589
rect 61872 24201 61930 24213
rect 61990 24589 62048 24601
rect 61990 24213 62002 24589
rect 62036 24213 62048 24589
rect 61990 24201 62048 24213
rect 62108 24589 62166 24601
rect 62108 24213 62120 24589
rect 62154 24213 62166 24589
rect 62108 24201 62166 24213
rect 62226 24589 62284 24601
rect 62226 24213 62238 24589
rect 62272 24213 62284 24589
rect 62226 24201 62284 24213
rect 62660 24593 62718 24605
rect 62660 24217 62672 24593
rect 62706 24217 62718 24593
rect 62660 24205 62718 24217
rect 62778 24593 62836 24605
rect 62778 24217 62790 24593
rect 62824 24217 62836 24593
rect 62778 24205 62836 24217
rect 62896 24593 62954 24605
rect 62896 24217 62908 24593
rect 62942 24217 62954 24593
rect 62896 24205 62954 24217
rect 63014 24593 63072 24605
rect 63014 24217 63026 24593
rect 63060 24217 63072 24593
rect 63014 24205 63072 24217
rect 63132 24593 63190 24605
rect 63132 24217 63144 24593
rect 63178 24217 63190 24593
rect 63132 24205 63190 24217
rect 63250 24593 63308 24605
rect 63250 24217 63262 24593
rect 63296 24217 63308 24593
rect 63250 24205 63308 24217
rect 63368 24593 63426 24605
rect 63368 24217 63380 24593
rect 63414 24217 63426 24593
rect 63368 24205 63426 24217
rect 50351 23623 50409 23635
rect 55389 23802 55447 23814
rect 55389 23626 55401 23802
rect 55435 23626 55447 23802
rect 55389 23614 55447 23626
rect 55507 23802 55565 23814
rect 55507 23626 55519 23802
rect 55553 23626 55565 23802
rect 55507 23614 55565 23626
rect 55625 23802 55683 23814
rect 55625 23626 55637 23802
rect 55671 23626 55683 23802
rect 55625 23614 55683 23626
rect 55743 23802 55801 23814
rect 55743 23626 55755 23802
rect 55789 23626 55801 23802
rect 55743 23614 55801 23626
rect 56531 23806 56589 23818
rect 56531 23630 56543 23806
rect 56577 23630 56589 23806
rect 56531 23618 56589 23630
rect 56649 23806 56707 23818
rect 56649 23630 56661 23806
rect 56695 23630 56707 23806
rect 56649 23618 56707 23630
rect 56767 23806 56825 23818
rect 56767 23630 56779 23806
rect 56813 23630 56825 23806
rect 56767 23618 56825 23630
rect 56885 23806 56943 23818
rect 56885 23630 56897 23806
rect 56931 23630 56943 23806
rect 56885 23618 56943 23630
rect 61947 23806 62005 23818
rect 61947 23630 61959 23806
rect 61993 23630 62005 23806
rect 61947 23618 62005 23630
rect 62065 23806 62123 23818
rect 62065 23630 62077 23806
rect 62111 23630 62123 23806
rect 62065 23618 62123 23630
rect 62183 23806 62241 23818
rect 62183 23630 62195 23806
rect 62229 23630 62241 23806
rect 62183 23618 62241 23630
rect 62301 23806 62359 23818
rect 62301 23630 62313 23806
rect 62347 23630 62359 23806
rect 62301 23618 62359 23630
rect 63089 23810 63147 23822
rect 63089 23634 63101 23810
rect 63135 23634 63147 23810
rect 63089 23622 63147 23634
rect 63207 23810 63265 23822
rect 63207 23634 63219 23810
rect 63253 23634 63265 23810
rect 63207 23622 63265 23634
rect 63325 23810 63383 23822
rect 63325 23634 63337 23810
rect 63371 23634 63383 23810
rect 63325 23622 63383 23634
rect 63443 23810 63501 23822
rect 63443 23634 63455 23810
rect 63489 23634 63501 23810
rect 63443 23622 63501 23634
rect 39602 22871 39660 22883
rect 39602 22695 39614 22871
rect 39648 22695 39660 22871
rect 39602 22683 39660 22695
rect 39720 22871 39778 22883
rect 39720 22695 39732 22871
rect 39766 22695 39778 22871
rect 39720 22683 39778 22695
rect 39838 22871 39896 22883
rect 39838 22695 39850 22871
rect 39884 22695 39896 22871
rect 39838 22683 39896 22695
rect 39956 22871 40014 22883
rect 39956 22695 39968 22871
rect 40002 22695 40014 22871
rect 39956 22683 40014 22695
rect 40074 22871 40132 22883
rect 40074 22695 40086 22871
rect 40120 22695 40132 22871
rect 40074 22683 40132 22695
rect 40192 22871 40250 22883
rect 40192 22695 40204 22871
rect 40238 22695 40250 22871
rect 40192 22683 40250 22695
rect 40310 22871 40368 22883
rect 40310 22695 40322 22871
rect 40356 22695 40368 22871
rect 40310 22683 40368 22695
rect 40428 22871 40486 22883
rect 40428 22695 40440 22871
rect 40474 22695 40486 22871
rect 40428 22683 40486 22695
rect 40546 22871 40604 22883
rect 40546 22695 40558 22871
rect 40592 22695 40604 22871
rect 40546 22683 40604 22695
rect 40664 22871 40722 22883
rect 40664 22695 40676 22871
rect 40710 22695 40722 22871
rect 46115 22868 46173 22880
rect 40664 22683 40722 22695
rect 46115 22692 46127 22868
rect 46161 22692 46173 22868
rect 46115 22680 46173 22692
rect 46233 22868 46291 22880
rect 46233 22692 46245 22868
rect 46279 22692 46291 22868
rect 46233 22680 46291 22692
rect 46351 22868 46409 22880
rect 46351 22692 46363 22868
rect 46397 22692 46409 22868
rect 46351 22680 46409 22692
rect 46469 22868 46527 22880
rect 46469 22692 46481 22868
rect 46515 22692 46527 22868
rect 46469 22680 46527 22692
rect 46587 22868 46645 22880
rect 46587 22692 46599 22868
rect 46633 22692 46645 22868
rect 46587 22680 46645 22692
rect 46705 22868 46763 22880
rect 46705 22692 46717 22868
rect 46751 22692 46763 22868
rect 46705 22680 46763 22692
rect 46823 22868 46881 22880
rect 46823 22692 46835 22868
rect 46869 22692 46881 22868
rect 46823 22680 46881 22692
rect 46941 22868 46999 22880
rect 46941 22692 46953 22868
rect 46987 22692 46999 22868
rect 46941 22680 46999 22692
rect 47059 22868 47117 22880
rect 47059 22692 47071 22868
rect 47105 22692 47117 22868
rect 47059 22680 47117 22692
rect 47177 22868 47235 22880
rect 47177 22692 47189 22868
rect 47223 22692 47235 22868
rect 52649 22863 52707 22875
rect 47177 22680 47235 22692
rect 52649 22687 52661 22863
rect 52695 22687 52707 22863
rect 41550 22454 41608 22466
rect 3473 21984 3531 21996
rect 3000 21784 3058 21796
rect 3000 21608 3012 21784
rect 3046 21608 3058 21784
rect 3000 21596 3058 21608
rect 3118 21784 3176 21796
rect 3118 21608 3130 21784
rect 3164 21608 3176 21784
rect 3118 21596 3176 21608
rect 3236 21784 3294 21796
rect 3236 21608 3248 21784
rect 3282 21608 3294 21784
rect 3236 21596 3294 21608
rect 3354 21784 3412 21796
rect 3354 21608 3366 21784
rect 3400 21608 3412 21784
rect 3354 21596 3412 21608
rect 3473 21608 3485 21984
rect 3519 21608 3531 21984
rect 3473 21596 3531 21608
rect 3591 21984 3649 21996
rect 3591 21608 3603 21984
rect 3637 21608 3649 21984
rect 3591 21596 3649 21608
rect 3709 21984 3767 21996
rect 3709 21608 3721 21984
rect 3755 21608 3767 21984
rect 3709 21596 3767 21608
rect 3827 21984 3885 21996
rect 3827 21608 3839 21984
rect 3873 21608 3885 21984
rect 3827 21596 3885 21608
rect 3946 21984 4004 21996
rect 3946 21608 3958 21984
rect 3992 21608 4004 21984
rect 3946 21596 4004 21608
rect 4064 21984 4122 21996
rect 4064 21608 4076 21984
rect 4110 21608 4122 21984
rect 4064 21596 4122 21608
rect 4182 21984 4240 21996
rect 4182 21608 4194 21984
rect 4228 21608 4240 21984
rect 4182 21596 4240 21608
rect 4300 21984 4358 21996
rect 4300 21608 4312 21984
rect 4346 21608 4358 21984
rect 4300 21596 4358 21608
rect 4418 21984 4476 21996
rect 4418 21608 4430 21984
rect 4464 21608 4476 21984
rect 4418 21596 4476 21608
rect 4536 21984 4594 21996
rect 4536 21608 4548 21984
rect 4582 21608 4594 21984
rect 4536 21596 4594 21608
rect 4654 21984 4712 21996
rect 4654 21608 4666 21984
rect 4700 21608 4712 21984
rect 4654 21596 4712 21608
rect 4767 21984 4825 21996
rect 4767 21608 4779 21984
rect 4813 21608 4825 21984
rect 4767 21596 4825 21608
rect 4885 21984 4943 21996
rect 4885 21608 4897 21984
rect 4931 21608 4943 21984
rect 4885 21596 4943 21608
rect 5003 21984 5061 21996
rect 5003 21608 5015 21984
rect 5049 21608 5061 21984
rect 5003 21596 5061 21608
rect 5121 21984 5179 21996
rect 5121 21608 5133 21984
rect 5167 21796 5179 21984
rect 6617 21984 6675 21996
rect 5167 21784 5266 21796
rect 5167 21608 5220 21784
rect 5254 21608 5266 21784
rect 5121 21596 5266 21608
rect 5326 21784 5384 21796
rect 5326 21608 5338 21784
rect 5372 21608 5384 21784
rect 5326 21596 5384 21608
rect 5444 21784 5502 21796
rect 5444 21608 5456 21784
rect 5490 21608 5502 21784
rect 5444 21596 5502 21608
rect 5562 21784 5620 21796
rect 5562 21608 5574 21784
rect 5608 21608 5620 21784
rect 5562 21596 5620 21608
rect 6144 21784 6202 21796
rect 6144 21608 6156 21784
rect 6190 21608 6202 21784
rect 6144 21596 6202 21608
rect 6262 21784 6320 21796
rect 6262 21608 6274 21784
rect 6308 21608 6320 21784
rect 6262 21596 6320 21608
rect 6380 21784 6438 21796
rect 6380 21608 6392 21784
rect 6426 21608 6438 21784
rect 6380 21596 6438 21608
rect 6498 21784 6556 21796
rect 6498 21608 6510 21784
rect 6544 21608 6556 21784
rect 6498 21596 6556 21608
rect 6617 21608 6629 21984
rect 6663 21608 6675 21984
rect 6617 21596 6675 21608
rect 6735 21984 6793 21996
rect 6735 21608 6747 21984
rect 6781 21608 6793 21984
rect 6735 21596 6793 21608
rect 6853 21984 6911 21996
rect 6853 21608 6865 21984
rect 6899 21608 6911 21984
rect 6853 21596 6911 21608
rect 6971 21984 7029 21996
rect 6971 21608 6983 21984
rect 7017 21608 7029 21984
rect 6971 21596 7029 21608
rect 7090 21984 7148 21996
rect 7090 21608 7102 21984
rect 7136 21608 7148 21984
rect 7090 21596 7148 21608
rect 7208 21984 7266 21996
rect 7208 21608 7220 21984
rect 7254 21608 7266 21984
rect 7208 21596 7266 21608
rect 7326 21984 7384 21996
rect 7326 21608 7338 21984
rect 7372 21608 7384 21984
rect 7326 21596 7384 21608
rect 7444 21984 7502 21996
rect 7444 21608 7456 21984
rect 7490 21608 7502 21984
rect 7444 21596 7502 21608
rect 7562 21984 7620 21996
rect 7562 21608 7574 21984
rect 7608 21608 7620 21984
rect 7562 21596 7620 21608
rect 7680 21984 7738 21996
rect 7680 21608 7692 21984
rect 7726 21608 7738 21984
rect 7680 21596 7738 21608
rect 7798 21984 7856 21996
rect 7798 21608 7810 21984
rect 7844 21608 7856 21984
rect 7798 21596 7856 21608
rect 7911 21984 7969 21996
rect 7911 21608 7923 21984
rect 7957 21608 7969 21984
rect 7911 21596 7969 21608
rect 8029 21984 8087 21996
rect 8029 21608 8041 21984
rect 8075 21608 8087 21984
rect 8029 21596 8087 21608
rect 8147 21984 8205 21996
rect 8147 21608 8159 21984
rect 8193 21608 8205 21984
rect 8147 21596 8205 21608
rect 8265 21984 8323 21996
rect 41066 22254 41124 22266
rect 8265 21608 8277 21984
rect 8311 21796 8323 21984
rect 9749 21980 9807 21992
rect 8311 21784 8410 21796
rect 8311 21608 8364 21784
rect 8398 21608 8410 21784
rect 8265 21596 8410 21608
rect 8470 21784 8528 21796
rect 8470 21608 8482 21784
rect 8516 21608 8528 21784
rect 8470 21596 8528 21608
rect 8588 21784 8646 21796
rect 8588 21608 8600 21784
rect 8634 21608 8646 21784
rect 8588 21596 8646 21608
rect 8706 21784 8764 21796
rect 8706 21608 8718 21784
rect 8752 21608 8764 21784
rect 8706 21596 8764 21608
rect 9276 21780 9334 21792
rect 9276 21604 9288 21780
rect 9322 21604 9334 21780
rect 9276 21592 9334 21604
rect 9394 21780 9452 21792
rect 9394 21604 9406 21780
rect 9440 21604 9452 21780
rect 9394 21592 9452 21604
rect 9512 21780 9570 21792
rect 9512 21604 9524 21780
rect 9558 21604 9570 21780
rect 9512 21592 9570 21604
rect 9630 21780 9688 21792
rect 9630 21604 9642 21780
rect 9676 21604 9688 21780
rect 9630 21592 9688 21604
rect 9749 21604 9761 21980
rect 9795 21604 9807 21980
rect 9749 21592 9807 21604
rect 9867 21980 9925 21992
rect 9867 21604 9879 21980
rect 9913 21604 9925 21980
rect 9867 21592 9925 21604
rect 9985 21980 10043 21992
rect 9985 21604 9997 21980
rect 10031 21604 10043 21980
rect 9985 21592 10043 21604
rect 10103 21980 10161 21992
rect 10103 21604 10115 21980
rect 10149 21604 10161 21980
rect 10103 21592 10161 21604
rect 10222 21980 10280 21992
rect 10222 21604 10234 21980
rect 10268 21604 10280 21980
rect 10222 21592 10280 21604
rect 10340 21980 10398 21992
rect 10340 21604 10352 21980
rect 10386 21604 10398 21980
rect 10340 21592 10398 21604
rect 10458 21980 10516 21992
rect 10458 21604 10470 21980
rect 10504 21604 10516 21980
rect 10458 21592 10516 21604
rect 10576 21980 10634 21992
rect 10576 21604 10588 21980
rect 10622 21604 10634 21980
rect 10576 21592 10634 21604
rect 10694 21980 10752 21992
rect 10694 21604 10706 21980
rect 10740 21604 10752 21980
rect 10694 21592 10752 21604
rect 10812 21980 10870 21992
rect 10812 21604 10824 21980
rect 10858 21604 10870 21980
rect 10812 21592 10870 21604
rect 10930 21980 10988 21992
rect 10930 21604 10942 21980
rect 10976 21604 10988 21980
rect 10930 21592 10988 21604
rect 11043 21980 11101 21992
rect 11043 21604 11055 21980
rect 11089 21604 11101 21980
rect 11043 21592 11101 21604
rect 11161 21980 11219 21992
rect 11161 21604 11173 21980
rect 11207 21604 11219 21980
rect 11161 21592 11219 21604
rect 11279 21980 11337 21992
rect 11279 21604 11291 21980
rect 11325 21604 11337 21980
rect 11279 21592 11337 21604
rect 11397 21980 11455 21992
rect 11397 21604 11409 21980
rect 11443 21792 11455 21980
rect 12893 21980 12951 21992
rect 11443 21780 11542 21792
rect 11443 21604 11496 21780
rect 11530 21604 11542 21780
rect 11397 21592 11542 21604
rect 11602 21780 11660 21792
rect 11602 21604 11614 21780
rect 11648 21604 11660 21780
rect 11602 21592 11660 21604
rect 11720 21780 11778 21792
rect 11720 21604 11732 21780
rect 11766 21604 11778 21780
rect 11720 21592 11778 21604
rect 11838 21780 11896 21792
rect 11838 21604 11850 21780
rect 11884 21604 11896 21780
rect 11838 21592 11896 21604
rect 12420 21780 12478 21792
rect 12420 21604 12432 21780
rect 12466 21604 12478 21780
rect 12420 21592 12478 21604
rect 12538 21780 12596 21792
rect 12538 21604 12550 21780
rect 12584 21604 12596 21780
rect 12538 21592 12596 21604
rect 12656 21780 12714 21792
rect 12656 21604 12668 21780
rect 12702 21604 12714 21780
rect 12656 21592 12714 21604
rect 12774 21780 12832 21792
rect 12774 21604 12786 21780
rect 12820 21604 12832 21780
rect 12774 21592 12832 21604
rect 12893 21604 12905 21980
rect 12939 21604 12951 21980
rect 12893 21592 12951 21604
rect 13011 21980 13069 21992
rect 13011 21604 13023 21980
rect 13057 21604 13069 21980
rect 13011 21592 13069 21604
rect 13129 21980 13187 21992
rect 13129 21604 13141 21980
rect 13175 21604 13187 21980
rect 13129 21592 13187 21604
rect 13247 21980 13305 21992
rect 13247 21604 13259 21980
rect 13293 21604 13305 21980
rect 13247 21592 13305 21604
rect 13366 21980 13424 21992
rect 13366 21604 13378 21980
rect 13412 21604 13424 21980
rect 13366 21592 13424 21604
rect 13484 21980 13542 21992
rect 13484 21604 13496 21980
rect 13530 21604 13542 21980
rect 13484 21592 13542 21604
rect 13602 21980 13660 21992
rect 13602 21604 13614 21980
rect 13648 21604 13660 21980
rect 13602 21592 13660 21604
rect 13720 21980 13778 21992
rect 13720 21604 13732 21980
rect 13766 21604 13778 21980
rect 13720 21592 13778 21604
rect 13838 21980 13896 21992
rect 13838 21604 13850 21980
rect 13884 21604 13896 21980
rect 13838 21592 13896 21604
rect 13956 21980 14014 21992
rect 13956 21604 13968 21980
rect 14002 21604 14014 21980
rect 13956 21592 14014 21604
rect 14074 21980 14132 21992
rect 14074 21604 14086 21980
rect 14120 21604 14132 21980
rect 14074 21592 14132 21604
rect 14187 21980 14245 21992
rect 14187 21604 14199 21980
rect 14233 21604 14245 21980
rect 14187 21592 14245 21604
rect 14305 21980 14363 21992
rect 14305 21604 14317 21980
rect 14351 21604 14363 21980
rect 14305 21592 14363 21604
rect 14423 21980 14481 21992
rect 14423 21604 14435 21980
rect 14469 21604 14481 21980
rect 14423 21592 14481 21604
rect 14541 21980 14599 21992
rect 14541 21604 14553 21980
rect 14587 21792 14599 21980
rect 16095 21984 16153 21996
rect 14587 21780 14686 21792
rect 14587 21604 14640 21780
rect 14674 21604 14686 21780
rect 14541 21592 14686 21604
rect 14746 21780 14804 21792
rect 14746 21604 14758 21780
rect 14792 21604 14804 21780
rect 14746 21592 14804 21604
rect 14864 21780 14922 21792
rect 14864 21604 14876 21780
rect 14910 21604 14922 21780
rect 14864 21592 14922 21604
rect 14982 21780 15040 21792
rect 14982 21604 14994 21780
rect 15028 21604 15040 21780
rect 14982 21592 15040 21604
rect 15622 21784 15680 21796
rect 15622 21608 15634 21784
rect 15668 21608 15680 21784
rect 15622 21596 15680 21608
rect 15740 21784 15798 21796
rect 15740 21608 15752 21784
rect 15786 21608 15798 21784
rect 15740 21596 15798 21608
rect 15858 21784 15916 21796
rect 15858 21608 15870 21784
rect 15904 21608 15916 21784
rect 15858 21596 15916 21608
rect 15976 21784 16034 21796
rect 15976 21608 15988 21784
rect 16022 21608 16034 21784
rect 15976 21596 16034 21608
rect 16095 21608 16107 21984
rect 16141 21608 16153 21984
rect 16095 21596 16153 21608
rect 16213 21984 16271 21996
rect 16213 21608 16225 21984
rect 16259 21608 16271 21984
rect 16213 21596 16271 21608
rect 16331 21984 16389 21996
rect 16331 21608 16343 21984
rect 16377 21608 16389 21984
rect 16331 21596 16389 21608
rect 16449 21984 16507 21996
rect 16449 21608 16461 21984
rect 16495 21608 16507 21984
rect 16449 21596 16507 21608
rect 16568 21984 16626 21996
rect 16568 21608 16580 21984
rect 16614 21608 16626 21984
rect 16568 21596 16626 21608
rect 16686 21984 16744 21996
rect 16686 21608 16698 21984
rect 16732 21608 16744 21984
rect 16686 21596 16744 21608
rect 16804 21984 16862 21996
rect 16804 21608 16816 21984
rect 16850 21608 16862 21984
rect 16804 21596 16862 21608
rect 16922 21984 16980 21996
rect 16922 21608 16934 21984
rect 16968 21608 16980 21984
rect 16922 21596 16980 21608
rect 17040 21984 17098 21996
rect 17040 21608 17052 21984
rect 17086 21608 17098 21984
rect 17040 21596 17098 21608
rect 17158 21984 17216 21996
rect 17158 21608 17170 21984
rect 17204 21608 17216 21984
rect 17158 21596 17216 21608
rect 17276 21984 17334 21996
rect 17276 21608 17288 21984
rect 17322 21608 17334 21984
rect 17276 21596 17334 21608
rect 17389 21984 17447 21996
rect 17389 21608 17401 21984
rect 17435 21608 17447 21984
rect 17389 21596 17447 21608
rect 17507 21984 17565 21996
rect 17507 21608 17519 21984
rect 17553 21608 17565 21984
rect 17507 21596 17565 21608
rect 17625 21984 17683 21996
rect 17625 21608 17637 21984
rect 17671 21608 17683 21984
rect 17625 21596 17683 21608
rect 17743 21984 17801 21996
rect 17743 21608 17755 21984
rect 17789 21796 17801 21984
rect 19239 21984 19297 21996
rect 17789 21784 17888 21796
rect 17789 21608 17842 21784
rect 17876 21608 17888 21784
rect 17743 21596 17888 21608
rect 17948 21784 18006 21796
rect 17948 21608 17960 21784
rect 17994 21608 18006 21784
rect 17948 21596 18006 21608
rect 18066 21784 18124 21796
rect 18066 21608 18078 21784
rect 18112 21608 18124 21784
rect 18066 21596 18124 21608
rect 18184 21784 18242 21796
rect 18184 21608 18196 21784
rect 18230 21608 18242 21784
rect 18184 21596 18242 21608
rect 18766 21784 18824 21796
rect 18766 21608 18778 21784
rect 18812 21608 18824 21784
rect 18766 21596 18824 21608
rect 18884 21784 18942 21796
rect 18884 21608 18896 21784
rect 18930 21608 18942 21784
rect 18884 21596 18942 21608
rect 19002 21784 19060 21796
rect 19002 21608 19014 21784
rect 19048 21608 19060 21784
rect 19002 21596 19060 21608
rect 19120 21784 19178 21796
rect 19120 21608 19132 21784
rect 19166 21608 19178 21784
rect 19120 21596 19178 21608
rect 19239 21608 19251 21984
rect 19285 21608 19297 21984
rect 19239 21596 19297 21608
rect 19357 21984 19415 21996
rect 19357 21608 19369 21984
rect 19403 21608 19415 21984
rect 19357 21596 19415 21608
rect 19475 21984 19533 21996
rect 19475 21608 19487 21984
rect 19521 21608 19533 21984
rect 19475 21596 19533 21608
rect 19593 21984 19651 21996
rect 19593 21608 19605 21984
rect 19639 21608 19651 21984
rect 19593 21596 19651 21608
rect 19712 21984 19770 21996
rect 19712 21608 19724 21984
rect 19758 21608 19770 21984
rect 19712 21596 19770 21608
rect 19830 21984 19888 21996
rect 19830 21608 19842 21984
rect 19876 21608 19888 21984
rect 19830 21596 19888 21608
rect 19948 21984 20006 21996
rect 19948 21608 19960 21984
rect 19994 21608 20006 21984
rect 19948 21596 20006 21608
rect 20066 21984 20124 21996
rect 20066 21608 20078 21984
rect 20112 21608 20124 21984
rect 20066 21596 20124 21608
rect 20184 21984 20242 21996
rect 20184 21608 20196 21984
rect 20230 21608 20242 21984
rect 20184 21596 20242 21608
rect 20302 21984 20360 21996
rect 20302 21608 20314 21984
rect 20348 21608 20360 21984
rect 20302 21596 20360 21608
rect 20420 21984 20478 21996
rect 20420 21608 20432 21984
rect 20466 21608 20478 21984
rect 20420 21596 20478 21608
rect 20533 21984 20591 21996
rect 20533 21608 20545 21984
rect 20579 21608 20591 21984
rect 20533 21596 20591 21608
rect 20651 21984 20709 21996
rect 20651 21608 20663 21984
rect 20697 21608 20709 21984
rect 20651 21596 20709 21608
rect 20769 21984 20827 21996
rect 20769 21608 20781 21984
rect 20815 21608 20827 21984
rect 20769 21596 20827 21608
rect 20887 21984 20945 21996
rect 20887 21608 20899 21984
rect 20933 21796 20945 21984
rect 22371 21980 22429 21992
rect 20933 21784 21032 21796
rect 20933 21608 20986 21784
rect 21020 21608 21032 21784
rect 20887 21596 21032 21608
rect 21092 21784 21150 21796
rect 21092 21608 21104 21784
rect 21138 21608 21150 21784
rect 21092 21596 21150 21608
rect 21210 21784 21268 21796
rect 21210 21608 21222 21784
rect 21256 21608 21268 21784
rect 21210 21596 21268 21608
rect 21328 21784 21386 21796
rect 21328 21608 21340 21784
rect 21374 21608 21386 21784
rect 21328 21596 21386 21608
rect 21898 21780 21956 21792
rect 21898 21604 21910 21780
rect 21944 21604 21956 21780
rect 21898 21592 21956 21604
rect 22016 21780 22074 21792
rect 22016 21604 22028 21780
rect 22062 21604 22074 21780
rect 22016 21592 22074 21604
rect 22134 21780 22192 21792
rect 22134 21604 22146 21780
rect 22180 21604 22192 21780
rect 22134 21592 22192 21604
rect 22252 21780 22310 21792
rect 22252 21604 22264 21780
rect 22298 21604 22310 21780
rect 22252 21592 22310 21604
rect 22371 21604 22383 21980
rect 22417 21604 22429 21980
rect 22371 21592 22429 21604
rect 22489 21980 22547 21992
rect 22489 21604 22501 21980
rect 22535 21604 22547 21980
rect 22489 21592 22547 21604
rect 22607 21980 22665 21992
rect 22607 21604 22619 21980
rect 22653 21604 22665 21980
rect 22607 21592 22665 21604
rect 22725 21980 22783 21992
rect 22725 21604 22737 21980
rect 22771 21604 22783 21980
rect 22725 21592 22783 21604
rect 22844 21980 22902 21992
rect 22844 21604 22856 21980
rect 22890 21604 22902 21980
rect 22844 21592 22902 21604
rect 22962 21980 23020 21992
rect 22962 21604 22974 21980
rect 23008 21604 23020 21980
rect 22962 21592 23020 21604
rect 23080 21980 23138 21992
rect 23080 21604 23092 21980
rect 23126 21604 23138 21980
rect 23080 21592 23138 21604
rect 23198 21980 23256 21992
rect 23198 21604 23210 21980
rect 23244 21604 23256 21980
rect 23198 21592 23256 21604
rect 23316 21980 23374 21992
rect 23316 21604 23328 21980
rect 23362 21604 23374 21980
rect 23316 21592 23374 21604
rect 23434 21980 23492 21992
rect 23434 21604 23446 21980
rect 23480 21604 23492 21980
rect 23434 21592 23492 21604
rect 23552 21980 23610 21992
rect 23552 21604 23564 21980
rect 23598 21604 23610 21980
rect 23552 21592 23610 21604
rect 23665 21980 23723 21992
rect 23665 21604 23677 21980
rect 23711 21604 23723 21980
rect 23665 21592 23723 21604
rect 23783 21980 23841 21992
rect 23783 21604 23795 21980
rect 23829 21604 23841 21980
rect 23783 21592 23841 21604
rect 23901 21980 23959 21992
rect 23901 21604 23913 21980
rect 23947 21604 23959 21980
rect 23901 21592 23959 21604
rect 24019 21980 24077 21992
rect 24019 21604 24031 21980
rect 24065 21792 24077 21980
rect 25515 21980 25573 21992
rect 24065 21780 24164 21792
rect 24065 21604 24118 21780
rect 24152 21604 24164 21780
rect 24019 21592 24164 21604
rect 24224 21780 24282 21792
rect 24224 21604 24236 21780
rect 24270 21604 24282 21780
rect 24224 21592 24282 21604
rect 24342 21780 24400 21792
rect 24342 21604 24354 21780
rect 24388 21604 24400 21780
rect 24342 21592 24400 21604
rect 24460 21780 24518 21792
rect 24460 21604 24472 21780
rect 24506 21604 24518 21780
rect 24460 21592 24518 21604
rect 25042 21780 25100 21792
rect 25042 21604 25054 21780
rect 25088 21604 25100 21780
rect 25042 21592 25100 21604
rect 25160 21780 25218 21792
rect 25160 21604 25172 21780
rect 25206 21604 25218 21780
rect 25160 21592 25218 21604
rect 25278 21780 25336 21792
rect 25278 21604 25290 21780
rect 25324 21604 25336 21780
rect 25278 21592 25336 21604
rect 25396 21780 25454 21792
rect 25396 21604 25408 21780
rect 25442 21604 25454 21780
rect 25396 21592 25454 21604
rect 25515 21604 25527 21980
rect 25561 21604 25573 21980
rect 25515 21592 25573 21604
rect 25633 21980 25691 21992
rect 25633 21604 25645 21980
rect 25679 21604 25691 21980
rect 25633 21592 25691 21604
rect 25751 21980 25809 21992
rect 25751 21604 25763 21980
rect 25797 21604 25809 21980
rect 25751 21592 25809 21604
rect 25869 21980 25927 21992
rect 25869 21604 25881 21980
rect 25915 21604 25927 21980
rect 25869 21592 25927 21604
rect 25988 21980 26046 21992
rect 25988 21604 26000 21980
rect 26034 21604 26046 21980
rect 25988 21592 26046 21604
rect 26106 21980 26164 21992
rect 26106 21604 26118 21980
rect 26152 21604 26164 21980
rect 26106 21592 26164 21604
rect 26224 21980 26282 21992
rect 26224 21604 26236 21980
rect 26270 21604 26282 21980
rect 26224 21592 26282 21604
rect 26342 21980 26400 21992
rect 26342 21604 26354 21980
rect 26388 21604 26400 21980
rect 26342 21592 26400 21604
rect 26460 21980 26518 21992
rect 26460 21604 26472 21980
rect 26506 21604 26518 21980
rect 26460 21592 26518 21604
rect 26578 21980 26636 21992
rect 26578 21604 26590 21980
rect 26624 21604 26636 21980
rect 26578 21592 26636 21604
rect 26696 21980 26754 21992
rect 26696 21604 26708 21980
rect 26742 21604 26754 21980
rect 26696 21592 26754 21604
rect 26809 21980 26867 21992
rect 26809 21604 26821 21980
rect 26855 21604 26867 21980
rect 26809 21592 26867 21604
rect 26927 21980 26985 21992
rect 26927 21604 26939 21980
rect 26973 21604 26985 21980
rect 26927 21592 26985 21604
rect 27045 21980 27103 21992
rect 27045 21604 27057 21980
rect 27091 21604 27103 21980
rect 27045 21592 27103 21604
rect 27163 21980 27221 21992
rect 27163 21604 27175 21980
rect 27209 21792 27221 21980
rect 41066 22078 41078 22254
rect 41112 22078 41124 22254
rect 41066 22066 41124 22078
rect 41184 22254 41242 22266
rect 41184 22078 41196 22254
rect 41230 22078 41242 22254
rect 41184 22066 41242 22078
rect 41302 22254 41360 22266
rect 41302 22078 41314 22254
rect 41348 22078 41360 22254
rect 41302 22066 41360 22078
rect 41420 22254 41478 22266
rect 41420 22078 41432 22254
rect 41466 22078 41478 22254
rect 41420 22066 41478 22078
rect 41550 22078 41562 22454
rect 41596 22078 41608 22454
rect 41550 22066 41608 22078
rect 41668 22454 41726 22466
rect 41668 22078 41680 22454
rect 41714 22078 41726 22454
rect 41668 22066 41726 22078
rect 41786 22454 41844 22466
rect 41786 22078 41798 22454
rect 41832 22078 41844 22454
rect 41786 22066 41844 22078
rect 41904 22454 41962 22466
rect 41904 22078 41916 22454
rect 41950 22078 41962 22454
rect 41904 22066 41962 22078
rect 42022 22454 42080 22466
rect 42022 22078 42034 22454
rect 42068 22078 42080 22454
rect 42022 22066 42080 22078
rect 42140 22454 42198 22466
rect 42140 22078 42152 22454
rect 42186 22078 42198 22454
rect 42140 22066 42198 22078
rect 42258 22454 42316 22466
rect 42258 22078 42270 22454
rect 42304 22078 42316 22454
rect 43448 22454 43506 22466
rect 42258 22066 42316 22078
rect 42387 22254 42445 22266
rect 42387 22078 42399 22254
rect 42433 22078 42445 22254
rect 42387 22066 42445 22078
rect 42505 22254 42563 22266
rect 42505 22078 42517 22254
rect 42551 22078 42563 22254
rect 42505 22066 42563 22078
rect 42623 22254 42681 22266
rect 42623 22078 42635 22254
rect 42669 22078 42681 22254
rect 42623 22066 42681 22078
rect 42741 22254 42799 22266
rect 42741 22078 42753 22254
rect 42787 22078 42799 22254
rect 42741 22066 42799 22078
rect 42964 22254 43022 22266
rect 42964 22078 42976 22254
rect 43010 22078 43022 22254
rect 42964 22066 43022 22078
rect 43082 22254 43140 22266
rect 43082 22078 43094 22254
rect 43128 22078 43140 22254
rect 43082 22066 43140 22078
rect 43200 22254 43258 22266
rect 43200 22078 43212 22254
rect 43246 22078 43258 22254
rect 43200 22066 43258 22078
rect 43318 22254 43376 22266
rect 43318 22078 43330 22254
rect 43364 22078 43376 22254
rect 43318 22066 43376 22078
rect 43448 22078 43460 22454
rect 43494 22078 43506 22454
rect 43448 22066 43506 22078
rect 43566 22454 43624 22466
rect 43566 22078 43578 22454
rect 43612 22078 43624 22454
rect 43566 22066 43624 22078
rect 43684 22454 43742 22466
rect 43684 22078 43696 22454
rect 43730 22078 43742 22454
rect 43684 22066 43742 22078
rect 43802 22454 43860 22466
rect 43802 22078 43814 22454
rect 43848 22078 43860 22454
rect 43802 22066 43860 22078
rect 43920 22454 43978 22466
rect 43920 22078 43932 22454
rect 43966 22078 43978 22454
rect 43920 22066 43978 22078
rect 44038 22454 44096 22466
rect 44038 22078 44050 22454
rect 44084 22078 44096 22454
rect 44038 22066 44096 22078
rect 44156 22454 44214 22466
rect 44156 22078 44168 22454
rect 44202 22078 44214 22454
rect 52649 22675 52707 22687
rect 52767 22863 52825 22875
rect 52767 22687 52779 22863
rect 52813 22687 52825 22863
rect 52767 22675 52825 22687
rect 52885 22863 52943 22875
rect 52885 22687 52897 22863
rect 52931 22687 52943 22863
rect 52885 22675 52943 22687
rect 53003 22863 53061 22875
rect 53003 22687 53015 22863
rect 53049 22687 53061 22863
rect 53003 22675 53061 22687
rect 53121 22863 53179 22875
rect 53121 22687 53133 22863
rect 53167 22687 53179 22863
rect 53121 22675 53179 22687
rect 53239 22863 53297 22875
rect 53239 22687 53251 22863
rect 53285 22687 53297 22863
rect 53239 22675 53297 22687
rect 53357 22863 53415 22875
rect 53357 22687 53369 22863
rect 53403 22687 53415 22863
rect 53357 22675 53415 22687
rect 53475 22863 53533 22875
rect 53475 22687 53487 22863
rect 53521 22687 53533 22863
rect 53475 22675 53533 22687
rect 53593 22863 53651 22875
rect 53593 22687 53605 22863
rect 53639 22687 53651 22863
rect 53593 22675 53651 22687
rect 53711 22863 53769 22875
rect 53711 22687 53723 22863
rect 53757 22687 53769 22863
rect 59207 22867 59265 22879
rect 53711 22675 53769 22687
rect 59207 22691 59219 22867
rect 59253 22691 59265 22867
rect 59207 22679 59265 22691
rect 59325 22867 59383 22879
rect 59325 22691 59337 22867
rect 59371 22691 59383 22867
rect 59325 22679 59383 22691
rect 59443 22867 59501 22879
rect 59443 22691 59455 22867
rect 59489 22691 59501 22867
rect 59443 22679 59501 22691
rect 59561 22867 59619 22879
rect 59561 22691 59573 22867
rect 59607 22691 59619 22867
rect 59561 22679 59619 22691
rect 59679 22867 59737 22879
rect 59679 22691 59691 22867
rect 59725 22691 59737 22867
rect 59679 22679 59737 22691
rect 59797 22867 59855 22879
rect 59797 22691 59809 22867
rect 59843 22691 59855 22867
rect 59797 22679 59855 22691
rect 59915 22867 59973 22879
rect 59915 22691 59927 22867
rect 59961 22691 59973 22867
rect 59915 22679 59973 22691
rect 60033 22867 60091 22879
rect 60033 22691 60045 22867
rect 60079 22691 60091 22867
rect 60033 22679 60091 22691
rect 60151 22867 60209 22879
rect 60151 22691 60163 22867
rect 60197 22691 60209 22867
rect 60151 22679 60209 22691
rect 60269 22867 60327 22879
rect 60269 22691 60281 22867
rect 60315 22691 60327 22867
rect 60269 22679 60327 22691
rect 48063 22451 48121 22463
rect 44156 22066 44214 22078
rect 44285 22254 44343 22266
rect 44285 22078 44297 22254
rect 44331 22078 44343 22254
rect 44285 22066 44343 22078
rect 44403 22254 44461 22266
rect 44403 22078 44415 22254
rect 44449 22078 44461 22254
rect 44403 22066 44461 22078
rect 44521 22254 44579 22266
rect 44521 22078 44533 22254
rect 44567 22078 44579 22254
rect 44521 22066 44579 22078
rect 44639 22254 44697 22266
rect 44639 22078 44651 22254
rect 44685 22078 44697 22254
rect 44639 22066 44697 22078
rect 27209 21780 27308 21792
rect 27209 21604 27262 21780
rect 27296 21604 27308 21780
rect 27163 21592 27308 21604
rect 27368 21780 27426 21792
rect 27368 21604 27380 21780
rect 27414 21604 27426 21780
rect 27368 21592 27426 21604
rect 27486 21780 27544 21792
rect 27486 21604 27498 21780
rect 27532 21604 27544 21780
rect 27486 21592 27544 21604
rect 27604 21780 27662 21792
rect 27604 21604 27616 21780
rect 27650 21604 27662 21780
rect 27604 21592 27662 21604
rect 39597 21267 39655 21279
rect 39597 21091 39609 21267
rect 39643 21091 39655 21267
rect 39597 21079 39655 21091
rect 39715 21267 39773 21279
rect 39715 21091 39727 21267
rect 39761 21091 39773 21267
rect 39715 21079 39773 21091
rect 39833 21267 39891 21279
rect 39833 21091 39845 21267
rect 39879 21091 39891 21267
rect 39833 21079 39891 21091
rect 39951 21267 40009 21279
rect 39951 21091 39963 21267
rect 39997 21091 40009 21267
rect 39951 21079 40009 21091
rect 40069 21267 40127 21279
rect 40069 21091 40081 21267
rect 40115 21091 40127 21267
rect 40069 21079 40127 21091
rect 40187 21267 40245 21279
rect 40187 21091 40199 21267
rect 40233 21091 40245 21267
rect 40187 21079 40245 21091
rect 40305 21267 40363 21279
rect 40305 21091 40317 21267
rect 40351 21091 40363 21267
rect 40305 21079 40363 21091
rect 40423 21267 40481 21279
rect 40423 21091 40435 21267
rect 40469 21091 40481 21267
rect 40423 21079 40481 21091
rect 40541 21267 40599 21279
rect 40541 21091 40553 21267
rect 40587 21091 40599 21267
rect 40541 21079 40599 21091
rect 40659 21267 40717 21279
rect 40659 21091 40671 21267
rect 40705 21091 40717 21267
rect 40659 21079 40717 21091
rect 41493 21761 41551 21773
rect 41493 21385 41505 21761
rect 41539 21385 41551 21761
rect 41493 21373 41551 21385
rect 41611 21761 41669 21773
rect 41611 21385 41623 21761
rect 41657 21385 41669 21761
rect 41611 21373 41669 21385
rect 41729 21761 41787 21773
rect 41729 21385 41741 21761
rect 41775 21385 41787 21761
rect 41729 21373 41787 21385
rect 41847 21761 41905 21773
rect 41847 21385 41859 21761
rect 41893 21385 41905 21761
rect 41847 21373 41905 21385
rect 41965 21761 42023 21773
rect 41965 21385 41977 21761
rect 42011 21385 42023 21761
rect 41965 21373 42023 21385
rect 42083 21761 42141 21773
rect 42083 21385 42095 21761
rect 42129 21385 42141 21761
rect 42083 21373 42141 21385
rect 42201 21761 42259 21773
rect 42201 21385 42213 21761
rect 42247 21385 42259 21761
rect 42201 21373 42259 21385
rect 47579 22251 47637 22263
rect 47579 22075 47591 22251
rect 47625 22075 47637 22251
rect 47579 22063 47637 22075
rect 47697 22251 47755 22263
rect 47697 22075 47709 22251
rect 47743 22075 47755 22251
rect 47697 22063 47755 22075
rect 47815 22251 47873 22263
rect 47815 22075 47827 22251
rect 47861 22075 47873 22251
rect 47815 22063 47873 22075
rect 47933 22251 47991 22263
rect 47933 22075 47945 22251
rect 47979 22075 47991 22251
rect 47933 22063 47991 22075
rect 48063 22075 48075 22451
rect 48109 22075 48121 22451
rect 48063 22063 48121 22075
rect 48181 22451 48239 22463
rect 48181 22075 48193 22451
rect 48227 22075 48239 22451
rect 48181 22063 48239 22075
rect 48299 22451 48357 22463
rect 48299 22075 48311 22451
rect 48345 22075 48357 22451
rect 48299 22063 48357 22075
rect 48417 22451 48475 22463
rect 48417 22075 48429 22451
rect 48463 22075 48475 22451
rect 48417 22063 48475 22075
rect 48535 22451 48593 22463
rect 48535 22075 48547 22451
rect 48581 22075 48593 22451
rect 48535 22063 48593 22075
rect 48653 22451 48711 22463
rect 48653 22075 48665 22451
rect 48699 22075 48711 22451
rect 48653 22063 48711 22075
rect 48771 22451 48829 22463
rect 48771 22075 48783 22451
rect 48817 22075 48829 22451
rect 49961 22451 50019 22463
rect 48771 22063 48829 22075
rect 48900 22251 48958 22263
rect 48900 22075 48912 22251
rect 48946 22075 48958 22251
rect 48900 22063 48958 22075
rect 49018 22251 49076 22263
rect 49018 22075 49030 22251
rect 49064 22075 49076 22251
rect 49018 22063 49076 22075
rect 49136 22251 49194 22263
rect 49136 22075 49148 22251
rect 49182 22075 49194 22251
rect 49136 22063 49194 22075
rect 49254 22251 49312 22263
rect 49254 22075 49266 22251
rect 49300 22075 49312 22251
rect 49254 22063 49312 22075
rect 49477 22251 49535 22263
rect 49477 22075 49489 22251
rect 49523 22075 49535 22251
rect 49477 22063 49535 22075
rect 49595 22251 49653 22263
rect 49595 22075 49607 22251
rect 49641 22075 49653 22251
rect 49595 22063 49653 22075
rect 49713 22251 49771 22263
rect 49713 22075 49725 22251
rect 49759 22075 49771 22251
rect 49713 22063 49771 22075
rect 49831 22251 49889 22263
rect 49831 22075 49843 22251
rect 49877 22075 49889 22251
rect 49831 22063 49889 22075
rect 49961 22075 49973 22451
rect 50007 22075 50019 22451
rect 49961 22063 50019 22075
rect 50079 22451 50137 22463
rect 50079 22075 50091 22451
rect 50125 22075 50137 22451
rect 50079 22063 50137 22075
rect 50197 22451 50255 22463
rect 50197 22075 50209 22451
rect 50243 22075 50255 22451
rect 50197 22063 50255 22075
rect 50315 22451 50373 22463
rect 50315 22075 50327 22451
rect 50361 22075 50373 22451
rect 50315 22063 50373 22075
rect 50433 22451 50491 22463
rect 50433 22075 50445 22451
rect 50479 22075 50491 22451
rect 50433 22063 50491 22075
rect 50551 22451 50609 22463
rect 50551 22075 50563 22451
rect 50597 22075 50609 22451
rect 50551 22063 50609 22075
rect 50669 22451 50727 22463
rect 50669 22075 50681 22451
rect 50715 22075 50727 22451
rect 54597 22446 54655 22458
rect 50669 22063 50727 22075
rect 50798 22251 50856 22263
rect 50798 22075 50810 22251
rect 50844 22075 50856 22251
rect 50798 22063 50856 22075
rect 50916 22251 50974 22263
rect 50916 22075 50928 22251
rect 50962 22075 50974 22251
rect 50916 22063 50974 22075
rect 51034 22251 51092 22263
rect 51034 22075 51046 22251
rect 51080 22075 51092 22251
rect 51034 22063 51092 22075
rect 51152 22251 51210 22263
rect 51152 22075 51164 22251
rect 51198 22075 51210 22251
rect 51152 22063 51210 22075
rect 43391 21761 43449 21773
rect 43391 21385 43403 21761
rect 43437 21385 43449 21761
rect 43391 21373 43449 21385
rect 43509 21761 43567 21773
rect 43509 21385 43521 21761
rect 43555 21385 43567 21761
rect 43509 21373 43567 21385
rect 43627 21761 43685 21773
rect 43627 21385 43639 21761
rect 43673 21385 43685 21761
rect 43627 21373 43685 21385
rect 43745 21761 43803 21773
rect 43745 21385 43757 21761
rect 43791 21385 43803 21761
rect 43745 21373 43803 21385
rect 43863 21761 43921 21773
rect 43863 21385 43875 21761
rect 43909 21385 43921 21761
rect 43863 21373 43921 21385
rect 43981 21761 44039 21773
rect 43981 21385 43993 21761
rect 44027 21385 44039 21761
rect 43981 21373 44039 21385
rect 44099 21761 44157 21773
rect 44099 21385 44111 21761
rect 44145 21385 44157 21761
rect 44099 21373 44157 21385
rect 46110 21264 46168 21276
rect 46110 21088 46122 21264
rect 46156 21088 46168 21264
rect 46110 21076 46168 21088
rect 46228 21264 46286 21276
rect 46228 21088 46240 21264
rect 46274 21088 46286 21264
rect 46228 21076 46286 21088
rect 46346 21264 46404 21276
rect 46346 21088 46358 21264
rect 46392 21088 46404 21264
rect 46346 21076 46404 21088
rect 46464 21264 46522 21276
rect 46464 21088 46476 21264
rect 46510 21088 46522 21264
rect 46464 21076 46522 21088
rect 46582 21264 46640 21276
rect 46582 21088 46594 21264
rect 46628 21088 46640 21264
rect 46582 21076 46640 21088
rect 46700 21264 46758 21276
rect 46700 21088 46712 21264
rect 46746 21088 46758 21264
rect 46700 21076 46758 21088
rect 46818 21264 46876 21276
rect 46818 21088 46830 21264
rect 46864 21088 46876 21264
rect 46818 21076 46876 21088
rect 46936 21264 46994 21276
rect 46936 21088 46948 21264
rect 46982 21088 46994 21264
rect 46936 21076 46994 21088
rect 47054 21264 47112 21276
rect 47054 21088 47066 21264
rect 47100 21088 47112 21264
rect 47054 21076 47112 21088
rect 47172 21264 47230 21276
rect 47172 21088 47184 21264
rect 47218 21088 47230 21264
rect 47172 21076 47230 21088
rect 48006 21758 48064 21770
rect 48006 21382 48018 21758
rect 48052 21382 48064 21758
rect 48006 21370 48064 21382
rect 48124 21758 48182 21770
rect 48124 21382 48136 21758
rect 48170 21382 48182 21758
rect 48124 21370 48182 21382
rect 48242 21758 48300 21770
rect 48242 21382 48254 21758
rect 48288 21382 48300 21758
rect 48242 21370 48300 21382
rect 48360 21758 48418 21770
rect 48360 21382 48372 21758
rect 48406 21382 48418 21758
rect 48360 21370 48418 21382
rect 48478 21758 48536 21770
rect 48478 21382 48490 21758
rect 48524 21382 48536 21758
rect 48478 21370 48536 21382
rect 48596 21758 48654 21770
rect 48596 21382 48608 21758
rect 48642 21382 48654 21758
rect 48596 21370 48654 21382
rect 48714 21758 48772 21770
rect 48714 21382 48726 21758
rect 48760 21382 48772 21758
rect 48714 21370 48772 21382
rect 54113 22246 54171 22258
rect 54113 22070 54125 22246
rect 54159 22070 54171 22246
rect 54113 22058 54171 22070
rect 54231 22246 54289 22258
rect 54231 22070 54243 22246
rect 54277 22070 54289 22246
rect 54231 22058 54289 22070
rect 54349 22246 54407 22258
rect 54349 22070 54361 22246
rect 54395 22070 54407 22246
rect 54349 22058 54407 22070
rect 54467 22246 54525 22258
rect 54467 22070 54479 22246
rect 54513 22070 54525 22246
rect 54467 22058 54525 22070
rect 54597 22070 54609 22446
rect 54643 22070 54655 22446
rect 54597 22058 54655 22070
rect 54715 22446 54773 22458
rect 54715 22070 54727 22446
rect 54761 22070 54773 22446
rect 54715 22058 54773 22070
rect 54833 22446 54891 22458
rect 54833 22070 54845 22446
rect 54879 22070 54891 22446
rect 54833 22058 54891 22070
rect 54951 22446 55009 22458
rect 54951 22070 54963 22446
rect 54997 22070 55009 22446
rect 54951 22058 55009 22070
rect 55069 22446 55127 22458
rect 55069 22070 55081 22446
rect 55115 22070 55127 22446
rect 55069 22058 55127 22070
rect 55187 22446 55245 22458
rect 55187 22070 55199 22446
rect 55233 22070 55245 22446
rect 55187 22058 55245 22070
rect 55305 22446 55363 22458
rect 55305 22070 55317 22446
rect 55351 22070 55363 22446
rect 56495 22446 56553 22458
rect 55305 22058 55363 22070
rect 55434 22246 55492 22258
rect 55434 22070 55446 22246
rect 55480 22070 55492 22246
rect 55434 22058 55492 22070
rect 55552 22246 55610 22258
rect 55552 22070 55564 22246
rect 55598 22070 55610 22246
rect 55552 22058 55610 22070
rect 55670 22246 55728 22258
rect 55670 22070 55682 22246
rect 55716 22070 55728 22246
rect 55670 22058 55728 22070
rect 55788 22246 55846 22258
rect 55788 22070 55800 22246
rect 55834 22070 55846 22246
rect 55788 22058 55846 22070
rect 56011 22246 56069 22258
rect 56011 22070 56023 22246
rect 56057 22070 56069 22246
rect 56011 22058 56069 22070
rect 56129 22246 56187 22258
rect 56129 22070 56141 22246
rect 56175 22070 56187 22246
rect 56129 22058 56187 22070
rect 56247 22246 56305 22258
rect 56247 22070 56259 22246
rect 56293 22070 56305 22246
rect 56247 22058 56305 22070
rect 56365 22246 56423 22258
rect 56365 22070 56377 22246
rect 56411 22070 56423 22246
rect 56365 22058 56423 22070
rect 56495 22070 56507 22446
rect 56541 22070 56553 22446
rect 56495 22058 56553 22070
rect 56613 22446 56671 22458
rect 56613 22070 56625 22446
rect 56659 22070 56671 22446
rect 56613 22058 56671 22070
rect 56731 22446 56789 22458
rect 56731 22070 56743 22446
rect 56777 22070 56789 22446
rect 56731 22058 56789 22070
rect 56849 22446 56907 22458
rect 56849 22070 56861 22446
rect 56895 22070 56907 22446
rect 56849 22058 56907 22070
rect 56967 22446 57025 22458
rect 56967 22070 56979 22446
rect 57013 22070 57025 22446
rect 56967 22058 57025 22070
rect 57085 22446 57143 22458
rect 57085 22070 57097 22446
rect 57131 22070 57143 22446
rect 57085 22058 57143 22070
rect 57203 22446 57261 22458
rect 57203 22070 57215 22446
rect 57249 22070 57261 22446
rect 61155 22450 61213 22462
rect 57203 22058 57261 22070
rect 57332 22246 57390 22258
rect 57332 22070 57344 22246
rect 57378 22070 57390 22246
rect 57332 22058 57390 22070
rect 57450 22246 57508 22258
rect 57450 22070 57462 22246
rect 57496 22070 57508 22246
rect 57450 22058 57508 22070
rect 57568 22246 57626 22258
rect 57568 22070 57580 22246
rect 57614 22070 57626 22246
rect 57568 22058 57626 22070
rect 57686 22246 57744 22258
rect 57686 22070 57698 22246
rect 57732 22070 57744 22246
rect 57686 22058 57744 22070
rect 49904 21758 49962 21770
rect 49904 21382 49916 21758
rect 49950 21382 49962 21758
rect 49904 21370 49962 21382
rect 50022 21758 50080 21770
rect 50022 21382 50034 21758
rect 50068 21382 50080 21758
rect 50022 21370 50080 21382
rect 50140 21758 50198 21770
rect 50140 21382 50152 21758
rect 50186 21382 50198 21758
rect 50140 21370 50198 21382
rect 50258 21758 50316 21770
rect 50258 21382 50270 21758
rect 50304 21382 50316 21758
rect 50258 21370 50316 21382
rect 50376 21758 50434 21770
rect 50376 21382 50388 21758
rect 50422 21382 50434 21758
rect 50376 21370 50434 21382
rect 50494 21758 50552 21770
rect 50494 21382 50506 21758
rect 50540 21382 50552 21758
rect 50494 21370 50552 21382
rect 50612 21758 50670 21770
rect 50612 21382 50624 21758
rect 50658 21382 50670 21758
rect 50612 21370 50670 21382
rect 52644 21259 52702 21271
rect 52644 21083 52656 21259
rect 52690 21083 52702 21259
rect 52644 21071 52702 21083
rect 52762 21259 52820 21271
rect 52762 21083 52774 21259
rect 52808 21083 52820 21259
rect 52762 21071 52820 21083
rect 52880 21259 52938 21271
rect 52880 21083 52892 21259
rect 52926 21083 52938 21259
rect 52880 21071 52938 21083
rect 52998 21259 53056 21271
rect 52998 21083 53010 21259
rect 53044 21083 53056 21259
rect 52998 21071 53056 21083
rect 53116 21259 53174 21271
rect 53116 21083 53128 21259
rect 53162 21083 53174 21259
rect 53116 21071 53174 21083
rect 53234 21259 53292 21271
rect 53234 21083 53246 21259
rect 53280 21083 53292 21259
rect 53234 21071 53292 21083
rect 53352 21259 53410 21271
rect 53352 21083 53364 21259
rect 53398 21083 53410 21259
rect 53352 21071 53410 21083
rect 53470 21259 53528 21271
rect 53470 21083 53482 21259
rect 53516 21083 53528 21259
rect 53470 21071 53528 21083
rect 53588 21259 53646 21271
rect 53588 21083 53600 21259
rect 53634 21083 53646 21259
rect 53588 21071 53646 21083
rect 53706 21259 53764 21271
rect 53706 21083 53718 21259
rect 53752 21083 53764 21259
rect 53706 21071 53764 21083
rect 54540 21753 54598 21765
rect 54540 21377 54552 21753
rect 54586 21377 54598 21753
rect 54540 21365 54598 21377
rect 54658 21753 54716 21765
rect 54658 21377 54670 21753
rect 54704 21377 54716 21753
rect 54658 21365 54716 21377
rect 54776 21753 54834 21765
rect 54776 21377 54788 21753
rect 54822 21377 54834 21753
rect 54776 21365 54834 21377
rect 54894 21753 54952 21765
rect 54894 21377 54906 21753
rect 54940 21377 54952 21753
rect 54894 21365 54952 21377
rect 55012 21753 55070 21765
rect 55012 21377 55024 21753
rect 55058 21377 55070 21753
rect 55012 21365 55070 21377
rect 55130 21753 55188 21765
rect 55130 21377 55142 21753
rect 55176 21377 55188 21753
rect 55130 21365 55188 21377
rect 55248 21753 55306 21765
rect 55248 21377 55260 21753
rect 55294 21377 55306 21753
rect 55248 21365 55306 21377
rect 60671 22250 60729 22262
rect 60671 22074 60683 22250
rect 60717 22074 60729 22250
rect 60671 22062 60729 22074
rect 60789 22250 60847 22262
rect 60789 22074 60801 22250
rect 60835 22074 60847 22250
rect 60789 22062 60847 22074
rect 60907 22250 60965 22262
rect 60907 22074 60919 22250
rect 60953 22074 60965 22250
rect 60907 22062 60965 22074
rect 61025 22250 61083 22262
rect 61025 22074 61037 22250
rect 61071 22074 61083 22250
rect 61025 22062 61083 22074
rect 61155 22074 61167 22450
rect 61201 22074 61213 22450
rect 61155 22062 61213 22074
rect 61273 22450 61331 22462
rect 61273 22074 61285 22450
rect 61319 22074 61331 22450
rect 61273 22062 61331 22074
rect 61391 22450 61449 22462
rect 61391 22074 61403 22450
rect 61437 22074 61449 22450
rect 61391 22062 61449 22074
rect 61509 22450 61567 22462
rect 61509 22074 61521 22450
rect 61555 22074 61567 22450
rect 61509 22062 61567 22074
rect 61627 22450 61685 22462
rect 61627 22074 61639 22450
rect 61673 22074 61685 22450
rect 61627 22062 61685 22074
rect 61745 22450 61803 22462
rect 61745 22074 61757 22450
rect 61791 22074 61803 22450
rect 61745 22062 61803 22074
rect 61863 22450 61921 22462
rect 61863 22074 61875 22450
rect 61909 22074 61921 22450
rect 63053 22450 63111 22462
rect 61863 22062 61921 22074
rect 61992 22250 62050 22262
rect 61992 22074 62004 22250
rect 62038 22074 62050 22250
rect 61992 22062 62050 22074
rect 62110 22250 62168 22262
rect 62110 22074 62122 22250
rect 62156 22074 62168 22250
rect 62110 22062 62168 22074
rect 62228 22250 62286 22262
rect 62228 22074 62240 22250
rect 62274 22074 62286 22250
rect 62228 22062 62286 22074
rect 62346 22250 62404 22262
rect 62346 22074 62358 22250
rect 62392 22074 62404 22250
rect 62346 22062 62404 22074
rect 62569 22250 62627 22262
rect 62569 22074 62581 22250
rect 62615 22074 62627 22250
rect 62569 22062 62627 22074
rect 62687 22250 62745 22262
rect 62687 22074 62699 22250
rect 62733 22074 62745 22250
rect 62687 22062 62745 22074
rect 62805 22250 62863 22262
rect 62805 22074 62817 22250
rect 62851 22074 62863 22250
rect 62805 22062 62863 22074
rect 62923 22250 62981 22262
rect 62923 22074 62935 22250
rect 62969 22074 62981 22250
rect 62923 22062 62981 22074
rect 63053 22074 63065 22450
rect 63099 22074 63111 22450
rect 63053 22062 63111 22074
rect 63171 22450 63229 22462
rect 63171 22074 63183 22450
rect 63217 22074 63229 22450
rect 63171 22062 63229 22074
rect 63289 22450 63347 22462
rect 63289 22074 63301 22450
rect 63335 22074 63347 22450
rect 63289 22062 63347 22074
rect 63407 22450 63465 22462
rect 63407 22074 63419 22450
rect 63453 22074 63465 22450
rect 63407 22062 63465 22074
rect 63525 22450 63583 22462
rect 63525 22074 63537 22450
rect 63571 22074 63583 22450
rect 63525 22062 63583 22074
rect 63643 22450 63701 22462
rect 63643 22074 63655 22450
rect 63689 22074 63701 22450
rect 63643 22062 63701 22074
rect 63761 22450 63819 22462
rect 63761 22074 63773 22450
rect 63807 22074 63819 22450
rect 63761 22062 63819 22074
rect 63890 22250 63948 22262
rect 63890 22074 63902 22250
rect 63936 22074 63948 22250
rect 63890 22062 63948 22074
rect 64008 22250 64066 22262
rect 64008 22074 64020 22250
rect 64054 22074 64066 22250
rect 64008 22062 64066 22074
rect 64126 22250 64184 22262
rect 64126 22074 64138 22250
rect 64172 22074 64184 22250
rect 64126 22062 64184 22074
rect 64244 22250 64302 22262
rect 64244 22074 64256 22250
rect 64290 22074 64302 22250
rect 64244 22062 64302 22074
rect 56438 21753 56496 21765
rect 56438 21377 56450 21753
rect 56484 21377 56496 21753
rect 56438 21365 56496 21377
rect 56556 21753 56614 21765
rect 56556 21377 56568 21753
rect 56602 21377 56614 21753
rect 56556 21365 56614 21377
rect 56674 21753 56732 21765
rect 56674 21377 56686 21753
rect 56720 21377 56732 21753
rect 56674 21365 56732 21377
rect 56792 21753 56850 21765
rect 56792 21377 56804 21753
rect 56838 21377 56850 21753
rect 56792 21365 56850 21377
rect 56910 21753 56968 21765
rect 56910 21377 56922 21753
rect 56956 21377 56968 21753
rect 56910 21365 56968 21377
rect 57028 21753 57086 21765
rect 57028 21377 57040 21753
rect 57074 21377 57086 21753
rect 57028 21365 57086 21377
rect 57146 21753 57204 21765
rect 57146 21377 57158 21753
rect 57192 21377 57204 21753
rect 57146 21365 57204 21377
rect 59202 21263 59260 21275
rect 59202 21087 59214 21263
rect 59248 21087 59260 21263
rect 59202 21075 59260 21087
rect 59320 21263 59378 21275
rect 59320 21087 59332 21263
rect 59366 21087 59378 21263
rect 59320 21075 59378 21087
rect 59438 21263 59496 21275
rect 59438 21087 59450 21263
rect 59484 21087 59496 21263
rect 59438 21075 59496 21087
rect 59556 21263 59614 21275
rect 59556 21087 59568 21263
rect 59602 21087 59614 21263
rect 59556 21075 59614 21087
rect 59674 21263 59732 21275
rect 59674 21087 59686 21263
rect 59720 21087 59732 21263
rect 59674 21075 59732 21087
rect 59792 21263 59850 21275
rect 59792 21087 59804 21263
rect 59838 21087 59850 21263
rect 59792 21075 59850 21087
rect 59910 21263 59968 21275
rect 59910 21087 59922 21263
rect 59956 21087 59968 21263
rect 59910 21075 59968 21087
rect 60028 21263 60086 21275
rect 60028 21087 60040 21263
rect 60074 21087 60086 21263
rect 60028 21075 60086 21087
rect 60146 21263 60204 21275
rect 60146 21087 60158 21263
rect 60192 21087 60204 21263
rect 60146 21075 60204 21087
rect 60264 21263 60322 21275
rect 60264 21087 60276 21263
rect 60310 21087 60322 21263
rect 60264 21075 60322 21087
rect 61098 21757 61156 21769
rect 61098 21381 61110 21757
rect 61144 21381 61156 21757
rect 61098 21369 61156 21381
rect 61216 21757 61274 21769
rect 61216 21381 61228 21757
rect 61262 21381 61274 21757
rect 61216 21369 61274 21381
rect 61334 21757 61392 21769
rect 61334 21381 61346 21757
rect 61380 21381 61392 21757
rect 61334 21369 61392 21381
rect 61452 21757 61510 21769
rect 61452 21381 61464 21757
rect 61498 21381 61510 21757
rect 61452 21369 61510 21381
rect 61570 21757 61628 21769
rect 61570 21381 61582 21757
rect 61616 21381 61628 21757
rect 61570 21369 61628 21381
rect 61688 21757 61746 21769
rect 61688 21381 61700 21757
rect 61734 21381 61746 21757
rect 61688 21369 61746 21381
rect 61806 21757 61864 21769
rect 61806 21381 61818 21757
rect 61852 21381 61864 21757
rect 61806 21369 61864 21381
rect 70713 22061 70913 22073
rect 70713 22027 70725 22061
rect 70901 22027 70913 22061
rect 70713 22015 70913 22027
rect 70713 21943 70913 21955
rect 70713 21909 70725 21943
rect 70901 21909 70913 21943
rect 70713 21897 70913 21909
rect 62996 21757 63054 21769
rect 62996 21381 63008 21757
rect 63042 21381 63054 21757
rect 62996 21369 63054 21381
rect 63114 21757 63172 21769
rect 63114 21381 63126 21757
rect 63160 21381 63172 21757
rect 63114 21369 63172 21381
rect 63232 21757 63290 21769
rect 63232 21381 63244 21757
rect 63278 21381 63290 21757
rect 63232 21369 63290 21381
rect 63350 21757 63408 21769
rect 63350 21381 63362 21757
rect 63396 21381 63408 21757
rect 63350 21369 63408 21381
rect 63468 21757 63526 21769
rect 63468 21381 63480 21757
rect 63514 21381 63526 21757
rect 63468 21369 63526 21381
rect 63586 21757 63644 21769
rect 63586 21381 63598 21757
rect 63632 21381 63644 21757
rect 63586 21369 63644 21381
rect 63704 21757 63762 21769
rect 63704 21381 63716 21757
rect 63750 21381 63762 21757
rect 63704 21369 63762 21381
rect 70713 21825 70913 21837
rect 70713 21791 70725 21825
rect 70901 21791 70913 21825
rect 70713 21779 70913 21791
rect 70713 21707 70913 21719
rect 70713 21673 70725 21707
rect 70901 21673 70913 21707
rect 70713 21632 70913 21673
rect 70513 21620 70913 21632
rect 70513 21586 70525 21620
rect 70901 21586 70913 21620
rect 70513 21574 70913 21586
rect 70513 21502 70913 21514
rect 70513 21468 70525 21502
rect 70901 21468 70913 21502
rect 70513 21456 70913 21468
rect 70513 21384 70913 21396
rect 70513 21350 70525 21384
rect 70901 21350 70913 21384
rect 70513 21338 70913 21350
rect 70513 21266 70913 21278
rect 70513 21232 70525 21266
rect 70901 21232 70913 21266
rect 70513 21220 70913 21232
rect 70513 21153 70913 21165
rect 70513 21119 70525 21153
rect 70901 21119 70913 21153
rect 70513 21107 70913 21119
rect 70513 21035 70913 21047
rect 70513 21001 70525 21035
rect 70901 21001 70913 21035
rect 70513 20989 70913 21001
rect 70513 20917 70913 20929
rect 70513 20883 70525 20917
rect 70901 20883 70913 20917
rect 70513 20871 70913 20883
rect 70513 20799 70913 20811
rect 70513 20765 70525 20799
rect 70901 20765 70913 20799
rect 70513 20753 70913 20765
rect 70513 20681 70913 20693
rect 70513 20647 70525 20681
rect 70901 20647 70913 20681
rect 70513 20635 70913 20647
rect 70513 20563 70913 20575
rect 70513 20529 70525 20563
rect 70901 20529 70913 20563
rect 70513 20517 70913 20529
rect 70513 20445 70913 20457
rect 70513 20411 70525 20445
rect 70901 20411 70913 20445
rect 70513 20399 70913 20411
rect 70513 20326 70913 20338
rect 70513 20292 70525 20326
rect 70901 20292 70913 20326
rect 70513 20280 70913 20292
rect 70513 20208 70913 20220
rect 70513 20174 70525 20208
rect 70901 20174 70913 20208
rect 70513 20162 70913 20174
rect 70513 20090 70913 20102
rect 70513 20056 70525 20090
rect 70901 20056 70913 20090
rect 70513 20044 70913 20056
rect 70513 19972 70913 19984
rect 70513 19938 70525 19972
rect 70901 19938 70913 19972
rect 70513 19926 70913 19938
rect 70713 19853 70913 19865
rect 70713 19819 70725 19853
rect 70901 19819 70913 19853
rect 70713 19807 70913 19819
rect 70713 19735 70913 19747
rect 70713 19701 70725 19735
rect 70901 19701 70913 19735
rect 70713 19689 70913 19701
rect 70713 19617 70913 19629
rect 70713 19583 70725 19617
rect 70901 19583 70913 19617
rect 70713 19571 70913 19583
rect 70713 19499 70913 19511
rect 70713 19465 70725 19499
rect 70901 19465 70913 19499
rect 70713 19453 70913 19465
rect 39599 18989 39657 19001
rect 39599 18613 39611 18989
rect 39645 18613 39657 18989
rect 39599 18601 39657 18613
rect 39717 18989 39775 19001
rect 39717 18613 39729 18989
rect 39763 18613 39775 18989
rect 39717 18601 39775 18613
rect 39835 18989 39893 19001
rect 39835 18613 39847 18989
rect 39881 18613 39893 18989
rect 39835 18601 39893 18613
rect 39953 18989 40011 19001
rect 39953 18613 39965 18989
rect 39999 18613 40011 18989
rect 39953 18601 40011 18613
rect 40071 18989 40129 19001
rect 40071 18613 40083 18989
rect 40117 18613 40129 18989
rect 40071 18601 40129 18613
rect 40189 18989 40247 19001
rect 40189 18613 40201 18989
rect 40235 18613 40247 18989
rect 40189 18601 40247 18613
rect 40307 18989 40365 19001
rect 40307 18613 40319 18989
rect 40353 18613 40365 18989
rect 40307 18601 40365 18613
rect 40741 18985 40799 18997
rect 40741 18609 40753 18985
rect 40787 18609 40799 18985
rect 40741 18597 40799 18609
rect 40859 18985 40917 18997
rect 40859 18609 40871 18985
rect 40905 18609 40917 18985
rect 40859 18597 40917 18609
rect 40977 18985 41035 18997
rect 40977 18609 40989 18985
rect 41023 18609 41035 18985
rect 40977 18597 41035 18609
rect 41095 18985 41153 18997
rect 41095 18609 41107 18985
rect 41141 18609 41153 18985
rect 41095 18597 41153 18609
rect 41213 18985 41271 18997
rect 41213 18609 41225 18985
rect 41259 18609 41271 18985
rect 41213 18597 41271 18609
rect 41331 18985 41389 18997
rect 41331 18609 41343 18985
rect 41377 18609 41389 18985
rect 41331 18597 41389 18609
rect 41449 18985 41507 18997
rect 41449 18609 41461 18985
rect 41495 18609 41507 18985
rect 46157 18985 46215 18997
rect 42712 18913 42770 18925
rect 42712 18737 42724 18913
rect 42758 18737 42770 18913
rect 42712 18725 42770 18737
rect 42830 18913 42888 18925
rect 42830 18737 42842 18913
rect 42876 18737 42888 18913
rect 42830 18725 42888 18737
rect 42948 18913 43006 18925
rect 42948 18737 42960 18913
rect 42994 18737 43006 18913
rect 42948 18725 43006 18737
rect 43066 18913 43124 18925
rect 43066 18737 43078 18913
rect 43112 18737 43124 18913
rect 43066 18725 43124 18737
rect 43184 18913 43242 18925
rect 43184 18737 43196 18913
rect 43230 18737 43242 18913
rect 43184 18725 43242 18737
rect 43302 18913 43360 18925
rect 43302 18737 43314 18913
rect 43348 18737 43360 18913
rect 43302 18725 43360 18737
rect 43420 18913 43478 18925
rect 43420 18737 43432 18913
rect 43466 18737 43478 18913
rect 43420 18725 43478 18737
rect 43538 18913 43596 18925
rect 43538 18737 43550 18913
rect 43584 18737 43596 18913
rect 43538 18725 43596 18737
rect 43656 18913 43714 18925
rect 43656 18737 43668 18913
rect 43702 18737 43714 18913
rect 43656 18725 43714 18737
rect 43774 18913 43832 18925
rect 43774 18737 43786 18913
rect 43820 18737 43832 18913
rect 43774 18725 43832 18737
rect 41449 18597 41507 18609
rect 46157 18609 46169 18985
rect 46203 18609 46215 18985
rect 46157 18597 46215 18609
rect 46275 18985 46333 18997
rect 46275 18609 46287 18985
rect 46321 18609 46333 18985
rect 46275 18597 46333 18609
rect 46393 18985 46451 18997
rect 46393 18609 46405 18985
rect 46439 18609 46451 18985
rect 46393 18597 46451 18609
rect 46511 18985 46569 18997
rect 46511 18609 46523 18985
rect 46557 18609 46569 18985
rect 46511 18597 46569 18609
rect 46629 18985 46687 18997
rect 46629 18609 46641 18985
rect 46675 18609 46687 18985
rect 46629 18597 46687 18609
rect 46747 18985 46805 18997
rect 46747 18609 46759 18985
rect 46793 18609 46805 18985
rect 46747 18597 46805 18609
rect 46865 18985 46923 18997
rect 46865 18609 46877 18985
rect 46911 18609 46923 18985
rect 46865 18597 46923 18609
rect 47299 18981 47357 18993
rect 47299 18605 47311 18981
rect 47345 18605 47357 18981
rect 39524 18206 39582 18218
rect 39524 18030 39536 18206
rect 39570 18030 39582 18206
rect 39524 18018 39582 18030
rect 39642 18206 39700 18218
rect 39642 18030 39654 18206
rect 39688 18030 39700 18206
rect 39642 18018 39700 18030
rect 39760 18206 39818 18218
rect 39760 18030 39772 18206
rect 39806 18030 39818 18206
rect 39760 18018 39818 18030
rect 39878 18206 39936 18218
rect 39878 18030 39890 18206
rect 39924 18030 39936 18206
rect 39878 18018 39936 18030
rect 40666 18202 40724 18214
rect 40666 18026 40678 18202
rect 40712 18026 40724 18202
rect 40666 18014 40724 18026
rect 40784 18202 40842 18214
rect 40784 18026 40796 18202
rect 40830 18026 40842 18202
rect 40784 18014 40842 18026
rect 40902 18202 40960 18214
rect 40902 18026 40914 18202
rect 40948 18026 40960 18202
rect 40902 18014 40960 18026
rect 41020 18202 41078 18214
rect 41020 18026 41032 18202
rect 41066 18026 41078 18202
rect 41020 18014 41078 18026
rect 47299 18593 47357 18605
rect 47417 18981 47475 18993
rect 47417 18605 47429 18981
rect 47463 18605 47475 18981
rect 47417 18593 47475 18605
rect 47535 18981 47593 18993
rect 47535 18605 47547 18981
rect 47581 18605 47593 18981
rect 47535 18593 47593 18605
rect 47653 18981 47711 18993
rect 47653 18605 47665 18981
rect 47699 18605 47711 18981
rect 47653 18593 47711 18605
rect 47771 18981 47829 18993
rect 47771 18605 47783 18981
rect 47817 18605 47829 18981
rect 47771 18593 47829 18605
rect 47889 18981 47947 18993
rect 47889 18605 47901 18981
rect 47935 18605 47947 18981
rect 47889 18593 47947 18605
rect 48007 18981 48065 18993
rect 52691 18990 52749 19002
rect 48007 18605 48019 18981
rect 48053 18605 48065 18981
rect 49270 18909 49328 18921
rect 49270 18733 49282 18909
rect 49316 18733 49328 18909
rect 49270 18721 49328 18733
rect 49388 18909 49446 18921
rect 49388 18733 49400 18909
rect 49434 18733 49446 18909
rect 49388 18721 49446 18733
rect 49506 18909 49564 18921
rect 49506 18733 49518 18909
rect 49552 18733 49564 18909
rect 49506 18721 49564 18733
rect 49624 18909 49682 18921
rect 49624 18733 49636 18909
rect 49670 18733 49682 18909
rect 49624 18721 49682 18733
rect 49742 18909 49800 18921
rect 49742 18733 49754 18909
rect 49788 18733 49800 18909
rect 49742 18721 49800 18733
rect 49860 18909 49918 18921
rect 49860 18733 49872 18909
rect 49906 18733 49918 18909
rect 49860 18721 49918 18733
rect 49978 18909 50036 18921
rect 49978 18733 49990 18909
rect 50024 18733 50036 18909
rect 49978 18721 50036 18733
rect 50096 18909 50154 18921
rect 50096 18733 50108 18909
rect 50142 18733 50154 18909
rect 50096 18721 50154 18733
rect 50214 18909 50272 18921
rect 50214 18733 50226 18909
rect 50260 18733 50272 18909
rect 50214 18721 50272 18733
rect 50332 18909 50390 18921
rect 50332 18733 50344 18909
rect 50378 18733 50390 18909
rect 50332 18721 50390 18733
rect 48007 18593 48065 18605
rect 52691 18614 52703 18990
rect 52737 18614 52749 18990
rect 52691 18602 52749 18614
rect 52809 18990 52867 19002
rect 52809 18614 52821 18990
rect 52855 18614 52867 18990
rect 52809 18602 52867 18614
rect 52927 18990 52985 19002
rect 52927 18614 52939 18990
rect 52973 18614 52985 18990
rect 52927 18602 52985 18614
rect 53045 18990 53103 19002
rect 53045 18614 53057 18990
rect 53091 18614 53103 18990
rect 53045 18602 53103 18614
rect 53163 18990 53221 19002
rect 53163 18614 53175 18990
rect 53209 18614 53221 18990
rect 53163 18602 53221 18614
rect 53281 18990 53339 19002
rect 53281 18614 53293 18990
rect 53327 18614 53339 18990
rect 53281 18602 53339 18614
rect 53399 18990 53457 19002
rect 53399 18614 53411 18990
rect 53445 18614 53457 18990
rect 53399 18602 53457 18614
rect 53833 18986 53891 18998
rect 53833 18610 53845 18986
rect 53879 18610 53891 18986
rect 46082 18202 46140 18214
rect 46082 18026 46094 18202
rect 46128 18026 46140 18202
rect 46082 18014 46140 18026
rect 46200 18202 46258 18214
rect 46200 18026 46212 18202
rect 46246 18026 46258 18202
rect 46200 18014 46258 18026
rect 46318 18202 46376 18214
rect 46318 18026 46330 18202
rect 46364 18026 46376 18202
rect 46318 18014 46376 18026
rect 46436 18202 46494 18214
rect 46436 18026 46448 18202
rect 46482 18026 46494 18202
rect 46436 18014 46494 18026
rect 47224 18198 47282 18210
rect 47224 18022 47236 18198
rect 47270 18022 47282 18198
rect 47224 18010 47282 18022
rect 47342 18198 47400 18210
rect 47342 18022 47354 18198
rect 47388 18022 47400 18198
rect 47342 18010 47400 18022
rect 47460 18198 47518 18210
rect 47460 18022 47472 18198
rect 47506 18022 47518 18198
rect 47460 18010 47518 18022
rect 47578 18198 47636 18210
rect 47578 18022 47590 18198
rect 47624 18022 47636 18198
rect 47578 18010 47636 18022
rect 53833 18598 53891 18610
rect 53951 18986 54009 18998
rect 53951 18610 53963 18986
rect 53997 18610 54009 18986
rect 53951 18598 54009 18610
rect 54069 18986 54127 18998
rect 54069 18610 54081 18986
rect 54115 18610 54127 18986
rect 54069 18598 54127 18610
rect 54187 18986 54245 18998
rect 54187 18610 54199 18986
rect 54233 18610 54245 18986
rect 54187 18598 54245 18610
rect 54305 18986 54363 18998
rect 54305 18610 54317 18986
rect 54351 18610 54363 18986
rect 54305 18598 54363 18610
rect 54423 18986 54481 18998
rect 54423 18610 54435 18986
rect 54469 18610 54481 18986
rect 54423 18598 54481 18610
rect 54541 18986 54599 18998
rect 54541 18610 54553 18986
rect 54587 18610 54599 18986
rect 59204 18993 59262 19005
rect 55804 18914 55862 18926
rect 55804 18738 55816 18914
rect 55850 18738 55862 18914
rect 55804 18726 55862 18738
rect 55922 18914 55980 18926
rect 55922 18738 55934 18914
rect 55968 18738 55980 18914
rect 55922 18726 55980 18738
rect 56040 18914 56098 18926
rect 56040 18738 56052 18914
rect 56086 18738 56098 18914
rect 56040 18726 56098 18738
rect 56158 18914 56216 18926
rect 56158 18738 56170 18914
rect 56204 18738 56216 18914
rect 56158 18726 56216 18738
rect 56276 18914 56334 18926
rect 56276 18738 56288 18914
rect 56322 18738 56334 18914
rect 56276 18726 56334 18738
rect 56394 18914 56452 18926
rect 56394 18738 56406 18914
rect 56440 18738 56452 18914
rect 56394 18726 56452 18738
rect 56512 18914 56570 18926
rect 56512 18738 56524 18914
rect 56558 18738 56570 18914
rect 56512 18726 56570 18738
rect 56630 18914 56688 18926
rect 56630 18738 56642 18914
rect 56676 18738 56688 18914
rect 56630 18726 56688 18738
rect 56748 18914 56806 18926
rect 56748 18738 56760 18914
rect 56794 18738 56806 18914
rect 56748 18726 56806 18738
rect 56866 18914 56924 18926
rect 56866 18738 56878 18914
rect 56912 18738 56924 18914
rect 56866 18726 56924 18738
rect 54541 18598 54599 18610
rect 59204 18617 59216 18993
rect 59250 18617 59262 18993
rect 59204 18605 59262 18617
rect 59322 18993 59380 19005
rect 59322 18617 59334 18993
rect 59368 18617 59380 18993
rect 59322 18605 59380 18617
rect 59440 18993 59498 19005
rect 59440 18617 59452 18993
rect 59486 18617 59498 18993
rect 59440 18605 59498 18617
rect 59558 18993 59616 19005
rect 59558 18617 59570 18993
rect 59604 18617 59616 18993
rect 59558 18605 59616 18617
rect 59676 18993 59734 19005
rect 59676 18617 59688 18993
rect 59722 18617 59734 18993
rect 59676 18605 59734 18617
rect 59794 18993 59852 19005
rect 59794 18617 59806 18993
rect 59840 18617 59852 18993
rect 59794 18605 59852 18617
rect 59912 18993 59970 19005
rect 59912 18617 59924 18993
rect 59958 18617 59970 18993
rect 59912 18605 59970 18617
rect 60346 18989 60404 19001
rect 60346 18613 60358 18989
rect 60392 18613 60404 18989
rect 52616 18207 52674 18219
rect 52616 18031 52628 18207
rect 52662 18031 52674 18207
rect 52616 18019 52674 18031
rect 52734 18207 52792 18219
rect 52734 18031 52746 18207
rect 52780 18031 52792 18207
rect 52734 18019 52792 18031
rect 52852 18207 52910 18219
rect 52852 18031 52864 18207
rect 52898 18031 52910 18207
rect 52852 18019 52910 18031
rect 52970 18207 53028 18219
rect 52970 18031 52982 18207
rect 53016 18031 53028 18207
rect 52970 18019 53028 18031
rect 53758 18203 53816 18215
rect 53758 18027 53770 18203
rect 53804 18027 53816 18203
rect 53758 18015 53816 18027
rect 53876 18203 53934 18215
rect 53876 18027 53888 18203
rect 53922 18027 53934 18203
rect 53876 18015 53934 18027
rect 53994 18203 54052 18215
rect 53994 18027 54006 18203
rect 54040 18027 54052 18203
rect 53994 18015 54052 18027
rect 54112 18203 54170 18215
rect 54112 18027 54124 18203
rect 54158 18027 54170 18203
rect 54112 18015 54170 18027
rect 60346 18601 60404 18613
rect 60464 18989 60522 19001
rect 60464 18613 60476 18989
rect 60510 18613 60522 18989
rect 60464 18601 60522 18613
rect 60582 18989 60640 19001
rect 60582 18613 60594 18989
rect 60628 18613 60640 18989
rect 60582 18601 60640 18613
rect 60700 18989 60758 19001
rect 60700 18613 60712 18989
rect 60746 18613 60758 18989
rect 60700 18601 60758 18613
rect 60818 18989 60876 19001
rect 60818 18613 60830 18989
rect 60864 18613 60876 18989
rect 60818 18601 60876 18613
rect 60936 18989 60994 19001
rect 60936 18613 60948 18989
rect 60982 18613 60994 18989
rect 60936 18601 60994 18613
rect 61054 18989 61112 19001
rect 61054 18613 61066 18989
rect 61100 18613 61112 18989
rect 62317 18917 62375 18929
rect 62317 18741 62329 18917
rect 62363 18741 62375 18917
rect 62317 18729 62375 18741
rect 62435 18917 62493 18929
rect 62435 18741 62447 18917
rect 62481 18741 62493 18917
rect 62435 18729 62493 18741
rect 62553 18917 62611 18929
rect 62553 18741 62565 18917
rect 62599 18741 62611 18917
rect 62553 18729 62611 18741
rect 62671 18917 62729 18929
rect 62671 18741 62683 18917
rect 62717 18741 62729 18917
rect 62671 18729 62729 18741
rect 62789 18917 62847 18929
rect 62789 18741 62801 18917
rect 62835 18741 62847 18917
rect 62789 18729 62847 18741
rect 62907 18917 62965 18929
rect 62907 18741 62919 18917
rect 62953 18741 62965 18917
rect 62907 18729 62965 18741
rect 63025 18917 63083 18929
rect 63025 18741 63037 18917
rect 63071 18741 63083 18917
rect 63025 18729 63083 18741
rect 63143 18917 63201 18929
rect 63143 18741 63155 18917
rect 63189 18741 63201 18917
rect 63143 18729 63201 18741
rect 63261 18917 63319 18929
rect 63261 18741 63273 18917
rect 63307 18741 63319 18917
rect 63261 18729 63319 18741
rect 63379 18917 63437 18929
rect 63379 18741 63391 18917
rect 63425 18741 63437 18917
rect 70713 18917 70913 18929
rect 70713 18883 70725 18917
rect 70901 18883 70913 18917
rect 70713 18871 70913 18883
rect 63379 18729 63437 18741
rect 70713 18799 70913 18811
rect 70713 18765 70725 18799
rect 70901 18765 70913 18799
rect 70713 18753 70913 18765
rect 61054 18601 61112 18613
rect 70713 18681 70913 18693
rect 70713 18647 70725 18681
rect 70901 18647 70913 18681
rect 70713 18635 70913 18647
rect 70713 18563 70913 18575
rect 70713 18529 70725 18563
rect 70901 18529 70913 18563
rect 59129 18210 59187 18222
rect 59129 18034 59141 18210
rect 59175 18034 59187 18210
rect 59129 18022 59187 18034
rect 59247 18210 59305 18222
rect 59247 18034 59259 18210
rect 59293 18034 59305 18210
rect 59247 18022 59305 18034
rect 59365 18210 59423 18222
rect 59365 18034 59377 18210
rect 59411 18034 59423 18210
rect 59365 18022 59423 18034
rect 59483 18210 59541 18222
rect 59483 18034 59495 18210
rect 59529 18034 59541 18210
rect 59483 18022 59541 18034
rect 60271 18206 60329 18218
rect 60271 18030 60283 18206
rect 60317 18030 60329 18206
rect 60271 18018 60329 18030
rect 60389 18206 60447 18218
rect 60389 18030 60401 18206
rect 60435 18030 60447 18206
rect 60389 18018 60447 18030
rect 60507 18206 60565 18218
rect 60507 18030 60519 18206
rect 60553 18030 60565 18206
rect 60507 18018 60565 18030
rect 60625 18206 60683 18218
rect 60625 18030 60637 18206
rect 60671 18030 60683 18206
rect 60625 18018 60683 18030
rect 70713 18488 70913 18529
rect 70513 18476 70913 18488
rect 70513 18442 70525 18476
rect 70901 18442 70913 18476
rect 70513 18430 70913 18442
rect 70513 18358 70913 18370
rect 70513 18324 70525 18358
rect 70901 18324 70913 18358
rect 70513 18312 70913 18324
rect 70513 18240 70913 18252
rect 70513 18206 70525 18240
rect 70901 18206 70913 18240
rect 70513 18194 70913 18206
rect 70513 18122 70913 18134
rect 70513 18088 70525 18122
rect 70901 18088 70913 18122
rect 70513 18076 70913 18088
rect 70513 18009 70913 18021
rect 70513 17975 70525 18009
rect 70901 17975 70913 18009
rect 70513 17963 70913 17975
rect 70513 17891 70913 17903
rect 70513 17857 70525 17891
rect 70901 17857 70913 17891
rect 70513 17845 70913 17857
rect 70513 17773 70913 17785
rect 70513 17739 70525 17773
rect 70901 17739 70913 17773
rect 70513 17727 70913 17739
rect 70513 17655 70913 17667
rect 70513 17621 70525 17655
rect 70901 17621 70913 17655
rect 70513 17609 70913 17621
rect 70513 17537 70913 17549
rect 70513 17503 70525 17537
rect 70901 17503 70913 17537
rect 70513 17491 70913 17503
rect 42698 17263 42756 17275
rect 42698 17087 42710 17263
rect 42744 17087 42756 17263
rect 4508 16796 4566 16808
rect 4508 16420 4520 16796
rect 4554 16420 4566 16796
rect 4508 16408 4566 16420
rect 4626 16796 4684 16808
rect 4626 16420 4638 16796
rect 4672 16420 4684 16796
rect 4626 16408 4684 16420
rect 4744 16796 4802 16808
rect 4744 16420 4756 16796
rect 4790 16420 4802 16796
rect 4744 16408 4802 16420
rect 4862 16796 4920 16808
rect 4862 16420 4874 16796
rect 4908 16420 4920 16796
rect 4862 16408 4920 16420
rect 4980 16796 5038 16808
rect 4980 16420 4992 16796
rect 5026 16420 5038 16796
rect 4980 16408 5038 16420
rect 5098 16796 5156 16808
rect 5098 16420 5110 16796
rect 5144 16420 5156 16796
rect 5098 16408 5156 16420
rect 5216 16796 5274 16808
rect 5216 16420 5228 16796
rect 5262 16420 5274 16796
rect 5216 16408 5274 16420
rect 5676 16798 5734 16810
rect 5676 16422 5688 16798
rect 5722 16422 5734 16798
rect 5676 16410 5734 16422
rect 5794 16798 5852 16810
rect 5794 16422 5806 16798
rect 5840 16422 5852 16798
rect 5794 16410 5852 16422
rect 5912 16798 5970 16810
rect 5912 16422 5924 16798
rect 5958 16422 5970 16798
rect 5912 16410 5970 16422
rect 6030 16798 6088 16810
rect 6030 16422 6042 16798
rect 6076 16422 6088 16798
rect 6030 16410 6088 16422
rect 6148 16798 6206 16810
rect 6148 16422 6160 16798
rect 6194 16422 6206 16798
rect 6148 16410 6206 16422
rect 6266 16798 6324 16810
rect 6266 16422 6278 16798
rect 6312 16422 6324 16798
rect 6266 16410 6324 16422
rect 6384 16798 6442 16810
rect 42698 17075 42756 17087
rect 42816 17263 42874 17275
rect 42816 17087 42828 17263
rect 42862 17087 42874 17263
rect 42816 17075 42874 17087
rect 42934 17263 42992 17275
rect 42934 17087 42946 17263
rect 42980 17087 42992 17263
rect 42934 17075 42992 17087
rect 43052 17263 43110 17275
rect 43052 17087 43064 17263
rect 43098 17087 43110 17263
rect 43052 17075 43110 17087
rect 43170 17263 43228 17275
rect 43170 17087 43182 17263
rect 43216 17087 43228 17263
rect 43170 17075 43228 17087
rect 43288 17263 43346 17275
rect 43288 17087 43300 17263
rect 43334 17087 43346 17263
rect 43288 17075 43346 17087
rect 43406 17263 43464 17275
rect 43406 17087 43418 17263
rect 43452 17087 43464 17263
rect 43406 17075 43464 17087
rect 43524 17263 43582 17275
rect 43524 17087 43536 17263
rect 43570 17087 43582 17263
rect 43524 17075 43582 17087
rect 43642 17263 43700 17275
rect 43642 17087 43654 17263
rect 43688 17087 43700 17263
rect 43642 17075 43700 17087
rect 43760 17263 43818 17275
rect 43760 17087 43772 17263
rect 43806 17087 43818 17263
rect 49256 17259 49314 17271
rect 43760 17075 43818 17087
rect 49256 17083 49268 17259
rect 49302 17083 49314 17259
rect 49256 17071 49314 17083
rect 49374 17259 49432 17271
rect 49374 17083 49386 17259
rect 49420 17083 49432 17259
rect 49374 17071 49432 17083
rect 49492 17259 49550 17271
rect 49492 17083 49504 17259
rect 49538 17083 49550 17259
rect 49492 17071 49550 17083
rect 49610 17259 49668 17271
rect 49610 17083 49622 17259
rect 49656 17083 49668 17259
rect 49610 17071 49668 17083
rect 49728 17259 49786 17271
rect 49728 17083 49740 17259
rect 49774 17083 49786 17259
rect 49728 17071 49786 17083
rect 49846 17259 49904 17271
rect 49846 17083 49858 17259
rect 49892 17083 49904 17259
rect 49846 17071 49904 17083
rect 49964 17259 50022 17271
rect 49964 17083 49976 17259
rect 50010 17083 50022 17259
rect 49964 17071 50022 17083
rect 50082 17259 50140 17271
rect 50082 17083 50094 17259
rect 50128 17083 50140 17259
rect 50082 17071 50140 17083
rect 50200 17259 50258 17271
rect 50200 17083 50212 17259
rect 50246 17083 50258 17259
rect 50200 17071 50258 17083
rect 50318 17259 50376 17271
rect 50318 17083 50330 17259
rect 50364 17083 50376 17259
rect 55790 17264 55848 17276
rect 50318 17071 50376 17083
rect 55790 17088 55802 17264
rect 55836 17088 55848 17264
rect 55790 17076 55848 17088
rect 55908 17264 55966 17276
rect 55908 17088 55920 17264
rect 55954 17088 55966 17264
rect 55908 17076 55966 17088
rect 56026 17264 56084 17276
rect 56026 17088 56038 17264
rect 56072 17088 56084 17264
rect 56026 17076 56084 17088
rect 56144 17264 56202 17276
rect 56144 17088 56156 17264
rect 56190 17088 56202 17264
rect 56144 17076 56202 17088
rect 56262 17264 56320 17276
rect 56262 17088 56274 17264
rect 56308 17088 56320 17264
rect 56262 17076 56320 17088
rect 56380 17264 56438 17276
rect 56380 17088 56392 17264
rect 56426 17088 56438 17264
rect 56380 17076 56438 17088
rect 56498 17264 56556 17276
rect 56498 17088 56510 17264
rect 56544 17088 56556 17264
rect 56498 17076 56556 17088
rect 56616 17264 56674 17276
rect 56616 17088 56628 17264
rect 56662 17088 56674 17264
rect 56616 17076 56674 17088
rect 56734 17264 56792 17276
rect 56734 17088 56746 17264
rect 56780 17088 56792 17264
rect 56734 17076 56792 17088
rect 56852 17264 56910 17276
rect 56852 17088 56864 17264
rect 56898 17088 56910 17264
rect 70513 17419 70913 17431
rect 70513 17385 70525 17419
rect 70901 17385 70913 17419
rect 70513 17373 70913 17385
rect 70513 17301 70913 17313
rect 62303 17267 62361 17279
rect 56852 17076 56910 17088
rect 62303 17091 62315 17267
rect 62349 17091 62361 17267
rect 62303 17079 62361 17091
rect 62421 17267 62479 17279
rect 62421 17091 62433 17267
rect 62467 17091 62479 17267
rect 62421 17079 62479 17091
rect 62539 17267 62597 17279
rect 62539 17091 62551 17267
rect 62585 17091 62597 17267
rect 62539 17079 62597 17091
rect 62657 17267 62715 17279
rect 62657 17091 62669 17267
rect 62703 17091 62715 17267
rect 62657 17079 62715 17091
rect 62775 17267 62833 17279
rect 62775 17091 62787 17267
rect 62821 17091 62833 17267
rect 62775 17079 62833 17091
rect 62893 17267 62951 17279
rect 62893 17091 62905 17267
rect 62939 17091 62951 17267
rect 62893 17079 62951 17091
rect 63011 17267 63069 17279
rect 63011 17091 63023 17267
rect 63057 17091 63069 17267
rect 63011 17079 63069 17091
rect 63129 17267 63187 17279
rect 63129 17091 63141 17267
rect 63175 17091 63187 17267
rect 63129 17079 63187 17091
rect 63247 17267 63305 17279
rect 63247 17091 63259 17267
rect 63293 17091 63305 17267
rect 63247 17079 63305 17091
rect 63365 17267 63423 17279
rect 63365 17091 63377 17267
rect 63411 17091 63423 17267
rect 70513 17267 70525 17301
rect 70901 17267 70913 17301
rect 70513 17255 70913 17267
rect 70513 17182 70913 17194
rect 70513 17148 70525 17182
rect 70901 17148 70913 17182
rect 70513 17136 70913 17148
rect 63365 17079 63423 17091
rect 6384 16422 6396 16798
rect 6430 16422 6442 16798
rect 6384 16410 6442 16422
rect 6844 16796 6902 16808
rect 6844 16420 6856 16796
rect 6890 16420 6902 16796
rect 6844 16408 6902 16420
rect 6962 16796 7020 16808
rect 6962 16420 6974 16796
rect 7008 16420 7020 16796
rect 6962 16408 7020 16420
rect 7080 16796 7138 16808
rect 7080 16420 7092 16796
rect 7126 16420 7138 16796
rect 7080 16408 7138 16420
rect 7198 16796 7256 16808
rect 7198 16420 7210 16796
rect 7244 16420 7256 16796
rect 7198 16408 7256 16420
rect 7316 16796 7374 16808
rect 7316 16420 7328 16796
rect 7362 16420 7374 16796
rect 7316 16408 7374 16420
rect 7434 16796 7492 16808
rect 7434 16420 7446 16796
rect 7480 16420 7492 16796
rect 7434 16408 7492 16420
rect 7552 16796 7610 16808
rect 7552 16420 7564 16796
rect 7598 16420 7610 16796
rect 7552 16408 7610 16420
rect 8012 16798 8070 16810
rect 8012 16422 8024 16798
rect 8058 16422 8070 16798
rect 8012 16410 8070 16422
rect 8130 16798 8188 16810
rect 8130 16422 8142 16798
rect 8176 16422 8188 16798
rect 8130 16410 8188 16422
rect 8248 16798 8306 16810
rect 8248 16422 8260 16798
rect 8294 16422 8306 16798
rect 8248 16410 8306 16422
rect 8366 16798 8424 16810
rect 8366 16422 8378 16798
rect 8412 16422 8424 16798
rect 8366 16410 8424 16422
rect 8484 16798 8542 16810
rect 8484 16422 8496 16798
rect 8530 16422 8542 16798
rect 8484 16410 8542 16422
rect 8602 16798 8660 16810
rect 8602 16422 8614 16798
rect 8648 16422 8660 16798
rect 8602 16410 8660 16422
rect 8720 16798 8778 16810
rect 8720 16422 8732 16798
rect 8766 16422 8778 16798
rect 8720 16410 8778 16422
rect 9186 16796 9244 16808
rect 9186 16420 9198 16796
rect 9232 16420 9244 16796
rect 4433 16008 4491 16020
rect 4433 15832 4445 16008
rect 4479 15832 4491 16008
rect 4433 15820 4491 15832
rect 4551 16008 4609 16020
rect 4551 15832 4563 16008
rect 4597 15832 4609 16008
rect 4551 15820 4609 15832
rect 4669 16008 4727 16020
rect 4669 15832 4681 16008
rect 4715 15832 4727 16008
rect 4669 15820 4727 15832
rect 4787 16008 4845 16020
rect 4787 15832 4799 16008
rect 4833 15832 4845 16008
rect 4787 15820 4845 15832
rect 5601 16007 5659 16019
rect 5601 15831 5613 16007
rect 5647 15831 5659 16007
rect 5601 15819 5659 15831
rect 5719 16007 5777 16019
rect 5719 15831 5731 16007
rect 5765 15831 5777 16007
rect 5719 15819 5777 15831
rect 5837 16007 5895 16019
rect 5837 15831 5849 16007
rect 5883 15831 5895 16007
rect 5837 15819 5895 15831
rect 5955 16007 6013 16019
rect 5955 15831 5967 16007
rect 6001 15831 6013 16007
rect 5955 15819 6013 15831
rect 9186 16408 9244 16420
rect 9304 16796 9362 16808
rect 9304 16420 9316 16796
rect 9350 16420 9362 16796
rect 9304 16408 9362 16420
rect 9422 16796 9480 16808
rect 9422 16420 9434 16796
rect 9468 16420 9480 16796
rect 9422 16408 9480 16420
rect 9540 16796 9598 16808
rect 9540 16420 9552 16796
rect 9586 16420 9598 16796
rect 9540 16408 9598 16420
rect 9658 16796 9716 16808
rect 9658 16420 9670 16796
rect 9704 16420 9716 16796
rect 9658 16408 9716 16420
rect 9776 16796 9834 16808
rect 9776 16420 9788 16796
rect 9822 16420 9834 16796
rect 9776 16408 9834 16420
rect 9894 16796 9952 16808
rect 9894 16420 9906 16796
rect 9940 16420 9952 16796
rect 9894 16408 9952 16420
rect 10354 16794 10412 16806
rect 10354 16418 10366 16794
rect 10400 16418 10412 16794
rect 6769 16007 6827 16019
rect 6769 15831 6781 16007
rect 6815 15831 6827 16007
rect 6769 15819 6827 15831
rect 6887 16007 6945 16019
rect 6887 15831 6899 16007
rect 6933 15831 6945 16007
rect 6887 15819 6945 15831
rect 7005 16007 7063 16019
rect 7005 15831 7017 16007
rect 7051 15831 7063 16007
rect 7005 15819 7063 15831
rect 7123 16007 7181 16019
rect 7123 15831 7135 16007
rect 7169 15831 7181 16007
rect 7123 15819 7181 15831
rect 10354 16406 10412 16418
rect 10472 16794 10530 16806
rect 10472 16418 10484 16794
rect 10518 16418 10530 16794
rect 10472 16406 10530 16418
rect 10590 16794 10648 16806
rect 10590 16418 10602 16794
rect 10636 16418 10648 16794
rect 10590 16406 10648 16418
rect 10708 16794 10766 16806
rect 10708 16418 10720 16794
rect 10754 16418 10766 16794
rect 10708 16406 10766 16418
rect 10826 16794 10884 16806
rect 10826 16418 10838 16794
rect 10872 16418 10884 16794
rect 10826 16406 10884 16418
rect 10944 16794 11002 16806
rect 10944 16418 10956 16794
rect 10990 16418 11002 16794
rect 10944 16406 11002 16418
rect 11062 16794 11120 16806
rect 11062 16418 11074 16794
rect 11108 16418 11120 16794
rect 11062 16406 11120 16418
rect 11522 16796 11580 16808
rect 11522 16420 11534 16796
rect 11568 16420 11580 16796
rect 11522 16408 11580 16420
rect 11640 16796 11698 16808
rect 11640 16420 11652 16796
rect 11686 16420 11698 16796
rect 11640 16408 11698 16420
rect 11758 16796 11816 16808
rect 11758 16420 11770 16796
rect 11804 16420 11816 16796
rect 11758 16408 11816 16420
rect 11876 16796 11934 16808
rect 11876 16420 11888 16796
rect 11922 16420 11934 16796
rect 11876 16408 11934 16420
rect 11994 16796 12052 16808
rect 11994 16420 12006 16796
rect 12040 16420 12052 16796
rect 11994 16408 12052 16420
rect 12112 16796 12170 16808
rect 12112 16420 12124 16796
rect 12158 16420 12170 16796
rect 12112 16408 12170 16420
rect 12230 16796 12288 16808
rect 12230 16420 12242 16796
rect 12276 16420 12288 16796
rect 12230 16408 12288 16420
rect 12690 16796 12748 16808
rect 12690 16420 12702 16796
rect 12736 16420 12748 16796
rect 12690 16408 12748 16420
rect 12808 16796 12866 16808
rect 12808 16420 12820 16796
rect 12854 16420 12866 16796
rect 12808 16408 12866 16420
rect 12926 16796 12984 16808
rect 12926 16420 12938 16796
rect 12972 16420 12984 16796
rect 12926 16408 12984 16420
rect 13044 16796 13102 16808
rect 13044 16420 13056 16796
rect 13090 16420 13102 16796
rect 13044 16408 13102 16420
rect 13162 16796 13220 16808
rect 13162 16420 13174 16796
rect 13208 16420 13220 16796
rect 13162 16408 13220 16420
rect 13280 16796 13338 16808
rect 13280 16420 13292 16796
rect 13326 16420 13338 16796
rect 13280 16408 13338 16420
rect 13398 16796 13456 16808
rect 13398 16420 13410 16796
rect 13444 16420 13456 16796
rect 39206 16846 39264 16858
rect 13398 16408 13456 16420
rect 13791 16601 13849 16613
rect 13791 16425 13803 16601
rect 13837 16425 13849 16601
rect 13791 16413 13849 16425
rect 13909 16601 13967 16613
rect 13909 16425 13921 16601
rect 13955 16425 13967 16601
rect 13909 16413 13967 16425
rect 14027 16601 14085 16613
rect 14027 16425 14039 16601
rect 14073 16425 14085 16601
rect 14027 16413 14085 16425
rect 14145 16601 14203 16613
rect 14145 16425 14157 16601
rect 14191 16425 14203 16601
rect 14145 16413 14203 16425
rect 14263 16601 14321 16613
rect 14263 16425 14275 16601
rect 14309 16425 14321 16601
rect 14263 16413 14321 16425
rect 14381 16601 14439 16613
rect 14381 16425 14393 16601
rect 14427 16425 14439 16601
rect 14381 16413 14439 16425
rect 14499 16601 14557 16613
rect 14499 16425 14511 16601
rect 14545 16425 14557 16601
rect 14499 16413 14557 16425
rect 14617 16601 14675 16613
rect 14617 16425 14629 16601
rect 14663 16425 14675 16601
rect 14617 16413 14675 16425
rect 14735 16601 14793 16613
rect 14735 16425 14747 16601
rect 14781 16425 14793 16601
rect 14735 16413 14793 16425
rect 14853 16601 14911 16613
rect 14853 16425 14865 16601
rect 14899 16425 14911 16601
rect 14853 16413 14911 16425
rect 15239 16601 15297 16613
rect 15239 16425 15251 16601
rect 15285 16425 15297 16601
rect 15239 16413 15297 16425
rect 15357 16601 15415 16613
rect 15357 16425 15369 16601
rect 15403 16425 15415 16601
rect 15357 16413 15415 16425
rect 15475 16601 15533 16613
rect 15475 16425 15487 16601
rect 15521 16425 15533 16601
rect 15475 16413 15533 16425
rect 15593 16601 15651 16613
rect 15593 16425 15605 16601
rect 15639 16425 15651 16601
rect 15593 16413 15651 16425
rect 15711 16601 15769 16613
rect 15711 16425 15723 16601
rect 15757 16425 15769 16601
rect 15711 16413 15769 16425
rect 15829 16601 15887 16613
rect 15829 16425 15841 16601
rect 15875 16425 15887 16601
rect 15829 16413 15887 16425
rect 15947 16601 16005 16613
rect 15947 16425 15959 16601
rect 15993 16425 16005 16601
rect 15947 16413 16005 16425
rect 16065 16601 16123 16613
rect 16065 16425 16077 16601
rect 16111 16425 16123 16601
rect 16065 16413 16123 16425
rect 16183 16601 16241 16613
rect 16183 16425 16195 16601
rect 16229 16425 16241 16601
rect 16183 16413 16241 16425
rect 16301 16601 16359 16613
rect 16301 16425 16313 16601
rect 16347 16425 16359 16601
rect 16301 16413 16359 16425
rect 16737 16599 16795 16611
rect 16737 16423 16749 16599
rect 16783 16423 16795 16599
rect 7938 16008 7996 16020
rect 7938 15832 7950 16008
rect 7984 15832 7996 16008
rect 7938 15820 7996 15832
rect 8056 16008 8114 16020
rect 8056 15832 8068 16008
rect 8102 15832 8114 16008
rect 8056 15820 8114 15832
rect 8174 16008 8232 16020
rect 8174 15832 8186 16008
rect 8220 15832 8232 16008
rect 8174 15820 8232 15832
rect 8292 16008 8350 16020
rect 8292 15832 8304 16008
rect 8338 15832 8350 16008
rect 8292 15820 8350 15832
rect 9110 16012 9168 16024
rect 9110 15836 9122 16012
rect 9156 15836 9168 16012
rect 9110 15824 9168 15836
rect 9228 16012 9286 16024
rect 9228 15836 9240 16012
rect 9274 15836 9286 16012
rect 9228 15824 9286 15836
rect 9346 16012 9404 16024
rect 9346 15836 9358 16012
rect 9392 15836 9404 16012
rect 9346 15824 9404 15836
rect 9464 16012 9522 16024
rect 9464 15836 9476 16012
rect 9510 15836 9522 16012
rect 9464 15824 9522 15836
rect 10279 16012 10337 16024
rect 10279 15836 10291 16012
rect 10325 15836 10337 16012
rect 10279 15824 10337 15836
rect 10397 16012 10455 16024
rect 10397 15836 10409 16012
rect 10443 15836 10455 16012
rect 10397 15824 10455 15836
rect 10515 16012 10573 16024
rect 10515 15836 10527 16012
rect 10561 15836 10573 16012
rect 10515 15824 10573 15836
rect 10633 16012 10691 16024
rect 10633 15836 10645 16012
rect 10679 15836 10691 16012
rect 10633 15824 10691 15836
rect 11447 16012 11505 16024
rect 11447 15836 11459 16012
rect 11493 15836 11505 16012
rect 11447 15824 11505 15836
rect 11565 16012 11623 16024
rect 11565 15836 11577 16012
rect 11611 15836 11623 16012
rect 11565 15824 11623 15836
rect 11683 16012 11741 16024
rect 11683 15836 11695 16012
rect 11729 15836 11741 16012
rect 11683 15824 11741 15836
rect 11801 16012 11859 16024
rect 11801 15836 11813 16012
rect 11847 15836 11859 16012
rect 11801 15824 11859 15836
rect 16737 16411 16795 16423
rect 16855 16599 16913 16611
rect 16855 16423 16867 16599
rect 16901 16423 16913 16599
rect 16855 16411 16913 16423
rect 16973 16599 17031 16611
rect 16973 16423 16985 16599
rect 17019 16423 17031 16599
rect 16973 16411 17031 16423
rect 17091 16599 17149 16611
rect 17091 16423 17103 16599
rect 17137 16423 17149 16599
rect 17091 16411 17149 16423
rect 17209 16599 17267 16611
rect 17209 16423 17221 16599
rect 17255 16423 17267 16599
rect 17209 16411 17267 16423
rect 17327 16599 17385 16611
rect 17327 16423 17339 16599
rect 17373 16423 17385 16599
rect 17327 16411 17385 16423
rect 17445 16599 17503 16611
rect 17445 16423 17457 16599
rect 17491 16423 17503 16599
rect 17445 16411 17503 16423
rect 17563 16599 17621 16611
rect 17563 16423 17575 16599
rect 17609 16423 17621 16599
rect 17563 16411 17621 16423
rect 17681 16599 17739 16611
rect 17681 16423 17693 16599
rect 17727 16423 17739 16599
rect 17681 16411 17739 16423
rect 17799 16599 17857 16611
rect 17799 16423 17811 16599
rect 17845 16423 17857 16599
rect 17799 16411 17857 16423
rect 18185 16599 18243 16611
rect 18185 16423 18197 16599
rect 18231 16423 18243 16599
rect 18185 16411 18243 16423
rect 18303 16599 18361 16611
rect 18303 16423 18315 16599
rect 18349 16423 18361 16599
rect 18303 16411 18361 16423
rect 18421 16599 18479 16611
rect 18421 16423 18433 16599
rect 18467 16423 18479 16599
rect 18421 16411 18479 16423
rect 18539 16599 18597 16611
rect 18539 16423 18551 16599
rect 18585 16423 18597 16599
rect 18539 16411 18597 16423
rect 18657 16599 18715 16611
rect 18657 16423 18669 16599
rect 18703 16423 18715 16599
rect 18657 16411 18715 16423
rect 18775 16599 18833 16611
rect 18775 16423 18787 16599
rect 18821 16423 18833 16599
rect 18775 16411 18833 16423
rect 18893 16599 18951 16611
rect 18893 16423 18905 16599
rect 18939 16423 18951 16599
rect 18893 16411 18951 16423
rect 19011 16599 19069 16611
rect 19011 16423 19023 16599
rect 19057 16423 19069 16599
rect 19011 16411 19069 16423
rect 19129 16599 19187 16611
rect 19129 16423 19141 16599
rect 19175 16423 19187 16599
rect 19129 16411 19187 16423
rect 19247 16599 19305 16611
rect 19247 16423 19259 16599
rect 19293 16423 19305 16599
rect 19247 16411 19305 16423
rect 19705 16601 19763 16613
rect 19705 16425 19717 16601
rect 19751 16425 19763 16601
rect 19705 16413 19763 16425
rect 19823 16601 19881 16613
rect 19823 16425 19835 16601
rect 19869 16425 19881 16601
rect 19823 16413 19881 16425
rect 19941 16601 19999 16613
rect 19941 16425 19953 16601
rect 19987 16425 19999 16601
rect 19941 16413 19999 16425
rect 20059 16601 20117 16613
rect 20059 16425 20071 16601
rect 20105 16425 20117 16601
rect 20059 16413 20117 16425
rect 20177 16601 20235 16613
rect 20177 16425 20189 16601
rect 20223 16425 20235 16601
rect 20177 16413 20235 16425
rect 20295 16601 20353 16613
rect 20295 16425 20307 16601
rect 20341 16425 20353 16601
rect 20295 16413 20353 16425
rect 20413 16601 20471 16613
rect 20413 16425 20425 16601
rect 20459 16425 20471 16601
rect 20413 16413 20471 16425
rect 20531 16601 20589 16613
rect 20531 16425 20543 16601
rect 20577 16425 20589 16601
rect 20531 16413 20589 16425
rect 20649 16601 20707 16613
rect 20649 16425 20661 16601
rect 20695 16425 20707 16601
rect 20649 16413 20707 16425
rect 20767 16601 20825 16613
rect 20767 16425 20779 16601
rect 20813 16425 20825 16601
rect 20767 16413 20825 16425
rect 21153 16601 21211 16613
rect 21153 16425 21165 16601
rect 21199 16425 21211 16601
rect 21153 16413 21211 16425
rect 21271 16601 21329 16613
rect 21271 16425 21283 16601
rect 21317 16425 21329 16601
rect 21271 16413 21329 16425
rect 21389 16601 21447 16613
rect 21389 16425 21401 16601
rect 21435 16425 21447 16601
rect 21389 16413 21447 16425
rect 21507 16601 21565 16613
rect 21507 16425 21519 16601
rect 21553 16425 21565 16601
rect 21507 16413 21565 16425
rect 21625 16601 21683 16613
rect 21625 16425 21637 16601
rect 21671 16425 21683 16601
rect 21625 16413 21683 16425
rect 21743 16601 21801 16613
rect 21743 16425 21755 16601
rect 21789 16425 21801 16601
rect 21743 16413 21801 16425
rect 21861 16601 21919 16613
rect 21861 16425 21873 16601
rect 21907 16425 21919 16601
rect 21861 16413 21919 16425
rect 21979 16601 22037 16613
rect 21979 16425 21991 16601
rect 22025 16425 22037 16601
rect 21979 16413 22037 16425
rect 22097 16601 22155 16613
rect 22097 16425 22109 16601
rect 22143 16425 22155 16601
rect 22097 16413 22155 16425
rect 22215 16601 22273 16613
rect 38723 16646 38781 16658
rect 22215 16425 22227 16601
rect 22261 16425 22273 16601
rect 22215 16413 22273 16425
rect 22651 16599 22709 16611
rect 22651 16423 22663 16599
rect 22697 16423 22709 16599
rect 12614 16006 12672 16018
rect 12614 15830 12626 16006
rect 12660 15830 12672 16006
rect 12614 15818 12672 15830
rect 12732 16006 12790 16018
rect 12732 15830 12744 16006
rect 12778 15830 12790 16006
rect 12732 15818 12790 15830
rect 12850 16006 12908 16018
rect 12850 15830 12862 16006
rect 12896 15830 12908 16006
rect 12850 15818 12908 15830
rect 12968 16006 13026 16018
rect 12968 15830 12980 16006
rect 13014 15830 13026 16006
rect 12968 15818 13026 15830
rect 22651 16411 22709 16423
rect 22769 16599 22827 16611
rect 22769 16423 22781 16599
rect 22815 16423 22827 16599
rect 22769 16411 22827 16423
rect 22887 16599 22945 16611
rect 22887 16423 22899 16599
rect 22933 16423 22945 16599
rect 22887 16411 22945 16423
rect 23005 16599 23063 16611
rect 23005 16423 23017 16599
rect 23051 16423 23063 16599
rect 23005 16411 23063 16423
rect 23123 16599 23181 16611
rect 23123 16423 23135 16599
rect 23169 16423 23181 16599
rect 23123 16411 23181 16423
rect 23241 16599 23299 16611
rect 23241 16423 23253 16599
rect 23287 16423 23299 16599
rect 23241 16411 23299 16423
rect 23359 16599 23417 16611
rect 23359 16423 23371 16599
rect 23405 16423 23417 16599
rect 23359 16411 23417 16423
rect 23477 16599 23535 16611
rect 23477 16423 23489 16599
rect 23523 16423 23535 16599
rect 23477 16411 23535 16423
rect 23595 16599 23653 16611
rect 23595 16423 23607 16599
rect 23641 16423 23653 16599
rect 23595 16411 23653 16423
rect 23713 16599 23771 16611
rect 23713 16423 23725 16599
rect 23759 16423 23771 16599
rect 23713 16411 23771 16423
rect 24099 16599 24157 16611
rect 24099 16423 24111 16599
rect 24145 16423 24157 16599
rect 24099 16411 24157 16423
rect 24217 16599 24275 16611
rect 24217 16423 24229 16599
rect 24263 16423 24275 16599
rect 24217 16411 24275 16423
rect 24335 16599 24393 16611
rect 24335 16423 24347 16599
rect 24381 16423 24393 16599
rect 24335 16411 24393 16423
rect 24453 16599 24511 16611
rect 24453 16423 24465 16599
rect 24499 16423 24511 16599
rect 24453 16411 24511 16423
rect 24571 16599 24629 16611
rect 24571 16423 24583 16599
rect 24617 16423 24629 16599
rect 24571 16411 24629 16423
rect 24689 16599 24747 16611
rect 24689 16423 24701 16599
rect 24735 16423 24747 16599
rect 24689 16411 24747 16423
rect 24807 16599 24865 16611
rect 24807 16423 24819 16599
rect 24853 16423 24865 16599
rect 24807 16411 24865 16423
rect 24925 16599 24983 16611
rect 24925 16423 24937 16599
rect 24971 16423 24983 16599
rect 24925 16411 24983 16423
rect 25043 16599 25101 16611
rect 25043 16423 25055 16599
rect 25089 16423 25101 16599
rect 25043 16411 25101 16423
rect 25161 16599 25219 16611
rect 25161 16423 25173 16599
rect 25207 16423 25219 16599
rect 38723 16470 38735 16646
rect 38769 16470 38781 16646
rect 38723 16458 38781 16470
rect 38841 16646 38899 16658
rect 38841 16470 38853 16646
rect 38887 16470 38899 16646
rect 38841 16458 38899 16470
rect 38959 16646 39017 16658
rect 38959 16470 38971 16646
rect 39005 16470 39017 16646
rect 38959 16458 39017 16470
rect 39077 16646 39135 16658
rect 39077 16470 39089 16646
rect 39123 16470 39135 16646
rect 39077 16458 39135 16470
rect 39206 16470 39218 16846
rect 39252 16470 39264 16846
rect 39206 16458 39264 16470
rect 39324 16846 39382 16858
rect 39324 16470 39336 16846
rect 39370 16470 39382 16846
rect 39324 16458 39382 16470
rect 39442 16846 39500 16858
rect 39442 16470 39454 16846
rect 39488 16470 39500 16846
rect 39442 16458 39500 16470
rect 39560 16846 39618 16858
rect 39560 16470 39572 16846
rect 39606 16470 39618 16846
rect 39560 16458 39618 16470
rect 39678 16846 39736 16858
rect 39678 16470 39690 16846
rect 39724 16470 39736 16846
rect 39678 16458 39736 16470
rect 39796 16846 39854 16858
rect 39796 16470 39808 16846
rect 39842 16470 39854 16846
rect 39796 16458 39854 16470
rect 39914 16846 39972 16858
rect 39914 16470 39926 16846
rect 39960 16470 39972 16846
rect 41104 16846 41162 16858
rect 39914 16458 39972 16470
rect 40044 16646 40102 16658
rect 40044 16470 40056 16646
rect 40090 16470 40102 16646
rect 40044 16458 40102 16470
rect 40162 16646 40220 16658
rect 40162 16470 40174 16646
rect 40208 16470 40220 16646
rect 40162 16458 40220 16470
rect 40280 16646 40338 16658
rect 40280 16470 40292 16646
rect 40326 16470 40338 16646
rect 40280 16458 40338 16470
rect 40398 16646 40456 16658
rect 40398 16470 40410 16646
rect 40444 16470 40456 16646
rect 40398 16458 40456 16470
rect 40621 16646 40679 16658
rect 40621 16470 40633 16646
rect 40667 16470 40679 16646
rect 40621 16458 40679 16470
rect 40739 16646 40797 16658
rect 40739 16470 40751 16646
rect 40785 16470 40797 16646
rect 40739 16458 40797 16470
rect 40857 16646 40915 16658
rect 40857 16470 40869 16646
rect 40903 16470 40915 16646
rect 40857 16458 40915 16470
rect 40975 16646 41033 16658
rect 40975 16470 40987 16646
rect 41021 16470 41033 16646
rect 40975 16458 41033 16470
rect 41104 16470 41116 16846
rect 41150 16470 41162 16846
rect 41104 16458 41162 16470
rect 41222 16846 41280 16858
rect 41222 16470 41234 16846
rect 41268 16470 41280 16846
rect 41222 16458 41280 16470
rect 41340 16846 41398 16858
rect 41340 16470 41352 16846
rect 41386 16470 41398 16846
rect 41340 16458 41398 16470
rect 41458 16846 41516 16858
rect 41458 16470 41470 16846
rect 41504 16470 41516 16846
rect 41458 16458 41516 16470
rect 41576 16846 41634 16858
rect 41576 16470 41588 16846
rect 41622 16470 41634 16846
rect 41576 16458 41634 16470
rect 41694 16846 41752 16858
rect 41694 16470 41706 16846
rect 41740 16470 41752 16846
rect 41694 16458 41752 16470
rect 41812 16846 41870 16858
rect 41812 16470 41824 16846
rect 41858 16470 41870 16846
rect 45764 16842 45822 16854
rect 41812 16458 41870 16470
rect 41942 16646 42000 16658
rect 41942 16470 41954 16646
rect 41988 16470 42000 16646
rect 41942 16458 42000 16470
rect 42060 16646 42118 16658
rect 42060 16470 42072 16646
rect 42106 16470 42118 16646
rect 42060 16458 42118 16470
rect 42178 16646 42236 16658
rect 42178 16470 42190 16646
rect 42224 16470 42236 16646
rect 42178 16458 42236 16470
rect 42296 16646 42354 16658
rect 42296 16470 42308 16646
rect 42342 16470 42354 16646
rect 42296 16458 42354 16470
rect 25161 16411 25219 16423
rect 39263 16153 39321 16165
rect 39263 15777 39275 16153
rect 39309 15777 39321 16153
rect 39263 15765 39321 15777
rect 39381 16153 39439 16165
rect 39381 15777 39393 16153
rect 39427 15777 39439 16153
rect 39381 15765 39439 15777
rect 39499 16153 39557 16165
rect 39499 15777 39511 16153
rect 39545 15777 39557 16153
rect 39499 15765 39557 15777
rect 39617 16153 39675 16165
rect 39617 15777 39629 16153
rect 39663 15777 39675 16153
rect 39617 15765 39675 15777
rect 39735 16153 39793 16165
rect 39735 15777 39747 16153
rect 39781 15777 39793 16153
rect 39735 15765 39793 15777
rect 39853 16153 39911 16165
rect 39853 15777 39865 16153
rect 39899 15777 39911 16153
rect 39853 15765 39911 15777
rect 39971 16153 40029 16165
rect 39971 15777 39983 16153
rect 40017 15777 40029 16153
rect 39971 15765 40029 15777
rect 45281 16642 45339 16654
rect 45281 16466 45293 16642
rect 45327 16466 45339 16642
rect 45281 16454 45339 16466
rect 45399 16642 45457 16654
rect 45399 16466 45411 16642
rect 45445 16466 45457 16642
rect 45399 16454 45457 16466
rect 45517 16642 45575 16654
rect 45517 16466 45529 16642
rect 45563 16466 45575 16642
rect 45517 16454 45575 16466
rect 45635 16642 45693 16654
rect 45635 16466 45647 16642
rect 45681 16466 45693 16642
rect 45635 16454 45693 16466
rect 45764 16466 45776 16842
rect 45810 16466 45822 16842
rect 45764 16454 45822 16466
rect 45882 16842 45940 16854
rect 45882 16466 45894 16842
rect 45928 16466 45940 16842
rect 45882 16454 45940 16466
rect 46000 16842 46058 16854
rect 46000 16466 46012 16842
rect 46046 16466 46058 16842
rect 46000 16454 46058 16466
rect 46118 16842 46176 16854
rect 46118 16466 46130 16842
rect 46164 16466 46176 16842
rect 46118 16454 46176 16466
rect 46236 16842 46294 16854
rect 46236 16466 46248 16842
rect 46282 16466 46294 16842
rect 46236 16454 46294 16466
rect 46354 16842 46412 16854
rect 46354 16466 46366 16842
rect 46400 16466 46412 16842
rect 46354 16454 46412 16466
rect 46472 16842 46530 16854
rect 46472 16466 46484 16842
rect 46518 16466 46530 16842
rect 47662 16842 47720 16854
rect 46472 16454 46530 16466
rect 46602 16642 46660 16654
rect 46602 16466 46614 16642
rect 46648 16466 46660 16642
rect 46602 16454 46660 16466
rect 46720 16642 46778 16654
rect 46720 16466 46732 16642
rect 46766 16466 46778 16642
rect 46720 16454 46778 16466
rect 46838 16642 46896 16654
rect 46838 16466 46850 16642
rect 46884 16466 46896 16642
rect 46838 16454 46896 16466
rect 46956 16642 47014 16654
rect 46956 16466 46968 16642
rect 47002 16466 47014 16642
rect 46956 16454 47014 16466
rect 47179 16642 47237 16654
rect 47179 16466 47191 16642
rect 47225 16466 47237 16642
rect 47179 16454 47237 16466
rect 47297 16642 47355 16654
rect 47297 16466 47309 16642
rect 47343 16466 47355 16642
rect 47297 16454 47355 16466
rect 47415 16642 47473 16654
rect 47415 16466 47427 16642
rect 47461 16466 47473 16642
rect 47415 16454 47473 16466
rect 47533 16642 47591 16654
rect 47533 16466 47545 16642
rect 47579 16466 47591 16642
rect 47533 16454 47591 16466
rect 47662 16466 47674 16842
rect 47708 16466 47720 16842
rect 47662 16454 47720 16466
rect 47780 16842 47838 16854
rect 47780 16466 47792 16842
rect 47826 16466 47838 16842
rect 47780 16454 47838 16466
rect 47898 16842 47956 16854
rect 47898 16466 47910 16842
rect 47944 16466 47956 16842
rect 47898 16454 47956 16466
rect 48016 16842 48074 16854
rect 48016 16466 48028 16842
rect 48062 16466 48074 16842
rect 48016 16454 48074 16466
rect 48134 16842 48192 16854
rect 48134 16466 48146 16842
rect 48180 16466 48192 16842
rect 48134 16454 48192 16466
rect 48252 16842 48310 16854
rect 48252 16466 48264 16842
rect 48298 16466 48310 16842
rect 48252 16454 48310 16466
rect 48370 16842 48428 16854
rect 48370 16466 48382 16842
rect 48416 16466 48428 16842
rect 52298 16847 52356 16859
rect 48370 16454 48428 16466
rect 48500 16642 48558 16654
rect 48500 16466 48512 16642
rect 48546 16466 48558 16642
rect 48500 16454 48558 16466
rect 48618 16642 48676 16654
rect 48618 16466 48630 16642
rect 48664 16466 48676 16642
rect 48618 16454 48676 16466
rect 48736 16642 48794 16654
rect 48736 16466 48748 16642
rect 48782 16466 48794 16642
rect 48736 16454 48794 16466
rect 48854 16642 48912 16654
rect 48854 16466 48866 16642
rect 48900 16466 48912 16642
rect 48854 16454 48912 16466
rect 41161 16153 41219 16165
rect 41161 15777 41173 16153
rect 41207 15777 41219 16153
rect 41161 15765 41219 15777
rect 41279 16153 41337 16165
rect 41279 15777 41291 16153
rect 41325 15777 41337 16153
rect 41279 15765 41337 15777
rect 41397 16153 41455 16165
rect 41397 15777 41409 16153
rect 41443 15777 41455 16153
rect 41397 15765 41455 15777
rect 41515 16153 41573 16165
rect 41515 15777 41527 16153
rect 41561 15777 41573 16153
rect 41515 15765 41573 15777
rect 41633 16153 41691 16165
rect 41633 15777 41645 16153
rect 41679 15777 41691 16153
rect 41633 15765 41691 15777
rect 41751 16153 41809 16165
rect 41751 15777 41763 16153
rect 41797 15777 41809 16153
rect 41751 15765 41809 15777
rect 41869 16153 41927 16165
rect 41869 15777 41881 16153
rect 41915 15777 41927 16153
rect 41869 15765 41927 15777
rect 42703 15659 42761 15671
rect 42703 15483 42715 15659
rect 42749 15483 42761 15659
rect 42703 15471 42761 15483
rect 42821 15659 42879 15671
rect 42821 15483 42833 15659
rect 42867 15483 42879 15659
rect 42821 15471 42879 15483
rect 42939 15659 42997 15671
rect 42939 15483 42951 15659
rect 42985 15483 42997 15659
rect 42939 15471 42997 15483
rect 43057 15659 43115 15671
rect 43057 15483 43069 15659
rect 43103 15483 43115 15659
rect 43057 15471 43115 15483
rect 43175 15659 43233 15671
rect 43175 15483 43187 15659
rect 43221 15483 43233 15659
rect 43175 15471 43233 15483
rect 43293 15659 43351 15671
rect 43293 15483 43305 15659
rect 43339 15483 43351 15659
rect 43293 15471 43351 15483
rect 43411 15659 43469 15671
rect 43411 15483 43423 15659
rect 43457 15483 43469 15659
rect 43411 15471 43469 15483
rect 43529 15659 43587 15671
rect 43529 15483 43541 15659
rect 43575 15483 43587 15659
rect 43529 15471 43587 15483
rect 43647 15659 43705 15671
rect 43647 15483 43659 15659
rect 43693 15483 43705 15659
rect 43647 15471 43705 15483
rect 43765 15659 43823 15671
rect 43765 15483 43777 15659
rect 43811 15483 43823 15659
rect 43765 15471 43823 15483
rect 45821 16149 45879 16161
rect 45821 15773 45833 16149
rect 45867 15773 45879 16149
rect 45821 15761 45879 15773
rect 45939 16149 45997 16161
rect 45939 15773 45951 16149
rect 45985 15773 45997 16149
rect 45939 15761 45997 15773
rect 46057 16149 46115 16161
rect 46057 15773 46069 16149
rect 46103 15773 46115 16149
rect 46057 15761 46115 15773
rect 46175 16149 46233 16161
rect 46175 15773 46187 16149
rect 46221 15773 46233 16149
rect 46175 15761 46233 15773
rect 46293 16149 46351 16161
rect 46293 15773 46305 16149
rect 46339 15773 46351 16149
rect 46293 15761 46351 15773
rect 46411 16149 46469 16161
rect 46411 15773 46423 16149
rect 46457 15773 46469 16149
rect 46411 15761 46469 15773
rect 46529 16149 46587 16161
rect 46529 15773 46541 16149
rect 46575 15773 46587 16149
rect 46529 15761 46587 15773
rect 51815 16647 51873 16659
rect 51815 16471 51827 16647
rect 51861 16471 51873 16647
rect 51815 16459 51873 16471
rect 51933 16647 51991 16659
rect 51933 16471 51945 16647
rect 51979 16471 51991 16647
rect 51933 16459 51991 16471
rect 52051 16647 52109 16659
rect 52051 16471 52063 16647
rect 52097 16471 52109 16647
rect 52051 16459 52109 16471
rect 52169 16647 52227 16659
rect 52169 16471 52181 16647
rect 52215 16471 52227 16647
rect 52169 16459 52227 16471
rect 52298 16471 52310 16847
rect 52344 16471 52356 16847
rect 52298 16459 52356 16471
rect 52416 16847 52474 16859
rect 52416 16471 52428 16847
rect 52462 16471 52474 16847
rect 52416 16459 52474 16471
rect 52534 16847 52592 16859
rect 52534 16471 52546 16847
rect 52580 16471 52592 16847
rect 52534 16459 52592 16471
rect 52652 16847 52710 16859
rect 52652 16471 52664 16847
rect 52698 16471 52710 16847
rect 52652 16459 52710 16471
rect 52770 16847 52828 16859
rect 52770 16471 52782 16847
rect 52816 16471 52828 16847
rect 52770 16459 52828 16471
rect 52888 16847 52946 16859
rect 52888 16471 52900 16847
rect 52934 16471 52946 16847
rect 52888 16459 52946 16471
rect 53006 16847 53064 16859
rect 53006 16471 53018 16847
rect 53052 16471 53064 16847
rect 54196 16847 54254 16859
rect 53006 16459 53064 16471
rect 53136 16647 53194 16659
rect 53136 16471 53148 16647
rect 53182 16471 53194 16647
rect 53136 16459 53194 16471
rect 53254 16647 53312 16659
rect 53254 16471 53266 16647
rect 53300 16471 53312 16647
rect 53254 16459 53312 16471
rect 53372 16647 53430 16659
rect 53372 16471 53384 16647
rect 53418 16471 53430 16647
rect 53372 16459 53430 16471
rect 53490 16647 53548 16659
rect 53490 16471 53502 16647
rect 53536 16471 53548 16647
rect 53490 16459 53548 16471
rect 53713 16647 53771 16659
rect 53713 16471 53725 16647
rect 53759 16471 53771 16647
rect 53713 16459 53771 16471
rect 53831 16647 53889 16659
rect 53831 16471 53843 16647
rect 53877 16471 53889 16647
rect 53831 16459 53889 16471
rect 53949 16647 54007 16659
rect 53949 16471 53961 16647
rect 53995 16471 54007 16647
rect 53949 16459 54007 16471
rect 54067 16647 54125 16659
rect 54067 16471 54079 16647
rect 54113 16471 54125 16647
rect 54067 16459 54125 16471
rect 54196 16471 54208 16847
rect 54242 16471 54254 16847
rect 54196 16459 54254 16471
rect 54314 16847 54372 16859
rect 54314 16471 54326 16847
rect 54360 16471 54372 16847
rect 54314 16459 54372 16471
rect 54432 16847 54490 16859
rect 54432 16471 54444 16847
rect 54478 16471 54490 16847
rect 54432 16459 54490 16471
rect 54550 16847 54608 16859
rect 54550 16471 54562 16847
rect 54596 16471 54608 16847
rect 54550 16459 54608 16471
rect 54668 16847 54726 16859
rect 54668 16471 54680 16847
rect 54714 16471 54726 16847
rect 54668 16459 54726 16471
rect 54786 16847 54844 16859
rect 54786 16471 54798 16847
rect 54832 16471 54844 16847
rect 54786 16459 54844 16471
rect 54904 16847 54962 16859
rect 54904 16471 54916 16847
rect 54950 16471 54962 16847
rect 58811 16850 58869 16862
rect 54904 16459 54962 16471
rect 55034 16647 55092 16659
rect 55034 16471 55046 16647
rect 55080 16471 55092 16647
rect 55034 16459 55092 16471
rect 55152 16647 55210 16659
rect 55152 16471 55164 16647
rect 55198 16471 55210 16647
rect 55152 16459 55210 16471
rect 55270 16647 55328 16659
rect 55270 16471 55282 16647
rect 55316 16471 55328 16647
rect 55270 16459 55328 16471
rect 55388 16647 55446 16659
rect 55388 16471 55400 16647
rect 55434 16471 55446 16647
rect 55388 16459 55446 16471
rect 47719 16149 47777 16161
rect 47719 15773 47731 16149
rect 47765 15773 47777 16149
rect 47719 15761 47777 15773
rect 47837 16149 47895 16161
rect 47837 15773 47849 16149
rect 47883 15773 47895 16149
rect 47837 15761 47895 15773
rect 47955 16149 48013 16161
rect 47955 15773 47967 16149
rect 48001 15773 48013 16149
rect 47955 15761 48013 15773
rect 48073 16149 48131 16161
rect 48073 15773 48085 16149
rect 48119 15773 48131 16149
rect 48073 15761 48131 15773
rect 48191 16149 48249 16161
rect 48191 15773 48203 16149
rect 48237 15773 48249 16149
rect 48191 15761 48249 15773
rect 48309 16149 48367 16161
rect 48309 15773 48321 16149
rect 48355 15773 48367 16149
rect 48309 15761 48367 15773
rect 48427 16149 48485 16161
rect 48427 15773 48439 16149
rect 48473 15773 48485 16149
rect 48427 15761 48485 15773
rect 49261 15655 49319 15667
rect 49261 15479 49273 15655
rect 49307 15479 49319 15655
rect 49261 15467 49319 15479
rect 49379 15655 49437 15667
rect 49379 15479 49391 15655
rect 49425 15479 49437 15655
rect 49379 15467 49437 15479
rect 49497 15655 49555 15667
rect 49497 15479 49509 15655
rect 49543 15479 49555 15655
rect 49497 15467 49555 15479
rect 49615 15655 49673 15667
rect 49615 15479 49627 15655
rect 49661 15479 49673 15655
rect 49615 15467 49673 15479
rect 49733 15655 49791 15667
rect 49733 15479 49745 15655
rect 49779 15479 49791 15655
rect 49733 15467 49791 15479
rect 49851 15655 49909 15667
rect 49851 15479 49863 15655
rect 49897 15479 49909 15655
rect 49851 15467 49909 15479
rect 49969 15655 50027 15667
rect 49969 15479 49981 15655
rect 50015 15479 50027 15655
rect 49969 15467 50027 15479
rect 50087 15655 50145 15667
rect 50087 15479 50099 15655
rect 50133 15479 50145 15655
rect 50087 15467 50145 15479
rect 50205 15655 50263 15667
rect 50205 15479 50217 15655
rect 50251 15479 50263 15655
rect 50205 15467 50263 15479
rect 50323 15655 50381 15667
rect 50323 15479 50335 15655
rect 50369 15479 50381 15655
rect 50323 15467 50381 15479
rect 52355 16154 52413 16166
rect 52355 15778 52367 16154
rect 52401 15778 52413 16154
rect 52355 15766 52413 15778
rect 52473 16154 52531 16166
rect 52473 15778 52485 16154
rect 52519 15778 52531 16154
rect 52473 15766 52531 15778
rect 52591 16154 52649 16166
rect 52591 15778 52603 16154
rect 52637 15778 52649 16154
rect 52591 15766 52649 15778
rect 52709 16154 52767 16166
rect 52709 15778 52721 16154
rect 52755 15778 52767 16154
rect 52709 15766 52767 15778
rect 52827 16154 52885 16166
rect 52827 15778 52839 16154
rect 52873 15778 52885 16154
rect 52827 15766 52885 15778
rect 52945 16154 53003 16166
rect 52945 15778 52957 16154
rect 52991 15778 53003 16154
rect 52945 15766 53003 15778
rect 53063 16154 53121 16166
rect 53063 15778 53075 16154
rect 53109 15778 53121 16154
rect 53063 15766 53121 15778
rect 971 14846 1029 14858
rect 498 14646 556 14658
rect 498 14470 510 14646
rect 544 14470 556 14646
rect 498 14458 556 14470
rect 616 14646 674 14658
rect 616 14470 628 14646
rect 662 14470 674 14646
rect 616 14458 674 14470
rect 734 14646 792 14658
rect 734 14470 746 14646
rect 780 14470 792 14646
rect 734 14458 792 14470
rect 852 14646 910 14658
rect 852 14470 864 14646
rect 898 14470 910 14646
rect 852 14458 910 14470
rect 971 14470 983 14846
rect 1017 14470 1029 14846
rect 971 14458 1029 14470
rect 1089 14846 1147 14858
rect 1089 14470 1101 14846
rect 1135 14470 1147 14846
rect 1089 14458 1147 14470
rect 1207 14846 1265 14858
rect 1207 14470 1219 14846
rect 1253 14470 1265 14846
rect 1207 14458 1265 14470
rect 1325 14846 1383 14858
rect 1325 14470 1337 14846
rect 1371 14470 1383 14846
rect 1325 14458 1383 14470
rect 1444 14846 1502 14858
rect 1444 14470 1456 14846
rect 1490 14470 1502 14846
rect 1444 14458 1502 14470
rect 1562 14846 1620 14858
rect 1562 14470 1574 14846
rect 1608 14470 1620 14846
rect 1562 14458 1620 14470
rect 1680 14846 1738 14858
rect 1680 14470 1692 14846
rect 1726 14470 1738 14846
rect 1680 14458 1738 14470
rect 1798 14846 1856 14858
rect 1798 14470 1810 14846
rect 1844 14470 1856 14846
rect 1798 14458 1856 14470
rect 1916 14846 1974 14858
rect 1916 14470 1928 14846
rect 1962 14470 1974 14846
rect 1916 14458 1974 14470
rect 2034 14846 2092 14858
rect 2034 14470 2046 14846
rect 2080 14470 2092 14846
rect 2034 14458 2092 14470
rect 2152 14846 2210 14858
rect 2152 14470 2164 14846
rect 2198 14470 2210 14846
rect 2152 14458 2210 14470
rect 2265 14846 2323 14858
rect 2265 14470 2277 14846
rect 2311 14470 2323 14846
rect 2265 14458 2323 14470
rect 2383 14846 2441 14858
rect 2383 14470 2395 14846
rect 2429 14470 2441 14846
rect 2383 14458 2441 14470
rect 2501 14846 2559 14858
rect 2501 14470 2513 14846
rect 2547 14470 2559 14846
rect 2501 14458 2559 14470
rect 2619 14846 2677 14858
rect 2619 14470 2631 14846
rect 2665 14658 2677 14846
rect 4115 14846 4173 14858
rect 2665 14646 2764 14658
rect 2665 14470 2718 14646
rect 2752 14470 2764 14646
rect 2619 14458 2764 14470
rect 2824 14646 2882 14658
rect 2824 14470 2836 14646
rect 2870 14470 2882 14646
rect 2824 14458 2882 14470
rect 2942 14646 3000 14658
rect 2942 14470 2954 14646
rect 2988 14470 3000 14646
rect 2942 14458 3000 14470
rect 3060 14646 3118 14658
rect 3060 14470 3072 14646
rect 3106 14470 3118 14646
rect 3060 14458 3118 14470
rect 3642 14646 3700 14658
rect 3642 14470 3654 14646
rect 3688 14470 3700 14646
rect 3642 14458 3700 14470
rect 3760 14646 3818 14658
rect 3760 14470 3772 14646
rect 3806 14470 3818 14646
rect 3760 14458 3818 14470
rect 3878 14646 3936 14658
rect 3878 14470 3890 14646
rect 3924 14470 3936 14646
rect 3878 14458 3936 14470
rect 3996 14646 4054 14658
rect 3996 14470 4008 14646
rect 4042 14470 4054 14646
rect 3996 14458 4054 14470
rect 4115 14470 4127 14846
rect 4161 14470 4173 14846
rect 4115 14458 4173 14470
rect 4233 14846 4291 14858
rect 4233 14470 4245 14846
rect 4279 14470 4291 14846
rect 4233 14458 4291 14470
rect 4351 14846 4409 14858
rect 4351 14470 4363 14846
rect 4397 14470 4409 14846
rect 4351 14458 4409 14470
rect 4469 14846 4527 14858
rect 4469 14470 4481 14846
rect 4515 14470 4527 14846
rect 4469 14458 4527 14470
rect 4588 14846 4646 14858
rect 4588 14470 4600 14846
rect 4634 14470 4646 14846
rect 4588 14458 4646 14470
rect 4706 14846 4764 14858
rect 4706 14470 4718 14846
rect 4752 14470 4764 14846
rect 4706 14458 4764 14470
rect 4824 14846 4882 14858
rect 4824 14470 4836 14846
rect 4870 14470 4882 14846
rect 4824 14458 4882 14470
rect 4942 14846 5000 14858
rect 4942 14470 4954 14846
rect 4988 14470 5000 14846
rect 4942 14458 5000 14470
rect 5060 14846 5118 14858
rect 5060 14470 5072 14846
rect 5106 14470 5118 14846
rect 5060 14458 5118 14470
rect 5178 14846 5236 14858
rect 5178 14470 5190 14846
rect 5224 14470 5236 14846
rect 5178 14458 5236 14470
rect 5296 14846 5354 14858
rect 5296 14470 5308 14846
rect 5342 14470 5354 14846
rect 5296 14458 5354 14470
rect 5409 14846 5467 14858
rect 5409 14470 5421 14846
rect 5455 14470 5467 14846
rect 5409 14458 5467 14470
rect 5527 14846 5585 14858
rect 5527 14470 5539 14846
rect 5573 14470 5585 14846
rect 5527 14458 5585 14470
rect 5645 14846 5703 14858
rect 5645 14470 5657 14846
rect 5691 14470 5703 14846
rect 5645 14458 5703 14470
rect 5763 14846 5821 14858
rect 5763 14470 5775 14846
rect 5809 14658 5821 14846
rect 7247 14842 7305 14854
rect 5809 14646 5908 14658
rect 5809 14470 5862 14646
rect 5896 14470 5908 14646
rect 5763 14458 5908 14470
rect 5968 14646 6026 14658
rect 5968 14470 5980 14646
rect 6014 14470 6026 14646
rect 5968 14458 6026 14470
rect 6086 14646 6144 14658
rect 6086 14470 6098 14646
rect 6132 14470 6144 14646
rect 6086 14458 6144 14470
rect 6204 14646 6262 14658
rect 6204 14470 6216 14646
rect 6250 14470 6262 14646
rect 6204 14458 6262 14470
rect 6774 14642 6832 14654
rect 6774 14466 6786 14642
rect 6820 14466 6832 14642
rect 6774 14454 6832 14466
rect 6892 14642 6950 14654
rect 6892 14466 6904 14642
rect 6938 14466 6950 14642
rect 6892 14454 6950 14466
rect 7010 14642 7068 14654
rect 7010 14466 7022 14642
rect 7056 14466 7068 14642
rect 7010 14454 7068 14466
rect 7128 14642 7186 14654
rect 7128 14466 7140 14642
rect 7174 14466 7186 14642
rect 7128 14454 7186 14466
rect 7247 14466 7259 14842
rect 7293 14466 7305 14842
rect 7247 14454 7305 14466
rect 7365 14842 7423 14854
rect 7365 14466 7377 14842
rect 7411 14466 7423 14842
rect 7365 14454 7423 14466
rect 7483 14842 7541 14854
rect 7483 14466 7495 14842
rect 7529 14466 7541 14842
rect 7483 14454 7541 14466
rect 7601 14842 7659 14854
rect 7601 14466 7613 14842
rect 7647 14466 7659 14842
rect 7601 14454 7659 14466
rect 7720 14842 7778 14854
rect 7720 14466 7732 14842
rect 7766 14466 7778 14842
rect 7720 14454 7778 14466
rect 7838 14842 7896 14854
rect 7838 14466 7850 14842
rect 7884 14466 7896 14842
rect 7838 14454 7896 14466
rect 7956 14842 8014 14854
rect 7956 14466 7968 14842
rect 8002 14466 8014 14842
rect 7956 14454 8014 14466
rect 8074 14842 8132 14854
rect 8074 14466 8086 14842
rect 8120 14466 8132 14842
rect 8074 14454 8132 14466
rect 8192 14842 8250 14854
rect 8192 14466 8204 14842
rect 8238 14466 8250 14842
rect 8192 14454 8250 14466
rect 8310 14842 8368 14854
rect 8310 14466 8322 14842
rect 8356 14466 8368 14842
rect 8310 14454 8368 14466
rect 8428 14842 8486 14854
rect 8428 14466 8440 14842
rect 8474 14466 8486 14842
rect 8428 14454 8486 14466
rect 8541 14842 8599 14854
rect 8541 14466 8553 14842
rect 8587 14466 8599 14842
rect 8541 14454 8599 14466
rect 8659 14842 8717 14854
rect 8659 14466 8671 14842
rect 8705 14466 8717 14842
rect 8659 14454 8717 14466
rect 8777 14842 8835 14854
rect 8777 14466 8789 14842
rect 8823 14466 8835 14842
rect 8777 14454 8835 14466
rect 8895 14842 8953 14854
rect 8895 14466 8907 14842
rect 8941 14654 8953 14842
rect 10391 14842 10449 14854
rect 8941 14642 9040 14654
rect 8941 14466 8994 14642
rect 9028 14466 9040 14642
rect 8895 14454 9040 14466
rect 9100 14642 9158 14654
rect 9100 14466 9112 14642
rect 9146 14466 9158 14642
rect 9100 14454 9158 14466
rect 9218 14642 9276 14654
rect 9218 14466 9230 14642
rect 9264 14466 9276 14642
rect 9218 14454 9276 14466
rect 9336 14642 9394 14654
rect 9336 14466 9348 14642
rect 9382 14466 9394 14642
rect 9336 14454 9394 14466
rect 9918 14642 9976 14654
rect 9918 14466 9930 14642
rect 9964 14466 9976 14642
rect 9918 14454 9976 14466
rect 10036 14642 10094 14654
rect 10036 14466 10048 14642
rect 10082 14466 10094 14642
rect 10036 14454 10094 14466
rect 10154 14642 10212 14654
rect 10154 14466 10166 14642
rect 10200 14466 10212 14642
rect 10154 14454 10212 14466
rect 10272 14642 10330 14654
rect 10272 14466 10284 14642
rect 10318 14466 10330 14642
rect 10272 14454 10330 14466
rect 10391 14466 10403 14842
rect 10437 14466 10449 14842
rect 10391 14454 10449 14466
rect 10509 14842 10567 14854
rect 10509 14466 10521 14842
rect 10555 14466 10567 14842
rect 10509 14454 10567 14466
rect 10627 14842 10685 14854
rect 10627 14466 10639 14842
rect 10673 14466 10685 14842
rect 10627 14454 10685 14466
rect 10745 14842 10803 14854
rect 10745 14466 10757 14842
rect 10791 14466 10803 14842
rect 10745 14454 10803 14466
rect 10864 14842 10922 14854
rect 10864 14466 10876 14842
rect 10910 14466 10922 14842
rect 10864 14454 10922 14466
rect 10982 14842 11040 14854
rect 10982 14466 10994 14842
rect 11028 14466 11040 14842
rect 10982 14454 11040 14466
rect 11100 14842 11158 14854
rect 11100 14466 11112 14842
rect 11146 14466 11158 14842
rect 11100 14454 11158 14466
rect 11218 14842 11276 14854
rect 11218 14466 11230 14842
rect 11264 14466 11276 14842
rect 11218 14454 11276 14466
rect 11336 14842 11394 14854
rect 11336 14466 11348 14842
rect 11382 14466 11394 14842
rect 11336 14454 11394 14466
rect 11454 14842 11512 14854
rect 11454 14466 11466 14842
rect 11500 14466 11512 14842
rect 11454 14454 11512 14466
rect 11572 14842 11630 14854
rect 11572 14466 11584 14842
rect 11618 14466 11630 14842
rect 11572 14454 11630 14466
rect 11685 14842 11743 14854
rect 11685 14466 11697 14842
rect 11731 14466 11743 14842
rect 11685 14454 11743 14466
rect 11803 14842 11861 14854
rect 11803 14466 11815 14842
rect 11849 14466 11861 14842
rect 11803 14454 11861 14466
rect 11921 14842 11979 14854
rect 11921 14466 11933 14842
rect 11967 14466 11979 14842
rect 11921 14454 11979 14466
rect 12039 14842 12097 14854
rect 12039 14466 12051 14842
rect 12085 14654 12097 14842
rect 13593 14846 13651 14858
rect 12085 14642 12184 14654
rect 12085 14466 12138 14642
rect 12172 14466 12184 14642
rect 12039 14454 12184 14466
rect 12244 14642 12302 14654
rect 12244 14466 12256 14642
rect 12290 14466 12302 14642
rect 12244 14454 12302 14466
rect 12362 14642 12420 14654
rect 12362 14466 12374 14642
rect 12408 14466 12420 14642
rect 12362 14454 12420 14466
rect 12480 14642 12538 14654
rect 12480 14466 12492 14642
rect 12526 14466 12538 14642
rect 12480 14454 12538 14466
rect 13120 14646 13178 14658
rect 13120 14470 13132 14646
rect 13166 14470 13178 14646
rect 13120 14458 13178 14470
rect 13238 14646 13296 14658
rect 13238 14470 13250 14646
rect 13284 14470 13296 14646
rect 13238 14458 13296 14470
rect 13356 14646 13414 14658
rect 13356 14470 13368 14646
rect 13402 14470 13414 14646
rect 13356 14458 13414 14470
rect 13474 14646 13532 14658
rect 13474 14470 13486 14646
rect 13520 14470 13532 14646
rect 13474 14458 13532 14470
rect 13593 14470 13605 14846
rect 13639 14470 13651 14846
rect 13593 14458 13651 14470
rect 13711 14846 13769 14858
rect 13711 14470 13723 14846
rect 13757 14470 13769 14846
rect 13711 14458 13769 14470
rect 13829 14846 13887 14858
rect 13829 14470 13841 14846
rect 13875 14470 13887 14846
rect 13829 14458 13887 14470
rect 13947 14846 14005 14858
rect 13947 14470 13959 14846
rect 13993 14470 14005 14846
rect 13947 14458 14005 14470
rect 14066 14846 14124 14858
rect 14066 14470 14078 14846
rect 14112 14470 14124 14846
rect 14066 14458 14124 14470
rect 14184 14846 14242 14858
rect 14184 14470 14196 14846
rect 14230 14470 14242 14846
rect 14184 14458 14242 14470
rect 14302 14846 14360 14858
rect 14302 14470 14314 14846
rect 14348 14470 14360 14846
rect 14302 14458 14360 14470
rect 14420 14846 14478 14858
rect 14420 14470 14432 14846
rect 14466 14470 14478 14846
rect 14420 14458 14478 14470
rect 14538 14846 14596 14858
rect 14538 14470 14550 14846
rect 14584 14470 14596 14846
rect 14538 14458 14596 14470
rect 14656 14846 14714 14858
rect 14656 14470 14668 14846
rect 14702 14470 14714 14846
rect 14656 14458 14714 14470
rect 14774 14846 14832 14858
rect 14774 14470 14786 14846
rect 14820 14470 14832 14846
rect 14774 14458 14832 14470
rect 14887 14846 14945 14858
rect 14887 14470 14899 14846
rect 14933 14470 14945 14846
rect 14887 14458 14945 14470
rect 15005 14846 15063 14858
rect 15005 14470 15017 14846
rect 15051 14470 15063 14846
rect 15005 14458 15063 14470
rect 15123 14846 15181 14858
rect 15123 14470 15135 14846
rect 15169 14470 15181 14846
rect 15123 14458 15181 14470
rect 15241 14846 15299 14858
rect 15241 14470 15253 14846
rect 15287 14658 15299 14846
rect 16737 14846 16795 14858
rect 15287 14646 15386 14658
rect 15287 14470 15340 14646
rect 15374 14470 15386 14646
rect 15241 14458 15386 14470
rect 15446 14646 15504 14658
rect 15446 14470 15458 14646
rect 15492 14470 15504 14646
rect 15446 14458 15504 14470
rect 15564 14646 15622 14658
rect 15564 14470 15576 14646
rect 15610 14470 15622 14646
rect 15564 14458 15622 14470
rect 15682 14646 15740 14658
rect 15682 14470 15694 14646
rect 15728 14470 15740 14646
rect 15682 14458 15740 14470
rect 16264 14646 16322 14658
rect 16264 14470 16276 14646
rect 16310 14470 16322 14646
rect 16264 14458 16322 14470
rect 16382 14646 16440 14658
rect 16382 14470 16394 14646
rect 16428 14470 16440 14646
rect 16382 14458 16440 14470
rect 16500 14646 16558 14658
rect 16500 14470 16512 14646
rect 16546 14470 16558 14646
rect 16500 14458 16558 14470
rect 16618 14646 16676 14658
rect 16618 14470 16630 14646
rect 16664 14470 16676 14646
rect 16618 14458 16676 14470
rect 16737 14470 16749 14846
rect 16783 14470 16795 14846
rect 16737 14458 16795 14470
rect 16855 14846 16913 14858
rect 16855 14470 16867 14846
rect 16901 14470 16913 14846
rect 16855 14458 16913 14470
rect 16973 14846 17031 14858
rect 16973 14470 16985 14846
rect 17019 14470 17031 14846
rect 16973 14458 17031 14470
rect 17091 14846 17149 14858
rect 17091 14470 17103 14846
rect 17137 14470 17149 14846
rect 17091 14458 17149 14470
rect 17210 14846 17268 14858
rect 17210 14470 17222 14846
rect 17256 14470 17268 14846
rect 17210 14458 17268 14470
rect 17328 14846 17386 14858
rect 17328 14470 17340 14846
rect 17374 14470 17386 14846
rect 17328 14458 17386 14470
rect 17446 14846 17504 14858
rect 17446 14470 17458 14846
rect 17492 14470 17504 14846
rect 17446 14458 17504 14470
rect 17564 14846 17622 14858
rect 17564 14470 17576 14846
rect 17610 14470 17622 14846
rect 17564 14458 17622 14470
rect 17682 14846 17740 14858
rect 17682 14470 17694 14846
rect 17728 14470 17740 14846
rect 17682 14458 17740 14470
rect 17800 14846 17858 14858
rect 17800 14470 17812 14846
rect 17846 14470 17858 14846
rect 17800 14458 17858 14470
rect 17918 14846 17976 14858
rect 17918 14470 17930 14846
rect 17964 14470 17976 14846
rect 17918 14458 17976 14470
rect 18031 14846 18089 14858
rect 18031 14470 18043 14846
rect 18077 14470 18089 14846
rect 18031 14458 18089 14470
rect 18149 14846 18207 14858
rect 18149 14470 18161 14846
rect 18195 14470 18207 14846
rect 18149 14458 18207 14470
rect 18267 14846 18325 14858
rect 18267 14470 18279 14846
rect 18313 14470 18325 14846
rect 18267 14458 18325 14470
rect 18385 14846 18443 14858
rect 18385 14470 18397 14846
rect 18431 14658 18443 14846
rect 19869 14842 19927 14854
rect 18431 14646 18530 14658
rect 18431 14470 18484 14646
rect 18518 14470 18530 14646
rect 18385 14458 18530 14470
rect 18590 14646 18648 14658
rect 18590 14470 18602 14646
rect 18636 14470 18648 14646
rect 18590 14458 18648 14470
rect 18708 14646 18766 14658
rect 18708 14470 18720 14646
rect 18754 14470 18766 14646
rect 18708 14458 18766 14470
rect 18826 14646 18884 14658
rect 18826 14470 18838 14646
rect 18872 14470 18884 14646
rect 18826 14458 18884 14470
rect 19396 14642 19454 14654
rect 19396 14466 19408 14642
rect 19442 14466 19454 14642
rect 19396 14454 19454 14466
rect 19514 14642 19572 14654
rect 19514 14466 19526 14642
rect 19560 14466 19572 14642
rect 19514 14454 19572 14466
rect 19632 14642 19690 14654
rect 19632 14466 19644 14642
rect 19678 14466 19690 14642
rect 19632 14454 19690 14466
rect 19750 14642 19808 14654
rect 19750 14466 19762 14642
rect 19796 14466 19808 14642
rect 19750 14454 19808 14466
rect 19869 14466 19881 14842
rect 19915 14466 19927 14842
rect 19869 14454 19927 14466
rect 19987 14842 20045 14854
rect 19987 14466 19999 14842
rect 20033 14466 20045 14842
rect 19987 14454 20045 14466
rect 20105 14842 20163 14854
rect 20105 14466 20117 14842
rect 20151 14466 20163 14842
rect 20105 14454 20163 14466
rect 20223 14842 20281 14854
rect 20223 14466 20235 14842
rect 20269 14466 20281 14842
rect 20223 14454 20281 14466
rect 20342 14842 20400 14854
rect 20342 14466 20354 14842
rect 20388 14466 20400 14842
rect 20342 14454 20400 14466
rect 20460 14842 20518 14854
rect 20460 14466 20472 14842
rect 20506 14466 20518 14842
rect 20460 14454 20518 14466
rect 20578 14842 20636 14854
rect 20578 14466 20590 14842
rect 20624 14466 20636 14842
rect 20578 14454 20636 14466
rect 20696 14842 20754 14854
rect 20696 14466 20708 14842
rect 20742 14466 20754 14842
rect 20696 14454 20754 14466
rect 20814 14842 20872 14854
rect 20814 14466 20826 14842
rect 20860 14466 20872 14842
rect 20814 14454 20872 14466
rect 20932 14842 20990 14854
rect 20932 14466 20944 14842
rect 20978 14466 20990 14842
rect 20932 14454 20990 14466
rect 21050 14842 21108 14854
rect 21050 14466 21062 14842
rect 21096 14466 21108 14842
rect 21050 14454 21108 14466
rect 21163 14842 21221 14854
rect 21163 14466 21175 14842
rect 21209 14466 21221 14842
rect 21163 14454 21221 14466
rect 21281 14842 21339 14854
rect 21281 14466 21293 14842
rect 21327 14466 21339 14842
rect 21281 14454 21339 14466
rect 21399 14842 21457 14854
rect 21399 14466 21411 14842
rect 21445 14466 21457 14842
rect 21399 14454 21457 14466
rect 21517 14842 21575 14854
rect 21517 14466 21529 14842
rect 21563 14654 21575 14842
rect 23013 14842 23071 14854
rect 21563 14642 21662 14654
rect 21563 14466 21616 14642
rect 21650 14466 21662 14642
rect 21517 14454 21662 14466
rect 21722 14642 21780 14654
rect 21722 14466 21734 14642
rect 21768 14466 21780 14642
rect 21722 14454 21780 14466
rect 21840 14642 21898 14654
rect 21840 14466 21852 14642
rect 21886 14466 21898 14642
rect 21840 14454 21898 14466
rect 21958 14642 22016 14654
rect 21958 14466 21970 14642
rect 22004 14466 22016 14642
rect 21958 14454 22016 14466
rect 22540 14642 22598 14654
rect 22540 14466 22552 14642
rect 22586 14466 22598 14642
rect 22540 14454 22598 14466
rect 22658 14642 22716 14654
rect 22658 14466 22670 14642
rect 22704 14466 22716 14642
rect 22658 14454 22716 14466
rect 22776 14642 22834 14654
rect 22776 14466 22788 14642
rect 22822 14466 22834 14642
rect 22776 14454 22834 14466
rect 22894 14642 22952 14654
rect 22894 14466 22906 14642
rect 22940 14466 22952 14642
rect 22894 14454 22952 14466
rect 23013 14466 23025 14842
rect 23059 14466 23071 14842
rect 23013 14454 23071 14466
rect 23131 14842 23189 14854
rect 23131 14466 23143 14842
rect 23177 14466 23189 14842
rect 23131 14454 23189 14466
rect 23249 14842 23307 14854
rect 23249 14466 23261 14842
rect 23295 14466 23307 14842
rect 23249 14454 23307 14466
rect 23367 14842 23425 14854
rect 23367 14466 23379 14842
rect 23413 14466 23425 14842
rect 23367 14454 23425 14466
rect 23486 14842 23544 14854
rect 23486 14466 23498 14842
rect 23532 14466 23544 14842
rect 23486 14454 23544 14466
rect 23604 14842 23662 14854
rect 23604 14466 23616 14842
rect 23650 14466 23662 14842
rect 23604 14454 23662 14466
rect 23722 14842 23780 14854
rect 23722 14466 23734 14842
rect 23768 14466 23780 14842
rect 23722 14454 23780 14466
rect 23840 14842 23898 14854
rect 23840 14466 23852 14842
rect 23886 14466 23898 14842
rect 23840 14454 23898 14466
rect 23958 14842 24016 14854
rect 23958 14466 23970 14842
rect 24004 14466 24016 14842
rect 23958 14454 24016 14466
rect 24076 14842 24134 14854
rect 24076 14466 24088 14842
rect 24122 14466 24134 14842
rect 24076 14454 24134 14466
rect 24194 14842 24252 14854
rect 24194 14466 24206 14842
rect 24240 14466 24252 14842
rect 24194 14454 24252 14466
rect 24307 14842 24365 14854
rect 24307 14466 24319 14842
rect 24353 14466 24365 14842
rect 24307 14454 24365 14466
rect 24425 14842 24483 14854
rect 24425 14466 24437 14842
rect 24471 14466 24483 14842
rect 24425 14454 24483 14466
rect 24543 14842 24601 14854
rect 24543 14466 24555 14842
rect 24589 14466 24601 14842
rect 24543 14454 24601 14466
rect 24661 14842 24719 14854
rect 24661 14466 24673 14842
rect 24707 14654 24719 14842
rect 58328 16650 58386 16662
rect 58328 16474 58340 16650
rect 58374 16474 58386 16650
rect 58328 16462 58386 16474
rect 58446 16650 58504 16662
rect 58446 16474 58458 16650
rect 58492 16474 58504 16650
rect 58446 16462 58504 16474
rect 58564 16650 58622 16662
rect 58564 16474 58576 16650
rect 58610 16474 58622 16650
rect 58564 16462 58622 16474
rect 58682 16650 58740 16662
rect 58682 16474 58694 16650
rect 58728 16474 58740 16650
rect 58682 16462 58740 16474
rect 58811 16474 58823 16850
rect 58857 16474 58869 16850
rect 58811 16462 58869 16474
rect 58929 16850 58987 16862
rect 58929 16474 58941 16850
rect 58975 16474 58987 16850
rect 58929 16462 58987 16474
rect 59047 16850 59105 16862
rect 59047 16474 59059 16850
rect 59093 16474 59105 16850
rect 59047 16462 59105 16474
rect 59165 16850 59223 16862
rect 59165 16474 59177 16850
rect 59211 16474 59223 16850
rect 59165 16462 59223 16474
rect 59283 16850 59341 16862
rect 59283 16474 59295 16850
rect 59329 16474 59341 16850
rect 59283 16462 59341 16474
rect 59401 16850 59459 16862
rect 59401 16474 59413 16850
rect 59447 16474 59459 16850
rect 59401 16462 59459 16474
rect 59519 16850 59577 16862
rect 59519 16474 59531 16850
rect 59565 16474 59577 16850
rect 60709 16850 60767 16862
rect 59519 16462 59577 16474
rect 59649 16650 59707 16662
rect 59649 16474 59661 16650
rect 59695 16474 59707 16650
rect 59649 16462 59707 16474
rect 59767 16650 59825 16662
rect 59767 16474 59779 16650
rect 59813 16474 59825 16650
rect 59767 16462 59825 16474
rect 59885 16650 59943 16662
rect 59885 16474 59897 16650
rect 59931 16474 59943 16650
rect 59885 16462 59943 16474
rect 60003 16650 60061 16662
rect 60003 16474 60015 16650
rect 60049 16474 60061 16650
rect 60003 16462 60061 16474
rect 60226 16650 60284 16662
rect 60226 16474 60238 16650
rect 60272 16474 60284 16650
rect 60226 16462 60284 16474
rect 60344 16650 60402 16662
rect 60344 16474 60356 16650
rect 60390 16474 60402 16650
rect 60344 16462 60402 16474
rect 60462 16650 60520 16662
rect 60462 16474 60474 16650
rect 60508 16474 60520 16650
rect 60462 16462 60520 16474
rect 60580 16650 60638 16662
rect 60580 16474 60592 16650
rect 60626 16474 60638 16650
rect 60580 16462 60638 16474
rect 60709 16474 60721 16850
rect 60755 16474 60767 16850
rect 60709 16462 60767 16474
rect 60827 16850 60885 16862
rect 60827 16474 60839 16850
rect 60873 16474 60885 16850
rect 60827 16462 60885 16474
rect 60945 16850 61003 16862
rect 60945 16474 60957 16850
rect 60991 16474 61003 16850
rect 60945 16462 61003 16474
rect 61063 16850 61121 16862
rect 61063 16474 61075 16850
rect 61109 16474 61121 16850
rect 61063 16462 61121 16474
rect 61181 16850 61239 16862
rect 61181 16474 61193 16850
rect 61227 16474 61239 16850
rect 61181 16462 61239 16474
rect 61299 16850 61357 16862
rect 61299 16474 61311 16850
rect 61345 16474 61357 16850
rect 61299 16462 61357 16474
rect 61417 16850 61475 16862
rect 61417 16474 61429 16850
rect 61463 16474 61475 16850
rect 70513 17064 70913 17076
rect 70513 17030 70525 17064
rect 70901 17030 70913 17064
rect 70513 17018 70913 17030
rect 70513 16946 70913 16958
rect 70513 16912 70525 16946
rect 70901 16912 70913 16946
rect 70513 16900 70913 16912
rect 61417 16462 61475 16474
rect 61547 16650 61605 16662
rect 61547 16474 61559 16650
rect 61593 16474 61605 16650
rect 61547 16462 61605 16474
rect 61665 16650 61723 16662
rect 61665 16474 61677 16650
rect 61711 16474 61723 16650
rect 61665 16462 61723 16474
rect 61783 16650 61841 16662
rect 61783 16474 61795 16650
rect 61829 16474 61841 16650
rect 61783 16462 61841 16474
rect 61901 16650 61959 16662
rect 61901 16474 61913 16650
rect 61947 16474 61959 16650
rect 61901 16462 61959 16474
rect 54253 16154 54311 16166
rect 54253 15778 54265 16154
rect 54299 15778 54311 16154
rect 54253 15766 54311 15778
rect 54371 16154 54429 16166
rect 54371 15778 54383 16154
rect 54417 15778 54429 16154
rect 54371 15766 54429 15778
rect 54489 16154 54547 16166
rect 54489 15778 54501 16154
rect 54535 15778 54547 16154
rect 54489 15766 54547 15778
rect 54607 16154 54665 16166
rect 54607 15778 54619 16154
rect 54653 15778 54665 16154
rect 54607 15766 54665 15778
rect 54725 16154 54783 16166
rect 54725 15778 54737 16154
rect 54771 15778 54783 16154
rect 54725 15766 54783 15778
rect 54843 16154 54901 16166
rect 54843 15778 54855 16154
rect 54889 15778 54901 16154
rect 54843 15766 54901 15778
rect 54961 16154 55019 16166
rect 54961 15778 54973 16154
rect 55007 15778 55019 16154
rect 54961 15766 55019 15778
rect 55795 15660 55853 15672
rect 55795 15484 55807 15660
rect 55841 15484 55853 15660
rect 55795 15472 55853 15484
rect 55913 15660 55971 15672
rect 55913 15484 55925 15660
rect 55959 15484 55971 15660
rect 55913 15472 55971 15484
rect 56031 15660 56089 15672
rect 56031 15484 56043 15660
rect 56077 15484 56089 15660
rect 56031 15472 56089 15484
rect 56149 15660 56207 15672
rect 56149 15484 56161 15660
rect 56195 15484 56207 15660
rect 56149 15472 56207 15484
rect 56267 15660 56325 15672
rect 56267 15484 56279 15660
rect 56313 15484 56325 15660
rect 56267 15472 56325 15484
rect 56385 15660 56443 15672
rect 56385 15484 56397 15660
rect 56431 15484 56443 15660
rect 56385 15472 56443 15484
rect 56503 15660 56561 15672
rect 56503 15484 56515 15660
rect 56549 15484 56561 15660
rect 56503 15472 56561 15484
rect 56621 15660 56679 15672
rect 56621 15484 56633 15660
rect 56667 15484 56679 15660
rect 56621 15472 56679 15484
rect 56739 15660 56797 15672
rect 56739 15484 56751 15660
rect 56785 15484 56797 15660
rect 56739 15472 56797 15484
rect 56857 15660 56915 15672
rect 56857 15484 56869 15660
rect 56903 15484 56915 15660
rect 56857 15472 56915 15484
rect 58868 16157 58926 16169
rect 58868 15781 58880 16157
rect 58914 15781 58926 16157
rect 58868 15769 58926 15781
rect 58986 16157 59044 16169
rect 58986 15781 58998 16157
rect 59032 15781 59044 16157
rect 58986 15769 59044 15781
rect 59104 16157 59162 16169
rect 59104 15781 59116 16157
rect 59150 15781 59162 16157
rect 59104 15769 59162 15781
rect 59222 16157 59280 16169
rect 59222 15781 59234 16157
rect 59268 15781 59280 16157
rect 59222 15769 59280 15781
rect 59340 16157 59398 16169
rect 59340 15781 59352 16157
rect 59386 15781 59398 16157
rect 59340 15769 59398 15781
rect 59458 16157 59516 16169
rect 59458 15781 59470 16157
rect 59504 15781 59516 16157
rect 59458 15769 59516 15781
rect 59576 16157 59634 16169
rect 59576 15781 59588 16157
rect 59622 15781 59634 16157
rect 59576 15769 59634 15781
rect 70513 16828 70913 16840
rect 70513 16794 70525 16828
rect 70901 16794 70913 16828
rect 70513 16782 70913 16794
rect 70713 16709 70913 16721
rect 70713 16675 70725 16709
rect 70901 16675 70913 16709
rect 70713 16663 70913 16675
rect 70713 16591 70913 16603
rect 70713 16557 70725 16591
rect 70901 16557 70913 16591
rect 70713 16545 70913 16557
rect 70713 16473 70913 16485
rect 70713 16439 70725 16473
rect 70901 16439 70913 16473
rect 70713 16427 70913 16439
rect 70713 16355 70913 16367
rect 70713 16321 70725 16355
rect 70901 16321 70913 16355
rect 70713 16309 70913 16321
rect 60766 16157 60824 16169
rect 60766 15781 60778 16157
rect 60812 15781 60824 16157
rect 60766 15769 60824 15781
rect 60884 16157 60942 16169
rect 60884 15781 60896 16157
rect 60930 15781 60942 16157
rect 60884 15769 60942 15781
rect 61002 16157 61060 16169
rect 61002 15781 61014 16157
rect 61048 15781 61060 16157
rect 61002 15769 61060 15781
rect 61120 16157 61178 16169
rect 61120 15781 61132 16157
rect 61166 15781 61178 16157
rect 61120 15769 61178 15781
rect 61238 16157 61296 16169
rect 61238 15781 61250 16157
rect 61284 15781 61296 16157
rect 61238 15769 61296 15781
rect 61356 16157 61414 16169
rect 61356 15781 61368 16157
rect 61402 15781 61414 16157
rect 61356 15769 61414 15781
rect 61474 16157 61532 16169
rect 61474 15781 61486 16157
rect 61520 15781 61532 16157
rect 61474 15769 61532 15781
rect 70709 15785 70909 15797
rect 70709 15751 70721 15785
rect 70897 15751 70909 15785
rect 70709 15739 70909 15751
rect 62308 15663 62366 15675
rect 62308 15487 62320 15663
rect 62354 15487 62366 15663
rect 62308 15475 62366 15487
rect 62426 15663 62484 15675
rect 62426 15487 62438 15663
rect 62472 15487 62484 15663
rect 62426 15475 62484 15487
rect 62544 15663 62602 15675
rect 62544 15487 62556 15663
rect 62590 15487 62602 15663
rect 62544 15475 62602 15487
rect 62662 15663 62720 15675
rect 62662 15487 62674 15663
rect 62708 15487 62720 15663
rect 62662 15475 62720 15487
rect 62780 15663 62838 15675
rect 62780 15487 62792 15663
rect 62826 15487 62838 15663
rect 62780 15475 62838 15487
rect 62898 15663 62956 15675
rect 62898 15487 62910 15663
rect 62944 15487 62956 15663
rect 62898 15475 62956 15487
rect 63016 15663 63074 15675
rect 63016 15487 63028 15663
rect 63062 15487 63074 15663
rect 63016 15475 63074 15487
rect 63134 15663 63192 15675
rect 63134 15487 63146 15663
rect 63180 15487 63192 15663
rect 63134 15475 63192 15487
rect 63252 15663 63310 15675
rect 63252 15487 63264 15663
rect 63298 15487 63310 15663
rect 63252 15475 63310 15487
rect 63370 15663 63428 15675
rect 63370 15487 63382 15663
rect 63416 15487 63428 15663
rect 63370 15475 63428 15487
rect 70709 15667 70909 15679
rect 70709 15633 70721 15667
rect 70897 15633 70909 15667
rect 70709 15621 70909 15633
rect 70709 15549 70909 15561
rect 70709 15515 70721 15549
rect 70897 15515 70909 15549
rect 70709 15503 70909 15515
rect 24707 14642 24806 14654
rect 24707 14466 24760 14642
rect 24794 14466 24806 14642
rect 24661 14454 24806 14466
rect 24866 14642 24924 14654
rect 24866 14466 24878 14642
rect 24912 14466 24924 14642
rect 24866 14454 24924 14466
rect 24984 14642 25042 14654
rect 24984 14466 24996 14642
rect 25030 14466 25042 14642
rect 24984 14454 25042 14466
rect 25102 14642 25160 14654
rect 25102 14466 25114 14642
rect 25148 14466 25160 14642
rect 70709 15431 70909 15443
rect 70709 15397 70721 15431
rect 70897 15397 70909 15431
rect 70709 15356 70909 15397
rect 70509 15344 70909 15356
rect 70509 15310 70521 15344
rect 70897 15310 70909 15344
rect 70509 15298 70909 15310
rect 70509 15226 70909 15238
rect 70509 15192 70521 15226
rect 70897 15192 70909 15226
rect 70509 15180 70909 15192
rect 70509 15108 70909 15120
rect 70509 15074 70521 15108
rect 70897 15074 70909 15108
rect 70509 15062 70909 15074
rect 70509 14990 70909 15002
rect 70509 14956 70521 14990
rect 70897 14956 70909 14990
rect 70509 14944 70909 14956
rect 70509 14877 70909 14889
rect 70509 14843 70521 14877
rect 70897 14843 70909 14877
rect 70509 14831 70909 14843
rect 70509 14759 70909 14771
rect 70509 14725 70521 14759
rect 70897 14725 70909 14759
rect 70509 14713 70909 14725
rect 25102 14454 25160 14466
rect 70509 14641 70909 14653
rect 70509 14607 70521 14641
rect 70897 14607 70909 14641
rect 70509 14595 70909 14607
rect 70509 14523 70909 14535
rect 70509 14489 70521 14523
rect 70897 14489 70909 14523
rect 70509 14477 70909 14489
rect 70509 14405 70909 14417
rect 70509 14371 70521 14405
rect 70897 14371 70909 14405
rect 70509 14359 70909 14371
rect 70509 14287 70909 14299
rect 70509 14253 70521 14287
rect 70897 14253 70909 14287
rect 70509 14241 70909 14253
rect 70509 14169 70909 14181
rect 70509 14135 70521 14169
rect 70897 14135 70909 14169
rect 70509 14123 70909 14135
rect 70509 14050 70909 14062
rect 70509 14016 70521 14050
rect 70897 14016 70909 14050
rect 70509 14004 70909 14016
rect 70509 13932 70909 13944
rect 70509 13898 70521 13932
rect 70897 13898 70909 13932
rect 70509 13886 70909 13898
rect 70509 13814 70909 13826
rect 70509 13780 70521 13814
rect 70897 13780 70909 13814
rect 70509 13768 70909 13780
rect 70509 13696 70909 13708
rect 70509 13662 70521 13696
rect 70897 13662 70909 13696
rect 70509 13650 70909 13662
rect 70709 13577 70909 13589
rect 70709 13543 70721 13577
rect 70897 13543 70909 13577
rect 70709 13531 70909 13543
rect 70709 13459 70909 13471
rect 70709 13425 70721 13459
rect 70897 13425 70909 13459
rect 70709 13413 70909 13425
rect 70709 13341 70909 13353
rect 70709 13307 70721 13341
rect 70897 13307 70909 13341
rect 70709 13295 70909 13307
rect 70709 13223 70909 13235
rect 70709 13189 70721 13223
rect 70897 13189 70909 13223
rect 30154 13168 30354 13180
rect 70709 13177 70909 13189
rect 30154 13134 30166 13168
rect 30342 13134 30354 13168
rect 30154 13122 30354 13134
rect 30154 13050 30354 13062
rect 30154 13016 30166 13050
rect 30342 13016 30354 13050
rect 30154 13004 30354 13016
rect 30154 12932 30354 12944
rect 30154 12898 30166 12932
rect 30342 12898 30354 12932
rect 30154 12886 30354 12898
rect 30154 12814 30354 12826
rect 30154 12780 30166 12814
rect 30342 12780 30354 12814
rect 30154 12768 30354 12780
rect 29954 12684 30354 12696
rect 29954 12650 29966 12684
rect 30342 12650 30354 12684
rect 29954 12638 30354 12650
rect 30647 12741 31047 12753
rect 30647 12707 30659 12741
rect 31035 12707 31047 12741
rect 30647 12695 31047 12707
rect 29954 12566 30354 12578
rect 29954 12532 29966 12566
rect 30342 12532 30354 12566
rect 29954 12520 30354 12532
rect 30647 12623 31047 12635
rect 30647 12589 30659 12623
rect 31035 12589 31047 12623
rect 30647 12577 31047 12589
rect 70709 12641 70909 12653
rect 70709 12607 70721 12641
rect 70897 12607 70909 12641
rect 70709 12595 70909 12607
rect 29954 12448 30354 12460
rect 29954 12414 29966 12448
rect 30342 12414 30354 12448
rect 29954 12402 30354 12414
rect 30647 12505 31047 12517
rect 30647 12471 30659 12505
rect 31035 12471 31047 12505
rect 30647 12459 31047 12471
rect 70709 12523 70909 12535
rect 70709 12489 70721 12523
rect 70897 12489 70909 12523
rect 70709 12477 70909 12489
rect 30647 12387 31047 12399
rect 30647 12353 30659 12387
rect 31035 12353 31047 12387
rect 29954 12330 30354 12342
rect 30647 12341 31047 12353
rect 29954 12296 29966 12330
rect 30342 12296 30354 12330
rect 29954 12284 30354 12296
rect 971 12112 1029 12124
rect 498 11912 556 11924
rect 498 11736 510 11912
rect 544 11736 556 11912
rect 498 11724 556 11736
rect 616 11912 674 11924
rect 616 11736 628 11912
rect 662 11736 674 11912
rect 616 11724 674 11736
rect 734 11912 792 11924
rect 734 11736 746 11912
rect 780 11736 792 11912
rect 734 11724 792 11736
rect 852 11912 910 11924
rect 852 11736 864 11912
rect 898 11736 910 11912
rect 852 11724 910 11736
rect 971 11736 983 12112
rect 1017 11736 1029 12112
rect 971 11724 1029 11736
rect 1089 12112 1147 12124
rect 1089 11736 1101 12112
rect 1135 11736 1147 12112
rect 1089 11724 1147 11736
rect 1207 12112 1265 12124
rect 1207 11736 1219 12112
rect 1253 11736 1265 12112
rect 1207 11724 1265 11736
rect 1325 12112 1383 12124
rect 1325 11736 1337 12112
rect 1371 11736 1383 12112
rect 1325 11724 1383 11736
rect 1444 12112 1502 12124
rect 1444 11736 1456 12112
rect 1490 11736 1502 12112
rect 1444 11724 1502 11736
rect 1562 12112 1620 12124
rect 1562 11736 1574 12112
rect 1608 11736 1620 12112
rect 1562 11724 1620 11736
rect 1680 12112 1738 12124
rect 1680 11736 1692 12112
rect 1726 11736 1738 12112
rect 1680 11724 1738 11736
rect 1798 12112 1856 12124
rect 1798 11736 1810 12112
rect 1844 11736 1856 12112
rect 1798 11724 1856 11736
rect 1916 12112 1974 12124
rect 1916 11736 1928 12112
rect 1962 11736 1974 12112
rect 1916 11724 1974 11736
rect 2034 12112 2092 12124
rect 2034 11736 2046 12112
rect 2080 11736 2092 12112
rect 2034 11724 2092 11736
rect 2152 12112 2210 12124
rect 2152 11736 2164 12112
rect 2198 11736 2210 12112
rect 2152 11724 2210 11736
rect 2265 12112 2323 12124
rect 2265 11736 2277 12112
rect 2311 11736 2323 12112
rect 2265 11724 2323 11736
rect 2383 12112 2441 12124
rect 2383 11736 2395 12112
rect 2429 11736 2441 12112
rect 2383 11724 2441 11736
rect 2501 12112 2559 12124
rect 2501 11736 2513 12112
rect 2547 11736 2559 12112
rect 2501 11724 2559 11736
rect 2619 12112 2677 12124
rect 2619 11736 2631 12112
rect 2665 11924 2677 12112
rect 4115 12112 4173 12124
rect 2665 11912 2764 11924
rect 2665 11736 2718 11912
rect 2752 11736 2764 11912
rect 2619 11724 2764 11736
rect 2824 11912 2882 11924
rect 2824 11736 2836 11912
rect 2870 11736 2882 11912
rect 2824 11724 2882 11736
rect 2942 11912 3000 11924
rect 2942 11736 2954 11912
rect 2988 11736 3000 11912
rect 2942 11724 3000 11736
rect 3060 11912 3118 11924
rect 3060 11736 3072 11912
rect 3106 11736 3118 11912
rect 3060 11724 3118 11736
rect 3642 11912 3700 11924
rect 3642 11736 3654 11912
rect 3688 11736 3700 11912
rect 3642 11724 3700 11736
rect 3760 11912 3818 11924
rect 3760 11736 3772 11912
rect 3806 11736 3818 11912
rect 3760 11724 3818 11736
rect 3878 11912 3936 11924
rect 3878 11736 3890 11912
rect 3924 11736 3936 11912
rect 3878 11724 3936 11736
rect 3996 11912 4054 11924
rect 3996 11736 4008 11912
rect 4042 11736 4054 11912
rect 3996 11724 4054 11736
rect 4115 11736 4127 12112
rect 4161 11736 4173 12112
rect 4115 11724 4173 11736
rect 4233 12112 4291 12124
rect 4233 11736 4245 12112
rect 4279 11736 4291 12112
rect 4233 11724 4291 11736
rect 4351 12112 4409 12124
rect 4351 11736 4363 12112
rect 4397 11736 4409 12112
rect 4351 11724 4409 11736
rect 4469 12112 4527 12124
rect 4469 11736 4481 12112
rect 4515 11736 4527 12112
rect 4469 11724 4527 11736
rect 4588 12112 4646 12124
rect 4588 11736 4600 12112
rect 4634 11736 4646 12112
rect 4588 11724 4646 11736
rect 4706 12112 4764 12124
rect 4706 11736 4718 12112
rect 4752 11736 4764 12112
rect 4706 11724 4764 11736
rect 4824 12112 4882 12124
rect 4824 11736 4836 12112
rect 4870 11736 4882 12112
rect 4824 11724 4882 11736
rect 4942 12112 5000 12124
rect 4942 11736 4954 12112
rect 4988 11736 5000 12112
rect 4942 11724 5000 11736
rect 5060 12112 5118 12124
rect 5060 11736 5072 12112
rect 5106 11736 5118 12112
rect 5060 11724 5118 11736
rect 5178 12112 5236 12124
rect 5178 11736 5190 12112
rect 5224 11736 5236 12112
rect 5178 11724 5236 11736
rect 5296 12112 5354 12124
rect 5296 11736 5308 12112
rect 5342 11736 5354 12112
rect 5296 11724 5354 11736
rect 5409 12112 5467 12124
rect 5409 11736 5421 12112
rect 5455 11736 5467 12112
rect 5409 11724 5467 11736
rect 5527 12112 5585 12124
rect 5527 11736 5539 12112
rect 5573 11736 5585 12112
rect 5527 11724 5585 11736
rect 5645 12112 5703 12124
rect 5645 11736 5657 12112
rect 5691 11736 5703 12112
rect 5645 11724 5703 11736
rect 5763 12112 5821 12124
rect 5763 11736 5775 12112
rect 5809 11924 5821 12112
rect 7247 12108 7305 12120
rect 5809 11912 5908 11924
rect 5809 11736 5862 11912
rect 5896 11736 5908 11912
rect 5763 11724 5908 11736
rect 5968 11912 6026 11924
rect 5968 11736 5980 11912
rect 6014 11736 6026 11912
rect 5968 11724 6026 11736
rect 6086 11912 6144 11924
rect 6086 11736 6098 11912
rect 6132 11736 6144 11912
rect 6086 11724 6144 11736
rect 6204 11912 6262 11924
rect 6204 11736 6216 11912
rect 6250 11736 6262 11912
rect 6204 11724 6262 11736
rect 6774 11908 6832 11920
rect 6774 11732 6786 11908
rect 6820 11732 6832 11908
rect 6774 11720 6832 11732
rect 6892 11908 6950 11920
rect 6892 11732 6904 11908
rect 6938 11732 6950 11908
rect 6892 11720 6950 11732
rect 7010 11908 7068 11920
rect 7010 11732 7022 11908
rect 7056 11732 7068 11908
rect 7010 11720 7068 11732
rect 7128 11908 7186 11920
rect 7128 11732 7140 11908
rect 7174 11732 7186 11908
rect 7128 11720 7186 11732
rect 7247 11732 7259 12108
rect 7293 11732 7305 12108
rect 7247 11720 7305 11732
rect 7365 12108 7423 12120
rect 7365 11732 7377 12108
rect 7411 11732 7423 12108
rect 7365 11720 7423 11732
rect 7483 12108 7541 12120
rect 7483 11732 7495 12108
rect 7529 11732 7541 12108
rect 7483 11720 7541 11732
rect 7601 12108 7659 12120
rect 7601 11732 7613 12108
rect 7647 11732 7659 12108
rect 7601 11720 7659 11732
rect 7720 12108 7778 12120
rect 7720 11732 7732 12108
rect 7766 11732 7778 12108
rect 7720 11720 7778 11732
rect 7838 12108 7896 12120
rect 7838 11732 7850 12108
rect 7884 11732 7896 12108
rect 7838 11720 7896 11732
rect 7956 12108 8014 12120
rect 7956 11732 7968 12108
rect 8002 11732 8014 12108
rect 7956 11720 8014 11732
rect 8074 12108 8132 12120
rect 8074 11732 8086 12108
rect 8120 11732 8132 12108
rect 8074 11720 8132 11732
rect 8192 12108 8250 12120
rect 8192 11732 8204 12108
rect 8238 11732 8250 12108
rect 8192 11720 8250 11732
rect 8310 12108 8368 12120
rect 8310 11732 8322 12108
rect 8356 11732 8368 12108
rect 8310 11720 8368 11732
rect 8428 12108 8486 12120
rect 8428 11732 8440 12108
rect 8474 11732 8486 12108
rect 8428 11720 8486 11732
rect 8541 12108 8599 12120
rect 8541 11732 8553 12108
rect 8587 11732 8599 12108
rect 8541 11720 8599 11732
rect 8659 12108 8717 12120
rect 8659 11732 8671 12108
rect 8705 11732 8717 12108
rect 8659 11720 8717 11732
rect 8777 12108 8835 12120
rect 8777 11732 8789 12108
rect 8823 11732 8835 12108
rect 8777 11720 8835 11732
rect 8895 12108 8953 12120
rect 8895 11732 8907 12108
rect 8941 11920 8953 12108
rect 10391 12108 10449 12120
rect 8941 11908 9040 11920
rect 8941 11732 8994 11908
rect 9028 11732 9040 11908
rect 8895 11720 9040 11732
rect 9100 11908 9158 11920
rect 9100 11732 9112 11908
rect 9146 11732 9158 11908
rect 9100 11720 9158 11732
rect 9218 11908 9276 11920
rect 9218 11732 9230 11908
rect 9264 11732 9276 11908
rect 9218 11720 9276 11732
rect 9336 11908 9394 11920
rect 9336 11732 9348 11908
rect 9382 11732 9394 11908
rect 9336 11720 9394 11732
rect 9918 11908 9976 11920
rect 9918 11732 9930 11908
rect 9964 11732 9976 11908
rect 9918 11720 9976 11732
rect 10036 11908 10094 11920
rect 10036 11732 10048 11908
rect 10082 11732 10094 11908
rect 10036 11720 10094 11732
rect 10154 11908 10212 11920
rect 10154 11732 10166 11908
rect 10200 11732 10212 11908
rect 10154 11720 10212 11732
rect 10272 11908 10330 11920
rect 10272 11732 10284 11908
rect 10318 11732 10330 11908
rect 10272 11720 10330 11732
rect 10391 11732 10403 12108
rect 10437 11732 10449 12108
rect 10391 11720 10449 11732
rect 10509 12108 10567 12120
rect 10509 11732 10521 12108
rect 10555 11732 10567 12108
rect 10509 11720 10567 11732
rect 10627 12108 10685 12120
rect 10627 11732 10639 12108
rect 10673 11732 10685 12108
rect 10627 11720 10685 11732
rect 10745 12108 10803 12120
rect 10745 11732 10757 12108
rect 10791 11732 10803 12108
rect 10745 11720 10803 11732
rect 10864 12108 10922 12120
rect 10864 11732 10876 12108
rect 10910 11732 10922 12108
rect 10864 11720 10922 11732
rect 10982 12108 11040 12120
rect 10982 11732 10994 12108
rect 11028 11732 11040 12108
rect 10982 11720 11040 11732
rect 11100 12108 11158 12120
rect 11100 11732 11112 12108
rect 11146 11732 11158 12108
rect 11100 11720 11158 11732
rect 11218 12108 11276 12120
rect 11218 11732 11230 12108
rect 11264 11732 11276 12108
rect 11218 11720 11276 11732
rect 11336 12108 11394 12120
rect 11336 11732 11348 12108
rect 11382 11732 11394 12108
rect 11336 11720 11394 11732
rect 11454 12108 11512 12120
rect 11454 11732 11466 12108
rect 11500 11732 11512 12108
rect 11454 11720 11512 11732
rect 11572 12108 11630 12120
rect 11572 11732 11584 12108
rect 11618 11732 11630 12108
rect 11572 11720 11630 11732
rect 11685 12108 11743 12120
rect 11685 11732 11697 12108
rect 11731 11732 11743 12108
rect 11685 11720 11743 11732
rect 11803 12108 11861 12120
rect 11803 11732 11815 12108
rect 11849 11732 11861 12108
rect 11803 11720 11861 11732
rect 11921 12108 11979 12120
rect 11921 11732 11933 12108
rect 11967 11732 11979 12108
rect 11921 11720 11979 11732
rect 12039 12108 12097 12120
rect 12039 11732 12051 12108
rect 12085 11920 12097 12108
rect 13593 12112 13651 12124
rect 12085 11908 12184 11920
rect 12085 11732 12138 11908
rect 12172 11732 12184 11908
rect 12039 11720 12184 11732
rect 12244 11908 12302 11920
rect 12244 11732 12256 11908
rect 12290 11732 12302 11908
rect 12244 11720 12302 11732
rect 12362 11908 12420 11920
rect 12362 11732 12374 11908
rect 12408 11732 12420 11908
rect 12362 11720 12420 11732
rect 12480 11908 12538 11920
rect 12480 11732 12492 11908
rect 12526 11732 12538 11908
rect 12480 11720 12538 11732
rect 13120 11912 13178 11924
rect 13120 11736 13132 11912
rect 13166 11736 13178 11912
rect 13120 11724 13178 11736
rect 13238 11912 13296 11924
rect 13238 11736 13250 11912
rect 13284 11736 13296 11912
rect 13238 11724 13296 11736
rect 13356 11912 13414 11924
rect 13356 11736 13368 11912
rect 13402 11736 13414 11912
rect 13356 11724 13414 11736
rect 13474 11912 13532 11924
rect 13474 11736 13486 11912
rect 13520 11736 13532 11912
rect 13474 11724 13532 11736
rect 13593 11736 13605 12112
rect 13639 11736 13651 12112
rect 13593 11724 13651 11736
rect 13711 12112 13769 12124
rect 13711 11736 13723 12112
rect 13757 11736 13769 12112
rect 13711 11724 13769 11736
rect 13829 12112 13887 12124
rect 13829 11736 13841 12112
rect 13875 11736 13887 12112
rect 13829 11724 13887 11736
rect 13947 12112 14005 12124
rect 13947 11736 13959 12112
rect 13993 11736 14005 12112
rect 13947 11724 14005 11736
rect 14066 12112 14124 12124
rect 14066 11736 14078 12112
rect 14112 11736 14124 12112
rect 14066 11724 14124 11736
rect 14184 12112 14242 12124
rect 14184 11736 14196 12112
rect 14230 11736 14242 12112
rect 14184 11724 14242 11736
rect 14302 12112 14360 12124
rect 14302 11736 14314 12112
rect 14348 11736 14360 12112
rect 14302 11724 14360 11736
rect 14420 12112 14478 12124
rect 14420 11736 14432 12112
rect 14466 11736 14478 12112
rect 14420 11724 14478 11736
rect 14538 12112 14596 12124
rect 14538 11736 14550 12112
rect 14584 11736 14596 12112
rect 14538 11724 14596 11736
rect 14656 12112 14714 12124
rect 14656 11736 14668 12112
rect 14702 11736 14714 12112
rect 14656 11724 14714 11736
rect 14774 12112 14832 12124
rect 14774 11736 14786 12112
rect 14820 11736 14832 12112
rect 14774 11724 14832 11736
rect 14887 12112 14945 12124
rect 14887 11736 14899 12112
rect 14933 11736 14945 12112
rect 14887 11724 14945 11736
rect 15005 12112 15063 12124
rect 15005 11736 15017 12112
rect 15051 11736 15063 12112
rect 15005 11724 15063 11736
rect 15123 12112 15181 12124
rect 15123 11736 15135 12112
rect 15169 11736 15181 12112
rect 15123 11724 15181 11736
rect 15241 12112 15299 12124
rect 15241 11736 15253 12112
rect 15287 11924 15299 12112
rect 16737 12112 16795 12124
rect 15287 11912 15386 11924
rect 15287 11736 15340 11912
rect 15374 11736 15386 11912
rect 15241 11724 15386 11736
rect 15446 11912 15504 11924
rect 15446 11736 15458 11912
rect 15492 11736 15504 11912
rect 15446 11724 15504 11736
rect 15564 11912 15622 11924
rect 15564 11736 15576 11912
rect 15610 11736 15622 11912
rect 15564 11724 15622 11736
rect 15682 11912 15740 11924
rect 15682 11736 15694 11912
rect 15728 11736 15740 11912
rect 15682 11724 15740 11736
rect 16264 11912 16322 11924
rect 16264 11736 16276 11912
rect 16310 11736 16322 11912
rect 16264 11724 16322 11736
rect 16382 11912 16440 11924
rect 16382 11736 16394 11912
rect 16428 11736 16440 11912
rect 16382 11724 16440 11736
rect 16500 11912 16558 11924
rect 16500 11736 16512 11912
rect 16546 11736 16558 11912
rect 16500 11724 16558 11736
rect 16618 11912 16676 11924
rect 16618 11736 16630 11912
rect 16664 11736 16676 11912
rect 16618 11724 16676 11736
rect 16737 11736 16749 12112
rect 16783 11736 16795 12112
rect 16737 11724 16795 11736
rect 16855 12112 16913 12124
rect 16855 11736 16867 12112
rect 16901 11736 16913 12112
rect 16855 11724 16913 11736
rect 16973 12112 17031 12124
rect 16973 11736 16985 12112
rect 17019 11736 17031 12112
rect 16973 11724 17031 11736
rect 17091 12112 17149 12124
rect 17091 11736 17103 12112
rect 17137 11736 17149 12112
rect 17091 11724 17149 11736
rect 17210 12112 17268 12124
rect 17210 11736 17222 12112
rect 17256 11736 17268 12112
rect 17210 11724 17268 11736
rect 17328 12112 17386 12124
rect 17328 11736 17340 12112
rect 17374 11736 17386 12112
rect 17328 11724 17386 11736
rect 17446 12112 17504 12124
rect 17446 11736 17458 12112
rect 17492 11736 17504 12112
rect 17446 11724 17504 11736
rect 17564 12112 17622 12124
rect 17564 11736 17576 12112
rect 17610 11736 17622 12112
rect 17564 11724 17622 11736
rect 17682 12112 17740 12124
rect 17682 11736 17694 12112
rect 17728 11736 17740 12112
rect 17682 11724 17740 11736
rect 17800 12112 17858 12124
rect 17800 11736 17812 12112
rect 17846 11736 17858 12112
rect 17800 11724 17858 11736
rect 17918 12112 17976 12124
rect 17918 11736 17930 12112
rect 17964 11736 17976 12112
rect 17918 11724 17976 11736
rect 18031 12112 18089 12124
rect 18031 11736 18043 12112
rect 18077 11736 18089 12112
rect 18031 11724 18089 11736
rect 18149 12112 18207 12124
rect 18149 11736 18161 12112
rect 18195 11736 18207 12112
rect 18149 11724 18207 11736
rect 18267 12112 18325 12124
rect 18267 11736 18279 12112
rect 18313 11736 18325 12112
rect 18267 11724 18325 11736
rect 18385 12112 18443 12124
rect 18385 11736 18397 12112
rect 18431 11924 18443 12112
rect 19869 12108 19927 12120
rect 18431 11912 18530 11924
rect 18431 11736 18484 11912
rect 18518 11736 18530 11912
rect 18385 11724 18530 11736
rect 18590 11912 18648 11924
rect 18590 11736 18602 11912
rect 18636 11736 18648 11912
rect 18590 11724 18648 11736
rect 18708 11912 18766 11924
rect 18708 11736 18720 11912
rect 18754 11736 18766 11912
rect 18708 11724 18766 11736
rect 18826 11912 18884 11924
rect 18826 11736 18838 11912
rect 18872 11736 18884 11912
rect 18826 11724 18884 11736
rect 19396 11908 19454 11920
rect 19396 11732 19408 11908
rect 19442 11732 19454 11908
rect 19396 11720 19454 11732
rect 19514 11908 19572 11920
rect 19514 11732 19526 11908
rect 19560 11732 19572 11908
rect 19514 11720 19572 11732
rect 19632 11908 19690 11920
rect 19632 11732 19644 11908
rect 19678 11732 19690 11908
rect 19632 11720 19690 11732
rect 19750 11908 19808 11920
rect 19750 11732 19762 11908
rect 19796 11732 19808 11908
rect 19750 11720 19808 11732
rect 19869 11732 19881 12108
rect 19915 11732 19927 12108
rect 19869 11720 19927 11732
rect 19987 12108 20045 12120
rect 19987 11732 19999 12108
rect 20033 11732 20045 12108
rect 19987 11720 20045 11732
rect 20105 12108 20163 12120
rect 20105 11732 20117 12108
rect 20151 11732 20163 12108
rect 20105 11720 20163 11732
rect 20223 12108 20281 12120
rect 20223 11732 20235 12108
rect 20269 11732 20281 12108
rect 20223 11720 20281 11732
rect 20342 12108 20400 12120
rect 20342 11732 20354 12108
rect 20388 11732 20400 12108
rect 20342 11720 20400 11732
rect 20460 12108 20518 12120
rect 20460 11732 20472 12108
rect 20506 11732 20518 12108
rect 20460 11720 20518 11732
rect 20578 12108 20636 12120
rect 20578 11732 20590 12108
rect 20624 11732 20636 12108
rect 20578 11720 20636 11732
rect 20696 12108 20754 12120
rect 20696 11732 20708 12108
rect 20742 11732 20754 12108
rect 20696 11720 20754 11732
rect 20814 12108 20872 12120
rect 20814 11732 20826 12108
rect 20860 11732 20872 12108
rect 20814 11720 20872 11732
rect 20932 12108 20990 12120
rect 20932 11732 20944 12108
rect 20978 11732 20990 12108
rect 20932 11720 20990 11732
rect 21050 12108 21108 12120
rect 21050 11732 21062 12108
rect 21096 11732 21108 12108
rect 21050 11720 21108 11732
rect 21163 12108 21221 12120
rect 21163 11732 21175 12108
rect 21209 11732 21221 12108
rect 21163 11720 21221 11732
rect 21281 12108 21339 12120
rect 21281 11732 21293 12108
rect 21327 11732 21339 12108
rect 21281 11720 21339 11732
rect 21399 12108 21457 12120
rect 21399 11732 21411 12108
rect 21445 11732 21457 12108
rect 21399 11720 21457 11732
rect 21517 12108 21575 12120
rect 21517 11732 21529 12108
rect 21563 11920 21575 12108
rect 23013 12108 23071 12120
rect 21563 11908 21662 11920
rect 21563 11732 21616 11908
rect 21650 11732 21662 11908
rect 21517 11720 21662 11732
rect 21722 11908 21780 11920
rect 21722 11732 21734 11908
rect 21768 11732 21780 11908
rect 21722 11720 21780 11732
rect 21840 11908 21898 11920
rect 21840 11732 21852 11908
rect 21886 11732 21898 11908
rect 21840 11720 21898 11732
rect 21958 11908 22016 11920
rect 21958 11732 21970 11908
rect 22004 11732 22016 11908
rect 21958 11720 22016 11732
rect 22540 11908 22598 11920
rect 22540 11732 22552 11908
rect 22586 11732 22598 11908
rect 22540 11720 22598 11732
rect 22658 11908 22716 11920
rect 22658 11732 22670 11908
rect 22704 11732 22716 11908
rect 22658 11720 22716 11732
rect 22776 11908 22834 11920
rect 22776 11732 22788 11908
rect 22822 11732 22834 11908
rect 22776 11720 22834 11732
rect 22894 11908 22952 11920
rect 22894 11732 22906 11908
rect 22940 11732 22952 11908
rect 22894 11720 22952 11732
rect 23013 11732 23025 12108
rect 23059 11732 23071 12108
rect 23013 11720 23071 11732
rect 23131 12108 23189 12120
rect 23131 11732 23143 12108
rect 23177 11732 23189 12108
rect 23131 11720 23189 11732
rect 23249 12108 23307 12120
rect 23249 11732 23261 12108
rect 23295 11732 23307 12108
rect 23249 11720 23307 11732
rect 23367 12108 23425 12120
rect 23367 11732 23379 12108
rect 23413 11732 23425 12108
rect 23367 11720 23425 11732
rect 23486 12108 23544 12120
rect 23486 11732 23498 12108
rect 23532 11732 23544 12108
rect 23486 11720 23544 11732
rect 23604 12108 23662 12120
rect 23604 11732 23616 12108
rect 23650 11732 23662 12108
rect 23604 11720 23662 11732
rect 23722 12108 23780 12120
rect 23722 11732 23734 12108
rect 23768 11732 23780 12108
rect 23722 11720 23780 11732
rect 23840 12108 23898 12120
rect 23840 11732 23852 12108
rect 23886 11732 23898 12108
rect 23840 11720 23898 11732
rect 23958 12108 24016 12120
rect 23958 11732 23970 12108
rect 24004 11732 24016 12108
rect 23958 11720 24016 11732
rect 24076 12108 24134 12120
rect 24076 11732 24088 12108
rect 24122 11732 24134 12108
rect 24076 11720 24134 11732
rect 24194 12108 24252 12120
rect 24194 11732 24206 12108
rect 24240 11732 24252 12108
rect 24194 11720 24252 11732
rect 24307 12108 24365 12120
rect 24307 11732 24319 12108
rect 24353 11732 24365 12108
rect 24307 11720 24365 11732
rect 24425 12108 24483 12120
rect 24425 11732 24437 12108
rect 24471 11732 24483 12108
rect 24425 11720 24483 11732
rect 24543 12108 24601 12120
rect 24543 11732 24555 12108
rect 24589 11732 24601 12108
rect 24543 11720 24601 11732
rect 24661 12108 24719 12120
rect 24661 11732 24673 12108
rect 24707 11920 24719 12108
rect 29954 12212 30354 12224
rect 29954 12178 29966 12212
rect 30342 12178 30354 12212
rect 29954 12166 30354 12178
rect 29954 12094 30354 12106
rect 29954 12060 29966 12094
rect 30342 12060 30354 12094
rect 29954 12048 30354 12060
rect 30647 12269 31047 12281
rect 30647 12235 30659 12269
rect 31035 12235 31047 12269
rect 30647 12223 31047 12235
rect 70709 12405 70909 12417
rect 70709 12371 70721 12405
rect 70897 12371 70909 12405
rect 70709 12359 70909 12371
rect 30647 12151 31047 12163
rect 30647 12117 30659 12151
rect 31035 12117 31047 12151
rect 30647 12105 31047 12117
rect 41558 12137 41616 12149
rect 29954 11976 30354 11988
rect 29954 11942 29966 11976
rect 30342 11942 30354 11976
rect 29954 11930 30354 11942
rect 24707 11908 24806 11920
rect 24707 11732 24760 11908
rect 24794 11732 24806 11908
rect 24661 11720 24806 11732
rect 24866 11908 24924 11920
rect 24866 11732 24878 11908
rect 24912 11732 24924 11908
rect 24866 11720 24924 11732
rect 24984 11908 25042 11920
rect 24984 11732 24996 11908
rect 25030 11732 25042 11908
rect 24984 11720 25042 11732
rect 25102 11908 25160 11920
rect 25102 11732 25114 11908
rect 25148 11732 25160 11908
rect 30154 11847 30354 11859
rect 30154 11813 30166 11847
rect 30342 11813 30354 11847
rect 30154 11801 30354 11813
rect 30647 12033 31047 12045
rect 30647 11999 30659 12033
rect 31035 11999 31047 12033
rect 30647 11987 31047 11999
rect 41558 11961 41570 12137
rect 41604 11961 41616 12137
rect 41558 11949 41616 11961
rect 41676 12137 41734 12149
rect 41676 11961 41688 12137
rect 41722 11961 41734 12137
rect 41676 11949 41734 11961
rect 41794 12137 41852 12149
rect 41794 11961 41806 12137
rect 41840 11961 41852 12137
rect 41794 11949 41852 11961
rect 41912 12137 41970 12149
rect 41912 11961 41924 12137
rect 41958 11961 41970 12137
rect 41912 11949 41970 11961
rect 42030 12137 42088 12149
rect 42030 11961 42042 12137
rect 42076 11961 42088 12137
rect 42030 11949 42088 11961
rect 42148 12137 42206 12149
rect 42148 11961 42160 12137
rect 42194 11961 42206 12137
rect 42148 11949 42206 11961
rect 42266 12137 42324 12149
rect 42266 11961 42278 12137
rect 42312 11961 42324 12137
rect 42266 11949 42324 11961
rect 42384 12137 42442 12149
rect 42384 11961 42396 12137
rect 42430 11961 42442 12137
rect 42384 11949 42442 11961
rect 42502 12137 42560 12149
rect 42502 11961 42514 12137
rect 42548 11961 42560 12137
rect 42502 11949 42560 11961
rect 42620 12137 42678 12149
rect 54761 12157 54819 12169
rect 42620 11961 42632 12137
rect 42666 11961 42678 12137
rect 42620 11949 42678 11961
rect 48107 12136 48165 12148
rect 48107 11960 48119 12136
rect 48153 11960 48165 12136
rect 25102 11720 25160 11732
rect 30154 11729 30354 11741
rect 30154 11695 30166 11729
rect 30342 11695 30354 11729
rect 48107 11948 48165 11960
rect 48225 12136 48283 12148
rect 48225 11960 48237 12136
rect 48271 11960 48283 12136
rect 48225 11948 48283 11960
rect 48343 12136 48401 12148
rect 48343 11960 48355 12136
rect 48389 11960 48401 12136
rect 48343 11948 48401 11960
rect 48461 12136 48519 12148
rect 48461 11960 48473 12136
rect 48507 11960 48519 12136
rect 48461 11948 48519 11960
rect 48579 12136 48637 12148
rect 48579 11960 48591 12136
rect 48625 11960 48637 12136
rect 48579 11948 48637 11960
rect 48697 12136 48755 12148
rect 48697 11960 48709 12136
rect 48743 11960 48755 12136
rect 48697 11948 48755 11960
rect 48815 12136 48873 12148
rect 48815 11960 48827 12136
rect 48861 11960 48873 12136
rect 48815 11948 48873 11960
rect 48933 12136 48991 12148
rect 48933 11960 48945 12136
rect 48979 11960 48991 12136
rect 48933 11948 48991 11960
rect 49051 12136 49109 12148
rect 49051 11960 49063 12136
rect 49097 11960 49109 12136
rect 49051 11948 49109 11960
rect 49169 12136 49227 12148
rect 49169 11960 49181 12136
rect 49215 11960 49227 12136
rect 54761 11981 54773 12157
rect 54807 11981 54819 12157
rect 54761 11969 54819 11981
rect 54879 12157 54937 12169
rect 54879 11981 54891 12157
rect 54925 11981 54937 12157
rect 54879 11969 54937 11981
rect 54997 12157 55055 12169
rect 54997 11981 55009 12157
rect 55043 11981 55055 12157
rect 54997 11969 55055 11981
rect 55115 12157 55173 12169
rect 55115 11981 55127 12157
rect 55161 11981 55173 12157
rect 55115 11969 55173 11981
rect 55233 12157 55291 12169
rect 55233 11981 55245 12157
rect 55279 11981 55291 12157
rect 55233 11969 55291 11981
rect 55351 12157 55409 12169
rect 55351 11981 55363 12157
rect 55397 11981 55409 12157
rect 55351 11969 55409 11981
rect 55469 12157 55527 12169
rect 55469 11981 55481 12157
rect 55515 11981 55527 12157
rect 55469 11969 55527 11981
rect 55587 12157 55645 12169
rect 55587 11981 55599 12157
rect 55633 11981 55645 12157
rect 55587 11969 55645 11981
rect 55705 12157 55763 12169
rect 55705 11981 55717 12157
rect 55751 11981 55763 12157
rect 55705 11969 55763 11981
rect 55823 12157 55881 12169
rect 55823 11981 55835 12157
rect 55869 11981 55881 12157
rect 70709 12287 70909 12299
rect 70709 12253 70721 12287
rect 70897 12253 70909 12287
rect 70709 12212 70909 12253
rect 70509 12200 70909 12212
rect 70509 12166 70521 12200
rect 70897 12166 70909 12200
rect 70509 12154 70909 12166
rect 70509 12082 70909 12094
rect 70509 12048 70521 12082
rect 70897 12048 70909 12082
rect 70509 12036 70909 12048
rect 55823 11969 55881 11981
rect 63414 11990 63472 12002
rect 49169 11948 49227 11960
rect 30154 11683 30354 11695
rect 30154 11611 30354 11623
rect 30154 11577 30166 11611
rect 30342 11577 30354 11611
rect 30154 11565 30354 11577
rect 30154 11493 30354 11505
rect 30154 11459 30166 11493
rect 30342 11459 30354 11493
rect 30154 11447 30354 11459
rect 63414 11814 63426 11990
rect 63460 11814 63472 11990
rect 63414 11802 63472 11814
rect 63532 11990 63590 12002
rect 63532 11814 63544 11990
rect 63578 11814 63590 11990
rect 63532 11802 63590 11814
rect 63650 11990 63708 12002
rect 63650 11814 63662 11990
rect 63696 11814 63708 11990
rect 63650 11802 63708 11814
rect 63768 11990 63826 12002
rect 63768 11814 63780 11990
rect 63814 11814 63826 11990
rect 63768 11802 63826 11814
rect 63886 11990 63944 12002
rect 63886 11814 63898 11990
rect 63932 11814 63944 11990
rect 63886 11802 63944 11814
rect 64004 11990 64062 12002
rect 64004 11814 64016 11990
rect 64050 11814 64062 11990
rect 64004 11802 64062 11814
rect 64122 11990 64180 12002
rect 64122 11814 64134 11990
rect 64168 11814 64180 11990
rect 64122 11802 64180 11814
rect 64240 11990 64298 12002
rect 64240 11814 64252 11990
rect 64286 11814 64298 11990
rect 64240 11802 64298 11814
rect 64358 11990 64416 12002
rect 64358 11814 64370 11990
rect 64404 11814 64416 11990
rect 64358 11802 64416 11814
rect 64476 11990 64534 12002
rect 64476 11814 64488 11990
rect 64522 11814 64534 11990
rect 70509 11964 70909 11976
rect 70509 11930 70521 11964
rect 70897 11930 70909 11964
rect 70509 11918 70909 11930
rect 64476 11802 64534 11814
rect 65706 11785 65764 11797
rect 65222 11585 65280 11597
rect 30152 11100 30352 11112
rect 30152 11066 30164 11100
rect 30340 11066 30352 11100
rect 30152 11054 30352 11066
rect 65222 11409 65234 11585
rect 65268 11409 65280 11585
rect 65222 11397 65280 11409
rect 65340 11585 65398 11597
rect 65340 11409 65352 11585
rect 65386 11409 65398 11585
rect 65340 11397 65398 11409
rect 65458 11585 65516 11597
rect 65458 11409 65470 11585
rect 65504 11409 65516 11585
rect 65458 11397 65516 11409
rect 65576 11585 65634 11597
rect 65576 11409 65588 11585
rect 65622 11409 65634 11585
rect 65576 11397 65634 11409
rect 65706 11409 65718 11785
rect 65752 11409 65764 11785
rect 65706 11397 65764 11409
rect 65824 11785 65882 11797
rect 65824 11409 65836 11785
rect 65870 11409 65882 11785
rect 65824 11397 65882 11409
rect 65942 11785 66000 11797
rect 65942 11409 65954 11785
rect 65988 11409 66000 11785
rect 65942 11397 66000 11409
rect 66060 11785 66118 11797
rect 66060 11409 66072 11785
rect 66106 11409 66118 11785
rect 66060 11397 66118 11409
rect 66178 11785 66236 11797
rect 66178 11409 66190 11785
rect 66224 11409 66236 11785
rect 66178 11397 66236 11409
rect 66296 11785 66354 11797
rect 66296 11409 66308 11785
rect 66342 11409 66354 11785
rect 66296 11397 66354 11409
rect 66414 11785 66472 11797
rect 66414 11409 66426 11785
rect 66460 11409 66472 11785
rect 70509 11846 70909 11858
rect 70509 11812 70521 11846
rect 70897 11812 70909 11846
rect 70509 11800 70909 11812
rect 70509 11733 70909 11745
rect 70509 11699 70521 11733
rect 70897 11699 70909 11733
rect 70509 11687 70909 11699
rect 66414 11397 66472 11409
rect 66543 11585 66601 11597
rect 66543 11409 66555 11585
rect 66589 11409 66601 11585
rect 66543 11397 66601 11409
rect 66661 11585 66719 11597
rect 66661 11409 66673 11585
rect 66707 11409 66719 11585
rect 66661 11397 66719 11409
rect 66779 11585 66837 11597
rect 66779 11409 66791 11585
rect 66825 11409 66837 11585
rect 66779 11397 66837 11409
rect 66897 11585 66955 11597
rect 66897 11409 66909 11585
rect 66943 11409 66955 11585
rect 66897 11397 66955 11409
rect 67015 11582 67073 11594
rect 67015 11406 67027 11582
rect 67061 11406 67073 11582
rect 67015 11394 67073 11406
rect 67133 11582 67191 11594
rect 67133 11406 67145 11582
rect 67179 11406 67191 11582
rect 67133 11394 67191 11406
rect 67251 11582 67309 11594
rect 67251 11406 67263 11582
rect 67297 11406 67309 11582
rect 67251 11394 67309 11406
rect 67369 11582 67427 11594
rect 67369 11406 67381 11582
rect 67415 11406 67427 11582
rect 67369 11394 67427 11406
rect 67487 11582 67545 11594
rect 67487 11406 67499 11582
rect 67533 11406 67545 11582
rect 67487 11394 67545 11406
rect 67605 11582 67663 11594
rect 67605 11406 67617 11582
rect 67651 11406 67663 11582
rect 67605 11394 67663 11406
rect 67723 11582 67781 11594
rect 67723 11406 67735 11582
rect 67769 11406 67781 11582
rect 67723 11394 67781 11406
rect 67841 11582 67899 11594
rect 67841 11406 67853 11582
rect 67887 11406 67899 11582
rect 67841 11394 67899 11406
rect 67959 11582 68017 11594
rect 67959 11406 67971 11582
rect 68005 11406 68017 11582
rect 67959 11394 68017 11406
rect 68077 11582 68135 11594
rect 68077 11406 68089 11582
rect 68123 11406 68135 11582
rect 70509 11615 70909 11627
rect 70509 11581 70521 11615
rect 70897 11581 70909 11615
rect 70509 11569 70909 11581
rect 68077 11394 68135 11406
rect 30152 10982 30352 10994
rect 30152 10948 30164 10982
rect 30340 10948 30352 10982
rect 30152 10936 30352 10948
rect 65649 11092 65707 11104
rect 30152 10864 30352 10876
rect 30152 10830 30164 10864
rect 30340 10830 30352 10864
rect 30152 10818 30352 10830
rect 30152 10746 30352 10758
rect 30152 10712 30164 10746
rect 30340 10712 30352 10746
rect 30152 10700 30352 10712
rect 29952 10616 30352 10628
rect 29952 10582 29964 10616
rect 30340 10582 30352 10616
rect 29952 10570 30352 10582
rect 30645 10673 31045 10685
rect 30645 10639 30657 10673
rect 31033 10639 31045 10673
rect 30645 10627 31045 10639
rect 29952 10498 30352 10510
rect 29952 10464 29964 10498
rect 30340 10464 30352 10498
rect 29952 10452 30352 10464
rect 30645 10555 31045 10567
rect 30645 10521 30657 10555
rect 31033 10521 31045 10555
rect 30645 10509 31045 10521
rect 29952 10380 30352 10392
rect 29952 10346 29964 10380
rect 30340 10346 30352 10380
rect 29952 10334 30352 10346
rect 30645 10437 31045 10449
rect 30645 10403 30657 10437
rect 31033 10403 31045 10437
rect 30645 10391 31045 10403
rect 30645 10319 31045 10331
rect 30645 10285 30657 10319
rect 31033 10285 31045 10319
rect 29952 10262 30352 10274
rect 30645 10273 31045 10285
rect 29952 10228 29964 10262
rect 30340 10228 30352 10262
rect 29952 10216 30352 10228
rect 29952 10144 30352 10156
rect 29952 10110 29964 10144
rect 30340 10110 30352 10144
rect 29952 10098 30352 10110
rect 29952 10026 30352 10038
rect 29952 9992 29964 10026
rect 30340 9992 30352 10026
rect 29952 9980 30352 9992
rect 30645 10201 31045 10213
rect 30645 10167 30657 10201
rect 31033 10167 31045 10201
rect 30645 10155 31045 10167
rect 34894 10237 34952 10249
rect 30645 10083 31045 10095
rect 30645 10049 30657 10083
rect 31033 10049 31045 10083
rect 30645 10037 31045 10049
rect 34894 10061 34906 10237
rect 34940 10061 34952 10237
rect 34894 10049 34952 10061
rect 35012 10237 35070 10249
rect 35012 10061 35024 10237
rect 35058 10061 35070 10237
rect 35012 10049 35070 10061
rect 35130 10237 35188 10249
rect 35130 10061 35142 10237
rect 35176 10061 35188 10237
rect 35130 10049 35188 10061
rect 35248 10237 35306 10249
rect 35248 10061 35260 10237
rect 35294 10061 35306 10237
rect 35248 10049 35306 10061
rect 35366 10237 35424 10249
rect 35366 10061 35378 10237
rect 35412 10061 35424 10237
rect 35366 10049 35424 10061
rect 35484 10237 35542 10249
rect 35484 10061 35496 10237
rect 35530 10061 35542 10237
rect 35484 10049 35542 10061
rect 35602 10237 35660 10249
rect 35602 10061 35614 10237
rect 35648 10061 35660 10237
rect 35602 10049 35660 10061
rect 35720 10237 35778 10249
rect 35720 10061 35732 10237
rect 35766 10061 35778 10237
rect 35720 10049 35778 10061
rect 35838 10237 35896 10249
rect 35838 10061 35850 10237
rect 35884 10061 35896 10237
rect 35838 10049 35896 10061
rect 35956 10237 36014 10249
rect 35956 10061 35968 10237
rect 36002 10061 36014 10237
rect 65649 10716 65661 11092
rect 65695 10716 65707 11092
rect 65649 10704 65707 10716
rect 65767 11092 65825 11104
rect 65767 10716 65779 11092
rect 65813 10716 65825 11092
rect 65767 10704 65825 10716
rect 65885 11092 65943 11104
rect 65885 10716 65897 11092
rect 65931 10716 65943 11092
rect 65885 10704 65943 10716
rect 66003 11092 66061 11104
rect 66003 10716 66015 11092
rect 66049 10716 66061 11092
rect 66003 10704 66061 10716
rect 66121 11092 66179 11104
rect 66121 10716 66133 11092
rect 66167 10716 66179 11092
rect 66121 10704 66179 10716
rect 66239 11092 66297 11104
rect 66239 10716 66251 11092
rect 66285 10716 66297 11092
rect 66239 10704 66297 10716
rect 66357 11092 66415 11104
rect 66357 10716 66369 11092
rect 66403 10716 66415 11092
rect 66357 10704 66415 10716
rect 70509 11497 70909 11509
rect 70509 11463 70521 11497
rect 70897 11463 70909 11497
rect 70509 11451 70909 11463
rect 70509 11379 70909 11391
rect 70509 11345 70521 11379
rect 70897 11345 70909 11379
rect 70509 11333 70909 11345
rect 70509 11261 70909 11273
rect 70509 11227 70521 11261
rect 70897 11227 70909 11261
rect 70509 11215 70909 11227
rect 70509 11143 70909 11155
rect 70509 11109 70521 11143
rect 70897 11109 70909 11143
rect 70509 11097 70909 11109
rect 70509 11025 70909 11037
rect 70509 10991 70521 11025
rect 70897 10991 70909 11025
rect 70509 10979 70909 10991
rect 70509 10906 70909 10918
rect 70509 10872 70521 10906
rect 70897 10872 70909 10906
rect 70509 10860 70909 10872
rect 70509 10788 70909 10800
rect 70509 10754 70521 10788
rect 70897 10754 70909 10788
rect 70509 10742 70909 10754
rect 70509 10670 70909 10682
rect 70509 10636 70521 10670
rect 70897 10636 70909 10670
rect 70509 10624 70909 10636
rect 70509 10552 70909 10564
rect 70509 10518 70521 10552
rect 70897 10518 70909 10552
rect 70509 10506 70909 10518
rect 70709 10433 70909 10445
rect 70709 10399 70721 10433
rect 70897 10399 70909 10433
rect 70709 10387 70909 10399
rect 46658 10130 46716 10142
rect 35956 10049 36014 10061
rect 44333 10058 44391 10070
rect 29952 9908 30352 9920
rect 29952 9874 29964 9908
rect 30340 9874 30352 9908
rect 29952 9862 30352 9874
rect 30152 9779 30352 9791
rect 30152 9745 30164 9779
rect 30340 9745 30352 9779
rect 30152 9733 30352 9745
rect 30645 9965 31045 9977
rect 30645 9931 30657 9965
rect 31033 9931 31045 9965
rect 30645 9919 31045 9931
rect 40109 10042 40167 10054
rect 37784 9970 37842 9982
rect 30152 9661 30352 9673
rect 30152 9627 30164 9661
rect 30340 9627 30352 9661
rect 30152 9615 30352 9627
rect 30152 9543 30352 9555
rect 30152 9509 30164 9543
rect 30340 9509 30352 9543
rect 30152 9497 30352 9509
rect 981 9380 1039 9392
rect 508 9180 566 9192
rect 508 9004 520 9180
rect 554 9004 566 9180
rect 508 8992 566 9004
rect 626 9180 684 9192
rect 626 9004 638 9180
rect 672 9004 684 9180
rect 626 8992 684 9004
rect 744 9180 802 9192
rect 744 9004 756 9180
rect 790 9004 802 9180
rect 744 8992 802 9004
rect 862 9180 920 9192
rect 862 9004 874 9180
rect 908 9004 920 9180
rect 862 8992 920 9004
rect 981 9004 993 9380
rect 1027 9004 1039 9380
rect 981 8992 1039 9004
rect 1099 9380 1157 9392
rect 1099 9004 1111 9380
rect 1145 9004 1157 9380
rect 1099 8992 1157 9004
rect 1217 9380 1275 9392
rect 1217 9004 1229 9380
rect 1263 9004 1275 9380
rect 1217 8992 1275 9004
rect 1335 9380 1393 9392
rect 1335 9004 1347 9380
rect 1381 9004 1393 9380
rect 1335 8992 1393 9004
rect 1454 9380 1512 9392
rect 1454 9004 1466 9380
rect 1500 9004 1512 9380
rect 1454 8992 1512 9004
rect 1572 9380 1630 9392
rect 1572 9004 1584 9380
rect 1618 9004 1630 9380
rect 1572 8992 1630 9004
rect 1690 9380 1748 9392
rect 1690 9004 1702 9380
rect 1736 9004 1748 9380
rect 1690 8992 1748 9004
rect 1808 9380 1866 9392
rect 1808 9004 1820 9380
rect 1854 9004 1866 9380
rect 1808 8992 1866 9004
rect 1926 9380 1984 9392
rect 1926 9004 1938 9380
rect 1972 9004 1984 9380
rect 1926 8992 1984 9004
rect 2044 9380 2102 9392
rect 2044 9004 2056 9380
rect 2090 9004 2102 9380
rect 2044 8992 2102 9004
rect 2162 9380 2220 9392
rect 2162 9004 2174 9380
rect 2208 9004 2220 9380
rect 2162 8992 2220 9004
rect 2275 9380 2333 9392
rect 2275 9004 2287 9380
rect 2321 9004 2333 9380
rect 2275 8992 2333 9004
rect 2393 9380 2451 9392
rect 2393 9004 2405 9380
rect 2439 9004 2451 9380
rect 2393 8992 2451 9004
rect 2511 9380 2569 9392
rect 2511 9004 2523 9380
rect 2557 9004 2569 9380
rect 2511 8992 2569 9004
rect 2629 9380 2687 9392
rect 2629 9004 2641 9380
rect 2675 9192 2687 9380
rect 4125 9380 4183 9392
rect 2675 9180 2774 9192
rect 2675 9004 2728 9180
rect 2762 9004 2774 9180
rect 2629 8992 2774 9004
rect 2834 9180 2892 9192
rect 2834 9004 2846 9180
rect 2880 9004 2892 9180
rect 2834 8992 2892 9004
rect 2952 9180 3010 9192
rect 2952 9004 2964 9180
rect 2998 9004 3010 9180
rect 2952 8992 3010 9004
rect 3070 9180 3128 9192
rect 3070 9004 3082 9180
rect 3116 9004 3128 9180
rect 3070 8992 3128 9004
rect 3652 9180 3710 9192
rect 3652 9004 3664 9180
rect 3698 9004 3710 9180
rect 3652 8992 3710 9004
rect 3770 9180 3828 9192
rect 3770 9004 3782 9180
rect 3816 9004 3828 9180
rect 3770 8992 3828 9004
rect 3888 9180 3946 9192
rect 3888 9004 3900 9180
rect 3934 9004 3946 9180
rect 3888 8992 3946 9004
rect 4006 9180 4064 9192
rect 4006 9004 4018 9180
rect 4052 9004 4064 9180
rect 4006 8992 4064 9004
rect 4125 9004 4137 9380
rect 4171 9004 4183 9380
rect 4125 8992 4183 9004
rect 4243 9380 4301 9392
rect 4243 9004 4255 9380
rect 4289 9004 4301 9380
rect 4243 8992 4301 9004
rect 4361 9380 4419 9392
rect 4361 9004 4373 9380
rect 4407 9004 4419 9380
rect 4361 8992 4419 9004
rect 4479 9380 4537 9392
rect 4479 9004 4491 9380
rect 4525 9004 4537 9380
rect 4479 8992 4537 9004
rect 4598 9380 4656 9392
rect 4598 9004 4610 9380
rect 4644 9004 4656 9380
rect 4598 8992 4656 9004
rect 4716 9380 4774 9392
rect 4716 9004 4728 9380
rect 4762 9004 4774 9380
rect 4716 8992 4774 9004
rect 4834 9380 4892 9392
rect 4834 9004 4846 9380
rect 4880 9004 4892 9380
rect 4834 8992 4892 9004
rect 4952 9380 5010 9392
rect 4952 9004 4964 9380
rect 4998 9004 5010 9380
rect 4952 8992 5010 9004
rect 5070 9380 5128 9392
rect 5070 9004 5082 9380
rect 5116 9004 5128 9380
rect 5070 8992 5128 9004
rect 5188 9380 5246 9392
rect 5188 9004 5200 9380
rect 5234 9004 5246 9380
rect 5188 8992 5246 9004
rect 5306 9380 5364 9392
rect 5306 9004 5318 9380
rect 5352 9004 5364 9380
rect 5306 8992 5364 9004
rect 5419 9380 5477 9392
rect 5419 9004 5431 9380
rect 5465 9004 5477 9380
rect 5419 8992 5477 9004
rect 5537 9380 5595 9392
rect 5537 9004 5549 9380
rect 5583 9004 5595 9380
rect 5537 8992 5595 9004
rect 5655 9380 5713 9392
rect 5655 9004 5667 9380
rect 5701 9004 5713 9380
rect 5655 8992 5713 9004
rect 5773 9380 5831 9392
rect 5773 9004 5785 9380
rect 5819 9192 5831 9380
rect 7257 9376 7315 9388
rect 5819 9180 5918 9192
rect 5819 9004 5872 9180
rect 5906 9004 5918 9180
rect 5773 8992 5918 9004
rect 5978 9180 6036 9192
rect 5978 9004 5990 9180
rect 6024 9004 6036 9180
rect 5978 8992 6036 9004
rect 6096 9180 6154 9192
rect 6096 9004 6108 9180
rect 6142 9004 6154 9180
rect 6096 8992 6154 9004
rect 6214 9180 6272 9192
rect 6214 9004 6226 9180
rect 6260 9004 6272 9180
rect 6214 8992 6272 9004
rect 6784 9176 6842 9188
rect 6784 9000 6796 9176
rect 6830 9000 6842 9176
rect 6784 8988 6842 9000
rect 6902 9176 6960 9188
rect 6902 9000 6914 9176
rect 6948 9000 6960 9176
rect 6902 8988 6960 9000
rect 7020 9176 7078 9188
rect 7020 9000 7032 9176
rect 7066 9000 7078 9176
rect 7020 8988 7078 9000
rect 7138 9176 7196 9188
rect 7138 9000 7150 9176
rect 7184 9000 7196 9176
rect 7138 8988 7196 9000
rect 7257 9000 7269 9376
rect 7303 9000 7315 9376
rect 7257 8988 7315 9000
rect 7375 9376 7433 9388
rect 7375 9000 7387 9376
rect 7421 9000 7433 9376
rect 7375 8988 7433 9000
rect 7493 9376 7551 9388
rect 7493 9000 7505 9376
rect 7539 9000 7551 9376
rect 7493 8988 7551 9000
rect 7611 9376 7669 9388
rect 7611 9000 7623 9376
rect 7657 9000 7669 9376
rect 7611 8988 7669 9000
rect 7730 9376 7788 9388
rect 7730 9000 7742 9376
rect 7776 9000 7788 9376
rect 7730 8988 7788 9000
rect 7848 9376 7906 9388
rect 7848 9000 7860 9376
rect 7894 9000 7906 9376
rect 7848 8988 7906 9000
rect 7966 9376 8024 9388
rect 7966 9000 7978 9376
rect 8012 9000 8024 9376
rect 7966 8988 8024 9000
rect 8084 9376 8142 9388
rect 8084 9000 8096 9376
rect 8130 9000 8142 9376
rect 8084 8988 8142 9000
rect 8202 9376 8260 9388
rect 8202 9000 8214 9376
rect 8248 9000 8260 9376
rect 8202 8988 8260 9000
rect 8320 9376 8378 9388
rect 8320 9000 8332 9376
rect 8366 9000 8378 9376
rect 8320 8988 8378 9000
rect 8438 9376 8496 9388
rect 8438 9000 8450 9376
rect 8484 9000 8496 9376
rect 8438 8988 8496 9000
rect 8551 9376 8609 9388
rect 8551 9000 8563 9376
rect 8597 9000 8609 9376
rect 8551 8988 8609 9000
rect 8669 9376 8727 9388
rect 8669 9000 8681 9376
rect 8715 9000 8727 9376
rect 8669 8988 8727 9000
rect 8787 9376 8845 9388
rect 8787 9000 8799 9376
rect 8833 9000 8845 9376
rect 8787 8988 8845 9000
rect 8905 9376 8963 9388
rect 8905 9000 8917 9376
rect 8951 9188 8963 9376
rect 10401 9376 10459 9388
rect 8951 9176 9050 9188
rect 8951 9000 9004 9176
rect 9038 9000 9050 9176
rect 8905 8988 9050 9000
rect 9110 9176 9168 9188
rect 9110 9000 9122 9176
rect 9156 9000 9168 9176
rect 9110 8988 9168 9000
rect 9228 9176 9286 9188
rect 9228 9000 9240 9176
rect 9274 9000 9286 9176
rect 9228 8988 9286 9000
rect 9346 9176 9404 9188
rect 9346 9000 9358 9176
rect 9392 9000 9404 9176
rect 9346 8988 9404 9000
rect 9928 9176 9986 9188
rect 9928 9000 9940 9176
rect 9974 9000 9986 9176
rect 9928 8988 9986 9000
rect 10046 9176 10104 9188
rect 10046 9000 10058 9176
rect 10092 9000 10104 9176
rect 10046 8988 10104 9000
rect 10164 9176 10222 9188
rect 10164 9000 10176 9176
rect 10210 9000 10222 9176
rect 10164 8988 10222 9000
rect 10282 9176 10340 9188
rect 10282 9000 10294 9176
rect 10328 9000 10340 9176
rect 10282 8988 10340 9000
rect 10401 9000 10413 9376
rect 10447 9000 10459 9376
rect 10401 8988 10459 9000
rect 10519 9376 10577 9388
rect 10519 9000 10531 9376
rect 10565 9000 10577 9376
rect 10519 8988 10577 9000
rect 10637 9376 10695 9388
rect 10637 9000 10649 9376
rect 10683 9000 10695 9376
rect 10637 8988 10695 9000
rect 10755 9376 10813 9388
rect 10755 9000 10767 9376
rect 10801 9000 10813 9376
rect 10755 8988 10813 9000
rect 10874 9376 10932 9388
rect 10874 9000 10886 9376
rect 10920 9000 10932 9376
rect 10874 8988 10932 9000
rect 10992 9376 11050 9388
rect 10992 9000 11004 9376
rect 11038 9000 11050 9376
rect 10992 8988 11050 9000
rect 11110 9376 11168 9388
rect 11110 9000 11122 9376
rect 11156 9000 11168 9376
rect 11110 8988 11168 9000
rect 11228 9376 11286 9388
rect 11228 9000 11240 9376
rect 11274 9000 11286 9376
rect 11228 8988 11286 9000
rect 11346 9376 11404 9388
rect 11346 9000 11358 9376
rect 11392 9000 11404 9376
rect 11346 8988 11404 9000
rect 11464 9376 11522 9388
rect 11464 9000 11476 9376
rect 11510 9000 11522 9376
rect 11464 8988 11522 9000
rect 11582 9376 11640 9388
rect 11582 9000 11594 9376
rect 11628 9000 11640 9376
rect 11582 8988 11640 9000
rect 11695 9376 11753 9388
rect 11695 9000 11707 9376
rect 11741 9000 11753 9376
rect 11695 8988 11753 9000
rect 11813 9376 11871 9388
rect 11813 9000 11825 9376
rect 11859 9000 11871 9376
rect 11813 8988 11871 9000
rect 11931 9376 11989 9388
rect 11931 9000 11943 9376
rect 11977 9000 11989 9376
rect 11931 8988 11989 9000
rect 12049 9376 12107 9388
rect 12049 9000 12061 9376
rect 12095 9188 12107 9376
rect 13603 9380 13661 9392
rect 12095 9176 12194 9188
rect 12095 9000 12148 9176
rect 12182 9000 12194 9176
rect 12049 8988 12194 9000
rect 12254 9176 12312 9188
rect 12254 9000 12266 9176
rect 12300 9000 12312 9176
rect 12254 8988 12312 9000
rect 12372 9176 12430 9188
rect 12372 9000 12384 9176
rect 12418 9000 12430 9176
rect 12372 8988 12430 9000
rect 12490 9176 12548 9188
rect 12490 9000 12502 9176
rect 12536 9000 12548 9176
rect 12490 8988 12548 9000
rect 13130 9180 13188 9192
rect 13130 9004 13142 9180
rect 13176 9004 13188 9180
rect 13130 8992 13188 9004
rect 13248 9180 13306 9192
rect 13248 9004 13260 9180
rect 13294 9004 13306 9180
rect 13248 8992 13306 9004
rect 13366 9180 13424 9192
rect 13366 9004 13378 9180
rect 13412 9004 13424 9180
rect 13366 8992 13424 9004
rect 13484 9180 13542 9192
rect 13484 9004 13496 9180
rect 13530 9004 13542 9180
rect 13484 8992 13542 9004
rect 13603 9004 13615 9380
rect 13649 9004 13661 9380
rect 13603 8992 13661 9004
rect 13721 9380 13779 9392
rect 13721 9004 13733 9380
rect 13767 9004 13779 9380
rect 13721 8992 13779 9004
rect 13839 9380 13897 9392
rect 13839 9004 13851 9380
rect 13885 9004 13897 9380
rect 13839 8992 13897 9004
rect 13957 9380 14015 9392
rect 13957 9004 13969 9380
rect 14003 9004 14015 9380
rect 13957 8992 14015 9004
rect 14076 9380 14134 9392
rect 14076 9004 14088 9380
rect 14122 9004 14134 9380
rect 14076 8992 14134 9004
rect 14194 9380 14252 9392
rect 14194 9004 14206 9380
rect 14240 9004 14252 9380
rect 14194 8992 14252 9004
rect 14312 9380 14370 9392
rect 14312 9004 14324 9380
rect 14358 9004 14370 9380
rect 14312 8992 14370 9004
rect 14430 9380 14488 9392
rect 14430 9004 14442 9380
rect 14476 9004 14488 9380
rect 14430 8992 14488 9004
rect 14548 9380 14606 9392
rect 14548 9004 14560 9380
rect 14594 9004 14606 9380
rect 14548 8992 14606 9004
rect 14666 9380 14724 9392
rect 14666 9004 14678 9380
rect 14712 9004 14724 9380
rect 14666 8992 14724 9004
rect 14784 9380 14842 9392
rect 14784 9004 14796 9380
rect 14830 9004 14842 9380
rect 14784 8992 14842 9004
rect 14897 9380 14955 9392
rect 14897 9004 14909 9380
rect 14943 9004 14955 9380
rect 14897 8992 14955 9004
rect 15015 9380 15073 9392
rect 15015 9004 15027 9380
rect 15061 9004 15073 9380
rect 15015 8992 15073 9004
rect 15133 9380 15191 9392
rect 15133 9004 15145 9380
rect 15179 9004 15191 9380
rect 15133 8992 15191 9004
rect 15251 9380 15309 9392
rect 15251 9004 15263 9380
rect 15297 9192 15309 9380
rect 16747 9380 16805 9392
rect 15297 9180 15396 9192
rect 15297 9004 15350 9180
rect 15384 9004 15396 9180
rect 15251 8992 15396 9004
rect 15456 9180 15514 9192
rect 15456 9004 15468 9180
rect 15502 9004 15514 9180
rect 15456 8992 15514 9004
rect 15574 9180 15632 9192
rect 15574 9004 15586 9180
rect 15620 9004 15632 9180
rect 15574 8992 15632 9004
rect 15692 9180 15750 9192
rect 15692 9004 15704 9180
rect 15738 9004 15750 9180
rect 15692 8992 15750 9004
rect 16274 9180 16332 9192
rect 16274 9004 16286 9180
rect 16320 9004 16332 9180
rect 16274 8992 16332 9004
rect 16392 9180 16450 9192
rect 16392 9004 16404 9180
rect 16438 9004 16450 9180
rect 16392 8992 16450 9004
rect 16510 9180 16568 9192
rect 16510 9004 16522 9180
rect 16556 9004 16568 9180
rect 16510 8992 16568 9004
rect 16628 9180 16686 9192
rect 16628 9004 16640 9180
rect 16674 9004 16686 9180
rect 16628 8992 16686 9004
rect 16747 9004 16759 9380
rect 16793 9004 16805 9380
rect 16747 8992 16805 9004
rect 16865 9380 16923 9392
rect 16865 9004 16877 9380
rect 16911 9004 16923 9380
rect 16865 8992 16923 9004
rect 16983 9380 17041 9392
rect 16983 9004 16995 9380
rect 17029 9004 17041 9380
rect 16983 8992 17041 9004
rect 17101 9380 17159 9392
rect 17101 9004 17113 9380
rect 17147 9004 17159 9380
rect 17101 8992 17159 9004
rect 17220 9380 17278 9392
rect 17220 9004 17232 9380
rect 17266 9004 17278 9380
rect 17220 8992 17278 9004
rect 17338 9380 17396 9392
rect 17338 9004 17350 9380
rect 17384 9004 17396 9380
rect 17338 8992 17396 9004
rect 17456 9380 17514 9392
rect 17456 9004 17468 9380
rect 17502 9004 17514 9380
rect 17456 8992 17514 9004
rect 17574 9380 17632 9392
rect 17574 9004 17586 9380
rect 17620 9004 17632 9380
rect 17574 8992 17632 9004
rect 17692 9380 17750 9392
rect 17692 9004 17704 9380
rect 17738 9004 17750 9380
rect 17692 8992 17750 9004
rect 17810 9380 17868 9392
rect 17810 9004 17822 9380
rect 17856 9004 17868 9380
rect 17810 8992 17868 9004
rect 17928 9380 17986 9392
rect 17928 9004 17940 9380
rect 17974 9004 17986 9380
rect 17928 8992 17986 9004
rect 18041 9380 18099 9392
rect 18041 9004 18053 9380
rect 18087 9004 18099 9380
rect 18041 8992 18099 9004
rect 18159 9380 18217 9392
rect 18159 9004 18171 9380
rect 18205 9004 18217 9380
rect 18159 8992 18217 9004
rect 18277 9380 18335 9392
rect 18277 9004 18289 9380
rect 18323 9004 18335 9380
rect 18277 8992 18335 9004
rect 18395 9380 18453 9392
rect 30152 9425 30352 9437
rect 30152 9391 30164 9425
rect 30340 9391 30352 9425
rect 37784 9794 37796 9970
rect 37830 9794 37842 9970
rect 37784 9782 37842 9794
rect 37902 9970 37960 9982
rect 37902 9794 37914 9970
rect 37948 9794 37960 9970
rect 37902 9782 37960 9794
rect 38020 9970 38078 9982
rect 38020 9794 38032 9970
rect 38066 9794 38078 9970
rect 38020 9782 38078 9794
rect 38138 9970 38196 9982
rect 38138 9794 38150 9970
rect 38184 9794 38196 9970
rect 38138 9782 38196 9794
rect 38256 9970 38314 9982
rect 38256 9794 38268 9970
rect 38302 9794 38314 9970
rect 38256 9782 38314 9794
rect 38374 9970 38432 9982
rect 38374 9794 38386 9970
rect 38420 9794 38432 9970
rect 38374 9782 38432 9794
rect 38492 9970 38550 9982
rect 38492 9794 38504 9970
rect 38538 9794 38550 9970
rect 38492 9782 38550 9794
rect 38610 9970 38668 9982
rect 38610 9794 38622 9970
rect 38656 9794 38668 9970
rect 38610 9782 38668 9794
rect 38728 9970 38786 9982
rect 38728 9794 38740 9970
rect 38774 9794 38786 9970
rect 38728 9782 38786 9794
rect 38846 9970 38904 9982
rect 38846 9794 38858 9970
rect 38892 9794 38904 9970
rect 38846 9782 38904 9794
rect 40109 9666 40121 10042
rect 40155 9666 40167 10042
rect 40109 9654 40167 9666
rect 40227 10042 40285 10054
rect 40227 9666 40239 10042
rect 40273 9666 40285 10042
rect 40227 9654 40285 9666
rect 40345 10042 40403 10054
rect 40345 9666 40357 10042
rect 40391 9666 40403 10042
rect 40345 9654 40403 9666
rect 40463 10042 40521 10054
rect 40463 9666 40475 10042
rect 40509 9666 40521 10042
rect 40463 9654 40521 9666
rect 40581 10042 40639 10054
rect 40581 9666 40593 10042
rect 40627 9666 40639 10042
rect 40581 9654 40639 9666
rect 40699 10042 40757 10054
rect 40699 9666 40711 10042
rect 40745 9666 40757 10042
rect 40699 9654 40757 9666
rect 40817 10042 40875 10054
rect 40817 9666 40829 10042
rect 40863 9666 40875 10042
rect 40817 9654 40875 9666
rect 41251 10046 41309 10058
rect 41251 9670 41263 10046
rect 41297 9670 41309 10046
rect 41251 9658 41309 9670
rect 41369 10046 41427 10058
rect 41369 9670 41381 10046
rect 41415 9670 41427 10046
rect 41369 9658 41427 9670
rect 41487 10046 41545 10058
rect 41487 9670 41499 10046
rect 41533 9670 41545 10046
rect 41487 9658 41545 9670
rect 41605 10046 41663 10058
rect 41605 9670 41617 10046
rect 41651 9670 41663 10046
rect 41605 9658 41663 9670
rect 41723 10046 41781 10058
rect 41723 9670 41735 10046
rect 41769 9670 41781 10046
rect 41723 9658 41781 9670
rect 41841 10046 41899 10058
rect 41841 9670 41853 10046
rect 41887 9670 41899 10046
rect 41841 9658 41899 9670
rect 41959 10046 42017 10058
rect 41959 9670 41971 10046
rect 42005 9670 42017 10046
rect 44333 9882 44345 10058
rect 44379 9882 44391 10058
rect 44333 9870 44391 9882
rect 44451 10058 44509 10070
rect 44451 9882 44463 10058
rect 44497 9882 44509 10058
rect 44451 9870 44509 9882
rect 44569 10058 44627 10070
rect 44569 9882 44581 10058
rect 44615 9882 44627 10058
rect 44569 9870 44627 9882
rect 44687 10058 44745 10070
rect 44687 9882 44699 10058
rect 44733 9882 44745 10058
rect 44687 9870 44745 9882
rect 44805 10058 44863 10070
rect 44805 9882 44817 10058
rect 44851 9882 44863 10058
rect 44805 9870 44863 9882
rect 44923 10058 44981 10070
rect 44923 9882 44935 10058
rect 44969 9882 44981 10058
rect 44923 9870 44981 9882
rect 45041 10058 45099 10070
rect 45041 9882 45053 10058
rect 45087 9882 45099 10058
rect 45041 9870 45099 9882
rect 45159 10058 45217 10070
rect 45159 9882 45171 10058
rect 45205 9882 45217 10058
rect 45159 9870 45217 9882
rect 45277 10058 45335 10070
rect 45277 9882 45289 10058
rect 45323 9882 45335 10058
rect 45277 9870 45335 9882
rect 45395 10058 45453 10070
rect 45395 9882 45407 10058
rect 45441 9882 45453 10058
rect 45395 9870 45453 9882
rect 41959 9658 42017 9670
rect 18395 9004 18407 9380
rect 18441 9192 18453 9380
rect 19879 9376 19937 9388
rect 18441 9180 18540 9192
rect 18441 9004 18494 9180
rect 18528 9004 18540 9180
rect 18395 8992 18540 9004
rect 18600 9180 18658 9192
rect 18600 9004 18612 9180
rect 18646 9004 18658 9180
rect 18600 8992 18658 9004
rect 18718 9180 18776 9192
rect 18718 9004 18730 9180
rect 18764 9004 18776 9180
rect 18718 8992 18776 9004
rect 18836 9180 18894 9192
rect 18836 9004 18848 9180
rect 18882 9004 18894 9180
rect 18836 8992 18894 9004
rect 19406 9176 19464 9188
rect 19406 9000 19418 9176
rect 19452 9000 19464 9176
rect 19406 8988 19464 9000
rect 19524 9176 19582 9188
rect 19524 9000 19536 9176
rect 19570 9000 19582 9176
rect 19524 8988 19582 9000
rect 19642 9176 19700 9188
rect 19642 9000 19654 9176
rect 19688 9000 19700 9176
rect 19642 8988 19700 9000
rect 19760 9176 19818 9188
rect 19760 9000 19772 9176
rect 19806 9000 19818 9176
rect 19760 8988 19818 9000
rect 19879 9000 19891 9376
rect 19925 9000 19937 9376
rect 19879 8988 19937 9000
rect 19997 9376 20055 9388
rect 19997 9000 20009 9376
rect 20043 9000 20055 9376
rect 19997 8988 20055 9000
rect 20115 9376 20173 9388
rect 20115 9000 20127 9376
rect 20161 9000 20173 9376
rect 20115 8988 20173 9000
rect 20233 9376 20291 9388
rect 20233 9000 20245 9376
rect 20279 9000 20291 9376
rect 20233 8988 20291 9000
rect 20352 9376 20410 9388
rect 20352 9000 20364 9376
rect 20398 9000 20410 9376
rect 20352 8988 20410 9000
rect 20470 9376 20528 9388
rect 20470 9000 20482 9376
rect 20516 9000 20528 9376
rect 20470 8988 20528 9000
rect 20588 9376 20646 9388
rect 20588 9000 20600 9376
rect 20634 9000 20646 9376
rect 20588 8988 20646 9000
rect 20706 9376 20764 9388
rect 20706 9000 20718 9376
rect 20752 9000 20764 9376
rect 20706 8988 20764 9000
rect 20824 9376 20882 9388
rect 20824 9000 20836 9376
rect 20870 9000 20882 9376
rect 20824 8988 20882 9000
rect 20942 9376 21000 9388
rect 20942 9000 20954 9376
rect 20988 9000 21000 9376
rect 20942 8988 21000 9000
rect 21060 9376 21118 9388
rect 21060 9000 21072 9376
rect 21106 9000 21118 9376
rect 21060 8988 21118 9000
rect 21173 9376 21231 9388
rect 21173 9000 21185 9376
rect 21219 9000 21231 9376
rect 21173 8988 21231 9000
rect 21291 9376 21349 9388
rect 21291 9000 21303 9376
rect 21337 9000 21349 9376
rect 21291 8988 21349 9000
rect 21409 9376 21467 9388
rect 21409 9000 21421 9376
rect 21455 9000 21467 9376
rect 21409 8988 21467 9000
rect 21527 9376 21585 9388
rect 21527 9000 21539 9376
rect 21573 9188 21585 9376
rect 23023 9376 23081 9388
rect 21573 9176 21672 9188
rect 21573 9000 21626 9176
rect 21660 9000 21672 9176
rect 21527 8988 21672 9000
rect 21732 9176 21790 9188
rect 21732 9000 21744 9176
rect 21778 9000 21790 9176
rect 21732 8988 21790 9000
rect 21850 9176 21908 9188
rect 21850 9000 21862 9176
rect 21896 9000 21908 9176
rect 21850 8988 21908 9000
rect 21968 9176 22026 9188
rect 21968 9000 21980 9176
rect 22014 9000 22026 9176
rect 21968 8988 22026 9000
rect 22550 9176 22608 9188
rect 22550 9000 22562 9176
rect 22596 9000 22608 9176
rect 22550 8988 22608 9000
rect 22668 9176 22726 9188
rect 22668 9000 22680 9176
rect 22714 9000 22726 9176
rect 22668 8988 22726 9000
rect 22786 9176 22844 9188
rect 22786 9000 22798 9176
rect 22832 9000 22844 9176
rect 22786 8988 22844 9000
rect 22904 9176 22962 9188
rect 22904 9000 22916 9176
rect 22950 9000 22962 9176
rect 22904 8988 22962 9000
rect 23023 9000 23035 9376
rect 23069 9000 23081 9376
rect 23023 8988 23081 9000
rect 23141 9376 23199 9388
rect 23141 9000 23153 9376
rect 23187 9000 23199 9376
rect 23141 8988 23199 9000
rect 23259 9376 23317 9388
rect 23259 9000 23271 9376
rect 23305 9000 23317 9376
rect 23259 8988 23317 9000
rect 23377 9376 23435 9388
rect 23377 9000 23389 9376
rect 23423 9000 23435 9376
rect 23377 8988 23435 9000
rect 23496 9376 23554 9388
rect 23496 9000 23508 9376
rect 23542 9000 23554 9376
rect 23496 8988 23554 9000
rect 23614 9376 23672 9388
rect 23614 9000 23626 9376
rect 23660 9000 23672 9376
rect 23614 8988 23672 9000
rect 23732 9376 23790 9388
rect 23732 9000 23744 9376
rect 23778 9000 23790 9376
rect 23732 8988 23790 9000
rect 23850 9376 23908 9388
rect 23850 9000 23862 9376
rect 23896 9000 23908 9376
rect 23850 8988 23908 9000
rect 23968 9376 24026 9388
rect 23968 9000 23980 9376
rect 24014 9000 24026 9376
rect 23968 8988 24026 9000
rect 24086 9376 24144 9388
rect 24086 9000 24098 9376
rect 24132 9000 24144 9376
rect 24086 8988 24144 9000
rect 24204 9376 24262 9388
rect 24204 9000 24216 9376
rect 24250 9000 24262 9376
rect 24204 8988 24262 9000
rect 24317 9376 24375 9388
rect 24317 9000 24329 9376
rect 24363 9000 24375 9376
rect 24317 8988 24375 9000
rect 24435 9376 24493 9388
rect 24435 9000 24447 9376
rect 24481 9000 24493 9376
rect 24435 8988 24493 9000
rect 24553 9376 24611 9388
rect 24553 9000 24565 9376
rect 24599 9000 24611 9376
rect 24553 8988 24611 9000
rect 24671 9376 24729 9388
rect 30152 9379 30352 9391
rect 24671 9000 24683 9376
rect 24717 9188 24729 9376
rect 24717 9176 24816 9188
rect 24717 9000 24770 9176
rect 24804 9000 24816 9176
rect 24671 8988 24816 9000
rect 24876 9176 24934 9188
rect 24876 9000 24888 9176
rect 24922 9000 24934 9176
rect 24876 8988 24934 9000
rect 24994 9176 25052 9188
rect 24994 9000 25006 9176
rect 25040 9000 25052 9176
rect 24994 8988 25052 9000
rect 25112 9176 25170 9188
rect 25112 9000 25124 9176
rect 25158 9000 25170 9176
rect 46658 9754 46670 10130
rect 46704 9754 46716 10130
rect 46658 9742 46716 9754
rect 46776 10130 46834 10142
rect 46776 9754 46788 10130
rect 46822 9754 46834 10130
rect 46776 9742 46834 9754
rect 46894 10130 46952 10142
rect 46894 9754 46906 10130
rect 46940 9754 46952 10130
rect 46894 9742 46952 9754
rect 47012 10130 47070 10142
rect 47012 9754 47024 10130
rect 47058 9754 47070 10130
rect 47012 9742 47070 9754
rect 47130 10130 47188 10142
rect 47130 9754 47142 10130
rect 47176 9754 47188 10130
rect 47130 9742 47188 9754
rect 47248 10130 47306 10142
rect 47248 9754 47260 10130
rect 47294 9754 47306 10130
rect 47248 9742 47306 9754
rect 47366 10130 47424 10142
rect 47366 9754 47378 10130
rect 47412 9754 47424 10130
rect 47366 9742 47424 9754
rect 47800 10134 47858 10146
rect 47800 9758 47812 10134
rect 47846 9758 47858 10134
rect 47800 9746 47858 9758
rect 47918 10134 47976 10146
rect 47918 9758 47930 10134
rect 47964 9758 47976 10134
rect 47918 9746 47976 9758
rect 48036 10134 48094 10146
rect 48036 9758 48048 10134
rect 48082 9758 48094 10134
rect 48036 9746 48094 9758
rect 48154 10134 48212 10146
rect 48154 9758 48166 10134
rect 48200 9758 48212 10134
rect 48154 9746 48212 9758
rect 48272 10134 48330 10146
rect 48272 9758 48284 10134
rect 48318 9758 48330 10134
rect 48272 9746 48330 9758
rect 48390 10134 48448 10146
rect 48390 9758 48402 10134
rect 48436 9758 48448 10134
rect 48390 9746 48448 9758
rect 48508 10134 48566 10146
rect 48508 9758 48520 10134
rect 48554 9758 48566 10134
rect 59937 10130 59995 10142
rect 53312 10062 53370 10074
rect 50987 9990 51045 10002
rect 50987 9814 50999 9990
rect 51033 9814 51045 9990
rect 50987 9802 51045 9814
rect 51105 9990 51163 10002
rect 51105 9814 51117 9990
rect 51151 9814 51163 9990
rect 51105 9802 51163 9814
rect 51223 9990 51281 10002
rect 51223 9814 51235 9990
rect 51269 9814 51281 9990
rect 51223 9802 51281 9814
rect 51341 9990 51399 10002
rect 51341 9814 51353 9990
rect 51387 9814 51399 9990
rect 51341 9802 51399 9814
rect 51459 9990 51517 10002
rect 51459 9814 51471 9990
rect 51505 9814 51517 9990
rect 51459 9802 51517 9814
rect 51577 9990 51635 10002
rect 51577 9814 51589 9990
rect 51623 9814 51635 9990
rect 51577 9802 51635 9814
rect 51695 9990 51753 10002
rect 51695 9814 51707 9990
rect 51741 9814 51753 9990
rect 51695 9802 51753 9814
rect 51813 9990 51871 10002
rect 51813 9814 51825 9990
rect 51859 9814 51871 9990
rect 51813 9802 51871 9814
rect 51931 9990 51989 10002
rect 51931 9814 51943 9990
rect 51977 9814 51989 9990
rect 51931 9802 51989 9814
rect 52049 9990 52107 10002
rect 52049 9814 52061 9990
rect 52095 9814 52107 9990
rect 52049 9802 52107 9814
rect 48508 9746 48566 9758
rect 40538 9259 40596 9271
rect 40538 9083 40550 9259
rect 40584 9083 40596 9259
rect 40538 9071 40596 9083
rect 40656 9259 40714 9271
rect 40656 9083 40668 9259
rect 40702 9083 40714 9259
rect 40656 9071 40714 9083
rect 40774 9259 40832 9271
rect 40774 9083 40786 9259
rect 40820 9083 40832 9259
rect 40774 9071 40832 9083
rect 40892 9259 40950 9271
rect 40892 9083 40904 9259
rect 40938 9083 40950 9259
rect 40892 9071 40950 9083
rect 41680 9263 41738 9275
rect 41680 9087 41692 9263
rect 41726 9087 41738 9263
rect 41680 9075 41738 9087
rect 41798 9263 41856 9275
rect 41798 9087 41810 9263
rect 41844 9087 41856 9263
rect 41798 9075 41856 9087
rect 41916 9263 41974 9275
rect 41916 9087 41928 9263
rect 41962 9087 41974 9263
rect 41916 9075 41974 9087
rect 42034 9263 42092 9275
rect 42034 9087 42046 9263
rect 42080 9087 42092 9263
rect 53312 9686 53324 10062
rect 53358 9686 53370 10062
rect 53312 9674 53370 9686
rect 53430 10062 53488 10074
rect 53430 9686 53442 10062
rect 53476 9686 53488 10062
rect 53430 9674 53488 9686
rect 53548 10062 53606 10074
rect 53548 9686 53560 10062
rect 53594 9686 53606 10062
rect 53548 9674 53606 9686
rect 53666 10062 53724 10074
rect 53666 9686 53678 10062
rect 53712 9686 53724 10062
rect 53666 9674 53724 9686
rect 53784 10062 53842 10074
rect 53784 9686 53796 10062
rect 53830 9686 53842 10062
rect 53784 9674 53842 9686
rect 53902 10062 53960 10074
rect 53902 9686 53914 10062
rect 53948 9686 53960 10062
rect 53902 9674 53960 9686
rect 54020 10062 54078 10074
rect 54020 9686 54032 10062
rect 54066 9686 54078 10062
rect 54020 9674 54078 9686
rect 54454 10066 54512 10078
rect 54454 9690 54466 10066
rect 54500 9690 54512 10066
rect 54454 9678 54512 9690
rect 54572 10066 54630 10078
rect 54572 9690 54584 10066
rect 54618 9690 54630 10066
rect 54572 9678 54630 9690
rect 54690 10066 54748 10078
rect 54690 9690 54702 10066
rect 54736 9690 54748 10066
rect 54690 9678 54748 9690
rect 54808 10066 54866 10078
rect 54808 9690 54820 10066
rect 54854 9690 54866 10066
rect 54808 9678 54866 9690
rect 54926 10066 54984 10078
rect 54926 9690 54938 10066
rect 54972 9690 54984 10066
rect 54926 9678 54984 9690
rect 55044 10066 55102 10078
rect 55044 9690 55056 10066
rect 55090 9690 55102 10066
rect 55044 9678 55102 9690
rect 55162 10066 55220 10078
rect 55162 9690 55174 10066
rect 55208 9690 55220 10066
rect 57612 10058 57670 10070
rect 57612 9882 57624 10058
rect 57658 9882 57670 10058
rect 57612 9870 57670 9882
rect 57730 10058 57788 10070
rect 57730 9882 57742 10058
rect 57776 9882 57788 10058
rect 57730 9870 57788 9882
rect 57848 10058 57906 10070
rect 57848 9882 57860 10058
rect 57894 9882 57906 10058
rect 57848 9870 57906 9882
rect 57966 10058 58024 10070
rect 57966 9882 57978 10058
rect 58012 9882 58024 10058
rect 57966 9870 58024 9882
rect 58084 10058 58142 10070
rect 58084 9882 58096 10058
rect 58130 9882 58142 10058
rect 58084 9870 58142 9882
rect 58202 10058 58260 10070
rect 58202 9882 58214 10058
rect 58248 9882 58260 10058
rect 58202 9870 58260 9882
rect 58320 10058 58378 10070
rect 58320 9882 58332 10058
rect 58366 9882 58378 10058
rect 58320 9870 58378 9882
rect 58438 10058 58496 10070
rect 58438 9882 58450 10058
rect 58484 9882 58496 10058
rect 58438 9870 58496 9882
rect 58556 10058 58614 10070
rect 58556 9882 58568 10058
rect 58602 9882 58614 10058
rect 58556 9870 58614 9882
rect 58674 10058 58732 10070
rect 58674 9882 58686 10058
rect 58720 9882 58732 10058
rect 58674 9870 58732 9882
rect 55162 9678 55220 9690
rect 47087 9347 47145 9359
rect 47087 9171 47099 9347
rect 47133 9171 47145 9347
rect 47087 9159 47145 9171
rect 47205 9347 47263 9359
rect 47205 9171 47217 9347
rect 47251 9171 47263 9347
rect 47205 9159 47263 9171
rect 47323 9347 47381 9359
rect 47323 9171 47335 9347
rect 47369 9171 47381 9347
rect 47323 9159 47381 9171
rect 47441 9347 47499 9359
rect 47441 9171 47453 9347
rect 47487 9171 47499 9347
rect 47441 9159 47499 9171
rect 48229 9351 48287 9363
rect 48229 9175 48241 9351
rect 48275 9175 48287 9351
rect 48229 9163 48287 9175
rect 48347 9351 48405 9363
rect 48347 9175 48359 9351
rect 48393 9175 48405 9351
rect 48347 9163 48405 9175
rect 48465 9351 48523 9363
rect 48465 9175 48477 9351
rect 48511 9175 48523 9351
rect 48465 9163 48523 9175
rect 48583 9351 48641 9363
rect 48583 9175 48595 9351
rect 48629 9175 48641 9351
rect 48583 9163 48641 9175
rect 59937 9754 59949 10130
rect 59983 9754 59995 10130
rect 59937 9742 59995 9754
rect 60055 10130 60113 10142
rect 60055 9754 60067 10130
rect 60101 9754 60113 10130
rect 60055 9742 60113 9754
rect 60173 10130 60231 10142
rect 60173 9754 60185 10130
rect 60219 9754 60231 10130
rect 60173 9742 60231 9754
rect 60291 10130 60349 10142
rect 60291 9754 60303 10130
rect 60337 9754 60349 10130
rect 60291 9742 60349 9754
rect 60409 10130 60467 10142
rect 60409 9754 60421 10130
rect 60455 9754 60467 10130
rect 60409 9742 60467 9754
rect 60527 10130 60585 10142
rect 60527 9754 60539 10130
rect 60573 9754 60585 10130
rect 60527 9742 60585 9754
rect 60645 10130 60703 10142
rect 60645 9754 60657 10130
rect 60691 9754 60703 10130
rect 60645 9742 60703 9754
rect 61079 10134 61137 10146
rect 61079 9758 61091 10134
rect 61125 9758 61137 10134
rect 61079 9746 61137 9758
rect 61197 10134 61255 10146
rect 61197 9758 61209 10134
rect 61243 9758 61255 10134
rect 61197 9746 61255 9758
rect 61315 10134 61373 10146
rect 61315 9758 61327 10134
rect 61361 9758 61373 10134
rect 61315 9746 61373 9758
rect 61433 10134 61491 10146
rect 61433 9758 61445 10134
rect 61479 9758 61491 10134
rect 61433 9746 61491 9758
rect 61551 10134 61609 10146
rect 61551 9758 61563 10134
rect 61597 9758 61609 10134
rect 61551 9746 61609 9758
rect 61669 10134 61727 10146
rect 61669 9758 61681 10134
rect 61715 9758 61727 10134
rect 61669 9746 61727 9758
rect 61787 10134 61845 10146
rect 61787 9758 61799 10134
rect 61833 9758 61845 10134
rect 70709 10315 70909 10327
rect 70709 10281 70721 10315
rect 70897 10281 70909 10315
rect 70709 10269 70909 10281
rect 70709 10197 70909 10209
rect 70709 10163 70721 10197
rect 70897 10163 70909 10197
rect 70709 10151 70909 10163
rect 70709 10079 70909 10091
rect 70709 10045 70721 10079
rect 70897 10045 70909 10079
rect 70709 10033 70909 10045
rect 61787 9746 61845 9758
rect 42034 9075 42092 9087
rect 53741 9279 53799 9291
rect 53741 9103 53753 9279
rect 53787 9103 53799 9279
rect 53741 9091 53799 9103
rect 53859 9279 53917 9291
rect 53859 9103 53871 9279
rect 53905 9103 53917 9279
rect 53859 9091 53917 9103
rect 53977 9279 54035 9291
rect 53977 9103 53989 9279
rect 54023 9103 54035 9279
rect 53977 9091 54035 9103
rect 54095 9279 54153 9291
rect 54095 9103 54107 9279
rect 54141 9103 54153 9279
rect 54095 9091 54153 9103
rect 54883 9283 54941 9295
rect 54883 9107 54895 9283
rect 54929 9107 54941 9283
rect 54883 9095 54941 9107
rect 55001 9283 55059 9295
rect 55001 9107 55013 9283
rect 55047 9107 55059 9283
rect 55001 9095 55059 9107
rect 55119 9283 55177 9295
rect 55119 9107 55131 9283
rect 55165 9107 55177 9283
rect 55119 9095 55177 9107
rect 55237 9283 55295 9295
rect 55237 9107 55249 9283
rect 55283 9107 55295 9283
rect 70713 9439 70913 9451
rect 63409 9419 63467 9431
rect 60366 9347 60424 9359
rect 60366 9171 60378 9347
rect 60412 9171 60424 9347
rect 60366 9159 60424 9171
rect 60484 9347 60542 9359
rect 60484 9171 60496 9347
rect 60530 9171 60542 9347
rect 60484 9159 60542 9171
rect 60602 9347 60660 9359
rect 60602 9171 60614 9347
rect 60648 9171 60660 9347
rect 60602 9159 60660 9171
rect 60720 9347 60778 9359
rect 60720 9171 60732 9347
rect 60766 9171 60778 9347
rect 60720 9159 60778 9171
rect 61508 9351 61566 9363
rect 61508 9175 61520 9351
rect 61554 9175 61566 9351
rect 61508 9163 61566 9175
rect 61626 9351 61684 9363
rect 61626 9175 61638 9351
rect 61672 9175 61684 9351
rect 61626 9163 61684 9175
rect 61744 9351 61802 9363
rect 61744 9175 61756 9351
rect 61790 9175 61802 9351
rect 61744 9163 61802 9175
rect 61862 9351 61920 9363
rect 61862 9175 61874 9351
rect 61908 9175 61920 9351
rect 63409 9243 63421 9419
rect 63455 9243 63467 9419
rect 63409 9231 63467 9243
rect 63527 9419 63585 9431
rect 63527 9243 63539 9419
rect 63573 9243 63585 9419
rect 63527 9231 63585 9243
rect 63645 9419 63703 9431
rect 63645 9243 63657 9419
rect 63691 9243 63703 9419
rect 63645 9231 63703 9243
rect 63763 9419 63821 9431
rect 63763 9243 63775 9419
rect 63809 9243 63821 9419
rect 63763 9231 63821 9243
rect 63881 9419 63939 9431
rect 63881 9243 63893 9419
rect 63927 9243 63939 9419
rect 63881 9231 63939 9243
rect 63999 9419 64057 9431
rect 63999 9243 64011 9419
rect 64045 9243 64057 9419
rect 63999 9231 64057 9243
rect 64117 9419 64175 9431
rect 64117 9243 64129 9419
rect 64163 9243 64175 9419
rect 64117 9231 64175 9243
rect 64235 9419 64293 9431
rect 64235 9243 64247 9419
rect 64281 9243 64293 9419
rect 64235 9231 64293 9243
rect 64353 9419 64411 9431
rect 64353 9243 64365 9419
rect 64399 9243 64411 9419
rect 64353 9231 64411 9243
rect 64471 9419 64529 9431
rect 64471 9243 64483 9419
rect 64517 9243 64529 9419
rect 70713 9405 70725 9439
rect 70901 9405 70913 9439
rect 70713 9393 70913 9405
rect 64471 9231 64529 9243
rect 70713 9321 70913 9333
rect 70713 9287 70725 9321
rect 70901 9287 70913 9321
rect 70713 9275 70913 9287
rect 61862 9163 61920 9175
rect 55237 9095 55295 9107
rect 25112 8988 25170 9000
rect 30154 9031 30354 9043
rect 30154 8997 30166 9031
rect 30342 8997 30354 9031
rect 30154 8985 30354 8997
rect 30154 8913 30354 8925
rect 30154 8879 30166 8913
rect 30342 8879 30354 8913
rect 30154 8867 30354 8879
rect 70713 9203 70913 9215
rect 70713 9169 70725 9203
rect 70901 9169 70913 9203
rect 70713 9157 70913 9169
rect 70713 9085 70913 9097
rect 70713 9051 70725 9085
rect 70901 9051 70913 9085
rect 70713 9010 70913 9051
rect 70513 8998 70913 9010
rect 30154 8795 30354 8807
rect 30154 8761 30166 8795
rect 30342 8761 30354 8795
rect 30154 8749 30354 8761
rect 30154 8677 30354 8689
rect 30154 8643 30166 8677
rect 30342 8643 30354 8677
rect 30154 8631 30354 8643
rect 29954 8547 30354 8559
rect 29954 8513 29966 8547
rect 30342 8513 30354 8547
rect 29954 8501 30354 8513
rect 30647 8604 31047 8616
rect 30647 8570 30659 8604
rect 31035 8570 31047 8604
rect 30647 8558 31047 8570
rect 29954 8429 30354 8441
rect 29954 8395 29966 8429
rect 30342 8395 30354 8429
rect 29954 8383 30354 8395
rect 30647 8486 31047 8498
rect 30647 8452 30659 8486
rect 31035 8452 31047 8486
rect 30647 8440 31047 8452
rect 70513 8964 70525 8998
rect 70901 8964 70913 8998
rect 70513 8952 70913 8964
rect 70513 8880 70913 8892
rect 70513 8846 70525 8880
rect 70901 8846 70913 8880
rect 70513 8834 70913 8846
rect 70513 8762 70913 8774
rect 70513 8728 70525 8762
rect 70901 8728 70913 8762
rect 70513 8716 70913 8728
rect 70513 8644 70913 8656
rect 70513 8610 70525 8644
rect 70901 8610 70913 8644
rect 70513 8598 70913 8610
rect 29954 8311 30354 8323
rect 29954 8277 29966 8311
rect 30342 8277 30354 8311
rect 29954 8265 30354 8277
rect 30647 8368 31047 8380
rect 30647 8334 30659 8368
rect 31035 8334 31047 8368
rect 30647 8322 31047 8334
rect 30647 8250 31047 8262
rect 30647 8216 30659 8250
rect 31035 8216 31047 8250
rect 29954 8193 30354 8205
rect 30647 8204 31047 8216
rect 29954 8159 29966 8193
rect 30342 8159 30354 8193
rect 29954 8147 30354 8159
rect 29954 8075 30354 8087
rect 29954 8041 29966 8075
rect 30342 8041 30354 8075
rect 29954 8029 30354 8041
rect 29954 7957 30354 7969
rect 29954 7923 29966 7957
rect 30342 7923 30354 7957
rect 29954 7911 30354 7923
rect 30647 8132 31047 8144
rect 30647 8098 30659 8132
rect 31035 8098 31047 8132
rect 30647 8086 31047 8098
rect 37798 8320 37856 8332
rect 37798 8144 37810 8320
rect 37844 8144 37856 8320
rect 37798 8132 37856 8144
rect 37916 8320 37974 8332
rect 37916 8144 37928 8320
rect 37962 8144 37974 8320
rect 37916 8132 37974 8144
rect 38034 8320 38092 8332
rect 38034 8144 38046 8320
rect 38080 8144 38092 8320
rect 38034 8132 38092 8144
rect 38152 8320 38210 8332
rect 38152 8144 38164 8320
rect 38198 8144 38210 8320
rect 38152 8132 38210 8144
rect 38270 8320 38328 8332
rect 38270 8144 38282 8320
rect 38316 8144 38328 8320
rect 38270 8132 38328 8144
rect 38388 8320 38446 8332
rect 38388 8144 38400 8320
rect 38434 8144 38446 8320
rect 38388 8132 38446 8144
rect 38506 8320 38564 8332
rect 38506 8144 38518 8320
rect 38552 8144 38564 8320
rect 38506 8132 38564 8144
rect 38624 8320 38682 8332
rect 38624 8144 38636 8320
rect 38670 8144 38682 8320
rect 38624 8132 38682 8144
rect 38742 8320 38800 8332
rect 38742 8144 38754 8320
rect 38788 8144 38800 8320
rect 38742 8132 38800 8144
rect 38860 8320 38918 8332
rect 38860 8144 38872 8320
rect 38906 8144 38918 8320
rect 44347 8408 44405 8420
rect 44347 8232 44359 8408
rect 44393 8232 44405 8408
rect 44347 8220 44405 8232
rect 44465 8408 44523 8420
rect 44465 8232 44477 8408
rect 44511 8232 44523 8408
rect 44465 8220 44523 8232
rect 44583 8408 44641 8420
rect 44583 8232 44595 8408
rect 44629 8232 44641 8408
rect 44583 8220 44641 8232
rect 44701 8408 44759 8420
rect 44701 8232 44713 8408
rect 44747 8232 44759 8408
rect 44701 8220 44759 8232
rect 44819 8408 44877 8420
rect 44819 8232 44831 8408
rect 44865 8232 44877 8408
rect 44819 8220 44877 8232
rect 44937 8408 44995 8420
rect 44937 8232 44949 8408
rect 44983 8232 44995 8408
rect 44937 8220 44995 8232
rect 45055 8408 45113 8420
rect 45055 8232 45067 8408
rect 45101 8232 45113 8408
rect 45055 8220 45113 8232
rect 45173 8408 45231 8420
rect 45173 8232 45185 8408
rect 45219 8232 45231 8408
rect 45173 8220 45231 8232
rect 45291 8408 45349 8420
rect 45291 8232 45303 8408
rect 45337 8232 45349 8408
rect 45291 8220 45349 8232
rect 45409 8408 45467 8420
rect 45409 8232 45421 8408
rect 45455 8232 45467 8408
rect 70513 8531 70913 8543
rect 70513 8497 70525 8531
rect 70901 8497 70913 8531
rect 70513 8485 70913 8497
rect 51001 8340 51059 8352
rect 45409 8220 45467 8232
rect 38860 8132 38918 8144
rect 30647 8014 31047 8026
rect 30647 7980 30659 8014
rect 31035 7980 31047 8014
rect 30647 7968 31047 7980
rect 29954 7839 30354 7851
rect 29954 7805 29966 7839
rect 30342 7805 30354 7839
rect 29954 7793 30354 7805
rect 30154 7710 30354 7722
rect 30154 7676 30166 7710
rect 30342 7676 30354 7710
rect 30154 7664 30354 7676
rect 30647 7896 31047 7908
rect 30647 7862 30659 7896
rect 31035 7862 31047 7896
rect 51001 8164 51013 8340
rect 51047 8164 51059 8340
rect 51001 8152 51059 8164
rect 51119 8340 51177 8352
rect 51119 8164 51131 8340
rect 51165 8164 51177 8340
rect 51119 8152 51177 8164
rect 51237 8340 51295 8352
rect 51237 8164 51249 8340
rect 51283 8164 51295 8340
rect 51237 8152 51295 8164
rect 51355 8340 51413 8352
rect 51355 8164 51367 8340
rect 51401 8164 51413 8340
rect 51355 8152 51413 8164
rect 51473 8340 51531 8352
rect 51473 8164 51485 8340
rect 51519 8164 51531 8340
rect 51473 8152 51531 8164
rect 51591 8340 51649 8352
rect 51591 8164 51603 8340
rect 51637 8164 51649 8340
rect 51591 8152 51649 8164
rect 51709 8340 51767 8352
rect 51709 8164 51721 8340
rect 51755 8164 51767 8340
rect 51709 8152 51767 8164
rect 51827 8340 51885 8352
rect 51827 8164 51839 8340
rect 51873 8164 51885 8340
rect 51827 8152 51885 8164
rect 51945 8340 52003 8352
rect 51945 8164 51957 8340
rect 51991 8164 52003 8340
rect 51945 8152 52003 8164
rect 52063 8340 52121 8352
rect 52063 8164 52075 8340
rect 52109 8164 52121 8340
rect 57626 8408 57684 8420
rect 57626 8232 57638 8408
rect 57672 8232 57684 8408
rect 57626 8220 57684 8232
rect 57744 8408 57802 8420
rect 57744 8232 57756 8408
rect 57790 8232 57802 8408
rect 57744 8220 57802 8232
rect 57862 8408 57920 8420
rect 57862 8232 57874 8408
rect 57908 8232 57920 8408
rect 57862 8220 57920 8232
rect 57980 8408 58038 8420
rect 57980 8232 57992 8408
rect 58026 8232 58038 8408
rect 57980 8220 58038 8232
rect 58098 8408 58156 8420
rect 58098 8232 58110 8408
rect 58144 8232 58156 8408
rect 58098 8220 58156 8232
rect 58216 8408 58274 8420
rect 58216 8232 58228 8408
rect 58262 8232 58274 8408
rect 58216 8220 58274 8232
rect 58334 8408 58392 8420
rect 58334 8232 58346 8408
rect 58380 8232 58392 8408
rect 58334 8220 58392 8232
rect 58452 8408 58510 8420
rect 58452 8232 58464 8408
rect 58498 8232 58510 8408
rect 58452 8220 58510 8232
rect 58570 8408 58628 8420
rect 58570 8232 58582 8408
rect 58616 8232 58628 8408
rect 58570 8220 58628 8232
rect 58688 8408 58746 8420
rect 58688 8232 58700 8408
rect 58734 8232 58746 8408
rect 70513 8413 70913 8425
rect 70513 8379 70525 8413
rect 70901 8379 70913 8413
rect 70513 8367 70913 8379
rect 58688 8220 58746 8232
rect 52063 8152 52121 8164
rect 46295 7991 46353 8003
rect 39746 7903 39804 7915
rect 30647 7850 31047 7862
rect 34886 7652 34944 7664
rect 30154 7592 30354 7604
rect 30154 7558 30166 7592
rect 30342 7558 30354 7592
rect 30154 7546 30354 7558
rect 30154 7474 30354 7486
rect 30154 7440 30166 7474
rect 30342 7440 30354 7474
rect 34886 7476 34898 7652
rect 34932 7476 34944 7652
rect 34886 7464 34944 7476
rect 35004 7652 35062 7664
rect 35004 7476 35016 7652
rect 35050 7476 35062 7652
rect 35004 7464 35062 7476
rect 35122 7652 35180 7664
rect 35122 7476 35134 7652
rect 35168 7476 35180 7652
rect 35122 7464 35180 7476
rect 35240 7652 35298 7664
rect 35240 7476 35252 7652
rect 35286 7476 35298 7652
rect 35240 7464 35298 7476
rect 35358 7652 35416 7664
rect 35358 7476 35370 7652
rect 35404 7476 35416 7652
rect 35358 7464 35416 7476
rect 35476 7652 35534 7664
rect 35476 7476 35488 7652
rect 35522 7476 35534 7652
rect 35476 7464 35534 7476
rect 35594 7652 35652 7664
rect 35594 7476 35606 7652
rect 35640 7476 35652 7652
rect 35594 7464 35652 7476
rect 35712 7652 35770 7664
rect 35712 7476 35724 7652
rect 35758 7476 35770 7652
rect 35712 7464 35770 7476
rect 35830 7652 35888 7664
rect 35830 7476 35842 7652
rect 35876 7476 35888 7652
rect 35830 7464 35888 7476
rect 35948 7652 36006 7664
rect 35948 7476 35960 7652
rect 35994 7476 36006 7652
rect 39262 7703 39320 7715
rect 35948 7464 36006 7476
rect 30154 7428 30354 7440
rect 30154 7356 30354 7368
rect 30154 7322 30166 7356
rect 30342 7322 30354 7356
rect 30154 7310 30354 7322
rect 39262 7527 39274 7703
rect 39308 7527 39320 7703
rect 39262 7515 39320 7527
rect 39380 7703 39438 7715
rect 39380 7527 39392 7703
rect 39426 7527 39438 7703
rect 39380 7515 39438 7527
rect 39498 7703 39556 7715
rect 39498 7527 39510 7703
rect 39544 7527 39556 7703
rect 39498 7515 39556 7527
rect 39616 7703 39674 7715
rect 39616 7527 39628 7703
rect 39662 7527 39674 7703
rect 39616 7515 39674 7527
rect 39746 7527 39758 7903
rect 39792 7527 39804 7903
rect 39746 7515 39804 7527
rect 39864 7903 39922 7915
rect 39864 7527 39876 7903
rect 39910 7527 39922 7903
rect 39864 7515 39922 7527
rect 39982 7903 40040 7915
rect 39982 7527 39994 7903
rect 40028 7527 40040 7903
rect 39982 7515 40040 7527
rect 40100 7903 40158 7915
rect 40100 7527 40112 7903
rect 40146 7527 40158 7903
rect 40100 7515 40158 7527
rect 40218 7903 40276 7915
rect 40218 7527 40230 7903
rect 40264 7527 40276 7903
rect 40218 7515 40276 7527
rect 40336 7903 40394 7915
rect 40336 7527 40348 7903
rect 40382 7527 40394 7903
rect 40336 7515 40394 7527
rect 40454 7903 40512 7915
rect 40454 7527 40466 7903
rect 40500 7527 40512 7903
rect 41644 7903 41702 7915
rect 40454 7515 40512 7527
rect 40583 7703 40641 7715
rect 40583 7527 40595 7703
rect 40629 7527 40641 7703
rect 40583 7515 40641 7527
rect 40701 7703 40759 7715
rect 40701 7527 40713 7703
rect 40747 7527 40759 7703
rect 40701 7515 40759 7527
rect 40819 7703 40877 7715
rect 40819 7527 40831 7703
rect 40865 7527 40877 7703
rect 40819 7515 40877 7527
rect 40937 7703 40995 7715
rect 40937 7527 40949 7703
rect 40983 7527 40995 7703
rect 40937 7515 40995 7527
rect 41160 7703 41218 7715
rect 41160 7527 41172 7703
rect 41206 7527 41218 7703
rect 41160 7515 41218 7527
rect 41278 7703 41336 7715
rect 41278 7527 41290 7703
rect 41324 7527 41336 7703
rect 41278 7515 41336 7527
rect 41396 7703 41454 7715
rect 41396 7527 41408 7703
rect 41442 7527 41454 7703
rect 41396 7515 41454 7527
rect 41514 7703 41572 7715
rect 41514 7527 41526 7703
rect 41560 7527 41572 7703
rect 41514 7515 41572 7527
rect 41644 7527 41656 7903
rect 41690 7527 41702 7903
rect 41644 7515 41702 7527
rect 41762 7903 41820 7915
rect 41762 7527 41774 7903
rect 41808 7527 41820 7903
rect 41762 7515 41820 7527
rect 41880 7903 41938 7915
rect 41880 7527 41892 7903
rect 41926 7527 41938 7903
rect 41880 7515 41938 7527
rect 41998 7903 42056 7915
rect 41998 7527 42010 7903
rect 42044 7527 42056 7903
rect 41998 7515 42056 7527
rect 42116 7903 42174 7915
rect 42116 7527 42128 7903
rect 42162 7527 42174 7903
rect 42116 7515 42174 7527
rect 42234 7903 42292 7915
rect 42234 7527 42246 7903
rect 42280 7527 42292 7903
rect 42234 7515 42292 7527
rect 42352 7903 42410 7915
rect 42352 7527 42364 7903
rect 42398 7527 42410 7903
rect 42352 7515 42410 7527
rect 42481 7703 42539 7715
rect 42481 7527 42493 7703
rect 42527 7527 42539 7703
rect 42481 7515 42539 7527
rect 42599 7703 42657 7715
rect 42599 7527 42611 7703
rect 42645 7527 42657 7703
rect 42599 7515 42657 7527
rect 42717 7703 42775 7715
rect 42717 7527 42729 7703
rect 42763 7527 42775 7703
rect 42717 7515 42775 7527
rect 42835 7703 42893 7715
rect 42835 7527 42847 7703
rect 42881 7527 42893 7703
rect 45811 7791 45869 7803
rect 42835 7515 42893 7527
rect 30152 6963 30352 6975
rect 30152 6929 30164 6963
rect 30340 6929 30352 6963
rect 30152 6917 30352 6929
rect 30152 6845 30352 6857
rect 30152 6811 30164 6845
rect 30340 6811 30352 6845
rect 30152 6799 30352 6811
rect 30152 6727 30352 6739
rect 30152 6693 30164 6727
rect 30340 6693 30352 6727
rect 30152 6681 30352 6693
rect 37793 6716 37851 6728
rect 30152 6609 30352 6621
rect 3117 6545 3175 6557
rect 3117 6369 3129 6545
rect 3163 6369 3175 6545
rect 3117 6357 3175 6369
rect 3235 6545 3293 6557
rect 3235 6369 3247 6545
rect 3281 6369 3293 6545
rect 3235 6357 3293 6369
rect 3353 6545 3411 6557
rect 3353 6369 3365 6545
rect 3399 6369 3411 6545
rect 3353 6357 3411 6369
rect 3471 6545 3529 6557
rect 3471 6369 3483 6545
rect 3517 6369 3529 6545
rect 3471 6357 3529 6369
rect 3855 6545 3913 6557
rect 3855 6369 3867 6545
rect 3901 6369 3913 6545
rect 3855 6357 3913 6369
rect 3973 6545 4031 6557
rect 3973 6369 3985 6545
rect 4019 6369 4031 6545
rect 3973 6357 4031 6369
rect 4091 6545 4149 6557
rect 4091 6369 4103 6545
rect 4137 6369 4149 6545
rect 4091 6357 4149 6369
rect 4209 6545 4267 6557
rect 4209 6369 4221 6545
rect 4255 6369 4267 6545
rect 4209 6357 4267 6369
rect 4593 6545 4651 6557
rect 4593 6369 4605 6545
rect 4639 6369 4651 6545
rect 4593 6357 4651 6369
rect 4711 6545 4769 6557
rect 4711 6369 4723 6545
rect 4757 6369 4769 6545
rect 4711 6357 4769 6369
rect 4829 6545 4887 6557
rect 4829 6369 4841 6545
rect 4875 6369 4887 6545
rect 4829 6357 4887 6369
rect 4947 6545 5005 6557
rect 4947 6369 4959 6545
rect 4993 6369 5005 6545
rect 4947 6357 5005 6369
rect 5331 6545 5389 6557
rect 5331 6369 5343 6545
rect 5377 6369 5389 6545
rect 5331 6357 5389 6369
rect 5449 6545 5507 6557
rect 5449 6369 5461 6545
rect 5495 6369 5507 6545
rect 5449 6357 5507 6369
rect 5567 6545 5625 6557
rect 5567 6369 5579 6545
rect 5613 6369 5625 6545
rect 5567 6357 5625 6369
rect 5685 6545 5743 6557
rect 5685 6369 5697 6545
rect 5731 6369 5743 6545
rect 5685 6357 5743 6369
rect 6071 6545 6129 6557
rect 6071 6369 6083 6545
rect 6117 6369 6129 6545
rect 6071 6357 6129 6369
rect 6189 6545 6247 6557
rect 6189 6369 6201 6545
rect 6235 6369 6247 6545
rect 6189 6357 6247 6369
rect 6307 6545 6365 6557
rect 6307 6369 6319 6545
rect 6353 6369 6365 6545
rect 6307 6357 6365 6369
rect 6425 6545 6483 6557
rect 6425 6369 6437 6545
rect 6471 6369 6483 6545
rect 6425 6357 6483 6369
rect 6813 6547 6871 6559
rect 6813 6371 6825 6547
rect 6859 6371 6871 6547
rect 6813 6359 6871 6371
rect 6931 6547 6989 6559
rect 6931 6371 6943 6547
rect 6977 6371 6989 6547
rect 6931 6359 6989 6371
rect 7049 6547 7107 6559
rect 7049 6371 7061 6547
rect 7095 6371 7107 6547
rect 7049 6359 7107 6371
rect 7167 6547 7225 6559
rect 7167 6371 7179 6547
rect 7213 6371 7225 6547
rect 7167 6359 7225 6371
rect 7551 6551 7609 6563
rect 7551 6375 7563 6551
rect 7597 6375 7609 6551
rect 7551 6363 7609 6375
rect 7669 6551 7727 6563
rect 7669 6375 7681 6551
rect 7715 6375 7727 6551
rect 7669 6363 7727 6375
rect 7787 6551 7845 6563
rect 7787 6375 7799 6551
rect 7833 6375 7845 6551
rect 7787 6363 7845 6375
rect 7905 6551 7963 6563
rect 30152 6575 30164 6609
rect 30340 6575 30352 6609
rect 30152 6563 30352 6575
rect 7905 6375 7917 6551
rect 7951 6375 7963 6551
rect 7905 6363 7963 6375
rect 8289 6547 8347 6559
rect 8289 6371 8301 6547
rect 8335 6371 8347 6547
rect 8289 6359 8347 6371
rect 8407 6547 8465 6559
rect 8407 6371 8419 6547
rect 8453 6371 8465 6547
rect 8407 6359 8465 6371
rect 8525 6547 8583 6559
rect 8525 6371 8537 6547
rect 8571 6371 8583 6547
rect 8525 6359 8583 6371
rect 8643 6547 8701 6559
rect 8643 6371 8655 6547
rect 8689 6371 8701 6547
rect 8643 6359 8701 6371
rect 9704 6435 9762 6447
rect 9221 6235 9279 6247
rect 9221 6059 9233 6235
rect 9267 6059 9279 6235
rect 9221 6047 9279 6059
rect 9339 6235 9397 6247
rect 9339 6059 9351 6235
rect 9385 6059 9397 6235
rect 9339 6047 9397 6059
rect 9457 6235 9515 6247
rect 9457 6059 9469 6235
rect 9503 6059 9515 6235
rect 9457 6047 9515 6059
rect 9575 6235 9633 6247
rect 9575 6059 9587 6235
rect 9621 6059 9633 6235
rect 9575 6047 9633 6059
rect 9704 6059 9716 6435
rect 9750 6059 9762 6435
rect 9704 6047 9762 6059
rect 9822 6435 9880 6447
rect 9822 6059 9834 6435
rect 9868 6059 9880 6435
rect 9822 6047 9880 6059
rect 9940 6435 9998 6447
rect 9940 6059 9952 6435
rect 9986 6059 9998 6435
rect 9940 6047 9998 6059
rect 10058 6435 10116 6447
rect 10058 6059 10070 6435
rect 10104 6059 10116 6435
rect 10058 6047 10116 6059
rect 10176 6435 10234 6447
rect 10176 6059 10188 6435
rect 10222 6059 10234 6435
rect 10176 6047 10234 6059
rect 10294 6435 10352 6447
rect 10294 6059 10306 6435
rect 10340 6059 10352 6435
rect 10294 6047 10352 6059
rect 10412 6435 10470 6447
rect 10412 6059 10424 6435
rect 10458 6059 10470 6435
rect 11772 6433 11830 6445
rect 10412 6047 10470 6059
rect 10542 6235 10600 6247
rect 10542 6059 10554 6235
rect 10588 6059 10600 6235
rect 10542 6047 10600 6059
rect 10660 6235 10718 6247
rect 10660 6059 10672 6235
rect 10706 6059 10718 6235
rect 10660 6047 10718 6059
rect 10778 6235 10836 6247
rect 10778 6059 10790 6235
rect 10824 6059 10836 6235
rect 10778 6047 10836 6059
rect 10896 6235 10954 6247
rect 10896 6059 10908 6235
rect 10942 6059 10954 6235
rect 10896 6047 10954 6059
rect 11289 6233 11347 6245
rect 11289 6057 11301 6233
rect 11335 6057 11347 6233
rect 11289 6045 11347 6057
rect 11407 6233 11465 6245
rect 11407 6057 11419 6233
rect 11453 6057 11465 6233
rect 11407 6045 11465 6057
rect 11525 6233 11583 6245
rect 11525 6057 11537 6233
rect 11571 6057 11583 6233
rect 11525 6045 11583 6057
rect 11643 6233 11701 6245
rect 11643 6057 11655 6233
rect 11689 6057 11701 6233
rect 11643 6045 11701 6057
rect 11772 6057 11784 6433
rect 11818 6057 11830 6433
rect 11772 6045 11830 6057
rect 11890 6433 11948 6445
rect 11890 6057 11902 6433
rect 11936 6057 11948 6433
rect 11890 6045 11948 6057
rect 12008 6433 12066 6445
rect 12008 6057 12020 6433
rect 12054 6057 12066 6433
rect 12008 6045 12066 6057
rect 12126 6433 12184 6445
rect 12126 6057 12138 6433
rect 12172 6057 12184 6433
rect 12126 6045 12184 6057
rect 12244 6433 12302 6445
rect 12244 6057 12256 6433
rect 12290 6057 12302 6433
rect 12244 6045 12302 6057
rect 12362 6433 12420 6445
rect 12362 6057 12374 6433
rect 12408 6057 12420 6433
rect 12362 6045 12420 6057
rect 12480 6433 12538 6445
rect 12480 6057 12492 6433
rect 12526 6057 12538 6433
rect 13841 6435 13899 6447
rect 12480 6045 12538 6057
rect 12610 6233 12668 6245
rect 12610 6057 12622 6233
rect 12656 6057 12668 6233
rect 12610 6045 12668 6057
rect 12728 6233 12786 6245
rect 12728 6057 12740 6233
rect 12774 6057 12786 6233
rect 12728 6045 12786 6057
rect 12846 6233 12904 6245
rect 12846 6057 12858 6233
rect 12892 6057 12904 6233
rect 12846 6045 12904 6057
rect 12964 6233 13022 6245
rect 12964 6057 12976 6233
rect 13010 6057 13022 6233
rect 12964 6045 13022 6057
rect 13358 6235 13416 6247
rect 13358 6059 13370 6235
rect 13404 6059 13416 6235
rect 13358 6047 13416 6059
rect 13476 6235 13534 6247
rect 13476 6059 13488 6235
rect 13522 6059 13534 6235
rect 13476 6047 13534 6059
rect 13594 6235 13652 6247
rect 13594 6059 13606 6235
rect 13640 6059 13652 6235
rect 13594 6047 13652 6059
rect 13712 6235 13770 6247
rect 13712 6059 13724 6235
rect 13758 6059 13770 6235
rect 13712 6047 13770 6059
rect 13841 6059 13853 6435
rect 13887 6059 13899 6435
rect 13841 6047 13899 6059
rect 13959 6435 14017 6447
rect 13959 6059 13971 6435
rect 14005 6059 14017 6435
rect 13959 6047 14017 6059
rect 14077 6435 14135 6447
rect 14077 6059 14089 6435
rect 14123 6059 14135 6435
rect 14077 6047 14135 6059
rect 14195 6435 14253 6447
rect 14195 6059 14207 6435
rect 14241 6059 14253 6435
rect 14195 6047 14253 6059
rect 14313 6435 14371 6447
rect 14313 6059 14325 6435
rect 14359 6059 14371 6435
rect 14313 6047 14371 6059
rect 14431 6435 14489 6447
rect 14431 6059 14443 6435
rect 14477 6059 14489 6435
rect 14431 6047 14489 6059
rect 14549 6435 14607 6447
rect 14549 6059 14561 6435
rect 14595 6059 14607 6435
rect 15909 6433 15967 6445
rect 14549 6047 14607 6059
rect 14679 6235 14737 6247
rect 14679 6059 14691 6235
rect 14725 6059 14737 6235
rect 14679 6047 14737 6059
rect 14797 6235 14855 6247
rect 14797 6059 14809 6235
rect 14843 6059 14855 6235
rect 14797 6047 14855 6059
rect 14915 6235 14973 6247
rect 14915 6059 14927 6235
rect 14961 6059 14973 6235
rect 14915 6047 14973 6059
rect 15033 6235 15091 6247
rect 15033 6059 15045 6235
rect 15079 6059 15091 6235
rect 15033 6047 15091 6059
rect 15426 6233 15484 6245
rect 15426 6057 15438 6233
rect 15472 6057 15484 6233
rect 9761 5742 9819 5754
rect 9761 5366 9773 5742
rect 9807 5366 9819 5742
rect 9761 5354 9819 5366
rect 9879 5742 9937 5754
rect 9879 5366 9891 5742
rect 9925 5366 9937 5742
rect 9879 5354 9937 5366
rect 9997 5742 10055 5754
rect 9997 5366 10009 5742
rect 10043 5366 10055 5742
rect 9997 5354 10055 5366
rect 10115 5742 10173 5754
rect 10115 5366 10127 5742
rect 10161 5366 10173 5742
rect 10115 5354 10173 5366
rect 10233 5742 10291 5754
rect 10233 5366 10245 5742
rect 10279 5366 10291 5742
rect 10233 5354 10291 5366
rect 10351 5742 10409 5754
rect 10351 5366 10363 5742
rect 10397 5366 10409 5742
rect 10351 5354 10409 5366
rect 10469 5742 10527 5754
rect 10469 5366 10481 5742
rect 10515 5366 10527 5742
rect 10469 5354 10527 5366
rect 15426 6045 15484 6057
rect 15544 6233 15602 6245
rect 15544 6057 15556 6233
rect 15590 6057 15602 6233
rect 15544 6045 15602 6057
rect 15662 6233 15720 6245
rect 15662 6057 15674 6233
rect 15708 6057 15720 6233
rect 15662 6045 15720 6057
rect 15780 6233 15838 6245
rect 15780 6057 15792 6233
rect 15826 6057 15838 6233
rect 15780 6045 15838 6057
rect 15909 6057 15921 6433
rect 15955 6057 15967 6433
rect 15909 6045 15967 6057
rect 16027 6433 16085 6445
rect 16027 6057 16039 6433
rect 16073 6057 16085 6433
rect 16027 6045 16085 6057
rect 16145 6433 16203 6445
rect 16145 6057 16157 6433
rect 16191 6057 16203 6433
rect 16145 6045 16203 6057
rect 16263 6433 16321 6445
rect 16263 6057 16275 6433
rect 16309 6057 16321 6433
rect 16263 6045 16321 6057
rect 16381 6433 16439 6445
rect 16381 6057 16393 6433
rect 16427 6057 16439 6433
rect 16381 6045 16439 6057
rect 16499 6433 16557 6445
rect 16499 6057 16511 6433
rect 16545 6057 16557 6433
rect 16499 6045 16557 6057
rect 16617 6433 16675 6445
rect 16617 6057 16629 6433
rect 16663 6057 16675 6433
rect 17978 6433 18036 6445
rect 16617 6045 16675 6057
rect 16747 6233 16805 6245
rect 16747 6057 16759 6233
rect 16793 6057 16805 6233
rect 16747 6045 16805 6057
rect 16865 6233 16923 6245
rect 16865 6057 16877 6233
rect 16911 6057 16923 6233
rect 16865 6045 16923 6057
rect 16983 6233 17041 6245
rect 16983 6057 16995 6233
rect 17029 6057 17041 6233
rect 16983 6045 17041 6057
rect 17101 6233 17159 6245
rect 17101 6057 17113 6233
rect 17147 6057 17159 6233
rect 17101 6045 17159 6057
rect 17495 6233 17553 6245
rect 17495 6057 17507 6233
rect 17541 6057 17553 6233
rect 17495 6045 17553 6057
rect 17613 6233 17671 6245
rect 17613 6057 17625 6233
rect 17659 6057 17671 6233
rect 17613 6045 17671 6057
rect 17731 6233 17789 6245
rect 17731 6057 17743 6233
rect 17777 6057 17789 6233
rect 17731 6045 17789 6057
rect 17849 6233 17907 6245
rect 17849 6057 17861 6233
rect 17895 6057 17907 6233
rect 17849 6045 17907 6057
rect 17978 6057 17990 6433
rect 18024 6057 18036 6433
rect 17978 6045 18036 6057
rect 18096 6433 18154 6445
rect 18096 6057 18108 6433
rect 18142 6057 18154 6433
rect 18096 6045 18154 6057
rect 18214 6433 18272 6445
rect 18214 6057 18226 6433
rect 18260 6057 18272 6433
rect 18214 6045 18272 6057
rect 18332 6433 18390 6445
rect 18332 6057 18344 6433
rect 18378 6057 18390 6433
rect 18332 6045 18390 6057
rect 18450 6433 18508 6445
rect 18450 6057 18462 6433
rect 18496 6057 18508 6433
rect 18450 6045 18508 6057
rect 18568 6433 18626 6445
rect 18568 6057 18580 6433
rect 18614 6057 18626 6433
rect 18568 6045 18626 6057
rect 18686 6433 18744 6445
rect 18686 6057 18698 6433
rect 18732 6057 18744 6433
rect 20046 6431 20104 6443
rect 18686 6045 18744 6057
rect 18816 6233 18874 6245
rect 18816 6057 18828 6233
rect 18862 6057 18874 6233
rect 18816 6045 18874 6057
rect 18934 6233 18992 6245
rect 18934 6057 18946 6233
rect 18980 6057 18992 6233
rect 18934 6045 18992 6057
rect 19052 6233 19110 6245
rect 19052 6057 19064 6233
rect 19098 6057 19110 6233
rect 19052 6045 19110 6057
rect 19170 6233 19228 6245
rect 19170 6057 19182 6233
rect 19216 6057 19228 6233
rect 19170 6045 19228 6057
rect 19563 6231 19621 6243
rect 19563 6055 19575 6231
rect 19609 6055 19621 6231
rect 11829 5740 11887 5752
rect 11829 5364 11841 5740
rect 11875 5364 11887 5740
rect 11829 5352 11887 5364
rect 11947 5740 12005 5752
rect 11947 5364 11959 5740
rect 11993 5364 12005 5740
rect 11947 5352 12005 5364
rect 12065 5740 12123 5752
rect 12065 5364 12077 5740
rect 12111 5364 12123 5740
rect 12065 5352 12123 5364
rect 12183 5740 12241 5752
rect 12183 5364 12195 5740
rect 12229 5364 12241 5740
rect 12183 5352 12241 5364
rect 12301 5740 12359 5752
rect 12301 5364 12313 5740
rect 12347 5364 12359 5740
rect 12301 5352 12359 5364
rect 12419 5740 12477 5752
rect 12419 5364 12431 5740
rect 12465 5364 12477 5740
rect 12419 5352 12477 5364
rect 12537 5740 12595 5752
rect 12537 5364 12549 5740
rect 12583 5364 12595 5740
rect 12537 5352 12595 5364
rect 13898 5742 13956 5754
rect 13898 5366 13910 5742
rect 13944 5366 13956 5742
rect 13898 5354 13956 5366
rect 14016 5742 14074 5754
rect 14016 5366 14028 5742
rect 14062 5366 14074 5742
rect 14016 5354 14074 5366
rect 14134 5742 14192 5754
rect 14134 5366 14146 5742
rect 14180 5366 14192 5742
rect 14134 5354 14192 5366
rect 14252 5742 14310 5754
rect 14252 5366 14264 5742
rect 14298 5366 14310 5742
rect 14252 5354 14310 5366
rect 14370 5742 14428 5754
rect 14370 5366 14382 5742
rect 14416 5366 14428 5742
rect 14370 5354 14428 5366
rect 14488 5742 14546 5754
rect 14488 5366 14500 5742
rect 14534 5366 14546 5742
rect 14488 5354 14546 5366
rect 14606 5742 14664 5754
rect 14606 5366 14618 5742
rect 14652 5366 14664 5742
rect 14606 5354 14664 5366
rect 15966 5740 16024 5752
rect 15966 5364 15978 5740
rect 16012 5364 16024 5740
rect 15966 5352 16024 5364
rect 16084 5740 16142 5752
rect 16084 5364 16096 5740
rect 16130 5364 16142 5740
rect 16084 5352 16142 5364
rect 16202 5740 16260 5752
rect 16202 5364 16214 5740
rect 16248 5364 16260 5740
rect 16202 5352 16260 5364
rect 16320 5740 16378 5752
rect 16320 5364 16332 5740
rect 16366 5364 16378 5740
rect 16320 5352 16378 5364
rect 16438 5740 16496 5752
rect 16438 5364 16450 5740
rect 16484 5364 16496 5740
rect 16438 5352 16496 5364
rect 16556 5740 16614 5752
rect 16556 5364 16568 5740
rect 16602 5364 16614 5740
rect 16556 5352 16614 5364
rect 16674 5740 16732 5752
rect 16674 5364 16686 5740
rect 16720 5364 16732 5740
rect 16674 5352 16732 5364
rect 19563 6043 19621 6055
rect 19681 6231 19739 6243
rect 19681 6055 19693 6231
rect 19727 6055 19739 6231
rect 19681 6043 19739 6055
rect 19799 6231 19857 6243
rect 19799 6055 19811 6231
rect 19845 6055 19857 6231
rect 19799 6043 19857 6055
rect 19917 6231 19975 6243
rect 19917 6055 19929 6231
rect 19963 6055 19975 6231
rect 19917 6043 19975 6055
rect 20046 6055 20058 6431
rect 20092 6055 20104 6431
rect 20046 6043 20104 6055
rect 20164 6431 20222 6443
rect 20164 6055 20176 6431
rect 20210 6055 20222 6431
rect 20164 6043 20222 6055
rect 20282 6431 20340 6443
rect 20282 6055 20294 6431
rect 20328 6055 20340 6431
rect 20282 6043 20340 6055
rect 20400 6431 20458 6443
rect 20400 6055 20412 6431
rect 20446 6055 20458 6431
rect 20400 6043 20458 6055
rect 20518 6431 20576 6443
rect 20518 6055 20530 6431
rect 20564 6055 20576 6431
rect 20518 6043 20576 6055
rect 20636 6431 20694 6443
rect 20636 6055 20648 6431
rect 20682 6055 20694 6431
rect 20636 6043 20694 6055
rect 20754 6431 20812 6443
rect 20754 6055 20766 6431
rect 20800 6055 20812 6431
rect 22115 6433 22173 6445
rect 20754 6043 20812 6055
rect 20884 6231 20942 6243
rect 20884 6055 20896 6231
rect 20930 6055 20942 6231
rect 20884 6043 20942 6055
rect 21002 6231 21060 6243
rect 21002 6055 21014 6231
rect 21048 6055 21060 6231
rect 21002 6043 21060 6055
rect 21120 6231 21178 6243
rect 21120 6055 21132 6231
rect 21166 6055 21178 6231
rect 21120 6043 21178 6055
rect 21238 6231 21296 6243
rect 21238 6055 21250 6231
rect 21284 6055 21296 6231
rect 21238 6043 21296 6055
rect 21632 6233 21690 6245
rect 21632 6057 21644 6233
rect 21678 6057 21690 6233
rect 21632 6045 21690 6057
rect 21750 6233 21808 6245
rect 21750 6057 21762 6233
rect 21796 6057 21808 6233
rect 21750 6045 21808 6057
rect 21868 6233 21926 6245
rect 21868 6057 21880 6233
rect 21914 6057 21926 6233
rect 21868 6045 21926 6057
rect 21986 6233 22044 6245
rect 21986 6057 21998 6233
rect 22032 6057 22044 6233
rect 21986 6045 22044 6057
rect 22115 6057 22127 6433
rect 22161 6057 22173 6433
rect 22115 6045 22173 6057
rect 22233 6433 22291 6445
rect 22233 6057 22245 6433
rect 22279 6057 22291 6433
rect 22233 6045 22291 6057
rect 22351 6433 22409 6445
rect 22351 6057 22363 6433
rect 22397 6057 22409 6433
rect 22351 6045 22409 6057
rect 22469 6433 22527 6445
rect 22469 6057 22481 6433
rect 22515 6057 22527 6433
rect 22469 6045 22527 6057
rect 22587 6433 22645 6445
rect 22587 6057 22599 6433
rect 22633 6057 22645 6433
rect 22587 6045 22645 6057
rect 22705 6433 22763 6445
rect 22705 6057 22717 6433
rect 22751 6057 22763 6433
rect 22705 6045 22763 6057
rect 22823 6433 22881 6445
rect 29952 6479 30352 6491
rect 29952 6445 29964 6479
rect 30340 6445 30352 6479
rect 22823 6057 22835 6433
rect 22869 6057 22881 6433
rect 24183 6431 24241 6443
rect 22823 6045 22881 6057
rect 22953 6233 23011 6245
rect 22953 6057 22965 6233
rect 22999 6057 23011 6233
rect 22953 6045 23011 6057
rect 23071 6233 23129 6245
rect 23071 6057 23083 6233
rect 23117 6057 23129 6233
rect 23071 6045 23129 6057
rect 23189 6233 23247 6245
rect 23189 6057 23201 6233
rect 23235 6057 23247 6233
rect 23189 6045 23247 6057
rect 23307 6233 23365 6245
rect 23307 6057 23319 6233
rect 23353 6057 23365 6233
rect 23307 6045 23365 6057
rect 23700 6231 23758 6243
rect 23700 6055 23712 6231
rect 23746 6055 23758 6231
rect 18035 5740 18093 5752
rect 18035 5364 18047 5740
rect 18081 5364 18093 5740
rect 18035 5352 18093 5364
rect 18153 5740 18211 5752
rect 18153 5364 18165 5740
rect 18199 5364 18211 5740
rect 18153 5352 18211 5364
rect 18271 5740 18329 5752
rect 18271 5364 18283 5740
rect 18317 5364 18329 5740
rect 18271 5352 18329 5364
rect 18389 5740 18447 5752
rect 18389 5364 18401 5740
rect 18435 5364 18447 5740
rect 18389 5352 18447 5364
rect 18507 5740 18565 5752
rect 18507 5364 18519 5740
rect 18553 5364 18565 5740
rect 18507 5352 18565 5364
rect 18625 5740 18683 5752
rect 18625 5364 18637 5740
rect 18671 5364 18683 5740
rect 18625 5352 18683 5364
rect 18743 5740 18801 5752
rect 18743 5364 18755 5740
rect 18789 5364 18801 5740
rect 18743 5352 18801 5364
rect 23700 6043 23758 6055
rect 23818 6231 23876 6243
rect 23818 6055 23830 6231
rect 23864 6055 23876 6231
rect 23818 6043 23876 6055
rect 23936 6231 23994 6243
rect 23936 6055 23948 6231
rect 23982 6055 23994 6231
rect 23936 6043 23994 6055
rect 24054 6231 24112 6243
rect 24054 6055 24066 6231
rect 24100 6055 24112 6231
rect 24054 6043 24112 6055
rect 24183 6055 24195 6431
rect 24229 6055 24241 6431
rect 24183 6043 24241 6055
rect 24301 6431 24359 6443
rect 24301 6055 24313 6431
rect 24347 6055 24359 6431
rect 24301 6043 24359 6055
rect 24419 6431 24477 6443
rect 24419 6055 24431 6431
rect 24465 6055 24477 6431
rect 24419 6043 24477 6055
rect 24537 6431 24595 6443
rect 24537 6055 24549 6431
rect 24583 6055 24595 6431
rect 24537 6043 24595 6055
rect 24655 6431 24713 6443
rect 24655 6055 24667 6431
rect 24701 6055 24713 6431
rect 24655 6043 24713 6055
rect 24773 6431 24831 6443
rect 24773 6055 24785 6431
rect 24819 6055 24831 6431
rect 24773 6043 24831 6055
rect 24891 6431 24949 6443
rect 29952 6433 30352 6445
rect 30645 6536 31045 6548
rect 30645 6502 30657 6536
rect 31033 6502 31045 6536
rect 37793 6540 37805 6716
rect 37839 6540 37851 6716
rect 37793 6528 37851 6540
rect 37911 6716 37969 6728
rect 37911 6540 37923 6716
rect 37957 6540 37969 6716
rect 37911 6528 37969 6540
rect 38029 6716 38087 6728
rect 38029 6540 38041 6716
rect 38075 6540 38087 6716
rect 38029 6528 38087 6540
rect 38147 6716 38205 6728
rect 38147 6540 38159 6716
rect 38193 6540 38205 6716
rect 38147 6528 38205 6540
rect 38265 6716 38323 6728
rect 38265 6540 38277 6716
rect 38311 6540 38323 6716
rect 38265 6528 38323 6540
rect 38383 6716 38441 6728
rect 38383 6540 38395 6716
rect 38429 6540 38441 6716
rect 38383 6528 38441 6540
rect 38501 6716 38559 6728
rect 38501 6540 38513 6716
rect 38547 6540 38559 6716
rect 38501 6528 38559 6540
rect 38619 6716 38677 6728
rect 38619 6540 38631 6716
rect 38665 6540 38677 6716
rect 38619 6528 38677 6540
rect 38737 6716 38795 6728
rect 38737 6540 38749 6716
rect 38783 6540 38795 6716
rect 38737 6528 38795 6540
rect 38855 6716 38913 6728
rect 38855 6540 38867 6716
rect 38901 6540 38913 6716
rect 38855 6528 38913 6540
rect 39689 7210 39747 7222
rect 39689 6834 39701 7210
rect 39735 6834 39747 7210
rect 39689 6822 39747 6834
rect 39807 7210 39865 7222
rect 39807 6834 39819 7210
rect 39853 6834 39865 7210
rect 39807 6822 39865 6834
rect 39925 7210 39983 7222
rect 39925 6834 39937 7210
rect 39971 6834 39983 7210
rect 39925 6822 39983 6834
rect 40043 7210 40101 7222
rect 40043 6834 40055 7210
rect 40089 6834 40101 7210
rect 40043 6822 40101 6834
rect 40161 7210 40219 7222
rect 40161 6834 40173 7210
rect 40207 6834 40219 7210
rect 40161 6822 40219 6834
rect 40279 7210 40337 7222
rect 40279 6834 40291 7210
rect 40325 6834 40337 7210
rect 40279 6822 40337 6834
rect 40397 7210 40455 7222
rect 40397 6834 40409 7210
rect 40443 6834 40455 7210
rect 40397 6822 40455 6834
rect 30645 6490 31045 6502
rect 24891 6055 24903 6431
rect 24937 6055 24949 6431
rect 29952 6361 30352 6373
rect 29952 6327 29964 6361
rect 30340 6327 30352 6361
rect 29952 6315 30352 6327
rect 30645 6418 31045 6430
rect 30645 6384 30657 6418
rect 31033 6384 31045 6418
rect 30645 6372 31045 6384
rect 24891 6043 24949 6055
rect 25021 6231 25079 6243
rect 25021 6055 25033 6231
rect 25067 6055 25079 6231
rect 25021 6043 25079 6055
rect 25139 6231 25197 6243
rect 25139 6055 25151 6231
rect 25185 6055 25197 6231
rect 25139 6043 25197 6055
rect 25257 6231 25315 6243
rect 25257 6055 25269 6231
rect 25303 6055 25315 6231
rect 25257 6043 25315 6055
rect 25375 6231 25433 6243
rect 25375 6055 25387 6231
rect 25421 6055 25433 6231
rect 25375 6043 25433 6055
rect 29952 6243 30352 6255
rect 29952 6209 29964 6243
rect 30340 6209 30352 6243
rect 29952 6197 30352 6209
rect 30645 6300 31045 6312
rect 30645 6266 30657 6300
rect 31033 6266 31045 6300
rect 30645 6254 31045 6266
rect 45811 7615 45823 7791
rect 45857 7615 45869 7791
rect 45811 7603 45869 7615
rect 45929 7791 45987 7803
rect 45929 7615 45941 7791
rect 45975 7615 45987 7791
rect 45929 7603 45987 7615
rect 46047 7791 46105 7803
rect 46047 7615 46059 7791
rect 46093 7615 46105 7791
rect 46047 7603 46105 7615
rect 46165 7791 46223 7803
rect 46165 7615 46177 7791
rect 46211 7615 46223 7791
rect 46165 7603 46223 7615
rect 46295 7615 46307 7991
rect 46341 7615 46353 7991
rect 46295 7603 46353 7615
rect 46413 7991 46471 8003
rect 46413 7615 46425 7991
rect 46459 7615 46471 7991
rect 46413 7603 46471 7615
rect 46531 7991 46589 8003
rect 46531 7615 46543 7991
rect 46577 7615 46589 7991
rect 46531 7603 46589 7615
rect 46649 7991 46707 8003
rect 46649 7615 46661 7991
rect 46695 7615 46707 7991
rect 46649 7603 46707 7615
rect 46767 7991 46825 8003
rect 46767 7615 46779 7991
rect 46813 7615 46825 7991
rect 46767 7603 46825 7615
rect 46885 7991 46943 8003
rect 46885 7615 46897 7991
rect 46931 7615 46943 7991
rect 46885 7603 46943 7615
rect 47003 7991 47061 8003
rect 47003 7615 47015 7991
rect 47049 7615 47061 7991
rect 48193 7991 48251 8003
rect 47003 7603 47061 7615
rect 47132 7791 47190 7803
rect 47132 7615 47144 7791
rect 47178 7615 47190 7791
rect 47132 7603 47190 7615
rect 47250 7791 47308 7803
rect 47250 7615 47262 7791
rect 47296 7615 47308 7791
rect 47250 7603 47308 7615
rect 47368 7791 47426 7803
rect 47368 7615 47380 7791
rect 47414 7615 47426 7791
rect 47368 7603 47426 7615
rect 47486 7791 47544 7803
rect 47486 7615 47498 7791
rect 47532 7615 47544 7791
rect 47486 7603 47544 7615
rect 47709 7791 47767 7803
rect 47709 7615 47721 7791
rect 47755 7615 47767 7791
rect 47709 7603 47767 7615
rect 47827 7791 47885 7803
rect 47827 7615 47839 7791
rect 47873 7615 47885 7791
rect 47827 7603 47885 7615
rect 47945 7791 48003 7803
rect 47945 7615 47957 7791
rect 47991 7615 48003 7791
rect 47945 7603 48003 7615
rect 48063 7791 48121 7803
rect 48063 7615 48075 7791
rect 48109 7615 48121 7791
rect 48063 7603 48121 7615
rect 48193 7615 48205 7991
rect 48239 7615 48251 7991
rect 48193 7603 48251 7615
rect 48311 7991 48369 8003
rect 48311 7615 48323 7991
rect 48357 7615 48369 7991
rect 48311 7603 48369 7615
rect 48429 7991 48487 8003
rect 48429 7615 48441 7991
rect 48475 7615 48487 7991
rect 48429 7603 48487 7615
rect 48547 7991 48605 8003
rect 48547 7615 48559 7991
rect 48593 7615 48605 7991
rect 48547 7603 48605 7615
rect 48665 7991 48723 8003
rect 48665 7615 48677 7991
rect 48711 7615 48723 7991
rect 48665 7603 48723 7615
rect 48783 7991 48841 8003
rect 48783 7615 48795 7991
rect 48829 7615 48841 7991
rect 48783 7603 48841 7615
rect 48901 7991 48959 8003
rect 48901 7615 48913 7991
rect 48947 7615 48959 7991
rect 70513 8295 70913 8307
rect 70513 8261 70525 8295
rect 70901 8261 70913 8295
rect 70513 8249 70913 8261
rect 70513 8177 70913 8189
rect 70513 8143 70525 8177
rect 70901 8143 70913 8177
rect 70513 8131 70913 8143
rect 70513 8059 70913 8071
rect 70513 8025 70525 8059
rect 70901 8025 70913 8059
rect 70513 8013 70913 8025
rect 59574 7991 59632 8003
rect 52949 7923 53007 7935
rect 48901 7603 48959 7615
rect 49030 7791 49088 7803
rect 49030 7615 49042 7791
rect 49076 7615 49088 7791
rect 49030 7603 49088 7615
rect 49148 7791 49206 7803
rect 49148 7615 49160 7791
rect 49194 7615 49206 7791
rect 49148 7603 49206 7615
rect 49266 7791 49324 7803
rect 49266 7615 49278 7791
rect 49312 7615 49324 7791
rect 49266 7603 49324 7615
rect 49384 7791 49442 7803
rect 49384 7615 49396 7791
rect 49430 7615 49442 7791
rect 49384 7603 49442 7615
rect 41587 7210 41645 7222
rect 41587 6834 41599 7210
rect 41633 6834 41645 7210
rect 41587 6822 41645 6834
rect 41705 7210 41763 7222
rect 41705 6834 41717 7210
rect 41751 6834 41763 7210
rect 41705 6822 41763 6834
rect 41823 7210 41881 7222
rect 41823 6834 41835 7210
rect 41869 6834 41881 7210
rect 41823 6822 41881 6834
rect 41941 7210 41999 7222
rect 41941 6834 41953 7210
rect 41987 6834 41999 7210
rect 41941 6822 41999 6834
rect 42059 7210 42117 7222
rect 42059 6834 42071 7210
rect 42105 6834 42117 7210
rect 42059 6822 42117 6834
rect 42177 7210 42235 7222
rect 42177 6834 42189 7210
rect 42223 6834 42235 7210
rect 42177 6822 42235 6834
rect 42295 7210 42353 7222
rect 42295 6834 42307 7210
rect 42341 6834 42353 7210
rect 42295 6822 42353 6834
rect 44342 6804 44400 6816
rect 44342 6628 44354 6804
rect 44388 6628 44400 6804
rect 44342 6616 44400 6628
rect 44460 6804 44518 6816
rect 44460 6628 44472 6804
rect 44506 6628 44518 6804
rect 44460 6616 44518 6628
rect 44578 6804 44636 6816
rect 44578 6628 44590 6804
rect 44624 6628 44636 6804
rect 44578 6616 44636 6628
rect 44696 6804 44754 6816
rect 44696 6628 44708 6804
rect 44742 6628 44754 6804
rect 44696 6616 44754 6628
rect 44814 6804 44872 6816
rect 44814 6628 44826 6804
rect 44860 6628 44872 6804
rect 44814 6616 44872 6628
rect 44932 6804 44990 6816
rect 44932 6628 44944 6804
rect 44978 6628 44990 6804
rect 44932 6616 44990 6628
rect 45050 6804 45108 6816
rect 45050 6628 45062 6804
rect 45096 6628 45108 6804
rect 45050 6616 45108 6628
rect 45168 6804 45226 6816
rect 45168 6628 45180 6804
rect 45214 6628 45226 6804
rect 45168 6616 45226 6628
rect 45286 6804 45344 6816
rect 45286 6628 45298 6804
rect 45332 6628 45344 6804
rect 45286 6616 45344 6628
rect 45404 6804 45462 6816
rect 45404 6628 45416 6804
rect 45450 6628 45462 6804
rect 45404 6616 45462 6628
rect 46238 7298 46296 7310
rect 46238 6922 46250 7298
rect 46284 6922 46296 7298
rect 46238 6910 46296 6922
rect 46356 7298 46414 7310
rect 46356 6922 46368 7298
rect 46402 6922 46414 7298
rect 46356 6910 46414 6922
rect 46474 7298 46532 7310
rect 46474 6922 46486 7298
rect 46520 6922 46532 7298
rect 46474 6910 46532 6922
rect 46592 7298 46650 7310
rect 46592 6922 46604 7298
rect 46638 6922 46650 7298
rect 46592 6910 46650 6922
rect 46710 7298 46768 7310
rect 46710 6922 46722 7298
rect 46756 6922 46768 7298
rect 46710 6910 46768 6922
rect 46828 7298 46886 7310
rect 46828 6922 46840 7298
rect 46874 6922 46886 7298
rect 46828 6910 46886 6922
rect 46946 7298 47004 7310
rect 46946 6922 46958 7298
rect 46992 6922 47004 7298
rect 46946 6910 47004 6922
rect 30645 6182 31045 6194
rect 30645 6148 30657 6182
rect 31033 6148 31045 6182
rect 29952 6125 30352 6137
rect 30645 6136 31045 6148
rect 29952 6091 29964 6125
rect 30340 6091 30352 6125
rect 29952 6079 30352 6091
rect 20103 5738 20161 5750
rect 20103 5362 20115 5738
rect 20149 5362 20161 5738
rect 20103 5350 20161 5362
rect 20221 5738 20279 5750
rect 20221 5362 20233 5738
rect 20267 5362 20279 5738
rect 20221 5350 20279 5362
rect 20339 5738 20397 5750
rect 20339 5362 20351 5738
rect 20385 5362 20397 5738
rect 20339 5350 20397 5362
rect 20457 5738 20515 5750
rect 20457 5362 20469 5738
rect 20503 5362 20515 5738
rect 20457 5350 20515 5362
rect 20575 5738 20633 5750
rect 20575 5362 20587 5738
rect 20621 5362 20633 5738
rect 20575 5350 20633 5362
rect 20693 5738 20751 5750
rect 20693 5362 20705 5738
rect 20739 5362 20751 5738
rect 20693 5350 20751 5362
rect 20811 5738 20869 5750
rect 20811 5362 20823 5738
rect 20857 5362 20869 5738
rect 20811 5350 20869 5362
rect 22172 5740 22230 5752
rect 22172 5364 22184 5740
rect 22218 5364 22230 5740
rect 22172 5352 22230 5364
rect 22290 5740 22348 5752
rect 22290 5364 22302 5740
rect 22336 5364 22348 5740
rect 22290 5352 22348 5364
rect 22408 5740 22466 5752
rect 22408 5364 22420 5740
rect 22454 5364 22466 5740
rect 22408 5352 22466 5364
rect 22526 5740 22584 5752
rect 22526 5364 22538 5740
rect 22572 5364 22584 5740
rect 22526 5352 22584 5364
rect 22644 5740 22702 5752
rect 22644 5364 22656 5740
rect 22690 5364 22702 5740
rect 22644 5352 22702 5364
rect 22762 5740 22820 5752
rect 22762 5364 22774 5740
rect 22808 5364 22820 5740
rect 22762 5352 22820 5364
rect 22880 5740 22938 5752
rect 22880 5364 22892 5740
rect 22926 5364 22938 5740
rect 22880 5352 22938 5364
rect 24240 5738 24298 5750
rect 24240 5362 24252 5738
rect 24286 5362 24298 5738
rect 24240 5350 24298 5362
rect 24358 5738 24416 5750
rect 24358 5362 24370 5738
rect 24404 5362 24416 5738
rect 24358 5350 24416 5362
rect 24476 5738 24534 5750
rect 24476 5362 24488 5738
rect 24522 5362 24534 5738
rect 24476 5350 24534 5362
rect 24594 5738 24652 5750
rect 24594 5362 24606 5738
rect 24640 5362 24652 5738
rect 24594 5350 24652 5362
rect 24712 5738 24770 5750
rect 24712 5362 24724 5738
rect 24758 5362 24770 5738
rect 24712 5350 24770 5362
rect 24830 5738 24888 5750
rect 24830 5362 24842 5738
rect 24876 5362 24888 5738
rect 24830 5350 24888 5362
rect 24948 5738 25006 5750
rect 24948 5362 24960 5738
rect 24994 5362 25006 5738
rect 24948 5350 25006 5362
rect 29952 6007 30352 6019
rect 29952 5973 29964 6007
rect 30340 5973 30352 6007
rect 29952 5961 30352 5973
rect 29952 5889 30352 5901
rect 29952 5855 29964 5889
rect 30340 5855 30352 5889
rect 29952 5843 30352 5855
rect 30645 6064 31045 6076
rect 30645 6030 30657 6064
rect 31033 6030 31045 6064
rect 30645 6018 31045 6030
rect 30645 5946 31045 5958
rect 30645 5912 30657 5946
rect 31033 5912 31045 5946
rect 30645 5900 31045 5912
rect 52465 7723 52523 7735
rect 52465 7547 52477 7723
rect 52511 7547 52523 7723
rect 52465 7535 52523 7547
rect 52583 7723 52641 7735
rect 52583 7547 52595 7723
rect 52629 7547 52641 7723
rect 52583 7535 52641 7547
rect 52701 7723 52759 7735
rect 52701 7547 52713 7723
rect 52747 7547 52759 7723
rect 52701 7535 52759 7547
rect 52819 7723 52877 7735
rect 52819 7547 52831 7723
rect 52865 7547 52877 7723
rect 52819 7535 52877 7547
rect 52949 7547 52961 7923
rect 52995 7547 53007 7923
rect 52949 7535 53007 7547
rect 53067 7923 53125 7935
rect 53067 7547 53079 7923
rect 53113 7547 53125 7923
rect 53067 7535 53125 7547
rect 53185 7923 53243 7935
rect 53185 7547 53197 7923
rect 53231 7547 53243 7923
rect 53185 7535 53243 7547
rect 53303 7923 53361 7935
rect 53303 7547 53315 7923
rect 53349 7547 53361 7923
rect 53303 7535 53361 7547
rect 53421 7923 53479 7935
rect 53421 7547 53433 7923
rect 53467 7547 53479 7923
rect 53421 7535 53479 7547
rect 53539 7923 53597 7935
rect 53539 7547 53551 7923
rect 53585 7547 53597 7923
rect 53539 7535 53597 7547
rect 53657 7923 53715 7935
rect 53657 7547 53669 7923
rect 53703 7547 53715 7923
rect 54847 7923 54905 7935
rect 53657 7535 53715 7547
rect 53786 7723 53844 7735
rect 53786 7547 53798 7723
rect 53832 7547 53844 7723
rect 53786 7535 53844 7547
rect 53904 7723 53962 7735
rect 53904 7547 53916 7723
rect 53950 7547 53962 7723
rect 53904 7535 53962 7547
rect 54022 7723 54080 7735
rect 54022 7547 54034 7723
rect 54068 7547 54080 7723
rect 54022 7535 54080 7547
rect 54140 7723 54198 7735
rect 54140 7547 54152 7723
rect 54186 7547 54198 7723
rect 54140 7535 54198 7547
rect 54363 7723 54421 7735
rect 54363 7547 54375 7723
rect 54409 7547 54421 7723
rect 54363 7535 54421 7547
rect 54481 7723 54539 7735
rect 54481 7547 54493 7723
rect 54527 7547 54539 7723
rect 54481 7535 54539 7547
rect 54599 7723 54657 7735
rect 54599 7547 54611 7723
rect 54645 7547 54657 7723
rect 54599 7535 54657 7547
rect 54717 7723 54775 7735
rect 54717 7547 54729 7723
rect 54763 7547 54775 7723
rect 54717 7535 54775 7547
rect 54847 7547 54859 7923
rect 54893 7547 54905 7923
rect 54847 7535 54905 7547
rect 54965 7923 55023 7935
rect 54965 7547 54977 7923
rect 55011 7547 55023 7923
rect 54965 7535 55023 7547
rect 55083 7923 55141 7935
rect 55083 7547 55095 7923
rect 55129 7547 55141 7923
rect 55083 7535 55141 7547
rect 55201 7923 55259 7935
rect 55201 7547 55213 7923
rect 55247 7547 55259 7923
rect 55201 7535 55259 7547
rect 55319 7923 55377 7935
rect 55319 7547 55331 7923
rect 55365 7547 55377 7923
rect 55319 7535 55377 7547
rect 55437 7923 55495 7935
rect 55437 7547 55449 7923
rect 55483 7547 55495 7923
rect 55437 7535 55495 7547
rect 55555 7923 55613 7935
rect 55555 7547 55567 7923
rect 55601 7547 55613 7923
rect 55555 7535 55613 7547
rect 55684 7723 55742 7735
rect 55684 7547 55696 7723
rect 55730 7547 55742 7723
rect 55684 7535 55742 7547
rect 55802 7723 55860 7735
rect 55802 7547 55814 7723
rect 55848 7547 55860 7723
rect 55802 7535 55860 7547
rect 55920 7723 55978 7735
rect 55920 7547 55932 7723
rect 55966 7547 55978 7723
rect 55920 7535 55978 7547
rect 56038 7723 56096 7735
rect 56038 7547 56050 7723
rect 56084 7547 56096 7723
rect 59090 7791 59148 7803
rect 56038 7535 56096 7547
rect 48136 7298 48194 7310
rect 48136 6922 48148 7298
rect 48182 6922 48194 7298
rect 48136 6910 48194 6922
rect 48254 7298 48312 7310
rect 48254 6922 48266 7298
rect 48300 6922 48312 7298
rect 48254 6910 48312 6922
rect 48372 7298 48430 7310
rect 48372 6922 48384 7298
rect 48418 6922 48430 7298
rect 48372 6910 48430 6922
rect 48490 7298 48548 7310
rect 48490 6922 48502 7298
rect 48536 6922 48548 7298
rect 48490 6910 48548 6922
rect 48608 7298 48666 7310
rect 48608 6922 48620 7298
rect 48654 6922 48666 7298
rect 48608 6910 48666 6922
rect 48726 7298 48784 7310
rect 48726 6922 48738 7298
rect 48772 6922 48784 7298
rect 48726 6910 48784 6922
rect 48844 7298 48902 7310
rect 48844 6922 48856 7298
rect 48890 6922 48902 7298
rect 48844 6910 48902 6922
rect 50996 6736 51054 6748
rect 50996 6560 51008 6736
rect 51042 6560 51054 6736
rect 50996 6548 51054 6560
rect 51114 6736 51172 6748
rect 51114 6560 51126 6736
rect 51160 6560 51172 6736
rect 51114 6548 51172 6560
rect 51232 6736 51290 6748
rect 51232 6560 51244 6736
rect 51278 6560 51290 6736
rect 51232 6548 51290 6560
rect 51350 6736 51408 6748
rect 51350 6560 51362 6736
rect 51396 6560 51408 6736
rect 51350 6548 51408 6560
rect 51468 6736 51526 6748
rect 51468 6560 51480 6736
rect 51514 6560 51526 6736
rect 51468 6548 51526 6560
rect 51586 6736 51644 6748
rect 51586 6560 51598 6736
rect 51632 6560 51644 6736
rect 51586 6548 51644 6560
rect 51704 6736 51762 6748
rect 51704 6560 51716 6736
rect 51750 6560 51762 6736
rect 51704 6548 51762 6560
rect 51822 6736 51880 6748
rect 51822 6560 51834 6736
rect 51868 6560 51880 6736
rect 51822 6548 51880 6560
rect 51940 6736 51998 6748
rect 51940 6560 51952 6736
rect 51986 6560 51998 6736
rect 51940 6548 51998 6560
rect 52058 6736 52116 6748
rect 52058 6560 52070 6736
rect 52104 6560 52116 6736
rect 52058 6548 52116 6560
rect 52892 7230 52950 7242
rect 52892 6854 52904 7230
rect 52938 6854 52950 7230
rect 52892 6842 52950 6854
rect 53010 7230 53068 7242
rect 53010 6854 53022 7230
rect 53056 6854 53068 7230
rect 53010 6842 53068 6854
rect 53128 7230 53186 7242
rect 53128 6854 53140 7230
rect 53174 6854 53186 7230
rect 53128 6842 53186 6854
rect 53246 7230 53304 7242
rect 53246 6854 53258 7230
rect 53292 6854 53304 7230
rect 53246 6842 53304 6854
rect 53364 7230 53422 7242
rect 53364 6854 53376 7230
rect 53410 6854 53422 7230
rect 53364 6842 53422 6854
rect 53482 7230 53540 7242
rect 53482 6854 53494 7230
rect 53528 6854 53540 7230
rect 53482 6842 53540 6854
rect 53600 7230 53658 7242
rect 53600 6854 53612 7230
rect 53646 6854 53658 7230
rect 53600 6842 53658 6854
rect 59090 7615 59102 7791
rect 59136 7615 59148 7791
rect 59090 7603 59148 7615
rect 59208 7791 59266 7803
rect 59208 7615 59220 7791
rect 59254 7615 59266 7791
rect 59208 7603 59266 7615
rect 59326 7791 59384 7803
rect 59326 7615 59338 7791
rect 59372 7615 59384 7791
rect 59326 7603 59384 7615
rect 59444 7791 59502 7803
rect 59444 7615 59456 7791
rect 59490 7615 59502 7791
rect 59444 7603 59502 7615
rect 59574 7615 59586 7991
rect 59620 7615 59632 7991
rect 59574 7603 59632 7615
rect 59692 7991 59750 8003
rect 59692 7615 59704 7991
rect 59738 7615 59750 7991
rect 59692 7603 59750 7615
rect 59810 7991 59868 8003
rect 59810 7615 59822 7991
rect 59856 7615 59868 7991
rect 59810 7603 59868 7615
rect 59928 7991 59986 8003
rect 59928 7615 59940 7991
rect 59974 7615 59986 7991
rect 59928 7603 59986 7615
rect 60046 7991 60104 8003
rect 60046 7615 60058 7991
rect 60092 7615 60104 7991
rect 60046 7603 60104 7615
rect 60164 7991 60222 8003
rect 60164 7615 60176 7991
rect 60210 7615 60222 7991
rect 60164 7603 60222 7615
rect 60282 7991 60340 8003
rect 60282 7615 60294 7991
rect 60328 7615 60340 7991
rect 61472 7991 61530 8003
rect 60282 7603 60340 7615
rect 60411 7791 60469 7803
rect 60411 7615 60423 7791
rect 60457 7615 60469 7791
rect 60411 7603 60469 7615
rect 60529 7791 60587 7803
rect 60529 7615 60541 7791
rect 60575 7615 60587 7791
rect 60529 7603 60587 7615
rect 60647 7791 60705 7803
rect 60647 7615 60659 7791
rect 60693 7615 60705 7791
rect 60647 7603 60705 7615
rect 60765 7791 60823 7803
rect 60765 7615 60777 7791
rect 60811 7615 60823 7791
rect 60765 7603 60823 7615
rect 60988 7791 61046 7803
rect 60988 7615 61000 7791
rect 61034 7615 61046 7791
rect 60988 7603 61046 7615
rect 61106 7791 61164 7803
rect 61106 7615 61118 7791
rect 61152 7615 61164 7791
rect 61106 7603 61164 7615
rect 61224 7791 61282 7803
rect 61224 7615 61236 7791
rect 61270 7615 61282 7791
rect 61224 7603 61282 7615
rect 61342 7791 61400 7803
rect 61342 7615 61354 7791
rect 61388 7615 61400 7791
rect 61342 7603 61400 7615
rect 61472 7615 61484 7991
rect 61518 7615 61530 7991
rect 61472 7603 61530 7615
rect 61590 7991 61648 8003
rect 61590 7615 61602 7991
rect 61636 7615 61648 7991
rect 61590 7603 61648 7615
rect 61708 7991 61766 8003
rect 61708 7615 61720 7991
rect 61754 7615 61766 7991
rect 61708 7603 61766 7615
rect 61826 7991 61884 8003
rect 61826 7615 61838 7991
rect 61872 7615 61884 7991
rect 61826 7603 61884 7615
rect 61944 7991 62002 8003
rect 61944 7615 61956 7991
rect 61990 7615 62002 7991
rect 61944 7603 62002 7615
rect 62062 7991 62120 8003
rect 62062 7615 62074 7991
rect 62108 7615 62120 7991
rect 62062 7603 62120 7615
rect 62180 7991 62238 8003
rect 62180 7615 62192 7991
rect 62226 7615 62238 7991
rect 70513 7941 70913 7953
rect 70513 7907 70525 7941
rect 70901 7907 70913 7941
rect 70513 7895 70913 7907
rect 70513 7823 70913 7835
rect 62180 7603 62238 7615
rect 62309 7791 62367 7803
rect 62309 7615 62321 7791
rect 62355 7615 62367 7791
rect 62309 7603 62367 7615
rect 62427 7791 62485 7803
rect 62427 7615 62439 7791
rect 62473 7615 62485 7791
rect 62427 7603 62485 7615
rect 62545 7791 62603 7803
rect 62545 7615 62557 7791
rect 62591 7615 62603 7791
rect 62545 7603 62603 7615
rect 62663 7791 62721 7803
rect 62663 7615 62675 7791
rect 62709 7615 62721 7791
rect 70513 7789 70525 7823
rect 70901 7789 70913 7823
rect 70513 7777 70913 7789
rect 62663 7603 62721 7615
rect 65708 7694 65766 7706
rect 54790 7230 54848 7242
rect 54790 6854 54802 7230
rect 54836 6854 54848 7230
rect 54790 6842 54848 6854
rect 54908 7230 54966 7242
rect 54908 6854 54920 7230
rect 54954 6854 54966 7230
rect 54908 6842 54966 6854
rect 55026 7230 55084 7242
rect 55026 6854 55038 7230
rect 55072 6854 55084 7230
rect 55026 6842 55084 6854
rect 55144 7230 55202 7242
rect 55144 6854 55156 7230
rect 55190 6854 55202 7230
rect 55144 6842 55202 6854
rect 55262 7230 55320 7242
rect 55262 6854 55274 7230
rect 55308 6854 55320 7230
rect 55262 6842 55320 6854
rect 55380 7230 55438 7242
rect 55380 6854 55392 7230
rect 55426 6854 55438 7230
rect 55380 6842 55438 6854
rect 55498 7230 55556 7242
rect 55498 6854 55510 7230
rect 55544 6854 55556 7230
rect 55498 6842 55556 6854
rect 57621 6804 57679 6816
rect 57621 6628 57633 6804
rect 57667 6628 57679 6804
rect 57621 6616 57679 6628
rect 57739 6804 57797 6816
rect 57739 6628 57751 6804
rect 57785 6628 57797 6804
rect 57739 6616 57797 6628
rect 57857 6804 57915 6816
rect 57857 6628 57869 6804
rect 57903 6628 57915 6804
rect 57857 6616 57915 6628
rect 57975 6804 58033 6816
rect 57975 6628 57987 6804
rect 58021 6628 58033 6804
rect 57975 6616 58033 6628
rect 58093 6804 58151 6816
rect 58093 6628 58105 6804
rect 58139 6628 58151 6804
rect 58093 6616 58151 6628
rect 58211 6804 58269 6816
rect 58211 6628 58223 6804
rect 58257 6628 58269 6804
rect 58211 6616 58269 6628
rect 58329 6804 58387 6816
rect 58329 6628 58341 6804
rect 58375 6628 58387 6804
rect 58329 6616 58387 6628
rect 58447 6804 58505 6816
rect 58447 6628 58459 6804
rect 58493 6628 58505 6804
rect 58447 6616 58505 6628
rect 58565 6804 58623 6816
rect 58565 6628 58577 6804
rect 58611 6628 58623 6804
rect 58565 6616 58623 6628
rect 58683 6804 58741 6816
rect 58683 6628 58695 6804
rect 58729 6628 58741 6804
rect 58683 6616 58741 6628
rect 59517 7298 59575 7310
rect 59517 6922 59529 7298
rect 59563 6922 59575 7298
rect 59517 6910 59575 6922
rect 59635 7298 59693 7310
rect 59635 6922 59647 7298
rect 59681 6922 59693 7298
rect 59635 6910 59693 6922
rect 59753 7298 59811 7310
rect 59753 6922 59765 7298
rect 59799 6922 59811 7298
rect 59753 6910 59811 6922
rect 59871 7298 59929 7310
rect 59871 6922 59883 7298
rect 59917 6922 59929 7298
rect 59871 6910 59929 6922
rect 59989 7298 60047 7310
rect 59989 6922 60001 7298
rect 60035 6922 60047 7298
rect 59989 6910 60047 6922
rect 60107 7298 60165 7310
rect 60107 6922 60119 7298
rect 60153 6922 60165 7298
rect 60107 6910 60165 6922
rect 60225 7298 60283 7310
rect 60225 6922 60237 7298
rect 60271 6922 60283 7298
rect 60225 6910 60283 6922
rect 29952 5771 30352 5783
rect 29952 5737 29964 5771
rect 30340 5737 30352 5771
rect 29952 5725 30352 5737
rect 30152 5642 30352 5654
rect 30152 5608 30164 5642
rect 30340 5608 30352 5642
rect 30152 5596 30352 5608
rect 30645 5828 31045 5840
rect 30645 5794 30657 5828
rect 31033 5794 31045 5828
rect 65224 7494 65282 7506
rect 61415 7298 61473 7310
rect 61415 6922 61427 7298
rect 61461 6922 61473 7298
rect 61415 6910 61473 6922
rect 61533 7298 61591 7310
rect 61533 6922 61545 7298
rect 61579 6922 61591 7298
rect 61533 6910 61591 6922
rect 61651 7298 61709 7310
rect 61651 6922 61663 7298
rect 61697 6922 61709 7298
rect 61651 6910 61709 6922
rect 61769 7298 61827 7310
rect 61769 6922 61781 7298
rect 61815 6922 61827 7298
rect 61769 6910 61827 6922
rect 61887 7298 61945 7310
rect 61887 6922 61899 7298
rect 61933 6922 61945 7298
rect 61887 6910 61945 6922
rect 62005 7298 62063 7310
rect 62005 6922 62017 7298
rect 62051 6922 62063 7298
rect 62005 6910 62063 6922
rect 62123 7298 62181 7310
rect 62123 6922 62135 7298
rect 62169 6922 62181 7298
rect 62123 6910 62181 6922
rect 65224 7318 65236 7494
rect 65270 7318 65282 7494
rect 65224 7306 65282 7318
rect 65342 7494 65400 7506
rect 65342 7318 65354 7494
rect 65388 7318 65400 7494
rect 65342 7306 65400 7318
rect 65460 7494 65518 7506
rect 65460 7318 65472 7494
rect 65506 7318 65518 7494
rect 65460 7306 65518 7318
rect 65578 7494 65636 7506
rect 65578 7318 65590 7494
rect 65624 7318 65636 7494
rect 65578 7306 65636 7318
rect 65708 7318 65720 7694
rect 65754 7318 65766 7694
rect 65708 7306 65766 7318
rect 65826 7694 65884 7706
rect 65826 7318 65838 7694
rect 65872 7318 65884 7694
rect 65826 7306 65884 7318
rect 65944 7694 66002 7706
rect 65944 7318 65956 7694
rect 65990 7318 66002 7694
rect 65944 7306 66002 7318
rect 66062 7694 66120 7706
rect 66062 7318 66074 7694
rect 66108 7318 66120 7694
rect 66062 7306 66120 7318
rect 66180 7694 66238 7706
rect 66180 7318 66192 7694
rect 66226 7318 66238 7694
rect 66180 7306 66238 7318
rect 66298 7694 66356 7706
rect 66298 7318 66310 7694
rect 66344 7318 66356 7694
rect 66298 7306 66356 7318
rect 66416 7694 66474 7706
rect 66416 7318 66428 7694
rect 66462 7318 66474 7694
rect 70513 7704 70913 7716
rect 70513 7670 70525 7704
rect 70901 7670 70913 7704
rect 70513 7658 70913 7670
rect 66416 7306 66474 7318
rect 66545 7494 66603 7506
rect 66545 7318 66557 7494
rect 66591 7318 66603 7494
rect 66545 7306 66603 7318
rect 66663 7494 66721 7506
rect 66663 7318 66675 7494
rect 66709 7318 66721 7494
rect 66663 7306 66721 7318
rect 66781 7494 66839 7506
rect 66781 7318 66793 7494
rect 66827 7318 66839 7494
rect 66781 7306 66839 7318
rect 66899 7494 66957 7506
rect 70513 7586 70913 7598
rect 70513 7552 70525 7586
rect 70901 7552 70913 7586
rect 70513 7540 70913 7552
rect 66899 7318 66911 7494
rect 66945 7318 66957 7494
rect 66899 7306 66957 7318
rect 67017 7491 67075 7503
rect 67017 7315 67029 7491
rect 67063 7315 67075 7491
rect 67017 7303 67075 7315
rect 67135 7491 67193 7503
rect 67135 7315 67147 7491
rect 67181 7315 67193 7491
rect 67135 7303 67193 7315
rect 67253 7491 67311 7503
rect 67253 7315 67265 7491
rect 67299 7315 67311 7491
rect 67253 7303 67311 7315
rect 67371 7491 67429 7503
rect 67371 7315 67383 7491
rect 67417 7315 67429 7491
rect 67371 7303 67429 7315
rect 67489 7491 67547 7503
rect 67489 7315 67501 7491
rect 67535 7315 67547 7491
rect 67489 7303 67547 7315
rect 67607 7491 67665 7503
rect 67607 7315 67619 7491
rect 67653 7315 67665 7491
rect 67607 7303 67665 7315
rect 67725 7491 67783 7503
rect 67725 7315 67737 7491
rect 67771 7315 67783 7491
rect 67725 7303 67783 7315
rect 67843 7491 67901 7503
rect 67843 7315 67855 7491
rect 67889 7315 67901 7491
rect 67843 7303 67901 7315
rect 67961 7491 68019 7503
rect 67961 7315 67973 7491
rect 68007 7315 68019 7491
rect 67961 7303 68019 7315
rect 68079 7491 68137 7503
rect 68079 7315 68091 7491
rect 68125 7315 68137 7491
rect 70513 7468 70913 7480
rect 70513 7434 70525 7468
rect 70901 7434 70913 7468
rect 70513 7422 70913 7434
rect 68079 7303 68137 7315
rect 70513 7350 70913 7362
rect 70513 7316 70525 7350
rect 70901 7316 70913 7350
rect 70513 7304 70913 7316
rect 65651 7001 65709 7013
rect 63409 6386 63467 6398
rect 63409 6210 63421 6386
rect 63455 6210 63467 6386
rect 63409 6198 63467 6210
rect 63527 6386 63585 6398
rect 63527 6210 63539 6386
rect 63573 6210 63585 6386
rect 63527 6198 63585 6210
rect 63645 6386 63703 6398
rect 63645 6210 63657 6386
rect 63691 6210 63703 6386
rect 63645 6198 63703 6210
rect 63763 6386 63821 6398
rect 63763 6210 63775 6386
rect 63809 6210 63821 6386
rect 63763 6198 63821 6210
rect 63881 6386 63939 6398
rect 63881 6210 63893 6386
rect 63927 6210 63939 6386
rect 63881 6198 63939 6210
rect 63999 6386 64057 6398
rect 63999 6210 64011 6386
rect 64045 6210 64057 6386
rect 63999 6198 64057 6210
rect 64117 6386 64175 6398
rect 64117 6210 64129 6386
rect 64163 6210 64175 6386
rect 64117 6198 64175 6210
rect 64235 6386 64293 6398
rect 64235 6210 64247 6386
rect 64281 6210 64293 6386
rect 64235 6198 64293 6210
rect 64353 6386 64411 6398
rect 64353 6210 64365 6386
rect 64399 6210 64411 6386
rect 64353 6198 64411 6210
rect 64471 6386 64529 6398
rect 64471 6210 64483 6386
rect 64517 6210 64529 6386
rect 65651 6625 65663 7001
rect 65697 6625 65709 7001
rect 65651 6613 65709 6625
rect 65769 7001 65827 7013
rect 65769 6625 65781 7001
rect 65815 6625 65827 7001
rect 65769 6613 65827 6625
rect 65887 7001 65945 7013
rect 65887 6625 65899 7001
rect 65933 6625 65945 7001
rect 65887 6613 65945 6625
rect 66005 7001 66063 7013
rect 66005 6625 66017 7001
rect 66051 6625 66063 7001
rect 66005 6613 66063 6625
rect 66123 7001 66181 7013
rect 66123 6625 66135 7001
rect 66169 6625 66181 7001
rect 66123 6613 66181 6625
rect 66241 7001 66299 7013
rect 66241 6625 66253 7001
rect 66287 6625 66299 7001
rect 66241 6613 66299 6625
rect 66359 7001 66417 7013
rect 66359 6625 66371 7001
rect 66405 6625 66417 7001
rect 66359 6613 66417 6625
rect 70713 7231 70913 7243
rect 70713 7197 70725 7231
rect 70901 7197 70913 7231
rect 70713 7185 70913 7197
rect 70713 7113 70913 7125
rect 70713 7079 70725 7113
rect 70901 7079 70913 7113
rect 70713 7067 70913 7079
rect 70713 6995 70913 7007
rect 70713 6961 70725 6995
rect 70901 6961 70913 6995
rect 70713 6949 70913 6961
rect 70713 6877 70913 6889
rect 70713 6843 70725 6877
rect 70901 6843 70913 6877
rect 70713 6831 70913 6843
rect 70713 6295 70913 6307
rect 64471 6198 64529 6210
rect 30645 5782 31045 5794
rect 30152 5524 30352 5536
rect 30152 5490 30164 5524
rect 30340 5490 30352 5524
rect 70713 6261 70725 6295
rect 70901 6261 70913 6295
rect 70713 6249 70913 6261
rect 70713 6177 70913 6189
rect 70713 6143 70725 6177
rect 70901 6143 70913 6177
rect 70713 6131 70913 6143
rect 70713 6059 70913 6071
rect 70713 6025 70725 6059
rect 70901 6025 70913 6059
rect 70713 6013 70913 6025
rect 70713 5941 70913 5953
rect 70713 5907 70725 5941
rect 70901 5907 70913 5941
rect 70713 5866 70913 5907
rect 70513 5854 70913 5866
rect 70513 5820 70525 5854
rect 70901 5820 70913 5854
rect 70513 5808 70913 5820
rect 70513 5736 70913 5748
rect 70513 5702 70525 5736
rect 70901 5702 70913 5736
rect 70513 5690 70913 5702
rect 70513 5618 70913 5630
rect 70513 5584 70525 5618
rect 70901 5584 70913 5618
rect 70513 5572 70913 5584
rect 30152 5478 30352 5490
rect 70513 5500 70913 5512
rect 70513 5466 70525 5500
rect 70901 5466 70913 5500
rect 70513 5454 70913 5466
rect 30152 5406 30352 5418
rect 30152 5372 30164 5406
rect 30340 5372 30352 5406
rect 30152 5360 30352 5372
rect 70513 5387 70913 5399
rect 70513 5353 70525 5387
rect 70901 5353 70913 5387
rect 70513 5341 70913 5353
rect 30152 5288 30352 5300
rect 30152 5254 30164 5288
rect 30340 5254 30352 5288
rect 30152 5242 30352 5254
rect 70513 5269 70913 5281
rect 70513 5235 70525 5269
rect 70901 5235 70913 5269
rect 70513 5223 70913 5235
rect 70513 5151 70913 5163
rect 70513 5117 70525 5151
rect 70901 5117 70913 5151
rect 70513 5105 70913 5117
rect 70513 5033 70913 5045
rect 70513 4999 70525 5033
rect 70901 4999 70913 5033
rect 70513 4987 70913 4999
rect 30152 4894 30352 4906
rect 30152 4860 30164 4894
rect 30340 4860 30352 4894
rect 30152 4848 30352 4860
rect 30152 4776 30352 4788
rect 30152 4742 30164 4776
rect 30340 4742 30352 4776
rect 30152 4730 30352 4742
rect 70513 4915 70913 4927
rect 70513 4881 70525 4915
rect 70901 4881 70913 4915
rect 70513 4869 70913 4881
rect 70513 4797 70913 4809
rect 70513 4763 70525 4797
rect 70901 4763 70913 4797
rect 70513 4751 70913 4763
rect 30152 4658 30352 4670
rect 30152 4624 30164 4658
rect 30340 4624 30352 4658
rect 30152 4612 30352 4624
rect 30152 4540 30352 4552
rect 30152 4506 30164 4540
rect 30340 4506 30352 4540
rect 30152 4494 30352 4506
rect 29952 4410 30352 4422
rect 29952 4376 29964 4410
rect 30340 4376 30352 4410
rect 29952 4364 30352 4376
rect 30645 4467 31045 4479
rect 30645 4433 30657 4467
rect 31033 4433 31045 4467
rect 30645 4421 31045 4433
rect 29952 4292 30352 4304
rect 29952 4258 29964 4292
rect 30340 4258 30352 4292
rect 29952 4246 30352 4258
rect 30645 4349 31045 4361
rect 30645 4315 30657 4349
rect 31033 4315 31045 4349
rect 30645 4303 31045 4315
rect 34867 4374 34925 4386
rect 29952 4174 30352 4186
rect 29952 4140 29964 4174
rect 30340 4140 30352 4174
rect 29952 4128 30352 4140
rect 30645 4231 31045 4243
rect 30645 4197 30657 4231
rect 31033 4197 31045 4231
rect 30645 4185 31045 4197
rect 34867 4198 34879 4374
rect 34913 4198 34925 4374
rect 34867 4186 34925 4198
rect 34985 4374 35043 4386
rect 34985 4198 34997 4374
rect 35031 4198 35043 4374
rect 34985 4186 35043 4198
rect 35103 4374 35161 4386
rect 35103 4198 35115 4374
rect 35149 4198 35161 4374
rect 35103 4186 35161 4198
rect 35221 4374 35279 4386
rect 35221 4198 35233 4374
rect 35267 4198 35279 4374
rect 35221 4186 35279 4198
rect 35339 4374 35397 4386
rect 35339 4198 35351 4374
rect 35385 4198 35397 4374
rect 35339 4186 35397 4198
rect 35457 4374 35515 4386
rect 35457 4198 35469 4374
rect 35503 4198 35515 4374
rect 35457 4186 35515 4198
rect 35575 4374 35633 4386
rect 35575 4198 35587 4374
rect 35621 4198 35633 4374
rect 35575 4186 35633 4198
rect 35693 4374 35751 4386
rect 35693 4198 35705 4374
rect 35739 4198 35751 4374
rect 35693 4186 35751 4198
rect 35811 4374 35869 4386
rect 35811 4198 35823 4374
rect 35857 4198 35869 4374
rect 35811 4186 35869 4198
rect 35929 4374 35987 4386
rect 35929 4198 35941 4374
rect 35975 4198 35987 4374
rect 40101 4262 40159 4274
rect 35929 4186 35987 4198
rect 37776 4190 37834 4202
rect 30645 4113 31045 4125
rect 30645 4079 30657 4113
rect 31033 4079 31045 4113
rect 29952 4056 30352 4068
rect 30645 4067 31045 4079
rect 29952 4022 29964 4056
rect 30340 4022 30352 4056
rect 29952 4010 30352 4022
rect 29952 3938 30352 3950
rect 29952 3904 29964 3938
rect 30340 3904 30352 3938
rect 29952 3892 30352 3904
rect 29952 3820 30352 3832
rect 29952 3786 29964 3820
rect 30340 3786 30352 3820
rect 29952 3774 30352 3786
rect 30645 3995 31045 4007
rect 30645 3961 30657 3995
rect 31033 3961 31045 3995
rect 30645 3949 31045 3961
rect 37776 4014 37788 4190
rect 37822 4014 37834 4190
rect 37776 4002 37834 4014
rect 37894 4190 37952 4202
rect 37894 4014 37906 4190
rect 37940 4014 37952 4190
rect 37894 4002 37952 4014
rect 38012 4190 38070 4202
rect 38012 4014 38024 4190
rect 38058 4014 38070 4190
rect 38012 4002 38070 4014
rect 38130 4190 38188 4202
rect 38130 4014 38142 4190
rect 38176 4014 38188 4190
rect 38130 4002 38188 4014
rect 38248 4190 38306 4202
rect 38248 4014 38260 4190
rect 38294 4014 38306 4190
rect 38248 4002 38306 4014
rect 38366 4190 38424 4202
rect 38366 4014 38378 4190
rect 38412 4014 38424 4190
rect 38366 4002 38424 4014
rect 38484 4190 38542 4202
rect 38484 4014 38496 4190
rect 38530 4014 38542 4190
rect 38484 4002 38542 4014
rect 38602 4190 38660 4202
rect 38602 4014 38614 4190
rect 38648 4014 38660 4190
rect 38602 4002 38660 4014
rect 38720 4190 38778 4202
rect 38720 4014 38732 4190
rect 38766 4014 38778 4190
rect 38720 4002 38778 4014
rect 38838 4190 38896 4202
rect 38838 4014 38850 4190
rect 38884 4014 38896 4190
rect 38838 4002 38896 4014
rect 30645 3877 31045 3889
rect 30645 3843 30657 3877
rect 31033 3843 31045 3877
rect 30645 3831 31045 3843
rect 29952 3702 30352 3714
rect 29952 3668 29964 3702
rect 30340 3668 30352 3702
rect 29952 3656 30352 3668
rect 30152 3573 30352 3585
rect 30152 3539 30164 3573
rect 30340 3539 30352 3573
rect 30152 3527 30352 3539
rect 30645 3759 31045 3771
rect 30645 3725 30657 3759
rect 31033 3725 31045 3759
rect 30645 3713 31045 3725
rect 40101 3886 40113 4262
rect 40147 3886 40159 4262
rect 40101 3874 40159 3886
rect 40219 4262 40277 4274
rect 40219 3886 40231 4262
rect 40265 3886 40277 4262
rect 40219 3874 40277 3886
rect 40337 4262 40395 4274
rect 40337 3886 40349 4262
rect 40383 3886 40395 4262
rect 40337 3874 40395 3886
rect 40455 4262 40513 4274
rect 40455 3886 40467 4262
rect 40501 3886 40513 4262
rect 40455 3874 40513 3886
rect 40573 4262 40631 4274
rect 40573 3886 40585 4262
rect 40619 3886 40631 4262
rect 40573 3874 40631 3886
rect 40691 4262 40749 4274
rect 40691 3886 40703 4262
rect 40737 3886 40749 4262
rect 40691 3874 40749 3886
rect 40809 4262 40867 4274
rect 40809 3886 40821 4262
rect 40855 3886 40867 4262
rect 40809 3874 40867 3886
rect 41243 4266 41301 4278
rect 41243 3890 41255 4266
rect 41289 3890 41301 4266
rect 41243 3878 41301 3890
rect 41361 4266 41419 4278
rect 41361 3890 41373 4266
rect 41407 3890 41419 4266
rect 41361 3878 41419 3890
rect 41479 4266 41537 4278
rect 41479 3890 41491 4266
rect 41525 3890 41537 4266
rect 41479 3878 41537 3890
rect 41597 4266 41655 4278
rect 41597 3890 41609 4266
rect 41643 3890 41655 4266
rect 41597 3878 41655 3890
rect 41715 4266 41773 4278
rect 41715 3890 41727 4266
rect 41761 3890 41773 4266
rect 41715 3878 41773 3890
rect 41833 4266 41891 4278
rect 41833 3890 41845 4266
rect 41879 3890 41891 4266
rect 41833 3878 41891 3890
rect 41951 4266 42009 4278
rect 70513 4679 70913 4691
rect 70513 4645 70525 4679
rect 70901 4645 70913 4679
rect 70513 4633 70913 4645
rect 70513 4560 70913 4572
rect 70513 4526 70525 4560
rect 70901 4526 70913 4560
rect 70513 4514 70913 4526
rect 63480 4466 63538 4478
rect 41951 3890 41963 4266
rect 41997 3890 42009 4266
rect 46652 4260 46710 4272
rect 44327 4188 44385 4200
rect 44327 4012 44339 4188
rect 44373 4012 44385 4188
rect 44327 4000 44385 4012
rect 44445 4188 44503 4200
rect 44445 4012 44457 4188
rect 44491 4012 44503 4188
rect 44445 4000 44503 4012
rect 44563 4188 44621 4200
rect 44563 4012 44575 4188
rect 44609 4012 44621 4188
rect 44563 4000 44621 4012
rect 44681 4188 44739 4200
rect 44681 4012 44693 4188
rect 44727 4012 44739 4188
rect 44681 4000 44739 4012
rect 44799 4188 44857 4200
rect 44799 4012 44811 4188
rect 44845 4012 44857 4188
rect 44799 4000 44857 4012
rect 44917 4188 44975 4200
rect 44917 4012 44929 4188
rect 44963 4012 44975 4188
rect 44917 4000 44975 4012
rect 45035 4188 45093 4200
rect 45035 4012 45047 4188
rect 45081 4012 45093 4188
rect 45035 4000 45093 4012
rect 45153 4188 45211 4200
rect 45153 4012 45165 4188
rect 45199 4012 45211 4188
rect 45153 4000 45211 4012
rect 45271 4188 45329 4200
rect 45271 4012 45283 4188
rect 45317 4012 45329 4188
rect 45271 4000 45329 4012
rect 45389 4188 45447 4200
rect 45389 4012 45401 4188
rect 45435 4012 45447 4188
rect 45389 4000 45447 4012
rect 41951 3878 42009 3890
rect 30152 3455 30352 3467
rect 30152 3421 30164 3455
rect 30340 3421 30352 3455
rect 30152 3409 30352 3421
rect 30152 3337 30352 3349
rect 30152 3303 30164 3337
rect 30340 3303 30352 3337
rect 46652 3884 46664 4260
rect 46698 3884 46710 4260
rect 46652 3872 46710 3884
rect 46770 4260 46828 4272
rect 46770 3884 46782 4260
rect 46816 3884 46828 4260
rect 46770 3872 46828 3884
rect 46888 4260 46946 4272
rect 46888 3884 46900 4260
rect 46934 3884 46946 4260
rect 46888 3872 46946 3884
rect 47006 4260 47064 4272
rect 47006 3884 47018 4260
rect 47052 3884 47064 4260
rect 47006 3872 47064 3884
rect 47124 4260 47182 4272
rect 47124 3884 47136 4260
rect 47170 3884 47182 4260
rect 47124 3872 47182 3884
rect 47242 4260 47300 4272
rect 47242 3884 47254 4260
rect 47288 3884 47300 4260
rect 47242 3872 47300 3884
rect 47360 4260 47418 4272
rect 47360 3884 47372 4260
rect 47406 3884 47418 4260
rect 47360 3872 47418 3884
rect 47794 4264 47852 4276
rect 47794 3888 47806 4264
rect 47840 3888 47852 4264
rect 47794 3876 47852 3888
rect 47912 4264 47970 4276
rect 47912 3888 47924 4264
rect 47958 3888 47970 4264
rect 47912 3876 47970 3888
rect 48030 4264 48088 4276
rect 48030 3888 48042 4264
rect 48076 3888 48088 4264
rect 48030 3876 48088 3888
rect 48148 4264 48206 4276
rect 48148 3888 48160 4264
rect 48194 3888 48206 4264
rect 48148 3876 48206 3888
rect 48266 4264 48324 4276
rect 48266 3888 48278 4264
rect 48312 3888 48324 4264
rect 48266 3876 48324 3888
rect 48384 4264 48442 4276
rect 48384 3888 48396 4264
rect 48430 3888 48442 4264
rect 48384 3876 48442 3888
rect 48502 4264 48560 4276
rect 48502 3888 48514 4264
rect 48548 3888 48560 4264
rect 53307 4261 53365 4273
rect 50982 4189 51040 4201
rect 50982 4013 50994 4189
rect 51028 4013 51040 4189
rect 50982 4001 51040 4013
rect 51100 4189 51158 4201
rect 51100 4013 51112 4189
rect 51146 4013 51158 4189
rect 51100 4001 51158 4013
rect 51218 4189 51276 4201
rect 51218 4013 51230 4189
rect 51264 4013 51276 4189
rect 51218 4001 51276 4013
rect 51336 4189 51394 4201
rect 51336 4013 51348 4189
rect 51382 4013 51394 4189
rect 51336 4001 51394 4013
rect 51454 4189 51512 4201
rect 51454 4013 51466 4189
rect 51500 4013 51512 4189
rect 51454 4001 51512 4013
rect 51572 4189 51630 4201
rect 51572 4013 51584 4189
rect 51618 4013 51630 4189
rect 51572 4001 51630 4013
rect 51690 4189 51748 4201
rect 51690 4013 51702 4189
rect 51736 4013 51748 4189
rect 51690 4001 51748 4013
rect 51808 4189 51866 4201
rect 51808 4013 51820 4189
rect 51854 4013 51866 4189
rect 51808 4001 51866 4013
rect 51926 4189 51984 4201
rect 51926 4013 51938 4189
rect 51972 4013 51984 4189
rect 51926 4001 51984 4013
rect 52044 4189 52102 4201
rect 52044 4013 52056 4189
rect 52090 4013 52102 4189
rect 52044 4001 52102 4013
rect 48502 3876 48560 3888
rect 30152 3291 30352 3303
rect 40530 3479 40588 3491
rect 40530 3303 40542 3479
rect 40576 3303 40588 3479
rect 40530 3291 40588 3303
rect 40648 3479 40706 3491
rect 40648 3303 40660 3479
rect 40694 3303 40706 3479
rect 40648 3291 40706 3303
rect 40766 3479 40824 3491
rect 40766 3303 40778 3479
rect 40812 3303 40824 3479
rect 40766 3291 40824 3303
rect 40884 3479 40942 3491
rect 40884 3303 40896 3479
rect 40930 3303 40942 3479
rect 40884 3291 40942 3303
rect 41672 3483 41730 3495
rect 41672 3307 41684 3483
rect 41718 3307 41730 3483
rect 41672 3295 41730 3307
rect 41790 3483 41848 3495
rect 41790 3307 41802 3483
rect 41836 3307 41848 3483
rect 41790 3295 41848 3307
rect 41908 3483 41966 3495
rect 41908 3307 41920 3483
rect 41954 3307 41966 3483
rect 41908 3295 41966 3307
rect 42026 3483 42084 3495
rect 42026 3307 42038 3483
rect 42072 3307 42084 3483
rect 53307 3885 53319 4261
rect 53353 3885 53365 4261
rect 53307 3873 53365 3885
rect 53425 4261 53483 4273
rect 53425 3885 53437 4261
rect 53471 3885 53483 4261
rect 53425 3873 53483 3885
rect 53543 4261 53601 4273
rect 53543 3885 53555 4261
rect 53589 3885 53601 4261
rect 53543 3873 53601 3885
rect 53661 4261 53719 4273
rect 53661 3885 53673 4261
rect 53707 3885 53719 4261
rect 53661 3873 53719 3885
rect 53779 4261 53837 4273
rect 53779 3885 53791 4261
rect 53825 3885 53837 4261
rect 53779 3873 53837 3885
rect 53897 4261 53955 4273
rect 53897 3885 53909 4261
rect 53943 3885 53955 4261
rect 53897 3873 53955 3885
rect 54015 4261 54073 4273
rect 54015 3885 54027 4261
rect 54061 3885 54073 4261
rect 54015 3873 54073 3885
rect 54449 4265 54507 4277
rect 54449 3889 54461 4265
rect 54495 3889 54507 4265
rect 54449 3877 54507 3889
rect 54567 4265 54625 4277
rect 54567 3889 54579 4265
rect 54613 3889 54625 4265
rect 54567 3877 54625 3889
rect 54685 4265 54743 4277
rect 54685 3889 54697 4265
rect 54731 3889 54743 4265
rect 54685 3877 54743 3889
rect 54803 4265 54861 4277
rect 54803 3889 54815 4265
rect 54849 3889 54861 4265
rect 54803 3877 54861 3889
rect 54921 4265 54979 4277
rect 54921 3889 54933 4265
rect 54967 3889 54979 4265
rect 54921 3877 54979 3889
rect 55039 4265 55097 4277
rect 55039 3889 55051 4265
rect 55085 3889 55097 4265
rect 55039 3877 55097 3889
rect 55157 4265 55215 4277
rect 63480 4290 63492 4466
rect 63526 4290 63538 4466
rect 63480 4278 63538 4290
rect 63598 4466 63656 4478
rect 63598 4290 63610 4466
rect 63644 4290 63656 4466
rect 63598 4278 63656 4290
rect 63716 4466 63774 4478
rect 63716 4290 63728 4466
rect 63762 4290 63774 4466
rect 63716 4278 63774 4290
rect 63834 4466 63892 4478
rect 63834 4290 63846 4466
rect 63880 4290 63892 4466
rect 63834 4278 63892 4290
rect 63952 4466 64010 4478
rect 63952 4290 63964 4466
rect 63998 4290 64010 4466
rect 63952 4278 64010 4290
rect 64070 4466 64128 4478
rect 64070 4290 64082 4466
rect 64116 4290 64128 4466
rect 64070 4278 64128 4290
rect 64188 4466 64246 4478
rect 64188 4290 64200 4466
rect 64234 4290 64246 4466
rect 64188 4278 64246 4290
rect 64306 4466 64364 4478
rect 64306 4290 64318 4466
rect 64352 4290 64364 4466
rect 64306 4278 64364 4290
rect 64424 4466 64482 4478
rect 64424 4290 64436 4466
rect 64470 4290 64482 4466
rect 64424 4278 64482 4290
rect 64542 4466 64600 4478
rect 64542 4290 64554 4466
rect 64588 4290 64600 4466
rect 64542 4278 64600 4290
rect 70513 4442 70913 4454
rect 70513 4408 70525 4442
rect 70901 4408 70913 4442
rect 70513 4396 70913 4408
rect 70513 4324 70913 4336
rect 70513 4290 70525 4324
rect 70901 4290 70913 4324
rect 70513 4278 70913 4290
rect 55157 3889 55169 4265
rect 55203 3889 55215 4265
rect 59929 4262 59987 4274
rect 57604 4190 57662 4202
rect 57604 4014 57616 4190
rect 57650 4014 57662 4190
rect 57604 4002 57662 4014
rect 57722 4190 57780 4202
rect 57722 4014 57734 4190
rect 57768 4014 57780 4190
rect 57722 4002 57780 4014
rect 57840 4190 57898 4202
rect 57840 4014 57852 4190
rect 57886 4014 57898 4190
rect 57840 4002 57898 4014
rect 57958 4190 58016 4202
rect 57958 4014 57970 4190
rect 58004 4014 58016 4190
rect 57958 4002 58016 4014
rect 58076 4190 58134 4202
rect 58076 4014 58088 4190
rect 58122 4014 58134 4190
rect 58076 4002 58134 4014
rect 58194 4190 58252 4202
rect 58194 4014 58206 4190
rect 58240 4014 58252 4190
rect 58194 4002 58252 4014
rect 58312 4190 58370 4202
rect 58312 4014 58324 4190
rect 58358 4014 58370 4190
rect 58312 4002 58370 4014
rect 58430 4190 58488 4202
rect 58430 4014 58442 4190
rect 58476 4014 58488 4190
rect 58430 4002 58488 4014
rect 58548 4190 58606 4202
rect 58548 4014 58560 4190
rect 58594 4014 58606 4190
rect 58548 4002 58606 4014
rect 58666 4190 58724 4202
rect 58666 4014 58678 4190
rect 58712 4014 58724 4190
rect 58666 4002 58724 4014
rect 55157 3877 55215 3889
rect 42026 3295 42084 3307
rect 30152 3219 30352 3231
rect 30152 3185 30164 3219
rect 30340 3185 30352 3219
rect 47081 3477 47139 3489
rect 47081 3301 47093 3477
rect 47127 3301 47139 3477
rect 47081 3289 47139 3301
rect 47199 3477 47257 3489
rect 47199 3301 47211 3477
rect 47245 3301 47257 3477
rect 47199 3289 47257 3301
rect 47317 3477 47375 3489
rect 47317 3301 47329 3477
rect 47363 3301 47375 3477
rect 47317 3289 47375 3301
rect 47435 3477 47493 3489
rect 47435 3301 47447 3477
rect 47481 3301 47493 3477
rect 47435 3289 47493 3301
rect 48223 3481 48281 3493
rect 48223 3305 48235 3481
rect 48269 3305 48281 3481
rect 48223 3293 48281 3305
rect 48341 3481 48399 3493
rect 48341 3305 48353 3481
rect 48387 3305 48399 3481
rect 48341 3293 48399 3305
rect 48459 3481 48517 3493
rect 48459 3305 48471 3481
rect 48505 3305 48517 3481
rect 48459 3293 48517 3305
rect 48577 3481 48635 3493
rect 48577 3305 48589 3481
rect 48623 3305 48635 3481
rect 59929 3886 59941 4262
rect 59975 3886 59987 4262
rect 59929 3874 59987 3886
rect 60047 4262 60105 4274
rect 60047 3886 60059 4262
rect 60093 3886 60105 4262
rect 60047 3874 60105 3886
rect 60165 4262 60223 4274
rect 60165 3886 60177 4262
rect 60211 3886 60223 4262
rect 60165 3874 60223 3886
rect 60283 4262 60341 4274
rect 60283 3886 60295 4262
rect 60329 3886 60341 4262
rect 60283 3874 60341 3886
rect 60401 4262 60459 4274
rect 60401 3886 60413 4262
rect 60447 3886 60459 4262
rect 60401 3874 60459 3886
rect 60519 4262 60577 4274
rect 60519 3886 60531 4262
rect 60565 3886 60577 4262
rect 60519 3874 60577 3886
rect 60637 4262 60695 4274
rect 60637 3886 60649 4262
rect 60683 3886 60695 4262
rect 60637 3874 60695 3886
rect 61071 4266 61129 4278
rect 61071 3890 61083 4266
rect 61117 3890 61129 4266
rect 61071 3878 61129 3890
rect 61189 4266 61247 4278
rect 61189 3890 61201 4266
rect 61235 3890 61247 4266
rect 61189 3878 61247 3890
rect 61307 4266 61365 4278
rect 61307 3890 61319 4266
rect 61353 3890 61365 4266
rect 61307 3878 61365 3890
rect 61425 4266 61483 4278
rect 61425 3890 61437 4266
rect 61471 3890 61483 4266
rect 61425 3878 61483 3890
rect 61543 4266 61601 4278
rect 61543 3890 61555 4266
rect 61589 3890 61601 4266
rect 61543 3878 61601 3890
rect 61661 4266 61719 4278
rect 61661 3890 61673 4266
rect 61707 3890 61719 4266
rect 61661 3878 61719 3890
rect 61779 4266 61837 4278
rect 61779 3890 61791 4266
rect 61825 3890 61837 4266
rect 65708 4199 65766 4211
rect 61779 3878 61837 3890
rect 48577 3293 48635 3305
rect 53736 3478 53794 3490
rect 53736 3302 53748 3478
rect 53782 3302 53794 3478
rect 53736 3290 53794 3302
rect 53854 3478 53912 3490
rect 53854 3302 53866 3478
rect 53900 3302 53912 3478
rect 53854 3290 53912 3302
rect 53972 3478 54030 3490
rect 53972 3302 53984 3478
rect 54018 3302 54030 3478
rect 53972 3290 54030 3302
rect 54090 3478 54148 3490
rect 54090 3302 54102 3478
rect 54136 3302 54148 3478
rect 54090 3290 54148 3302
rect 54878 3482 54936 3494
rect 54878 3306 54890 3482
rect 54924 3306 54936 3482
rect 54878 3294 54936 3306
rect 54996 3482 55054 3494
rect 54996 3306 55008 3482
rect 55042 3306 55054 3482
rect 54996 3294 55054 3306
rect 55114 3482 55172 3494
rect 55114 3306 55126 3482
rect 55160 3306 55172 3482
rect 55114 3294 55172 3306
rect 55232 3482 55290 3494
rect 55232 3306 55244 3482
rect 55278 3306 55290 3482
rect 65224 3999 65282 4011
rect 65224 3823 65236 3999
rect 65270 3823 65282 3999
rect 65224 3811 65282 3823
rect 65342 3999 65400 4011
rect 65342 3823 65354 3999
rect 65388 3823 65400 3999
rect 65342 3811 65400 3823
rect 65460 3999 65518 4011
rect 65460 3823 65472 3999
rect 65506 3823 65518 3999
rect 65460 3811 65518 3823
rect 65578 3999 65636 4011
rect 65578 3823 65590 3999
rect 65624 3823 65636 3999
rect 65578 3811 65636 3823
rect 65708 3823 65720 4199
rect 65754 3823 65766 4199
rect 65708 3811 65766 3823
rect 65826 4199 65884 4211
rect 65826 3823 65838 4199
rect 65872 3823 65884 4199
rect 65826 3811 65884 3823
rect 65944 4199 66002 4211
rect 65944 3823 65956 4199
rect 65990 3823 66002 4199
rect 65944 3811 66002 3823
rect 66062 4199 66120 4211
rect 66062 3823 66074 4199
rect 66108 3823 66120 4199
rect 66062 3811 66120 3823
rect 66180 4199 66238 4211
rect 66180 3823 66192 4199
rect 66226 3823 66238 4199
rect 66180 3811 66238 3823
rect 66298 4199 66356 4211
rect 66298 3823 66310 4199
rect 66344 3823 66356 4199
rect 66298 3811 66356 3823
rect 66416 4199 66474 4211
rect 66416 3823 66428 4199
rect 66462 3823 66474 4199
rect 70513 4206 70913 4218
rect 70513 4172 70525 4206
rect 70901 4172 70913 4206
rect 70513 4160 70913 4172
rect 70713 4087 70913 4099
rect 66416 3811 66474 3823
rect 66545 3999 66603 4011
rect 66545 3823 66557 3999
rect 66591 3823 66603 3999
rect 66545 3811 66603 3823
rect 66663 3999 66721 4011
rect 66663 3823 66675 3999
rect 66709 3823 66721 3999
rect 66663 3811 66721 3823
rect 66781 3999 66839 4011
rect 66781 3823 66793 3999
rect 66827 3823 66839 3999
rect 66781 3811 66839 3823
rect 66899 3999 66957 4011
rect 70713 4053 70725 4087
rect 70901 4053 70913 4087
rect 70713 4041 70913 4053
rect 66899 3823 66911 3999
rect 66945 3823 66957 3999
rect 66899 3811 66957 3823
rect 67017 3996 67075 4008
rect 67017 3820 67029 3996
rect 67063 3820 67075 3996
rect 67017 3808 67075 3820
rect 67135 3996 67193 4008
rect 67135 3820 67147 3996
rect 67181 3820 67193 3996
rect 67135 3808 67193 3820
rect 67253 3996 67311 4008
rect 67253 3820 67265 3996
rect 67299 3820 67311 3996
rect 67253 3808 67311 3820
rect 67371 3996 67429 4008
rect 67371 3820 67383 3996
rect 67417 3820 67429 3996
rect 67371 3808 67429 3820
rect 67489 3996 67547 4008
rect 67489 3820 67501 3996
rect 67535 3820 67547 3996
rect 67489 3808 67547 3820
rect 67607 3996 67665 4008
rect 67607 3820 67619 3996
rect 67653 3820 67665 3996
rect 67607 3808 67665 3820
rect 67725 3996 67783 4008
rect 67725 3820 67737 3996
rect 67771 3820 67783 3996
rect 67725 3808 67783 3820
rect 67843 3996 67901 4008
rect 67843 3820 67855 3996
rect 67889 3820 67901 3996
rect 67843 3808 67901 3820
rect 67961 3996 68019 4008
rect 67961 3820 67973 3996
rect 68007 3820 68019 3996
rect 67961 3808 68019 3820
rect 68079 3996 68137 4008
rect 68079 3820 68091 3996
rect 68125 3820 68137 3996
rect 68079 3808 68137 3820
rect 70713 3969 70913 3981
rect 70713 3935 70725 3969
rect 70901 3935 70913 3969
rect 70713 3923 70913 3935
rect 55232 3294 55290 3306
rect 60358 3479 60416 3491
rect 60358 3303 60370 3479
rect 60404 3303 60416 3479
rect 60358 3291 60416 3303
rect 60476 3479 60534 3491
rect 60476 3303 60488 3479
rect 60522 3303 60534 3479
rect 60476 3291 60534 3303
rect 60594 3479 60652 3491
rect 60594 3303 60606 3479
rect 60640 3303 60652 3479
rect 60594 3291 60652 3303
rect 60712 3479 60770 3491
rect 60712 3303 60724 3479
rect 60758 3303 60770 3479
rect 60712 3291 60770 3303
rect 61500 3483 61558 3495
rect 61500 3307 61512 3483
rect 61546 3307 61558 3483
rect 61500 3295 61558 3307
rect 61618 3483 61676 3495
rect 61618 3307 61630 3483
rect 61664 3307 61676 3483
rect 61618 3295 61676 3307
rect 61736 3483 61794 3495
rect 61736 3307 61748 3483
rect 61782 3307 61794 3483
rect 61736 3295 61794 3307
rect 61854 3483 61912 3495
rect 61854 3307 61866 3483
rect 61900 3307 61912 3483
rect 65651 3506 65709 3518
rect 61854 3295 61912 3307
rect 30152 3173 30352 3185
rect 30150 2826 30350 2838
rect 30150 2792 30162 2826
rect 30338 2792 30350 2826
rect 30150 2780 30350 2792
rect 30150 2708 30350 2720
rect 30150 2674 30162 2708
rect 30338 2674 30350 2708
rect 30150 2662 30350 2674
rect 65651 3130 65663 3506
rect 65697 3130 65709 3506
rect 65651 3118 65709 3130
rect 65769 3506 65827 3518
rect 65769 3130 65781 3506
rect 65815 3130 65827 3506
rect 65769 3118 65827 3130
rect 65887 3506 65945 3518
rect 65887 3130 65899 3506
rect 65933 3130 65945 3506
rect 65887 3118 65945 3130
rect 66005 3506 66063 3518
rect 66005 3130 66017 3506
rect 66051 3130 66063 3506
rect 66005 3118 66063 3130
rect 66123 3506 66181 3518
rect 66123 3130 66135 3506
rect 66169 3130 66181 3506
rect 66123 3118 66181 3130
rect 66241 3506 66299 3518
rect 66241 3130 66253 3506
rect 66287 3130 66299 3506
rect 66241 3118 66299 3130
rect 66359 3506 66417 3518
rect 66359 3130 66371 3506
rect 66405 3130 66417 3506
rect 66359 3118 66417 3130
rect 70713 3851 70913 3863
rect 70713 3817 70725 3851
rect 70901 3817 70913 3851
rect 70713 3805 70913 3817
rect 70713 3733 70913 3745
rect 70713 3699 70725 3733
rect 70901 3699 70913 3733
rect 70713 3687 70913 3699
rect 70709 3163 70909 3175
rect 70709 3129 70721 3163
rect 70897 3129 70909 3163
rect 70709 3117 70909 3129
rect 70709 3045 70909 3057
rect 70709 3011 70721 3045
rect 70897 3011 70909 3045
rect 70709 2999 70909 3011
rect 70709 2927 70909 2939
rect 70709 2893 70721 2927
rect 70897 2893 70909 2927
rect 70709 2881 70909 2893
rect 70709 2809 70909 2821
rect 30150 2590 30350 2602
rect 30150 2556 30162 2590
rect 30338 2556 30350 2590
rect 30150 2544 30350 2556
rect 37790 2540 37848 2552
rect 30150 2472 30350 2484
rect 30150 2438 30162 2472
rect 30338 2438 30350 2472
rect 30150 2426 30350 2438
rect 29950 2342 30350 2354
rect 29950 2308 29962 2342
rect 30338 2308 30350 2342
rect 29950 2296 30350 2308
rect 30643 2399 31043 2411
rect 30643 2365 30655 2399
rect 31031 2365 31043 2399
rect 30643 2353 31043 2365
rect 37790 2364 37802 2540
rect 37836 2364 37848 2540
rect 37790 2352 37848 2364
rect 37908 2540 37966 2552
rect 37908 2364 37920 2540
rect 37954 2364 37966 2540
rect 37908 2352 37966 2364
rect 38026 2540 38084 2552
rect 38026 2364 38038 2540
rect 38072 2364 38084 2540
rect 38026 2352 38084 2364
rect 38144 2540 38202 2552
rect 38144 2364 38156 2540
rect 38190 2364 38202 2540
rect 38144 2352 38202 2364
rect 38262 2540 38320 2552
rect 38262 2364 38274 2540
rect 38308 2364 38320 2540
rect 38262 2352 38320 2364
rect 38380 2540 38438 2552
rect 38380 2364 38392 2540
rect 38426 2364 38438 2540
rect 38380 2352 38438 2364
rect 38498 2540 38556 2552
rect 38498 2364 38510 2540
rect 38544 2364 38556 2540
rect 38498 2352 38556 2364
rect 38616 2540 38674 2552
rect 38616 2364 38628 2540
rect 38662 2364 38674 2540
rect 38616 2352 38674 2364
rect 38734 2540 38792 2552
rect 38734 2364 38746 2540
rect 38780 2364 38792 2540
rect 38734 2352 38792 2364
rect 38852 2540 38910 2552
rect 38852 2364 38864 2540
rect 38898 2364 38910 2540
rect 44341 2538 44399 2550
rect 38852 2352 38910 2364
rect 44341 2362 44353 2538
rect 44387 2362 44399 2538
rect 689 2128 747 2140
rect 689 1940 701 2128
rect 248 1928 306 1940
rect 248 1752 260 1928
rect 294 1752 306 1928
rect 248 1740 306 1752
rect 366 1928 424 1940
rect 366 1752 378 1928
rect 412 1752 424 1928
rect 366 1740 424 1752
rect 484 1928 542 1940
rect 484 1752 496 1928
rect 530 1752 542 1928
rect 484 1740 542 1752
rect 602 1928 701 1940
rect 602 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 747 2128
rect 602 1740 747 1752
rect 807 2128 865 2140
rect 807 1752 819 2128
rect 853 1752 865 2128
rect 807 1740 865 1752
rect 925 2128 983 2140
rect 925 1752 937 2128
rect 971 1752 983 2128
rect 925 1740 983 1752
rect 1043 2128 1101 2140
rect 1043 1752 1055 2128
rect 1089 1752 1101 2128
rect 1043 1740 1101 1752
rect 1156 2128 1214 2140
rect 1156 1752 1168 2128
rect 1202 1752 1214 2128
rect 1156 1740 1214 1752
rect 1274 2128 1332 2140
rect 1274 1752 1286 2128
rect 1320 1752 1332 2128
rect 1274 1740 1332 1752
rect 1392 2128 1450 2140
rect 1392 1752 1404 2128
rect 1438 1752 1450 2128
rect 1392 1740 1450 1752
rect 1510 2128 1568 2140
rect 1510 1752 1522 2128
rect 1556 1752 1568 2128
rect 1510 1740 1568 1752
rect 1628 2128 1686 2140
rect 1628 1752 1640 2128
rect 1674 1752 1686 2128
rect 1628 1740 1686 1752
rect 1746 2128 1804 2140
rect 1746 1752 1758 2128
rect 1792 1752 1804 2128
rect 1746 1740 1804 1752
rect 1864 2128 1922 2140
rect 1864 1752 1876 2128
rect 1910 1752 1922 2128
rect 1864 1740 1922 1752
rect 1983 2128 2041 2140
rect 1983 1752 1995 2128
rect 2029 1752 2041 2128
rect 1983 1740 2041 1752
rect 2101 2128 2159 2140
rect 2101 1752 2113 2128
rect 2147 1752 2159 2128
rect 2101 1740 2159 1752
rect 2219 2128 2277 2140
rect 2219 1752 2231 2128
rect 2265 1752 2277 2128
rect 2219 1740 2277 1752
rect 2337 2128 2395 2140
rect 2337 1752 2349 2128
rect 2383 1752 2395 2128
rect 3833 2128 3891 2140
rect 3833 1940 3845 2128
rect 2337 1740 2395 1752
rect 2456 1928 2514 1940
rect 2456 1752 2468 1928
rect 2502 1752 2514 1928
rect 2456 1740 2514 1752
rect 2574 1928 2632 1940
rect 2574 1752 2586 1928
rect 2620 1752 2632 1928
rect 2574 1740 2632 1752
rect 2692 1928 2750 1940
rect 2692 1752 2704 1928
rect 2738 1752 2750 1928
rect 2692 1740 2750 1752
rect 2810 1928 2868 1940
rect 2810 1752 2822 1928
rect 2856 1752 2868 1928
rect 2810 1740 2868 1752
rect 3392 1928 3450 1940
rect 3392 1752 3404 1928
rect 3438 1752 3450 1928
rect 3392 1740 3450 1752
rect 3510 1928 3568 1940
rect 3510 1752 3522 1928
rect 3556 1752 3568 1928
rect 3510 1740 3568 1752
rect 3628 1928 3686 1940
rect 3628 1752 3640 1928
rect 3674 1752 3686 1928
rect 3628 1740 3686 1752
rect 3746 1928 3845 1940
rect 3746 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3891 2128
rect 3746 1740 3891 1752
rect 3951 2128 4009 2140
rect 3951 1752 3963 2128
rect 3997 1752 4009 2128
rect 3951 1740 4009 1752
rect 4069 2128 4127 2140
rect 4069 1752 4081 2128
rect 4115 1752 4127 2128
rect 4069 1740 4127 1752
rect 4187 2128 4245 2140
rect 4187 1752 4199 2128
rect 4233 1752 4245 2128
rect 4187 1740 4245 1752
rect 4300 2128 4358 2140
rect 4300 1752 4312 2128
rect 4346 1752 4358 2128
rect 4300 1740 4358 1752
rect 4418 2128 4476 2140
rect 4418 1752 4430 2128
rect 4464 1752 4476 2128
rect 4418 1740 4476 1752
rect 4536 2128 4594 2140
rect 4536 1752 4548 2128
rect 4582 1752 4594 2128
rect 4536 1740 4594 1752
rect 4654 2128 4712 2140
rect 4654 1752 4666 2128
rect 4700 1752 4712 2128
rect 4654 1740 4712 1752
rect 4772 2128 4830 2140
rect 4772 1752 4784 2128
rect 4818 1752 4830 2128
rect 4772 1740 4830 1752
rect 4890 2128 4948 2140
rect 4890 1752 4902 2128
rect 4936 1752 4948 2128
rect 4890 1740 4948 1752
rect 5008 2128 5066 2140
rect 5008 1752 5020 2128
rect 5054 1752 5066 2128
rect 5008 1740 5066 1752
rect 5127 2128 5185 2140
rect 5127 1752 5139 2128
rect 5173 1752 5185 2128
rect 5127 1740 5185 1752
rect 5245 2128 5303 2140
rect 5245 1752 5257 2128
rect 5291 1752 5303 2128
rect 5245 1740 5303 1752
rect 5363 2128 5421 2140
rect 5363 1752 5375 2128
rect 5409 1752 5421 2128
rect 5363 1740 5421 1752
rect 5481 2128 5539 2140
rect 5481 1752 5493 2128
rect 5527 1752 5539 2128
rect 6965 2132 7023 2144
rect 6965 1944 6977 2132
rect 5481 1740 5539 1752
rect 5600 1928 5658 1940
rect 5600 1752 5612 1928
rect 5646 1752 5658 1928
rect 5600 1740 5658 1752
rect 5718 1928 5776 1940
rect 5718 1752 5730 1928
rect 5764 1752 5776 1928
rect 5718 1740 5776 1752
rect 5836 1928 5894 1940
rect 5836 1752 5848 1928
rect 5882 1752 5894 1928
rect 5836 1740 5894 1752
rect 5954 1928 6012 1940
rect 5954 1752 5966 1928
rect 6000 1752 6012 1928
rect 5954 1740 6012 1752
rect 6524 1932 6582 1944
rect 6524 1756 6536 1932
rect 6570 1756 6582 1932
rect 6524 1744 6582 1756
rect 6642 1932 6700 1944
rect 6642 1756 6654 1932
rect 6688 1756 6700 1932
rect 6642 1744 6700 1756
rect 6760 1932 6818 1944
rect 6760 1756 6772 1932
rect 6806 1756 6818 1932
rect 6760 1744 6818 1756
rect 6878 1932 6977 1944
rect 6878 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7023 2132
rect 6878 1744 7023 1756
rect 7083 2132 7141 2144
rect 7083 1756 7095 2132
rect 7129 1756 7141 2132
rect 7083 1744 7141 1756
rect 7201 2132 7259 2144
rect 7201 1756 7213 2132
rect 7247 1756 7259 2132
rect 7201 1744 7259 1756
rect 7319 2132 7377 2144
rect 7319 1756 7331 2132
rect 7365 1756 7377 2132
rect 7319 1744 7377 1756
rect 7432 2132 7490 2144
rect 7432 1756 7444 2132
rect 7478 1756 7490 2132
rect 7432 1744 7490 1756
rect 7550 2132 7608 2144
rect 7550 1756 7562 2132
rect 7596 1756 7608 2132
rect 7550 1744 7608 1756
rect 7668 2132 7726 2144
rect 7668 1756 7680 2132
rect 7714 1756 7726 2132
rect 7668 1744 7726 1756
rect 7786 2132 7844 2144
rect 7786 1756 7798 2132
rect 7832 1756 7844 2132
rect 7786 1744 7844 1756
rect 7904 2132 7962 2144
rect 7904 1756 7916 2132
rect 7950 1756 7962 2132
rect 7904 1744 7962 1756
rect 8022 2132 8080 2144
rect 8022 1756 8034 2132
rect 8068 1756 8080 2132
rect 8022 1744 8080 1756
rect 8140 2132 8198 2144
rect 8140 1756 8152 2132
rect 8186 1756 8198 2132
rect 8140 1744 8198 1756
rect 8259 2132 8317 2144
rect 8259 1756 8271 2132
rect 8305 1756 8317 2132
rect 8259 1744 8317 1756
rect 8377 2132 8435 2144
rect 8377 1756 8389 2132
rect 8423 1756 8435 2132
rect 8377 1744 8435 1756
rect 8495 2132 8553 2144
rect 8495 1756 8507 2132
rect 8541 1756 8553 2132
rect 8495 1744 8553 1756
rect 8613 2132 8671 2144
rect 8613 1756 8625 2132
rect 8659 1756 8671 2132
rect 10109 2132 10167 2144
rect 10109 1944 10121 2132
rect 8613 1744 8671 1756
rect 8732 1932 8790 1944
rect 8732 1756 8744 1932
rect 8778 1756 8790 1932
rect 8732 1744 8790 1756
rect 8850 1932 8908 1944
rect 8850 1756 8862 1932
rect 8896 1756 8908 1932
rect 8850 1744 8908 1756
rect 8968 1932 9026 1944
rect 8968 1756 8980 1932
rect 9014 1756 9026 1932
rect 8968 1744 9026 1756
rect 9086 1932 9144 1944
rect 9086 1756 9098 1932
rect 9132 1756 9144 1932
rect 9086 1744 9144 1756
rect 9668 1932 9726 1944
rect 9668 1756 9680 1932
rect 9714 1756 9726 1932
rect 9668 1744 9726 1756
rect 9786 1932 9844 1944
rect 9786 1756 9798 1932
rect 9832 1756 9844 1932
rect 9786 1744 9844 1756
rect 9904 1932 9962 1944
rect 9904 1756 9916 1932
rect 9950 1756 9962 1932
rect 9904 1744 9962 1756
rect 10022 1932 10121 1944
rect 10022 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10167 2132
rect 10022 1744 10167 1756
rect 10227 2132 10285 2144
rect 10227 1756 10239 2132
rect 10273 1756 10285 2132
rect 10227 1744 10285 1756
rect 10345 2132 10403 2144
rect 10345 1756 10357 2132
rect 10391 1756 10403 2132
rect 10345 1744 10403 1756
rect 10463 2132 10521 2144
rect 10463 1756 10475 2132
rect 10509 1756 10521 2132
rect 10463 1744 10521 1756
rect 10576 2132 10634 2144
rect 10576 1756 10588 2132
rect 10622 1756 10634 2132
rect 10576 1744 10634 1756
rect 10694 2132 10752 2144
rect 10694 1756 10706 2132
rect 10740 1756 10752 2132
rect 10694 1744 10752 1756
rect 10812 2132 10870 2144
rect 10812 1756 10824 2132
rect 10858 1756 10870 2132
rect 10812 1744 10870 1756
rect 10930 2132 10988 2144
rect 10930 1756 10942 2132
rect 10976 1756 10988 2132
rect 10930 1744 10988 1756
rect 11048 2132 11106 2144
rect 11048 1756 11060 2132
rect 11094 1756 11106 2132
rect 11048 1744 11106 1756
rect 11166 2132 11224 2144
rect 11166 1756 11178 2132
rect 11212 1756 11224 2132
rect 11166 1744 11224 1756
rect 11284 2132 11342 2144
rect 11284 1756 11296 2132
rect 11330 1756 11342 2132
rect 11284 1744 11342 1756
rect 11403 2132 11461 2144
rect 11403 1756 11415 2132
rect 11449 1756 11461 2132
rect 11403 1744 11461 1756
rect 11521 2132 11579 2144
rect 11521 1756 11533 2132
rect 11567 1756 11579 2132
rect 11521 1744 11579 1756
rect 11639 2132 11697 2144
rect 11639 1756 11651 2132
rect 11685 1756 11697 2132
rect 11639 1744 11697 1756
rect 11757 2132 11815 2144
rect 29950 2224 30350 2236
rect 29950 2190 29962 2224
rect 30338 2190 30350 2224
rect 29950 2178 30350 2190
rect 30643 2281 31043 2293
rect 30643 2247 30655 2281
rect 31031 2247 31043 2281
rect 30643 2235 31043 2247
rect 11757 1756 11769 2132
rect 11803 1756 11815 2132
rect 13311 2128 13369 2140
rect 11757 1744 11815 1756
rect 11876 1932 11934 1944
rect 11876 1756 11888 1932
rect 11922 1756 11934 1932
rect 11876 1744 11934 1756
rect 11994 1932 12052 1944
rect 11994 1756 12006 1932
rect 12040 1756 12052 1932
rect 11994 1744 12052 1756
rect 12112 1932 12170 1944
rect 12112 1756 12124 1932
rect 12158 1756 12170 1932
rect 12112 1744 12170 1756
rect 12230 1932 12288 1944
rect 13311 1940 13323 2128
rect 12230 1756 12242 1932
rect 12276 1756 12288 1932
rect 12230 1744 12288 1756
rect 12870 1928 12928 1940
rect 12870 1752 12882 1928
rect 12916 1752 12928 1928
rect 12870 1740 12928 1752
rect 12988 1928 13046 1940
rect 12988 1752 13000 1928
rect 13034 1752 13046 1928
rect 12988 1740 13046 1752
rect 13106 1928 13164 1940
rect 13106 1752 13118 1928
rect 13152 1752 13164 1928
rect 13106 1740 13164 1752
rect 13224 1928 13323 1940
rect 13224 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13369 2128
rect 13224 1740 13369 1752
rect 13429 2128 13487 2140
rect 13429 1752 13441 2128
rect 13475 1752 13487 2128
rect 13429 1740 13487 1752
rect 13547 2128 13605 2140
rect 13547 1752 13559 2128
rect 13593 1752 13605 2128
rect 13547 1740 13605 1752
rect 13665 2128 13723 2140
rect 13665 1752 13677 2128
rect 13711 1752 13723 2128
rect 13665 1740 13723 1752
rect 13778 2128 13836 2140
rect 13778 1752 13790 2128
rect 13824 1752 13836 2128
rect 13778 1740 13836 1752
rect 13896 2128 13954 2140
rect 13896 1752 13908 2128
rect 13942 1752 13954 2128
rect 13896 1740 13954 1752
rect 14014 2128 14072 2140
rect 14014 1752 14026 2128
rect 14060 1752 14072 2128
rect 14014 1740 14072 1752
rect 14132 2128 14190 2140
rect 14132 1752 14144 2128
rect 14178 1752 14190 2128
rect 14132 1740 14190 1752
rect 14250 2128 14308 2140
rect 14250 1752 14262 2128
rect 14296 1752 14308 2128
rect 14250 1740 14308 1752
rect 14368 2128 14426 2140
rect 14368 1752 14380 2128
rect 14414 1752 14426 2128
rect 14368 1740 14426 1752
rect 14486 2128 14544 2140
rect 14486 1752 14498 2128
rect 14532 1752 14544 2128
rect 14486 1740 14544 1752
rect 14605 2128 14663 2140
rect 14605 1752 14617 2128
rect 14651 1752 14663 2128
rect 14605 1740 14663 1752
rect 14723 2128 14781 2140
rect 14723 1752 14735 2128
rect 14769 1752 14781 2128
rect 14723 1740 14781 1752
rect 14841 2128 14899 2140
rect 14841 1752 14853 2128
rect 14887 1752 14899 2128
rect 14841 1740 14899 1752
rect 14959 2128 15017 2140
rect 14959 1752 14971 2128
rect 15005 1752 15017 2128
rect 16455 2128 16513 2140
rect 16455 1940 16467 2128
rect 14959 1740 15017 1752
rect 15078 1928 15136 1940
rect 15078 1752 15090 1928
rect 15124 1752 15136 1928
rect 15078 1740 15136 1752
rect 15196 1928 15254 1940
rect 15196 1752 15208 1928
rect 15242 1752 15254 1928
rect 15196 1740 15254 1752
rect 15314 1928 15372 1940
rect 15314 1752 15326 1928
rect 15360 1752 15372 1928
rect 15314 1740 15372 1752
rect 15432 1928 15490 1940
rect 15432 1752 15444 1928
rect 15478 1752 15490 1928
rect 15432 1740 15490 1752
rect 16014 1928 16072 1940
rect 16014 1752 16026 1928
rect 16060 1752 16072 1928
rect 16014 1740 16072 1752
rect 16132 1928 16190 1940
rect 16132 1752 16144 1928
rect 16178 1752 16190 1928
rect 16132 1740 16190 1752
rect 16250 1928 16308 1940
rect 16250 1752 16262 1928
rect 16296 1752 16308 1928
rect 16250 1740 16308 1752
rect 16368 1928 16467 1940
rect 16368 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16513 2128
rect 16368 1740 16513 1752
rect 16573 2128 16631 2140
rect 16573 1752 16585 2128
rect 16619 1752 16631 2128
rect 16573 1740 16631 1752
rect 16691 2128 16749 2140
rect 16691 1752 16703 2128
rect 16737 1752 16749 2128
rect 16691 1740 16749 1752
rect 16809 2128 16867 2140
rect 16809 1752 16821 2128
rect 16855 1752 16867 2128
rect 16809 1740 16867 1752
rect 16922 2128 16980 2140
rect 16922 1752 16934 2128
rect 16968 1752 16980 2128
rect 16922 1740 16980 1752
rect 17040 2128 17098 2140
rect 17040 1752 17052 2128
rect 17086 1752 17098 2128
rect 17040 1740 17098 1752
rect 17158 2128 17216 2140
rect 17158 1752 17170 2128
rect 17204 1752 17216 2128
rect 17158 1740 17216 1752
rect 17276 2128 17334 2140
rect 17276 1752 17288 2128
rect 17322 1752 17334 2128
rect 17276 1740 17334 1752
rect 17394 2128 17452 2140
rect 17394 1752 17406 2128
rect 17440 1752 17452 2128
rect 17394 1740 17452 1752
rect 17512 2128 17570 2140
rect 17512 1752 17524 2128
rect 17558 1752 17570 2128
rect 17512 1740 17570 1752
rect 17630 2128 17688 2140
rect 17630 1752 17642 2128
rect 17676 1752 17688 2128
rect 17630 1740 17688 1752
rect 17749 2128 17807 2140
rect 17749 1752 17761 2128
rect 17795 1752 17807 2128
rect 17749 1740 17807 1752
rect 17867 2128 17925 2140
rect 17867 1752 17879 2128
rect 17913 1752 17925 2128
rect 17867 1740 17925 1752
rect 17985 2128 18043 2140
rect 17985 1752 17997 2128
rect 18031 1752 18043 2128
rect 17985 1740 18043 1752
rect 18103 2128 18161 2140
rect 18103 1752 18115 2128
rect 18149 1752 18161 2128
rect 19587 2132 19645 2144
rect 19587 1944 19599 2132
rect 18103 1740 18161 1752
rect 18222 1928 18280 1940
rect 18222 1752 18234 1928
rect 18268 1752 18280 1928
rect 18222 1740 18280 1752
rect 18340 1928 18398 1940
rect 18340 1752 18352 1928
rect 18386 1752 18398 1928
rect 18340 1740 18398 1752
rect 18458 1928 18516 1940
rect 18458 1752 18470 1928
rect 18504 1752 18516 1928
rect 18458 1740 18516 1752
rect 18576 1928 18634 1940
rect 18576 1752 18588 1928
rect 18622 1752 18634 1928
rect 18576 1740 18634 1752
rect 19146 1932 19204 1944
rect 19146 1756 19158 1932
rect 19192 1756 19204 1932
rect 19146 1744 19204 1756
rect 19264 1932 19322 1944
rect 19264 1756 19276 1932
rect 19310 1756 19322 1932
rect 19264 1744 19322 1756
rect 19382 1932 19440 1944
rect 19382 1756 19394 1932
rect 19428 1756 19440 1932
rect 19382 1744 19440 1756
rect 19500 1932 19599 1944
rect 19500 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19645 2132
rect 19500 1744 19645 1756
rect 19705 2132 19763 2144
rect 19705 1756 19717 2132
rect 19751 1756 19763 2132
rect 19705 1744 19763 1756
rect 19823 2132 19881 2144
rect 19823 1756 19835 2132
rect 19869 1756 19881 2132
rect 19823 1744 19881 1756
rect 19941 2132 19999 2144
rect 19941 1756 19953 2132
rect 19987 1756 19999 2132
rect 19941 1744 19999 1756
rect 20054 2132 20112 2144
rect 20054 1756 20066 2132
rect 20100 1756 20112 2132
rect 20054 1744 20112 1756
rect 20172 2132 20230 2144
rect 20172 1756 20184 2132
rect 20218 1756 20230 2132
rect 20172 1744 20230 1756
rect 20290 2132 20348 2144
rect 20290 1756 20302 2132
rect 20336 1756 20348 2132
rect 20290 1744 20348 1756
rect 20408 2132 20466 2144
rect 20408 1756 20420 2132
rect 20454 1756 20466 2132
rect 20408 1744 20466 1756
rect 20526 2132 20584 2144
rect 20526 1756 20538 2132
rect 20572 1756 20584 2132
rect 20526 1744 20584 1756
rect 20644 2132 20702 2144
rect 20644 1756 20656 2132
rect 20690 1756 20702 2132
rect 20644 1744 20702 1756
rect 20762 2132 20820 2144
rect 20762 1756 20774 2132
rect 20808 1756 20820 2132
rect 20762 1744 20820 1756
rect 20881 2132 20939 2144
rect 20881 1756 20893 2132
rect 20927 1756 20939 2132
rect 20881 1744 20939 1756
rect 20999 2132 21057 2144
rect 20999 1756 21011 2132
rect 21045 1756 21057 2132
rect 20999 1744 21057 1756
rect 21117 2132 21175 2144
rect 21117 1756 21129 2132
rect 21163 1756 21175 2132
rect 21117 1744 21175 1756
rect 21235 2132 21293 2144
rect 21235 1756 21247 2132
rect 21281 1756 21293 2132
rect 22731 2132 22789 2144
rect 22731 1944 22743 2132
rect 21235 1744 21293 1756
rect 21354 1932 21412 1944
rect 21354 1756 21366 1932
rect 21400 1756 21412 1932
rect 21354 1744 21412 1756
rect 21472 1932 21530 1944
rect 21472 1756 21484 1932
rect 21518 1756 21530 1932
rect 21472 1744 21530 1756
rect 21590 1932 21648 1944
rect 21590 1756 21602 1932
rect 21636 1756 21648 1932
rect 21590 1744 21648 1756
rect 21708 1932 21766 1944
rect 21708 1756 21720 1932
rect 21754 1756 21766 1932
rect 21708 1744 21766 1756
rect 22290 1932 22348 1944
rect 22290 1756 22302 1932
rect 22336 1756 22348 1932
rect 22290 1744 22348 1756
rect 22408 1932 22466 1944
rect 22408 1756 22420 1932
rect 22454 1756 22466 1932
rect 22408 1744 22466 1756
rect 22526 1932 22584 1944
rect 22526 1756 22538 1932
rect 22572 1756 22584 1932
rect 22526 1744 22584 1756
rect 22644 1932 22743 1944
rect 22644 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22789 2132
rect 22644 1744 22789 1756
rect 22849 2132 22907 2144
rect 22849 1756 22861 2132
rect 22895 1756 22907 2132
rect 22849 1744 22907 1756
rect 22967 2132 23025 2144
rect 22967 1756 22979 2132
rect 23013 1756 23025 2132
rect 22967 1744 23025 1756
rect 23085 2132 23143 2144
rect 23085 1756 23097 2132
rect 23131 1756 23143 2132
rect 23085 1744 23143 1756
rect 23198 2132 23256 2144
rect 23198 1756 23210 2132
rect 23244 1756 23256 2132
rect 23198 1744 23256 1756
rect 23316 2132 23374 2144
rect 23316 1756 23328 2132
rect 23362 1756 23374 2132
rect 23316 1744 23374 1756
rect 23434 2132 23492 2144
rect 23434 1756 23446 2132
rect 23480 1756 23492 2132
rect 23434 1744 23492 1756
rect 23552 2132 23610 2144
rect 23552 1756 23564 2132
rect 23598 1756 23610 2132
rect 23552 1744 23610 1756
rect 23670 2132 23728 2144
rect 23670 1756 23682 2132
rect 23716 1756 23728 2132
rect 23670 1744 23728 1756
rect 23788 2132 23846 2144
rect 23788 1756 23800 2132
rect 23834 1756 23846 2132
rect 23788 1744 23846 1756
rect 23906 2132 23964 2144
rect 23906 1756 23918 2132
rect 23952 1756 23964 2132
rect 23906 1744 23964 1756
rect 24025 2132 24083 2144
rect 24025 1756 24037 2132
rect 24071 1756 24083 2132
rect 24025 1744 24083 1756
rect 24143 2132 24201 2144
rect 24143 1756 24155 2132
rect 24189 1756 24201 2132
rect 24143 1744 24201 1756
rect 24261 2132 24319 2144
rect 24261 1756 24273 2132
rect 24307 1756 24319 2132
rect 24261 1744 24319 1756
rect 24379 2132 24437 2144
rect 24379 1756 24391 2132
rect 24425 1756 24437 2132
rect 24379 1744 24437 1756
rect 24498 1932 24556 1944
rect 24498 1756 24510 1932
rect 24544 1756 24556 1932
rect 24498 1744 24556 1756
rect 24616 1932 24674 1944
rect 24616 1756 24628 1932
rect 24662 1756 24674 1932
rect 24616 1744 24674 1756
rect 24734 1932 24792 1944
rect 24734 1756 24746 1932
rect 24780 1756 24792 1932
rect 24734 1744 24792 1756
rect 24852 1932 24910 1944
rect 24852 1756 24864 1932
rect 24898 1756 24910 1932
rect 29950 2106 30350 2118
rect 29950 2072 29962 2106
rect 30338 2072 30350 2106
rect 29950 2060 30350 2072
rect 30643 2163 31043 2175
rect 30643 2129 30655 2163
rect 31031 2129 31043 2163
rect 30643 2117 31043 2129
rect 44341 2350 44399 2362
rect 44459 2538 44517 2550
rect 44459 2362 44471 2538
rect 44505 2362 44517 2538
rect 44459 2350 44517 2362
rect 44577 2538 44635 2550
rect 44577 2362 44589 2538
rect 44623 2362 44635 2538
rect 44577 2350 44635 2362
rect 44695 2538 44753 2550
rect 44695 2362 44707 2538
rect 44741 2362 44753 2538
rect 44695 2350 44753 2362
rect 44813 2538 44871 2550
rect 44813 2362 44825 2538
rect 44859 2362 44871 2538
rect 44813 2350 44871 2362
rect 44931 2538 44989 2550
rect 44931 2362 44943 2538
rect 44977 2362 44989 2538
rect 44931 2350 44989 2362
rect 45049 2538 45107 2550
rect 45049 2362 45061 2538
rect 45095 2362 45107 2538
rect 45049 2350 45107 2362
rect 45167 2538 45225 2550
rect 45167 2362 45179 2538
rect 45213 2362 45225 2538
rect 45167 2350 45225 2362
rect 45285 2538 45343 2550
rect 45285 2362 45297 2538
rect 45331 2362 45343 2538
rect 45285 2350 45343 2362
rect 45403 2538 45461 2550
rect 45403 2362 45415 2538
rect 45449 2362 45461 2538
rect 50996 2539 51054 2551
rect 45403 2350 45461 2362
rect 50996 2363 51008 2539
rect 51042 2363 51054 2539
rect 50996 2351 51054 2363
rect 51114 2539 51172 2551
rect 51114 2363 51126 2539
rect 51160 2363 51172 2539
rect 51114 2351 51172 2363
rect 51232 2539 51290 2551
rect 51232 2363 51244 2539
rect 51278 2363 51290 2539
rect 51232 2351 51290 2363
rect 51350 2539 51408 2551
rect 51350 2363 51362 2539
rect 51396 2363 51408 2539
rect 51350 2351 51408 2363
rect 51468 2539 51526 2551
rect 51468 2363 51480 2539
rect 51514 2363 51526 2539
rect 51468 2351 51526 2363
rect 51586 2539 51644 2551
rect 51586 2363 51598 2539
rect 51632 2363 51644 2539
rect 51586 2351 51644 2363
rect 51704 2539 51762 2551
rect 51704 2363 51716 2539
rect 51750 2363 51762 2539
rect 51704 2351 51762 2363
rect 51822 2539 51880 2551
rect 51822 2363 51834 2539
rect 51868 2363 51880 2539
rect 51822 2351 51880 2363
rect 51940 2539 51998 2551
rect 51940 2363 51952 2539
rect 51986 2363 51998 2539
rect 51940 2351 51998 2363
rect 52058 2539 52116 2551
rect 52058 2363 52070 2539
rect 52104 2363 52116 2539
rect 57618 2540 57676 2552
rect 52058 2351 52116 2363
rect 57618 2364 57630 2540
rect 57664 2364 57676 2540
rect 57618 2352 57676 2364
rect 57736 2540 57794 2552
rect 57736 2364 57748 2540
rect 57782 2364 57794 2540
rect 57736 2352 57794 2364
rect 57854 2540 57912 2552
rect 57854 2364 57866 2540
rect 57900 2364 57912 2540
rect 57854 2352 57912 2364
rect 57972 2540 58030 2552
rect 57972 2364 57984 2540
rect 58018 2364 58030 2540
rect 57972 2352 58030 2364
rect 58090 2540 58148 2552
rect 58090 2364 58102 2540
rect 58136 2364 58148 2540
rect 58090 2352 58148 2364
rect 58208 2540 58266 2552
rect 58208 2364 58220 2540
rect 58254 2364 58266 2540
rect 58208 2352 58266 2364
rect 58326 2540 58384 2552
rect 58326 2364 58338 2540
rect 58372 2364 58384 2540
rect 58326 2352 58384 2364
rect 58444 2540 58502 2552
rect 58444 2364 58456 2540
rect 58490 2364 58502 2540
rect 58444 2352 58502 2364
rect 58562 2540 58620 2552
rect 58562 2364 58574 2540
rect 58608 2364 58620 2540
rect 58562 2352 58620 2364
rect 58680 2540 58738 2552
rect 58680 2364 58692 2540
rect 58726 2364 58738 2540
rect 70709 2775 70721 2809
rect 70897 2775 70909 2809
rect 70709 2734 70909 2775
rect 70509 2722 70909 2734
rect 70509 2688 70521 2722
rect 70897 2688 70909 2722
rect 70509 2676 70909 2688
rect 70509 2604 70909 2616
rect 70509 2570 70521 2604
rect 70897 2570 70909 2604
rect 70509 2558 70909 2570
rect 70509 2486 70909 2498
rect 70509 2452 70521 2486
rect 70897 2452 70909 2486
rect 70509 2440 70909 2452
rect 58680 2352 58738 2364
rect 70509 2368 70909 2380
rect 39738 2123 39796 2135
rect 30643 2045 31043 2057
rect 30643 2011 30655 2045
rect 31031 2011 31043 2045
rect 29950 1988 30350 2000
rect 30643 1999 31043 2011
rect 29950 1954 29962 1988
rect 30338 1954 30350 1988
rect 29950 1942 30350 1954
rect 29950 1870 30350 1882
rect 29950 1836 29962 1870
rect 30338 1836 30350 1870
rect 29950 1824 30350 1836
rect 24852 1744 24910 1756
rect 29950 1752 30350 1764
rect 29950 1718 29962 1752
rect 30338 1718 30350 1752
rect 29950 1706 30350 1718
rect 30643 1927 31043 1939
rect 30643 1893 30655 1927
rect 31031 1893 31043 1927
rect 30643 1881 31043 1893
rect 30643 1809 31043 1821
rect 30643 1775 30655 1809
rect 31031 1775 31043 1809
rect 30643 1763 31043 1775
rect 29950 1634 30350 1646
rect 29950 1600 29962 1634
rect 30338 1600 30350 1634
rect 29950 1588 30350 1600
rect 30150 1505 30350 1517
rect 30150 1471 30162 1505
rect 30338 1471 30350 1505
rect 30150 1459 30350 1471
rect 30643 1691 31043 1703
rect 30643 1657 30655 1691
rect 31031 1657 31043 1691
rect 39254 1923 39312 1935
rect 30643 1645 31043 1657
rect 39254 1747 39266 1923
rect 39300 1747 39312 1923
rect 39254 1735 39312 1747
rect 39372 1923 39430 1935
rect 39372 1747 39384 1923
rect 39418 1747 39430 1923
rect 39372 1735 39430 1747
rect 39490 1923 39548 1935
rect 39490 1747 39502 1923
rect 39536 1747 39548 1923
rect 39490 1735 39548 1747
rect 39608 1923 39666 1935
rect 39608 1747 39620 1923
rect 39654 1747 39666 1923
rect 39608 1735 39666 1747
rect 39738 1747 39750 2123
rect 39784 1747 39796 2123
rect 39738 1735 39796 1747
rect 39856 2123 39914 2135
rect 39856 1747 39868 2123
rect 39902 1747 39914 2123
rect 39856 1735 39914 1747
rect 39974 2123 40032 2135
rect 39974 1747 39986 2123
rect 40020 1747 40032 2123
rect 39974 1735 40032 1747
rect 40092 2123 40150 2135
rect 40092 1747 40104 2123
rect 40138 1747 40150 2123
rect 40092 1735 40150 1747
rect 40210 2123 40268 2135
rect 40210 1747 40222 2123
rect 40256 1747 40268 2123
rect 40210 1735 40268 1747
rect 40328 2123 40386 2135
rect 40328 1747 40340 2123
rect 40374 1747 40386 2123
rect 40328 1735 40386 1747
rect 40446 2123 40504 2135
rect 40446 1747 40458 2123
rect 40492 1747 40504 2123
rect 41636 2123 41694 2135
rect 40446 1735 40504 1747
rect 40575 1923 40633 1935
rect 40575 1747 40587 1923
rect 40621 1747 40633 1923
rect 40575 1735 40633 1747
rect 40693 1923 40751 1935
rect 40693 1747 40705 1923
rect 40739 1747 40751 1923
rect 40693 1735 40751 1747
rect 40811 1923 40869 1935
rect 40811 1747 40823 1923
rect 40857 1747 40869 1923
rect 40811 1735 40869 1747
rect 40929 1923 40987 1935
rect 40929 1747 40941 1923
rect 40975 1747 40987 1923
rect 40929 1735 40987 1747
rect 41152 1923 41210 1935
rect 41152 1747 41164 1923
rect 41198 1747 41210 1923
rect 41152 1735 41210 1747
rect 41270 1923 41328 1935
rect 41270 1747 41282 1923
rect 41316 1747 41328 1923
rect 41270 1735 41328 1747
rect 41388 1923 41446 1935
rect 41388 1747 41400 1923
rect 41434 1747 41446 1923
rect 41388 1735 41446 1747
rect 41506 1923 41564 1935
rect 41506 1747 41518 1923
rect 41552 1747 41564 1923
rect 41506 1735 41564 1747
rect 41636 1747 41648 2123
rect 41682 1747 41694 2123
rect 41636 1735 41694 1747
rect 41754 2123 41812 2135
rect 41754 1747 41766 2123
rect 41800 1747 41812 2123
rect 41754 1735 41812 1747
rect 41872 2123 41930 2135
rect 41872 1747 41884 2123
rect 41918 1747 41930 2123
rect 41872 1735 41930 1747
rect 41990 2123 42048 2135
rect 41990 1747 42002 2123
rect 42036 1747 42048 2123
rect 41990 1735 42048 1747
rect 42108 2123 42166 2135
rect 42108 1747 42120 2123
rect 42154 1747 42166 2123
rect 42108 1735 42166 1747
rect 42226 2123 42284 2135
rect 42226 1747 42238 2123
rect 42272 1747 42284 2123
rect 42226 1735 42284 1747
rect 42344 2123 42402 2135
rect 42344 1747 42356 2123
rect 42390 1747 42402 2123
rect 46289 2121 46347 2133
rect 42344 1735 42402 1747
rect 42473 1923 42531 1935
rect 42473 1747 42485 1923
rect 42519 1747 42531 1923
rect 42473 1735 42531 1747
rect 42591 1923 42649 1935
rect 42591 1747 42603 1923
rect 42637 1747 42649 1923
rect 42591 1735 42649 1747
rect 42709 1923 42767 1935
rect 42709 1747 42721 1923
rect 42755 1747 42767 1923
rect 42709 1735 42767 1747
rect 42827 1923 42885 1935
rect 42827 1747 42839 1923
rect 42873 1747 42885 1923
rect 42827 1735 42885 1747
rect 34883 1614 34941 1626
rect 30150 1387 30350 1399
rect 30150 1353 30162 1387
rect 30338 1353 30350 1387
rect 34883 1438 34895 1614
rect 34929 1438 34941 1614
rect 34883 1426 34941 1438
rect 35001 1614 35059 1626
rect 35001 1438 35013 1614
rect 35047 1438 35059 1614
rect 35001 1426 35059 1438
rect 35119 1614 35177 1626
rect 35119 1438 35131 1614
rect 35165 1438 35177 1614
rect 35119 1426 35177 1438
rect 35237 1614 35295 1626
rect 35237 1438 35249 1614
rect 35283 1438 35295 1614
rect 35237 1426 35295 1438
rect 35355 1614 35413 1626
rect 35355 1438 35367 1614
rect 35401 1438 35413 1614
rect 35355 1426 35413 1438
rect 35473 1614 35531 1626
rect 35473 1438 35485 1614
rect 35519 1438 35531 1614
rect 35473 1426 35531 1438
rect 35591 1614 35649 1626
rect 35591 1438 35603 1614
rect 35637 1438 35649 1614
rect 35591 1426 35649 1438
rect 35709 1614 35767 1626
rect 35709 1438 35721 1614
rect 35755 1438 35767 1614
rect 35709 1426 35767 1438
rect 35827 1614 35885 1626
rect 35827 1438 35839 1614
rect 35873 1438 35885 1614
rect 35827 1426 35885 1438
rect 35945 1614 36003 1626
rect 35945 1438 35957 1614
rect 35991 1438 36003 1614
rect 35945 1426 36003 1438
rect 30150 1341 30350 1353
rect 30150 1269 30350 1281
rect 30150 1235 30162 1269
rect 30338 1235 30350 1269
rect 30150 1223 30350 1235
rect 30150 1151 30350 1163
rect 30150 1117 30162 1151
rect 30338 1117 30350 1151
rect 30150 1105 30350 1117
rect 37785 936 37843 948
rect 30152 757 30352 769
rect 30152 723 30164 757
rect 30340 723 30352 757
rect 30152 711 30352 723
rect 30152 639 30352 651
rect 30152 605 30164 639
rect 30340 605 30352 639
rect 30152 593 30352 605
rect 37785 760 37797 936
rect 37831 760 37843 936
rect 37785 748 37843 760
rect 37903 936 37961 948
rect 37903 760 37915 936
rect 37949 760 37961 936
rect 37903 748 37961 760
rect 38021 936 38079 948
rect 38021 760 38033 936
rect 38067 760 38079 936
rect 38021 748 38079 760
rect 38139 936 38197 948
rect 38139 760 38151 936
rect 38185 760 38197 936
rect 38139 748 38197 760
rect 38257 936 38315 948
rect 38257 760 38269 936
rect 38303 760 38315 936
rect 38257 748 38315 760
rect 38375 936 38433 948
rect 38375 760 38387 936
rect 38421 760 38433 936
rect 38375 748 38433 760
rect 38493 936 38551 948
rect 38493 760 38505 936
rect 38539 760 38551 936
rect 38493 748 38551 760
rect 38611 936 38669 948
rect 38611 760 38623 936
rect 38657 760 38669 936
rect 38611 748 38669 760
rect 38729 936 38787 948
rect 38729 760 38741 936
rect 38775 760 38787 936
rect 38729 748 38787 760
rect 38847 936 38905 948
rect 38847 760 38859 936
rect 38893 760 38905 936
rect 38847 748 38905 760
rect 39681 1430 39739 1442
rect 39681 1054 39693 1430
rect 39727 1054 39739 1430
rect 39681 1042 39739 1054
rect 39799 1430 39857 1442
rect 39799 1054 39811 1430
rect 39845 1054 39857 1430
rect 39799 1042 39857 1054
rect 39917 1430 39975 1442
rect 39917 1054 39929 1430
rect 39963 1054 39975 1430
rect 39917 1042 39975 1054
rect 40035 1430 40093 1442
rect 40035 1054 40047 1430
rect 40081 1054 40093 1430
rect 40035 1042 40093 1054
rect 40153 1430 40211 1442
rect 40153 1054 40165 1430
rect 40199 1054 40211 1430
rect 40153 1042 40211 1054
rect 40271 1430 40329 1442
rect 40271 1054 40283 1430
rect 40317 1054 40329 1430
rect 40271 1042 40329 1054
rect 40389 1430 40447 1442
rect 40389 1054 40401 1430
rect 40435 1054 40447 1430
rect 40389 1042 40447 1054
rect 30152 521 30352 533
rect 30152 487 30164 521
rect 30340 487 30352 521
rect 30152 475 30352 487
rect 45805 1921 45863 1933
rect 45805 1745 45817 1921
rect 45851 1745 45863 1921
rect 45805 1733 45863 1745
rect 45923 1921 45981 1933
rect 45923 1745 45935 1921
rect 45969 1745 45981 1921
rect 45923 1733 45981 1745
rect 46041 1921 46099 1933
rect 46041 1745 46053 1921
rect 46087 1745 46099 1921
rect 46041 1733 46099 1745
rect 46159 1921 46217 1933
rect 46159 1745 46171 1921
rect 46205 1745 46217 1921
rect 46159 1733 46217 1745
rect 46289 1745 46301 2121
rect 46335 1745 46347 2121
rect 46289 1733 46347 1745
rect 46407 2121 46465 2133
rect 46407 1745 46419 2121
rect 46453 1745 46465 2121
rect 46407 1733 46465 1745
rect 46525 2121 46583 2133
rect 46525 1745 46537 2121
rect 46571 1745 46583 2121
rect 46525 1733 46583 1745
rect 46643 2121 46701 2133
rect 46643 1745 46655 2121
rect 46689 1745 46701 2121
rect 46643 1733 46701 1745
rect 46761 2121 46819 2133
rect 46761 1745 46773 2121
rect 46807 1745 46819 2121
rect 46761 1733 46819 1745
rect 46879 2121 46937 2133
rect 46879 1745 46891 2121
rect 46925 1745 46937 2121
rect 46879 1733 46937 1745
rect 46997 2121 47055 2133
rect 46997 1745 47009 2121
rect 47043 1745 47055 2121
rect 48187 2121 48245 2133
rect 46997 1733 47055 1745
rect 47126 1921 47184 1933
rect 47126 1745 47138 1921
rect 47172 1745 47184 1921
rect 47126 1733 47184 1745
rect 47244 1921 47302 1933
rect 47244 1745 47256 1921
rect 47290 1745 47302 1921
rect 47244 1733 47302 1745
rect 47362 1921 47420 1933
rect 47362 1745 47374 1921
rect 47408 1745 47420 1921
rect 47362 1733 47420 1745
rect 47480 1921 47538 1933
rect 47480 1745 47492 1921
rect 47526 1745 47538 1921
rect 47480 1733 47538 1745
rect 47703 1921 47761 1933
rect 47703 1745 47715 1921
rect 47749 1745 47761 1921
rect 47703 1733 47761 1745
rect 47821 1921 47879 1933
rect 47821 1745 47833 1921
rect 47867 1745 47879 1921
rect 47821 1733 47879 1745
rect 47939 1921 47997 1933
rect 47939 1745 47951 1921
rect 47985 1745 47997 1921
rect 47939 1733 47997 1745
rect 48057 1921 48115 1933
rect 48057 1745 48069 1921
rect 48103 1745 48115 1921
rect 48057 1733 48115 1745
rect 48187 1745 48199 2121
rect 48233 1745 48245 2121
rect 48187 1733 48245 1745
rect 48305 2121 48363 2133
rect 48305 1745 48317 2121
rect 48351 1745 48363 2121
rect 48305 1733 48363 1745
rect 48423 2121 48481 2133
rect 48423 1745 48435 2121
rect 48469 1745 48481 2121
rect 48423 1733 48481 1745
rect 48541 2121 48599 2133
rect 48541 1745 48553 2121
rect 48587 1745 48599 2121
rect 48541 1733 48599 1745
rect 48659 2121 48717 2133
rect 48659 1745 48671 2121
rect 48705 1745 48717 2121
rect 48659 1733 48717 1745
rect 48777 2121 48835 2133
rect 48777 1745 48789 2121
rect 48823 1745 48835 2121
rect 48777 1733 48835 1745
rect 48895 2121 48953 2133
rect 48895 1745 48907 2121
rect 48941 1745 48953 2121
rect 52944 2122 53002 2134
rect 48895 1733 48953 1745
rect 49024 1921 49082 1933
rect 49024 1745 49036 1921
rect 49070 1745 49082 1921
rect 49024 1733 49082 1745
rect 49142 1921 49200 1933
rect 49142 1745 49154 1921
rect 49188 1745 49200 1921
rect 49142 1733 49200 1745
rect 49260 1921 49318 1933
rect 49260 1745 49272 1921
rect 49306 1745 49318 1921
rect 49260 1733 49318 1745
rect 49378 1921 49436 1933
rect 49378 1745 49390 1921
rect 49424 1745 49436 1921
rect 49378 1733 49436 1745
rect 41579 1430 41637 1442
rect 41579 1054 41591 1430
rect 41625 1054 41637 1430
rect 41579 1042 41637 1054
rect 41697 1430 41755 1442
rect 41697 1054 41709 1430
rect 41743 1054 41755 1430
rect 41697 1042 41755 1054
rect 41815 1430 41873 1442
rect 41815 1054 41827 1430
rect 41861 1054 41873 1430
rect 41815 1042 41873 1054
rect 41933 1430 41991 1442
rect 41933 1054 41945 1430
rect 41979 1054 41991 1430
rect 41933 1042 41991 1054
rect 42051 1430 42109 1442
rect 42051 1054 42063 1430
rect 42097 1054 42109 1430
rect 42051 1042 42109 1054
rect 42169 1430 42227 1442
rect 42169 1054 42181 1430
rect 42215 1054 42227 1430
rect 42169 1042 42227 1054
rect 42287 1430 42345 1442
rect 42287 1054 42299 1430
rect 42333 1054 42345 1430
rect 42287 1042 42345 1054
rect 44336 934 44394 946
rect 44336 758 44348 934
rect 44382 758 44394 934
rect 44336 746 44394 758
rect 44454 934 44512 946
rect 44454 758 44466 934
rect 44500 758 44512 934
rect 44454 746 44512 758
rect 44572 934 44630 946
rect 44572 758 44584 934
rect 44618 758 44630 934
rect 44572 746 44630 758
rect 44690 934 44748 946
rect 44690 758 44702 934
rect 44736 758 44748 934
rect 44690 746 44748 758
rect 44808 934 44866 946
rect 44808 758 44820 934
rect 44854 758 44866 934
rect 44808 746 44866 758
rect 44926 934 44984 946
rect 44926 758 44938 934
rect 44972 758 44984 934
rect 44926 746 44984 758
rect 45044 934 45102 946
rect 45044 758 45056 934
rect 45090 758 45102 934
rect 45044 746 45102 758
rect 45162 934 45220 946
rect 45162 758 45174 934
rect 45208 758 45220 934
rect 45162 746 45220 758
rect 45280 934 45338 946
rect 45280 758 45292 934
rect 45326 758 45338 934
rect 45280 746 45338 758
rect 45398 934 45456 946
rect 45398 758 45410 934
rect 45444 758 45456 934
rect 45398 746 45456 758
rect 46232 1428 46290 1440
rect 46232 1052 46244 1428
rect 46278 1052 46290 1428
rect 46232 1040 46290 1052
rect 46350 1428 46408 1440
rect 46350 1052 46362 1428
rect 46396 1052 46408 1428
rect 46350 1040 46408 1052
rect 46468 1428 46526 1440
rect 46468 1052 46480 1428
rect 46514 1052 46526 1428
rect 46468 1040 46526 1052
rect 46586 1428 46644 1440
rect 46586 1052 46598 1428
rect 46632 1052 46644 1428
rect 46586 1040 46644 1052
rect 46704 1428 46762 1440
rect 46704 1052 46716 1428
rect 46750 1052 46762 1428
rect 46704 1040 46762 1052
rect 46822 1428 46880 1440
rect 46822 1052 46834 1428
rect 46868 1052 46880 1428
rect 46822 1040 46880 1052
rect 46940 1428 46998 1440
rect 46940 1052 46952 1428
rect 46986 1052 46998 1428
rect 46940 1040 46998 1052
rect 30152 403 30352 415
rect 30152 369 30164 403
rect 30340 369 30352 403
rect 30152 357 30352 369
rect 29952 273 30352 285
rect 29952 239 29964 273
rect 30340 239 30352 273
rect 29952 227 30352 239
rect 30645 330 31045 342
rect 30645 296 30657 330
rect 31033 296 31045 330
rect 30645 284 31045 296
rect 29952 155 30352 167
rect 29952 121 29964 155
rect 30340 121 30352 155
rect 29952 109 30352 121
rect 30645 212 31045 224
rect 30645 178 30657 212
rect 31033 178 31045 212
rect 30645 166 31045 178
rect 52460 1922 52518 1934
rect 52460 1746 52472 1922
rect 52506 1746 52518 1922
rect 52460 1734 52518 1746
rect 52578 1922 52636 1934
rect 52578 1746 52590 1922
rect 52624 1746 52636 1922
rect 52578 1734 52636 1746
rect 52696 1922 52754 1934
rect 52696 1746 52708 1922
rect 52742 1746 52754 1922
rect 52696 1734 52754 1746
rect 52814 1922 52872 1934
rect 52814 1746 52826 1922
rect 52860 1746 52872 1922
rect 52814 1734 52872 1746
rect 52944 1746 52956 2122
rect 52990 1746 53002 2122
rect 52944 1734 53002 1746
rect 53062 2122 53120 2134
rect 53062 1746 53074 2122
rect 53108 1746 53120 2122
rect 53062 1734 53120 1746
rect 53180 2122 53238 2134
rect 53180 1746 53192 2122
rect 53226 1746 53238 2122
rect 53180 1734 53238 1746
rect 53298 2122 53356 2134
rect 53298 1746 53310 2122
rect 53344 1746 53356 2122
rect 53298 1734 53356 1746
rect 53416 2122 53474 2134
rect 53416 1746 53428 2122
rect 53462 1746 53474 2122
rect 53416 1734 53474 1746
rect 53534 2122 53592 2134
rect 53534 1746 53546 2122
rect 53580 1746 53592 2122
rect 53534 1734 53592 1746
rect 53652 2122 53710 2134
rect 53652 1746 53664 2122
rect 53698 1746 53710 2122
rect 54842 2122 54900 2134
rect 53652 1734 53710 1746
rect 53781 1922 53839 1934
rect 53781 1746 53793 1922
rect 53827 1746 53839 1922
rect 53781 1734 53839 1746
rect 53899 1922 53957 1934
rect 53899 1746 53911 1922
rect 53945 1746 53957 1922
rect 53899 1734 53957 1746
rect 54017 1922 54075 1934
rect 54017 1746 54029 1922
rect 54063 1746 54075 1922
rect 54017 1734 54075 1746
rect 54135 1922 54193 1934
rect 54135 1746 54147 1922
rect 54181 1746 54193 1922
rect 54135 1734 54193 1746
rect 54358 1922 54416 1934
rect 54358 1746 54370 1922
rect 54404 1746 54416 1922
rect 54358 1734 54416 1746
rect 54476 1922 54534 1934
rect 54476 1746 54488 1922
rect 54522 1746 54534 1922
rect 54476 1734 54534 1746
rect 54594 1922 54652 1934
rect 54594 1746 54606 1922
rect 54640 1746 54652 1922
rect 54594 1734 54652 1746
rect 54712 1922 54770 1934
rect 54712 1746 54724 1922
rect 54758 1746 54770 1922
rect 54712 1734 54770 1746
rect 54842 1746 54854 2122
rect 54888 1746 54900 2122
rect 54842 1734 54900 1746
rect 54960 2122 55018 2134
rect 54960 1746 54972 2122
rect 55006 1746 55018 2122
rect 54960 1734 55018 1746
rect 55078 2122 55136 2134
rect 55078 1746 55090 2122
rect 55124 1746 55136 2122
rect 55078 1734 55136 1746
rect 55196 2122 55254 2134
rect 55196 1746 55208 2122
rect 55242 1746 55254 2122
rect 55196 1734 55254 1746
rect 55314 2122 55372 2134
rect 55314 1746 55326 2122
rect 55360 1746 55372 2122
rect 55314 1734 55372 1746
rect 55432 2122 55490 2134
rect 55432 1746 55444 2122
rect 55478 1746 55490 2122
rect 55432 1734 55490 1746
rect 55550 2122 55608 2134
rect 55550 1746 55562 2122
rect 55596 1746 55608 2122
rect 70509 2334 70521 2368
rect 70897 2334 70909 2368
rect 70509 2322 70909 2334
rect 70509 2255 70909 2267
rect 59566 2123 59624 2135
rect 55550 1734 55608 1746
rect 55679 1922 55737 1934
rect 55679 1746 55691 1922
rect 55725 1746 55737 1922
rect 55679 1734 55737 1746
rect 55797 1922 55855 1934
rect 55797 1746 55809 1922
rect 55843 1746 55855 1922
rect 55797 1734 55855 1746
rect 55915 1922 55973 1934
rect 55915 1746 55927 1922
rect 55961 1746 55973 1922
rect 55915 1734 55973 1746
rect 56033 1922 56091 1934
rect 56033 1746 56045 1922
rect 56079 1746 56091 1922
rect 56033 1734 56091 1746
rect 48130 1428 48188 1440
rect 48130 1052 48142 1428
rect 48176 1052 48188 1428
rect 48130 1040 48188 1052
rect 48248 1428 48306 1440
rect 48248 1052 48260 1428
rect 48294 1052 48306 1428
rect 48248 1040 48306 1052
rect 48366 1428 48424 1440
rect 48366 1052 48378 1428
rect 48412 1052 48424 1428
rect 48366 1040 48424 1052
rect 48484 1428 48542 1440
rect 48484 1052 48496 1428
rect 48530 1052 48542 1428
rect 48484 1040 48542 1052
rect 48602 1428 48660 1440
rect 48602 1052 48614 1428
rect 48648 1052 48660 1428
rect 48602 1040 48660 1052
rect 48720 1428 48778 1440
rect 48720 1052 48732 1428
rect 48766 1052 48778 1428
rect 48720 1040 48778 1052
rect 48838 1428 48896 1440
rect 48838 1052 48850 1428
rect 48884 1052 48896 1428
rect 48838 1040 48896 1052
rect 50991 935 51049 947
rect 50991 759 51003 935
rect 51037 759 51049 935
rect 50991 747 51049 759
rect 51109 935 51167 947
rect 51109 759 51121 935
rect 51155 759 51167 935
rect 51109 747 51167 759
rect 51227 935 51285 947
rect 51227 759 51239 935
rect 51273 759 51285 935
rect 51227 747 51285 759
rect 51345 935 51403 947
rect 51345 759 51357 935
rect 51391 759 51403 935
rect 51345 747 51403 759
rect 51463 935 51521 947
rect 51463 759 51475 935
rect 51509 759 51521 935
rect 51463 747 51521 759
rect 51581 935 51639 947
rect 51581 759 51593 935
rect 51627 759 51639 935
rect 51581 747 51639 759
rect 51699 935 51757 947
rect 51699 759 51711 935
rect 51745 759 51757 935
rect 51699 747 51757 759
rect 51817 935 51875 947
rect 51817 759 51829 935
rect 51863 759 51875 935
rect 51817 747 51875 759
rect 51935 935 51993 947
rect 51935 759 51947 935
rect 51981 759 51993 935
rect 51935 747 51993 759
rect 52053 935 52111 947
rect 52053 759 52065 935
rect 52099 759 52111 935
rect 52053 747 52111 759
rect 52887 1429 52945 1441
rect 52887 1053 52899 1429
rect 52933 1053 52945 1429
rect 52887 1041 52945 1053
rect 53005 1429 53063 1441
rect 53005 1053 53017 1429
rect 53051 1053 53063 1429
rect 53005 1041 53063 1053
rect 53123 1429 53181 1441
rect 53123 1053 53135 1429
rect 53169 1053 53181 1429
rect 53123 1041 53181 1053
rect 53241 1429 53299 1441
rect 53241 1053 53253 1429
rect 53287 1053 53299 1429
rect 53241 1041 53299 1053
rect 53359 1429 53417 1441
rect 53359 1053 53371 1429
rect 53405 1053 53417 1429
rect 53359 1041 53417 1053
rect 53477 1429 53535 1441
rect 53477 1053 53489 1429
rect 53523 1053 53535 1429
rect 53477 1041 53535 1053
rect 53595 1429 53653 1441
rect 53595 1053 53607 1429
rect 53641 1053 53653 1429
rect 53595 1041 53653 1053
rect 29952 37 30352 49
rect 29952 3 29964 37
rect 30340 3 30352 37
rect 29952 -9 30352 3
rect 30645 94 31045 106
rect 30645 60 30657 94
rect 31033 60 31045 94
rect 30645 48 31045 60
rect 59082 1923 59140 1935
rect 59082 1747 59094 1923
rect 59128 1747 59140 1923
rect 59082 1735 59140 1747
rect 59200 1923 59258 1935
rect 59200 1747 59212 1923
rect 59246 1747 59258 1923
rect 59200 1735 59258 1747
rect 59318 1923 59376 1935
rect 59318 1747 59330 1923
rect 59364 1747 59376 1923
rect 59318 1735 59376 1747
rect 59436 1923 59494 1935
rect 59436 1747 59448 1923
rect 59482 1747 59494 1923
rect 59436 1735 59494 1747
rect 59566 1747 59578 2123
rect 59612 1747 59624 2123
rect 59566 1735 59624 1747
rect 59684 2123 59742 2135
rect 59684 1747 59696 2123
rect 59730 1747 59742 2123
rect 59684 1735 59742 1747
rect 59802 2123 59860 2135
rect 59802 1747 59814 2123
rect 59848 1747 59860 2123
rect 59802 1735 59860 1747
rect 59920 2123 59978 2135
rect 59920 1747 59932 2123
rect 59966 1747 59978 2123
rect 59920 1735 59978 1747
rect 60038 2123 60096 2135
rect 60038 1747 60050 2123
rect 60084 1747 60096 2123
rect 60038 1735 60096 1747
rect 60156 2123 60214 2135
rect 60156 1747 60168 2123
rect 60202 1747 60214 2123
rect 60156 1735 60214 1747
rect 60274 2123 60332 2135
rect 60274 1747 60286 2123
rect 60320 1747 60332 2123
rect 61464 2123 61522 2135
rect 60274 1735 60332 1747
rect 60403 1923 60461 1935
rect 60403 1747 60415 1923
rect 60449 1747 60461 1923
rect 60403 1735 60461 1747
rect 60521 1923 60579 1935
rect 60521 1747 60533 1923
rect 60567 1747 60579 1923
rect 60521 1735 60579 1747
rect 60639 1923 60697 1935
rect 60639 1747 60651 1923
rect 60685 1747 60697 1923
rect 60639 1735 60697 1747
rect 60757 1923 60815 1935
rect 60757 1747 60769 1923
rect 60803 1747 60815 1923
rect 60757 1735 60815 1747
rect 60980 1923 61038 1935
rect 60980 1747 60992 1923
rect 61026 1747 61038 1923
rect 60980 1735 61038 1747
rect 61098 1923 61156 1935
rect 61098 1747 61110 1923
rect 61144 1747 61156 1923
rect 61098 1735 61156 1747
rect 61216 1923 61274 1935
rect 61216 1747 61228 1923
rect 61262 1747 61274 1923
rect 61216 1735 61274 1747
rect 61334 1923 61392 1935
rect 61334 1747 61346 1923
rect 61380 1747 61392 1923
rect 61334 1735 61392 1747
rect 61464 1747 61476 2123
rect 61510 1747 61522 2123
rect 61464 1735 61522 1747
rect 61582 2123 61640 2135
rect 61582 1747 61594 2123
rect 61628 1747 61640 2123
rect 61582 1735 61640 1747
rect 61700 2123 61758 2135
rect 61700 1747 61712 2123
rect 61746 1747 61758 2123
rect 61700 1735 61758 1747
rect 61818 2123 61876 2135
rect 61818 1747 61830 2123
rect 61864 1747 61876 2123
rect 61818 1735 61876 1747
rect 61936 2123 61994 2135
rect 61936 1747 61948 2123
rect 61982 1747 61994 2123
rect 61936 1735 61994 1747
rect 62054 2123 62112 2135
rect 62054 1747 62066 2123
rect 62100 1747 62112 2123
rect 62054 1735 62112 1747
rect 62172 2123 62230 2135
rect 62172 1747 62184 2123
rect 62218 1747 62230 2123
rect 70509 2221 70521 2255
rect 70897 2221 70909 2255
rect 70509 2209 70909 2221
rect 70509 2137 70909 2149
rect 70509 2103 70521 2137
rect 70897 2103 70909 2137
rect 70509 2091 70909 2103
rect 62172 1735 62230 1747
rect 62301 1923 62359 1935
rect 62301 1747 62313 1923
rect 62347 1747 62359 1923
rect 62301 1735 62359 1747
rect 62419 1923 62477 1935
rect 62419 1747 62431 1923
rect 62465 1747 62477 1923
rect 62419 1735 62477 1747
rect 62537 1923 62595 1935
rect 62537 1747 62549 1923
rect 62583 1747 62595 1923
rect 62537 1735 62595 1747
rect 62655 1923 62713 1935
rect 62655 1747 62667 1923
rect 62701 1747 62713 1923
rect 62655 1735 62713 1747
rect 70509 2019 70909 2031
rect 70509 1985 70521 2019
rect 70897 1985 70909 2019
rect 70509 1973 70909 1985
rect 70509 1901 70909 1913
rect 70509 1867 70521 1901
rect 70897 1867 70909 1901
rect 70509 1855 70909 1867
rect 54785 1429 54843 1441
rect 54785 1053 54797 1429
rect 54831 1053 54843 1429
rect 54785 1041 54843 1053
rect 54903 1429 54961 1441
rect 54903 1053 54915 1429
rect 54949 1053 54961 1429
rect 54903 1041 54961 1053
rect 55021 1429 55079 1441
rect 55021 1053 55033 1429
rect 55067 1053 55079 1429
rect 55021 1041 55079 1053
rect 55139 1429 55197 1441
rect 55139 1053 55151 1429
rect 55185 1053 55197 1429
rect 55139 1041 55197 1053
rect 55257 1429 55315 1441
rect 55257 1053 55269 1429
rect 55303 1053 55315 1429
rect 55257 1041 55315 1053
rect 55375 1429 55433 1441
rect 55375 1053 55387 1429
rect 55421 1053 55433 1429
rect 55375 1041 55433 1053
rect 55493 1429 55551 1441
rect 55493 1053 55505 1429
rect 55539 1053 55551 1429
rect 55493 1041 55551 1053
rect 57613 936 57671 948
rect 57613 760 57625 936
rect 57659 760 57671 936
rect 57613 748 57671 760
rect 57731 936 57789 948
rect 57731 760 57743 936
rect 57777 760 57789 936
rect 57731 748 57789 760
rect 57849 936 57907 948
rect 57849 760 57861 936
rect 57895 760 57907 936
rect 57849 748 57907 760
rect 57967 936 58025 948
rect 57967 760 57979 936
rect 58013 760 58025 936
rect 57967 748 58025 760
rect 58085 936 58143 948
rect 58085 760 58097 936
rect 58131 760 58143 936
rect 58085 748 58143 760
rect 58203 936 58261 948
rect 58203 760 58215 936
rect 58249 760 58261 936
rect 58203 748 58261 760
rect 58321 936 58379 948
rect 58321 760 58333 936
rect 58367 760 58379 936
rect 58321 748 58379 760
rect 58439 936 58497 948
rect 58439 760 58451 936
rect 58485 760 58497 936
rect 58439 748 58497 760
rect 58557 936 58615 948
rect 58557 760 58569 936
rect 58603 760 58615 936
rect 58557 748 58615 760
rect 58675 936 58733 948
rect 58675 760 58687 936
rect 58721 760 58733 936
rect 58675 748 58733 760
rect 59509 1430 59567 1442
rect 59509 1054 59521 1430
rect 59555 1054 59567 1430
rect 59509 1042 59567 1054
rect 59627 1430 59685 1442
rect 59627 1054 59639 1430
rect 59673 1054 59685 1430
rect 59627 1042 59685 1054
rect 59745 1430 59803 1442
rect 59745 1054 59757 1430
rect 59791 1054 59803 1430
rect 59745 1042 59803 1054
rect 59863 1430 59921 1442
rect 59863 1054 59875 1430
rect 59909 1054 59921 1430
rect 59863 1042 59921 1054
rect 59981 1430 60039 1442
rect 59981 1054 59993 1430
rect 60027 1054 60039 1430
rect 59981 1042 60039 1054
rect 60099 1430 60157 1442
rect 60099 1054 60111 1430
rect 60145 1054 60157 1430
rect 60099 1042 60157 1054
rect 60217 1430 60275 1442
rect 60217 1054 60229 1430
rect 60263 1054 60275 1430
rect 60217 1042 60275 1054
rect 30645 -24 31045 -12
rect 30645 -58 30657 -24
rect 31033 -58 31045 -24
rect 29952 -81 30352 -69
rect 30645 -70 31045 -58
rect 29952 -115 29964 -81
rect 30340 -115 30352 -81
rect 29952 -127 30352 -115
rect 29952 -199 30352 -187
rect 29952 -233 29964 -199
rect 30340 -233 30352 -199
rect 29952 -245 30352 -233
rect 29952 -317 30352 -305
rect 29952 -351 29964 -317
rect 30340 -351 30352 -317
rect 29952 -363 30352 -351
rect 30645 -142 31045 -130
rect 30645 -176 30657 -142
rect 31033 -176 31045 -142
rect 30645 -188 31045 -176
rect 70509 1783 70909 1795
rect 70509 1749 70521 1783
rect 70897 1749 70909 1783
rect 70509 1737 70909 1749
rect 70509 1665 70909 1677
rect 70509 1631 70521 1665
rect 70897 1631 70909 1665
rect 70509 1619 70909 1631
rect 70509 1547 70909 1559
rect 70509 1513 70521 1547
rect 70897 1513 70909 1547
rect 70509 1501 70909 1513
rect 61407 1430 61465 1442
rect 61407 1054 61419 1430
rect 61453 1054 61465 1430
rect 61407 1042 61465 1054
rect 61525 1430 61583 1442
rect 61525 1054 61537 1430
rect 61571 1054 61583 1430
rect 61525 1042 61583 1054
rect 61643 1430 61701 1442
rect 61643 1054 61655 1430
rect 61689 1054 61701 1430
rect 61643 1042 61701 1054
rect 61761 1430 61819 1442
rect 61761 1054 61773 1430
rect 61807 1054 61819 1430
rect 61761 1042 61819 1054
rect 61879 1430 61937 1442
rect 61879 1054 61891 1430
rect 61925 1054 61937 1430
rect 61879 1042 61937 1054
rect 61997 1430 62055 1442
rect 61997 1054 62009 1430
rect 62043 1054 62055 1430
rect 61997 1042 62055 1054
rect 62115 1430 62173 1442
rect 62115 1054 62127 1430
rect 62161 1054 62173 1430
rect 62115 1042 62173 1054
rect 70509 1428 70909 1440
rect 63477 1396 63535 1408
rect 63477 1220 63489 1396
rect 63523 1220 63535 1396
rect 63477 1208 63535 1220
rect 63595 1396 63653 1408
rect 63595 1220 63607 1396
rect 63641 1220 63653 1396
rect 63595 1208 63653 1220
rect 63713 1396 63771 1408
rect 63713 1220 63725 1396
rect 63759 1220 63771 1396
rect 63713 1208 63771 1220
rect 63831 1396 63889 1408
rect 63831 1220 63843 1396
rect 63877 1220 63889 1396
rect 63831 1208 63889 1220
rect 63949 1396 64007 1408
rect 63949 1220 63961 1396
rect 63995 1220 64007 1396
rect 63949 1208 64007 1220
rect 64067 1396 64125 1408
rect 64067 1220 64079 1396
rect 64113 1220 64125 1396
rect 64067 1208 64125 1220
rect 64185 1396 64243 1408
rect 64185 1220 64197 1396
rect 64231 1220 64243 1396
rect 64185 1208 64243 1220
rect 64303 1396 64361 1408
rect 64303 1220 64315 1396
rect 64349 1220 64361 1396
rect 64303 1208 64361 1220
rect 64421 1396 64479 1408
rect 64421 1220 64433 1396
rect 64467 1220 64479 1396
rect 64421 1208 64479 1220
rect 64539 1396 64597 1408
rect 64539 1220 64551 1396
rect 64585 1220 64597 1396
rect 70509 1394 70521 1428
rect 70897 1394 70909 1428
rect 70509 1382 70909 1394
rect 64539 1208 64597 1220
rect 70509 1310 70909 1322
rect 70509 1276 70521 1310
rect 70897 1276 70909 1310
rect 70509 1264 70909 1276
rect 70509 1192 70909 1204
rect 70509 1158 70521 1192
rect 70897 1158 70909 1192
rect 70509 1146 70909 1158
rect 70509 1074 70909 1086
rect 70509 1040 70521 1074
rect 70897 1040 70909 1074
rect 70509 1028 70909 1040
rect 70709 955 70909 967
rect 70709 921 70721 955
rect 70897 921 70909 955
rect 70709 909 70909 921
rect 70709 837 70909 849
rect 70709 803 70721 837
rect 70897 803 70909 837
rect 70709 791 70909 803
rect 70709 719 70909 731
rect 70709 685 70721 719
rect 70897 685 70909 719
rect 70709 673 70909 685
rect 70709 601 70909 613
rect 70709 567 70721 601
rect 70897 567 70909 601
rect 70709 555 70909 567
rect 70709 19 70909 31
rect 70709 -15 70721 19
rect 70897 -15 70909 19
rect 70709 -27 70909 -15
rect 65708 -149 65766 -137
rect 30645 -260 31045 -248
rect 30645 -294 30657 -260
rect 31033 -294 31045 -260
rect 30645 -306 31045 -294
rect 29952 -435 30352 -423
rect 29952 -469 29964 -435
rect 30340 -469 30352 -435
rect 29952 -481 30352 -469
rect 30152 -564 30352 -552
rect 30152 -598 30164 -564
rect 30340 -598 30352 -564
rect 30152 -610 30352 -598
rect 30645 -378 31045 -366
rect 30645 -412 30657 -378
rect 31033 -412 31045 -378
rect 65224 -349 65282 -337
rect 30645 -424 31045 -412
rect 65224 -525 65236 -349
rect 65270 -525 65282 -349
rect 65224 -537 65282 -525
rect 65342 -349 65400 -337
rect 65342 -525 65354 -349
rect 65388 -525 65400 -349
rect 65342 -537 65400 -525
rect 65460 -349 65518 -337
rect 65460 -525 65472 -349
rect 65506 -525 65518 -349
rect 65460 -537 65518 -525
rect 65578 -349 65636 -337
rect 65578 -525 65590 -349
rect 65624 -525 65636 -349
rect 65578 -537 65636 -525
rect 65708 -525 65720 -149
rect 65754 -525 65766 -149
rect 65708 -537 65766 -525
rect 65826 -149 65884 -137
rect 65826 -525 65838 -149
rect 65872 -525 65884 -149
rect 65826 -537 65884 -525
rect 65944 -149 66002 -137
rect 65944 -525 65956 -149
rect 65990 -525 66002 -149
rect 65944 -537 66002 -525
rect 66062 -149 66120 -137
rect 66062 -525 66074 -149
rect 66108 -525 66120 -149
rect 66062 -537 66120 -525
rect 66180 -149 66238 -137
rect 66180 -525 66192 -149
rect 66226 -525 66238 -149
rect 66180 -537 66238 -525
rect 66298 -149 66356 -137
rect 66298 -525 66310 -149
rect 66344 -525 66356 -149
rect 66298 -537 66356 -525
rect 66416 -149 66474 -137
rect 66416 -525 66428 -149
rect 66462 -525 66474 -149
rect 70709 -99 70909 -87
rect 70709 -133 70721 -99
rect 70897 -133 70909 -99
rect 70709 -145 70909 -133
rect 70709 -217 70909 -205
rect 70709 -251 70721 -217
rect 70897 -251 70909 -217
rect 70709 -263 70909 -251
rect 66416 -537 66474 -525
rect 66545 -349 66603 -337
rect 66545 -525 66557 -349
rect 66591 -525 66603 -349
rect 66545 -537 66603 -525
rect 66663 -349 66721 -337
rect 66663 -525 66675 -349
rect 66709 -525 66721 -349
rect 66663 -537 66721 -525
rect 66781 -349 66839 -337
rect 66781 -525 66793 -349
rect 66827 -525 66839 -349
rect 66781 -537 66839 -525
rect 66899 -349 66957 -337
rect 70709 -335 70909 -323
rect 66899 -525 66911 -349
rect 66945 -525 66957 -349
rect 66899 -537 66957 -525
rect 67017 -352 67075 -340
rect 67017 -528 67029 -352
rect 67063 -528 67075 -352
rect 30152 -682 30352 -670
rect 30152 -716 30164 -682
rect 30340 -716 30352 -682
rect 30152 -728 30352 -716
rect 30152 -800 30352 -788
rect 30152 -834 30164 -800
rect 30340 -834 30352 -800
rect 67017 -540 67075 -528
rect 67135 -352 67193 -340
rect 67135 -528 67147 -352
rect 67181 -528 67193 -352
rect 67135 -540 67193 -528
rect 67253 -352 67311 -340
rect 67253 -528 67265 -352
rect 67299 -528 67311 -352
rect 67253 -540 67311 -528
rect 67371 -352 67429 -340
rect 67371 -528 67383 -352
rect 67417 -528 67429 -352
rect 67371 -540 67429 -528
rect 67489 -352 67547 -340
rect 67489 -528 67501 -352
rect 67535 -528 67547 -352
rect 67489 -540 67547 -528
rect 67607 -352 67665 -340
rect 67607 -528 67619 -352
rect 67653 -528 67665 -352
rect 67607 -540 67665 -528
rect 67725 -352 67783 -340
rect 67725 -528 67737 -352
rect 67771 -528 67783 -352
rect 67725 -540 67783 -528
rect 67843 -352 67901 -340
rect 67843 -528 67855 -352
rect 67889 -528 67901 -352
rect 67843 -540 67901 -528
rect 67961 -352 68019 -340
rect 67961 -528 67973 -352
rect 68007 -528 68019 -352
rect 67961 -540 68019 -528
rect 68079 -352 68137 -340
rect 68079 -528 68091 -352
rect 68125 -528 68137 -352
rect 70709 -369 70721 -335
rect 70897 -369 70909 -335
rect 70709 -410 70909 -369
rect 70509 -422 70909 -410
rect 70509 -456 70521 -422
rect 70897 -456 70909 -422
rect 70509 -468 70909 -456
rect 68079 -540 68137 -528
rect 30152 -846 30352 -834
rect 30152 -918 30352 -906
rect 65651 -842 65709 -830
rect 30152 -952 30164 -918
rect 30340 -952 30352 -918
rect 30152 -964 30352 -952
rect 30150 -1311 30350 -1299
rect 30150 -1345 30162 -1311
rect 30338 -1345 30350 -1311
rect 30150 -1357 30350 -1345
rect 30150 -1429 30350 -1417
rect 30150 -1463 30162 -1429
rect 30338 -1463 30350 -1429
rect 30150 -1475 30350 -1463
rect 30150 -1547 30350 -1535
rect 30150 -1581 30162 -1547
rect 30338 -1581 30350 -1547
rect 30150 -1593 30350 -1581
rect 63484 -1449 63542 -1437
rect 41593 -1567 41651 -1555
rect 30150 -1665 30350 -1653
rect 721 -1764 779 -1752
rect 721 -1952 733 -1764
rect 280 -1964 338 -1952
rect 280 -2140 292 -1964
rect 326 -2140 338 -1964
rect 280 -2152 338 -2140
rect 398 -1964 456 -1952
rect 398 -2140 410 -1964
rect 444 -2140 456 -1964
rect 398 -2152 456 -2140
rect 516 -1964 574 -1952
rect 516 -2140 528 -1964
rect 562 -2140 574 -1964
rect 516 -2152 574 -2140
rect 634 -1964 733 -1952
rect 634 -2140 646 -1964
rect 680 -2140 733 -1964
rect 767 -2140 779 -1764
rect 634 -2152 779 -2140
rect 839 -1764 897 -1752
rect 839 -2140 851 -1764
rect 885 -2140 897 -1764
rect 839 -2152 897 -2140
rect 957 -1764 1015 -1752
rect 957 -2140 969 -1764
rect 1003 -2140 1015 -1764
rect 957 -2152 1015 -2140
rect 1075 -1764 1133 -1752
rect 1075 -2140 1087 -1764
rect 1121 -2140 1133 -1764
rect 1075 -2152 1133 -2140
rect 1188 -1764 1246 -1752
rect 1188 -2140 1200 -1764
rect 1234 -2140 1246 -1764
rect 1188 -2152 1246 -2140
rect 1306 -1764 1364 -1752
rect 1306 -2140 1318 -1764
rect 1352 -2140 1364 -1764
rect 1306 -2152 1364 -2140
rect 1424 -1764 1482 -1752
rect 1424 -2140 1436 -1764
rect 1470 -2140 1482 -1764
rect 1424 -2152 1482 -2140
rect 1542 -1764 1600 -1752
rect 1542 -2140 1554 -1764
rect 1588 -2140 1600 -1764
rect 1542 -2152 1600 -2140
rect 1660 -1764 1718 -1752
rect 1660 -2140 1672 -1764
rect 1706 -2140 1718 -1764
rect 1660 -2152 1718 -2140
rect 1778 -1764 1836 -1752
rect 1778 -2140 1790 -1764
rect 1824 -2140 1836 -1764
rect 1778 -2152 1836 -2140
rect 1896 -1764 1954 -1752
rect 1896 -2140 1908 -1764
rect 1942 -2140 1954 -1764
rect 1896 -2152 1954 -2140
rect 2015 -1764 2073 -1752
rect 2015 -2140 2027 -1764
rect 2061 -2140 2073 -1764
rect 2015 -2152 2073 -2140
rect 2133 -1764 2191 -1752
rect 2133 -2140 2145 -1764
rect 2179 -2140 2191 -1764
rect 2133 -2152 2191 -2140
rect 2251 -1764 2309 -1752
rect 2251 -2140 2263 -1764
rect 2297 -2140 2309 -1764
rect 2251 -2152 2309 -2140
rect 2369 -1764 2427 -1752
rect 2369 -2140 2381 -1764
rect 2415 -2140 2427 -1764
rect 3865 -1764 3923 -1752
rect 3865 -1952 3877 -1764
rect 2369 -2152 2427 -2140
rect 2488 -1964 2546 -1952
rect 2488 -2140 2500 -1964
rect 2534 -2140 2546 -1964
rect 2488 -2152 2546 -2140
rect 2606 -1964 2664 -1952
rect 2606 -2140 2618 -1964
rect 2652 -2140 2664 -1964
rect 2606 -2152 2664 -2140
rect 2724 -1964 2782 -1952
rect 2724 -2140 2736 -1964
rect 2770 -2140 2782 -1964
rect 2724 -2152 2782 -2140
rect 2842 -1964 2900 -1952
rect 2842 -2140 2854 -1964
rect 2888 -2140 2900 -1964
rect 2842 -2152 2900 -2140
rect 3424 -1964 3482 -1952
rect 3424 -2140 3436 -1964
rect 3470 -2140 3482 -1964
rect 3424 -2152 3482 -2140
rect 3542 -1964 3600 -1952
rect 3542 -2140 3554 -1964
rect 3588 -2140 3600 -1964
rect 3542 -2152 3600 -2140
rect 3660 -1964 3718 -1952
rect 3660 -2140 3672 -1964
rect 3706 -2140 3718 -1964
rect 3660 -2152 3718 -2140
rect 3778 -1964 3877 -1952
rect 3778 -2140 3790 -1964
rect 3824 -2140 3877 -1964
rect 3911 -2140 3923 -1764
rect 3778 -2152 3923 -2140
rect 3983 -1764 4041 -1752
rect 3983 -2140 3995 -1764
rect 4029 -2140 4041 -1764
rect 3983 -2152 4041 -2140
rect 4101 -1764 4159 -1752
rect 4101 -2140 4113 -1764
rect 4147 -2140 4159 -1764
rect 4101 -2152 4159 -2140
rect 4219 -1764 4277 -1752
rect 4219 -2140 4231 -1764
rect 4265 -2140 4277 -1764
rect 4219 -2152 4277 -2140
rect 4332 -1764 4390 -1752
rect 4332 -2140 4344 -1764
rect 4378 -2140 4390 -1764
rect 4332 -2152 4390 -2140
rect 4450 -1764 4508 -1752
rect 4450 -2140 4462 -1764
rect 4496 -2140 4508 -1764
rect 4450 -2152 4508 -2140
rect 4568 -1764 4626 -1752
rect 4568 -2140 4580 -1764
rect 4614 -2140 4626 -1764
rect 4568 -2152 4626 -2140
rect 4686 -1764 4744 -1752
rect 4686 -2140 4698 -1764
rect 4732 -2140 4744 -1764
rect 4686 -2152 4744 -2140
rect 4804 -1764 4862 -1752
rect 4804 -2140 4816 -1764
rect 4850 -2140 4862 -1764
rect 4804 -2152 4862 -2140
rect 4922 -1764 4980 -1752
rect 4922 -2140 4934 -1764
rect 4968 -2140 4980 -1764
rect 4922 -2152 4980 -2140
rect 5040 -1764 5098 -1752
rect 5040 -2140 5052 -1764
rect 5086 -2140 5098 -1764
rect 5040 -2152 5098 -2140
rect 5159 -1764 5217 -1752
rect 5159 -2140 5171 -1764
rect 5205 -2140 5217 -1764
rect 5159 -2152 5217 -2140
rect 5277 -1764 5335 -1752
rect 5277 -2140 5289 -1764
rect 5323 -2140 5335 -1764
rect 5277 -2152 5335 -2140
rect 5395 -1764 5453 -1752
rect 5395 -2140 5407 -1764
rect 5441 -2140 5453 -1764
rect 5395 -2152 5453 -2140
rect 5513 -1764 5571 -1752
rect 5513 -2140 5525 -1764
rect 5559 -2140 5571 -1764
rect 6997 -1760 7055 -1748
rect 6997 -1948 7009 -1760
rect 5513 -2152 5571 -2140
rect 5632 -1964 5690 -1952
rect 5632 -2140 5644 -1964
rect 5678 -2140 5690 -1964
rect 5632 -2152 5690 -2140
rect 5750 -1964 5808 -1952
rect 5750 -2140 5762 -1964
rect 5796 -2140 5808 -1964
rect 5750 -2152 5808 -2140
rect 5868 -1964 5926 -1952
rect 5868 -2140 5880 -1964
rect 5914 -2140 5926 -1964
rect 5868 -2152 5926 -2140
rect 5986 -1964 6044 -1952
rect 5986 -2140 5998 -1964
rect 6032 -2140 6044 -1964
rect 5986 -2152 6044 -2140
rect 6556 -1960 6614 -1948
rect 6556 -2136 6568 -1960
rect 6602 -2136 6614 -1960
rect 6556 -2148 6614 -2136
rect 6674 -1960 6732 -1948
rect 6674 -2136 6686 -1960
rect 6720 -2136 6732 -1960
rect 6674 -2148 6732 -2136
rect 6792 -1960 6850 -1948
rect 6792 -2136 6804 -1960
rect 6838 -2136 6850 -1960
rect 6792 -2148 6850 -2136
rect 6910 -1960 7009 -1948
rect 6910 -2136 6922 -1960
rect 6956 -2136 7009 -1960
rect 7043 -2136 7055 -1760
rect 6910 -2148 7055 -2136
rect 7115 -1760 7173 -1748
rect 7115 -2136 7127 -1760
rect 7161 -2136 7173 -1760
rect 7115 -2148 7173 -2136
rect 7233 -1760 7291 -1748
rect 7233 -2136 7245 -1760
rect 7279 -2136 7291 -1760
rect 7233 -2148 7291 -2136
rect 7351 -1760 7409 -1748
rect 7351 -2136 7363 -1760
rect 7397 -2136 7409 -1760
rect 7351 -2148 7409 -2136
rect 7464 -1760 7522 -1748
rect 7464 -2136 7476 -1760
rect 7510 -2136 7522 -1760
rect 7464 -2148 7522 -2136
rect 7582 -1760 7640 -1748
rect 7582 -2136 7594 -1760
rect 7628 -2136 7640 -1760
rect 7582 -2148 7640 -2136
rect 7700 -1760 7758 -1748
rect 7700 -2136 7712 -1760
rect 7746 -2136 7758 -1760
rect 7700 -2148 7758 -2136
rect 7818 -1760 7876 -1748
rect 7818 -2136 7830 -1760
rect 7864 -2136 7876 -1760
rect 7818 -2148 7876 -2136
rect 7936 -1760 7994 -1748
rect 7936 -2136 7948 -1760
rect 7982 -2136 7994 -1760
rect 7936 -2148 7994 -2136
rect 8054 -1760 8112 -1748
rect 8054 -2136 8066 -1760
rect 8100 -2136 8112 -1760
rect 8054 -2148 8112 -2136
rect 8172 -1760 8230 -1748
rect 8172 -2136 8184 -1760
rect 8218 -2136 8230 -1760
rect 8172 -2148 8230 -2136
rect 8291 -1760 8349 -1748
rect 8291 -2136 8303 -1760
rect 8337 -2136 8349 -1760
rect 8291 -2148 8349 -2136
rect 8409 -1760 8467 -1748
rect 8409 -2136 8421 -1760
rect 8455 -2136 8467 -1760
rect 8409 -2148 8467 -2136
rect 8527 -1760 8585 -1748
rect 8527 -2136 8539 -1760
rect 8573 -2136 8585 -1760
rect 8527 -2148 8585 -2136
rect 8645 -1760 8703 -1748
rect 8645 -2136 8657 -1760
rect 8691 -2136 8703 -1760
rect 10141 -1760 10199 -1748
rect 10141 -1948 10153 -1760
rect 8645 -2148 8703 -2136
rect 8764 -1960 8822 -1948
rect 8764 -2136 8776 -1960
rect 8810 -2136 8822 -1960
rect 8764 -2148 8822 -2136
rect 8882 -1960 8940 -1948
rect 8882 -2136 8894 -1960
rect 8928 -2136 8940 -1960
rect 8882 -2148 8940 -2136
rect 9000 -1960 9058 -1948
rect 9000 -2136 9012 -1960
rect 9046 -2136 9058 -1960
rect 9000 -2148 9058 -2136
rect 9118 -1960 9176 -1948
rect 9118 -2136 9130 -1960
rect 9164 -2136 9176 -1960
rect 9118 -2148 9176 -2136
rect 9700 -1960 9758 -1948
rect 9700 -2136 9712 -1960
rect 9746 -2136 9758 -1960
rect 9700 -2148 9758 -2136
rect 9818 -1960 9876 -1948
rect 9818 -2136 9830 -1960
rect 9864 -2136 9876 -1960
rect 9818 -2148 9876 -2136
rect 9936 -1960 9994 -1948
rect 9936 -2136 9948 -1960
rect 9982 -2136 9994 -1960
rect 9936 -2148 9994 -2136
rect 10054 -1960 10153 -1948
rect 10054 -2136 10066 -1960
rect 10100 -2136 10153 -1960
rect 10187 -2136 10199 -1760
rect 10054 -2148 10199 -2136
rect 10259 -1760 10317 -1748
rect 10259 -2136 10271 -1760
rect 10305 -2136 10317 -1760
rect 10259 -2148 10317 -2136
rect 10377 -1760 10435 -1748
rect 10377 -2136 10389 -1760
rect 10423 -2136 10435 -1760
rect 10377 -2148 10435 -2136
rect 10495 -1760 10553 -1748
rect 10495 -2136 10507 -1760
rect 10541 -2136 10553 -1760
rect 10495 -2148 10553 -2136
rect 10608 -1760 10666 -1748
rect 10608 -2136 10620 -1760
rect 10654 -2136 10666 -1760
rect 10608 -2148 10666 -2136
rect 10726 -1760 10784 -1748
rect 10726 -2136 10738 -1760
rect 10772 -2136 10784 -1760
rect 10726 -2148 10784 -2136
rect 10844 -1760 10902 -1748
rect 10844 -2136 10856 -1760
rect 10890 -2136 10902 -1760
rect 10844 -2148 10902 -2136
rect 10962 -1760 11020 -1748
rect 10962 -2136 10974 -1760
rect 11008 -2136 11020 -1760
rect 10962 -2148 11020 -2136
rect 11080 -1760 11138 -1748
rect 11080 -2136 11092 -1760
rect 11126 -2136 11138 -1760
rect 11080 -2148 11138 -2136
rect 11198 -1760 11256 -1748
rect 11198 -2136 11210 -1760
rect 11244 -2136 11256 -1760
rect 11198 -2148 11256 -2136
rect 11316 -1760 11374 -1748
rect 11316 -2136 11328 -1760
rect 11362 -2136 11374 -1760
rect 11316 -2148 11374 -2136
rect 11435 -1760 11493 -1748
rect 11435 -2136 11447 -1760
rect 11481 -2136 11493 -1760
rect 11435 -2148 11493 -2136
rect 11553 -1760 11611 -1748
rect 11553 -2136 11565 -1760
rect 11599 -2136 11611 -1760
rect 11553 -2148 11611 -2136
rect 11671 -1760 11729 -1748
rect 11671 -2136 11683 -1760
rect 11717 -2136 11729 -1760
rect 11671 -2148 11729 -2136
rect 11789 -1760 11847 -1748
rect 30150 -1699 30162 -1665
rect 30338 -1699 30350 -1665
rect 30150 -1711 30350 -1699
rect 11789 -2136 11801 -1760
rect 11835 -2136 11847 -1760
rect 13343 -1764 13401 -1752
rect 11789 -2148 11847 -2136
rect 11908 -1960 11966 -1948
rect 11908 -2136 11920 -1960
rect 11954 -2136 11966 -1960
rect 11908 -2148 11966 -2136
rect 12026 -1960 12084 -1948
rect 12026 -2136 12038 -1960
rect 12072 -2136 12084 -1960
rect 12026 -2148 12084 -2136
rect 12144 -1960 12202 -1948
rect 12144 -2136 12156 -1960
rect 12190 -2136 12202 -1960
rect 12144 -2148 12202 -2136
rect 12262 -1960 12320 -1948
rect 13343 -1952 13355 -1764
rect 12262 -2136 12274 -1960
rect 12308 -2136 12320 -1960
rect 12262 -2148 12320 -2136
rect 12902 -1964 12960 -1952
rect 12902 -2140 12914 -1964
rect 12948 -2140 12960 -1964
rect 12902 -2152 12960 -2140
rect 13020 -1964 13078 -1952
rect 13020 -2140 13032 -1964
rect 13066 -2140 13078 -1964
rect 13020 -2152 13078 -2140
rect 13138 -1964 13196 -1952
rect 13138 -2140 13150 -1964
rect 13184 -2140 13196 -1964
rect 13138 -2152 13196 -2140
rect 13256 -1964 13355 -1952
rect 13256 -2140 13268 -1964
rect 13302 -2140 13355 -1964
rect 13389 -2140 13401 -1764
rect 13256 -2152 13401 -2140
rect 13461 -1764 13519 -1752
rect 13461 -2140 13473 -1764
rect 13507 -2140 13519 -1764
rect 13461 -2152 13519 -2140
rect 13579 -1764 13637 -1752
rect 13579 -2140 13591 -1764
rect 13625 -2140 13637 -1764
rect 13579 -2152 13637 -2140
rect 13697 -1764 13755 -1752
rect 13697 -2140 13709 -1764
rect 13743 -2140 13755 -1764
rect 13697 -2152 13755 -2140
rect 13810 -1764 13868 -1752
rect 13810 -2140 13822 -1764
rect 13856 -2140 13868 -1764
rect 13810 -2152 13868 -2140
rect 13928 -1764 13986 -1752
rect 13928 -2140 13940 -1764
rect 13974 -2140 13986 -1764
rect 13928 -2152 13986 -2140
rect 14046 -1764 14104 -1752
rect 14046 -2140 14058 -1764
rect 14092 -2140 14104 -1764
rect 14046 -2152 14104 -2140
rect 14164 -1764 14222 -1752
rect 14164 -2140 14176 -1764
rect 14210 -2140 14222 -1764
rect 14164 -2152 14222 -2140
rect 14282 -1764 14340 -1752
rect 14282 -2140 14294 -1764
rect 14328 -2140 14340 -1764
rect 14282 -2152 14340 -2140
rect 14400 -1764 14458 -1752
rect 14400 -2140 14412 -1764
rect 14446 -2140 14458 -1764
rect 14400 -2152 14458 -2140
rect 14518 -1764 14576 -1752
rect 14518 -2140 14530 -1764
rect 14564 -2140 14576 -1764
rect 14518 -2152 14576 -2140
rect 14637 -1764 14695 -1752
rect 14637 -2140 14649 -1764
rect 14683 -2140 14695 -1764
rect 14637 -2152 14695 -2140
rect 14755 -1764 14813 -1752
rect 14755 -2140 14767 -1764
rect 14801 -2140 14813 -1764
rect 14755 -2152 14813 -2140
rect 14873 -1764 14931 -1752
rect 14873 -2140 14885 -1764
rect 14919 -2140 14931 -1764
rect 14873 -2152 14931 -2140
rect 14991 -1764 15049 -1752
rect 14991 -2140 15003 -1764
rect 15037 -2140 15049 -1764
rect 16487 -1764 16545 -1752
rect 16487 -1952 16499 -1764
rect 14991 -2152 15049 -2140
rect 15110 -1964 15168 -1952
rect 15110 -2140 15122 -1964
rect 15156 -2140 15168 -1964
rect 15110 -2152 15168 -2140
rect 15228 -1964 15286 -1952
rect 15228 -2140 15240 -1964
rect 15274 -2140 15286 -1964
rect 15228 -2152 15286 -2140
rect 15346 -1964 15404 -1952
rect 15346 -2140 15358 -1964
rect 15392 -2140 15404 -1964
rect 15346 -2152 15404 -2140
rect 15464 -1964 15522 -1952
rect 15464 -2140 15476 -1964
rect 15510 -2140 15522 -1964
rect 15464 -2152 15522 -2140
rect 16046 -1964 16104 -1952
rect 16046 -2140 16058 -1964
rect 16092 -2140 16104 -1964
rect 16046 -2152 16104 -2140
rect 16164 -1964 16222 -1952
rect 16164 -2140 16176 -1964
rect 16210 -2140 16222 -1964
rect 16164 -2152 16222 -2140
rect 16282 -1964 16340 -1952
rect 16282 -2140 16294 -1964
rect 16328 -2140 16340 -1964
rect 16282 -2152 16340 -2140
rect 16400 -1964 16499 -1952
rect 16400 -2140 16412 -1964
rect 16446 -2140 16499 -1964
rect 16533 -2140 16545 -1764
rect 16400 -2152 16545 -2140
rect 16605 -1764 16663 -1752
rect 16605 -2140 16617 -1764
rect 16651 -2140 16663 -1764
rect 16605 -2152 16663 -2140
rect 16723 -1764 16781 -1752
rect 16723 -2140 16735 -1764
rect 16769 -2140 16781 -1764
rect 16723 -2152 16781 -2140
rect 16841 -1764 16899 -1752
rect 16841 -2140 16853 -1764
rect 16887 -2140 16899 -1764
rect 16841 -2152 16899 -2140
rect 16954 -1764 17012 -1752
rect 16954 -2140 16966 -1764
rect 17000 -2140 17012 -1764
rect 16954 -2152 17012 -2140
rect 17072 -1764 17130 -1752
rect 17072 -2140 17084 -1764
rect 17118 -2140 17130 -1764
rect 17072 -2152 17130 -2140
rect 17190 -1764 17248 -1752
rect 17190 -2140 17202 -1764
rect 17236 -2140 17248 -1764
rect 17190 -2152 17248 -2140
rect 17308 -1764 17366 -1752
rect 17308 -2140 17320 -1764
rect 17354 -2140 17366 -1764
rect 17308 -2152 17366 -2140
rect 17426 -1764 17484 -1752
rect 17426 -2140 17438 -1764
rect 17472 -2140 17484 -1764
rect 17426 -2152 17484 -2140
rect 17544 -1764 17602 -1752
rect 17544 -2140 17556 -1764
rect 17590 -2140 17602 -1764
rect 17544 -2152 17602 -2140
rect 17662 -1764 17720 -1752
rect 17662 -2140 17674 -1764
rect 17708 -2140 17720 -1764
rect 17662 -2152 17720 -2140
rect 17781 -1764 17839 -1752
rect 17781 -2140 17793 -1764
rect 17827 -2140 17839 -1764
rect 17781 -2152 17839 -2140
rect 17899 -1764 17957 -1752
rect 17899 -2140 17911 -1764
rect 17945 -2140 17957 -1764
rect 17899 -2152 17957 -2140
rect 18017 -1764 18075 -1752
rect 18017 -2140 18029 -1764
rect 18063 -2140 18075 -1764
rect 18017 -2152 18075 -2140
rect 18135 -1764 18193 -1752
rect 18135 -2140 18147 -1764
rect 18181 -2140 18193 -1764
rect 19619 -1760 19677 -1748
rect 19619 -1948 19631 -1760
rect 18135 -2152 18193 -2140
rect 18254 -1964 18312 -1952
rect 18254 -2140 18266 -1964
rect 18300 -2140 18312 -1964
rect 18254 -2152 18312 -2140
rect 18372 -1964 18430 -1952
rect 18372 -2140 18384 -1964
rect 18418 -2140 18430 -1964
rect 18372 -2152 18430 -2140
rect 18490 -1964 18548 -1952
rect 18490 -2140 18502 -1964
rect 18536 -2140 18548 -1964
rect 18490 -2152 18548 -2140
rect 18608 -1964 18666 -1952
rect 18608 -2140 18620 -1964
rect 18654 -2140 18666 -1964
rect 18608 -2152 18666 -2140
rect 19178 -1960 19236 -1948
rect 19178 -2136 19190 -1960
rect 19224 -2136 19236 -1960
rect 19178 -2148 19236 -2136
rect 19296 -1960 19354 -1948
rect 19296 -2136 19308 -1960
rect 19342 -2136 19354 -1960
rect 19296 -2148 19354 -2136
rect 19414 -1960 19472 -1948
rect 19414 -2136 19426 -1960
rect 19460 -2136 19472 -1960
rect 19414 -2148 19472 -2136
rect 19532 -1960 19631 -1948
rect 19532 -2136 19544 -1960
rect 19578 -2136 19631 -1960
rect 19665 -2136 19677 -1760
rect 19532 -2148 19677 -2136
rect 19737 -1760 19795 -1748
rect 19737 -2136 19749 -1760
rect 19783 -2136 19795 -1760
rect 19737 -2148 19795 -2136
rect 19855 -1760 19913 -1748
rect 19855 -2136 19867 -1760
rect 19901 -2136 19913 -1760
rect 19855 -2148 19913 -2136
rect 19973 -1760 20031 -1748
rect 19973 -2136 19985 -1760
rect 20019 -2136 20031 -1760
rect 19973 -2148 20031 -2136
rect 20086 -1760 20144 -1748
rect 20086 -2136 20098 -1760
rect 20132 -2136 20144 -1760
rect 20086 -2148 20144 -2136
rect 20204 -1760 20262 -1748
rect 20204 -2136 20216 -1760
rect 20250 -2136 20262 -1760
rect 20204 -2148 20262 -2136
rect 20322 -1760 20380 -1748
rect 20322 -2136 20334 -1760
rect 20368 -2136 20380 -1760
rect 20322 -2148 20380 -2136
rect 20440 -1760 20498 -1748
rect 20440 -2136 20452 -1760
rect 20486 -2136 20498 -1760
rect 20440 -2148 20498 -2136
rect 20558 -1760 20616 -1748
rect 20558 -2136 20570 -1760
rect 20604 -2136 20616 -1760
rect 20558 -2148 20616 -2136
rect 20676 -1760 20734 -1748
rect 20676 -2136 20688 -1760
rect 20722 -2136 20734 -1760
rect 20676 -2148 20734 -2136
rect 20794 -1760 20852 -1748
rect 20794 -2136 20806 -1760
rect 20840 -2136 20852 -1760
rect 20794 -2148 20852 -2136
rect 20913 -1760 20971 -1748
rect 20913 -2136 20925 -1760
rect 20959 -2136 20971 -1760
rect 20913 -2148 20971 -2136
rect 21031 -1760 21089 -1748
rect 21031 -2136 21043 -1760
rect 21077 -2136 21089 -1760
rect 21031 -2148 21089 -2136
rect 21149 -1760 21207 -1748
rect 21149 -2136 21161 -1760
rect 21195 -2136 21207 -1760
rect 21149 -2148 21207 -2136
rect 21267 -1760 21325 -1748
rect 21267 -2136 21279 -1760
rect 21313 -2136 21325 -1760
rect 22763 -1760 22821 -1748
rect 22763 -1948 22775 -1760
rect 21267 -2148 21325 -2136
rect 21386 -1960 21444 -1948
rect 21386 -2136 21398 -1960
rect 21432 -2136 21444 -1960
rect 21386 -2148 21444 -2136
rect 21504 -1960 21562 -1948
rect 21504 -2136 21516 -1960
rect 21550 -2136 21562 -1960
rect 21504 -2148 21562 -2136
rect 21622 -1960 21680 -1948
rect 21622 -2136 21634 -1960
rect 21668 -2136 21680 -1960
rect 21622 -2148 21680 -2136
rect 21740 -1960 21798 -1948
rect 21740 -2136 21752 -1960
rect 21786 -2136 21798 -1960
rect 21740 -2148 21798 -2136
rect 22322 -1960 22380 -1948
rect 22322 -2136 22334 -1960
rect 22368 -2136 22380 -1960
rect 22322 -2148 22380 -2136
rect 22440 -1960 22498 -1948
rect 22440 -2136 22452 -1960
rect 22486 -2136 22498 -1960
rect 22440 -2148 22498 -2136
rect 22558 -1960 22616 -1948
rect 22558 -2136 22570 -1960
rect 22604 -2136 22616 -1960
rect 22558 -2148 22616 -2136
rect 22676 -1960 22775 -1948
rect 22676 -2136 22688 -1960
rect 22722 -2136 22775 -1960
rect 22809 -2136 22821 -1760
rect 22676 -2148 22821 -2136
rect 22881 -1760 22939 -1748
rect 22881 -2136 22893 -1760
rect 22927 -2136 22939 -1760
rect 22881 -2148 22939 -2136
rect 22999 -1760 23057 -1748
rect 22999 -2136 23011 -1760
rect 23045 -2136 23057 -1760
rect 22999 -2148 23057 -2136
rect 23117 -1760 23175 -1748
rect 23117 -2136 23129 -1760
rect 23163 -2136 23175 -1760
rect 23117 -2148 23175 -2136
rect 23230 -1760 23288 -1748
rect 23230 -2136 23242 -1760
rect 23276 -2136 23288 -1760
rect 23230 -2148 23288 -2136
rect 23348 -1760 23406 -1748
rect 23348 -2136 23360 -1760
rect 23394 -2136 23406 -1760
rect 23348 -2148 23406 -2136
rect 23466 -1760 23524 -1748
rect 23466 -2136 23478 -1760
rect 23512 -2136 23524 -1760
rect 23466 -2148 23524 -2136
rect 23584 -1760 23642 -1748
rect 23584 -2136 23596 -1760
rect 23630 -2136 23642 -1760
rect 23584 -2148 23642 -2136
rect 23702 -1760 23760 -1748
rect 23702 -2136 23714 -1760
rect 23748 -2136 23760 -1760
rect 23702 -2148 23760 -2136
rect 23820 -1760 23878 -1748
rect 23820 -2136 23832 -1760
rect 23866 -2136 23878 -1760
rect 23820 -2148 23878 -2136
rect 23938 -1760 23996 -1748
rect 23938 -2136 23950 -1760
rect 23984 -2136 23996 -1760
rect 23938 -2148 23996 -2136
rect 24057 -1760 24115 -1748
rect 24057 -2136 24069 -1760
rect 24103 -2136 24115 -1760
rect 24057 -2148 24115 -2136
rect 24175 -1760 24233 -1748
rect 24175 -2136 24187 -1760
rect 24221 -2136 24233 -1760
rect 24175 -2148 24233 -2136
rect 24293 -1760 24351 -1748
rect 24293 -2136 24305 -1760
rect 24339 -2136 24351 -1760
rect 24293 -2148 24351 -2136
rect 24411 -1760 24469 -1748
rect 24411 -2136 24423 -1760
rect 24457 -2136 24469 -1760
rect 29950 -1795 30350 -1783
rect 29950 -1829 29962 -1795
rect 30338 -1829 30350 -1795
rect 29950 -1841 30350 -1829
rect 30643 -1738 31043 -1726
rect 30643 -1772 30655 -1738
rect 31031 -1772 31043 -1738
rect 41593 -1743 41605 -1567
rect 41639 -1743 41651 -1567
rect 30643 -1784 31043 -1772
rect 41593 -1755 41651 -1743
rect 41711 -1567 41769 -1555
rect 41711 -1743 41723 -1567
rect 41757 -1743 41769 -1567
rect 41711 -1755 41769 -1743
rect 41829 -1567 41887 -1555
rect 41829 -1743 41841 -1567
rect 41875 -1743 41887 -1567
rect 41829 -1755 41887 -1743
rect 41947 -1567 42005 -1555
rect 41947 -1743 41959 -1567
rect 41993 -1743 42005 -1567
rect 41947 -1755 42005 -1743
rect 42065 -1567 42123 -1555
rect 42065 -1743 42077 -1567
rect 42111 -1743 42123 -1567
rect 42065 -1755 42123 -1743
rect 42183 -1567 42241 -1555
rect 42183 -1743 42195 -1567
rect 42229 -1743 42241 -1567
rect 42183 -1755 42241 -1743
rect 42301 -1567 42359 -1555
rect 42301 -1743 42313 -1567
rect 42347 -1743 42359 -1567
rect 42301 -1755 42359 -1743
rect 42419 -1567 42477 -1555
rect 42419 -1743 42431 -1567
rect 42465 -1743 42477 -1567
rect 42419 -1755 42477 -1743
rect 42537 -1567 42595 -1555
rect 42537 -1743 42549 -1567
rect 42583 -1743 42595 -1567
rect 42537 -1755 42595 -1743
rect 42655 -1567 42713 -1555
rect 42655 -1743 42667 -1567
rect 42701 -1743 42713 -1567
rect 42655 -1755 42713 -1743
rect 48147 -1562 48205 -1550
rect 48147 -1738 48159 -1562
rect 48193 -1738 48205 -1562
rect 48147 -1750 48205 -1738
rect 48265 -1562 48323 -1550
rect 48265 -1738 48277 -1562
rect 48311 -1738 48323 -1562
rect 48265 -1750 48323 -1738
rect 48383 -1562 48441 -1550
rect 48383 -1738 48395 -1562
rect 48429 -1738 48441 -1562
rect 48383 -1750 48441 -1738
rect 48501 -1562 48559 -1550
rect 48501 -1738 48513 -1562
rect 48547 -1738 48559 -1562
rect 48501 -1750 48559 -1738
rect 48619 -1562 48677 -1550
rect 48619 -1738 48631 -1562
rect 48665 -1738 48677 -1562
rect 48619 -1750 48677 -1738
rect 48737 -1562 48795 -1550
rect 48737 -1738 48749 -1562
rect 48783 -1738 48795 -1562
rect 48737 -1750 48795 -1738
rect 48855 -1562 48913 -1550
rect 48855 -1738 48867 -1562
rect 48901 -1738 48913 -1562
rect 48855 -1750 48913 -1738
rect 48973 -1562 49031 -1550
rect 48973 -1738 48985 -1562
rect 49019 -1738 49031 -1562
rect 48973 -1750 49031 -1738
rect 49091 -1562 49149 -1550
rect 49091 -1738 49103 -1562
rect 49137 -1738 49149 -1562
rect 49091 -1750 49149 -1738
rect 49209 -1562 49267 -1550
rect 49209 -1738 49221 -1562
rect 49255 -1738 49267 -1562
rect 49209 -1750 49267 -1738
rect 54796 -1574 54854 -1562
rect 54796 -1750 54808 -1574
rect 54842 -1750 54854 -1574
rect 54796 -1762 54854 -1750
rect 54914 -1574 54972 -1562
rect 54914 -1750 54926 -1574
rect 54960 -1750 54972 -1574
rect 54914 -1762 54972 -1750
rect 55032 -1574 55090 -1562
rect 55032 -1750 55044 -1574
rect 55078 -1750 55090 -1574
rect 55032 -1762 55090 -1750
rect 55150 -1574 55208 -1562
rect 55150 -1750 55162 -1574
rect 55196 -1750 55208 -1574
rect 55150 -1762 55208 -1750
rect 55268 -1574 55326 -1562
rect 55268 -1750 55280 -1574
rect 55314 -1750 55326 -1574
rect 55268 -1762 55326 -1750
rect 55386 -1574 55444 -1562
rect 55386 -1750 55398 -1574
rect 55432 -1750 55444 -1574
rect 55386 -1762 55444 -1750
rect 55504 -1574 55562 -1562
rect 55504 -1750 55516 -1574
rect 55550 -1750 55562 -1574
rect 55504 -1762 55562 -1750
rect 55622 -1574 55680 -1562
rect 55622 -1750 55634 -1574
rect 55668 -1750 55680 -1574
rect 55622 -1762 55680 -1750
rect 55740 -1574 55798 -1562
rect 55740 -1750 55752 -1574
rect 55786 -1750 55798 -1574
rect 55740 -1762 55798 -1750
rect 55858 -1574 55916 -1562
rect 55858 -1750 55870 -1574
rect 55904 -1750 55916 -1574
rect 63484 -1625 63496 -1449
rect 63530 -1625 63542 -1449
rect 63484 -1637 63542 -1625
rect 63602 -1449 63660 -1437
rect 63602 -1625 63614 -1449
rect 63648 -1625 63660 -1449
rect 63602 -1637 63660 -1625
rect 63720 -1449 63778 -1437
rect 63720 -1625 63732 -1449
rect 63766 -1625 63778 -1449
rect 63720 -1637 63778 -1625
rect 63838 -1449 63896 -1437
rect 63838 -1625 63850 -1449
rect 63884 -1625 63896 -1449
rect 63838 -1637 63896 -1625
rect 63956 -1449 64014 -1437
rect 63956 -1625 63968 -1449
rect 64002 -1625 64014 -1449
rect 63956 -1637 64014 -1625
rect 64074 -1449 64132 -1437
rect 64074 -1625 64086 -1449
rect 64120 -1625 64132 -1449
rect 64074 -1637 64132 -1625
rect 64192 -1449 64250 -1437
rect 64192 -1625 64204 -1449
rect 64238 -1625 64250 -1449
rect 64192 -1637 64250 -1625
rect 64310 -1449 64368 -1437
rect 64310 -1625 64322 -1449
rect 64356 -1625 64368 -1449
rect 64310 -1637 64368 -1625
rect 64428 -1449 64486 -1437
rect 64428 -1625 64440 -1449
rect 64474 -1625 64486 -1449
rect 64428 -1637 64486 -1625
rect 64546 -1449 64604 -1437
rect 64546 -1625 64558 -1449
rect 64592 -1625 64604 -1449
rect 65651 -1218 65663 -842
rect 65697 -1218 65709 -842
rect 65651 -1230 65709 -1218
rect 65769 -842 65827 -830
rect 65769 -1218 65781 -842
rect 65815 -1218 65827 -842
rect 65769 -1230 65827 -1218
rect 65887 -842 65945 -830
rect 65887 -1218 65899 -842
rect 65933 -1218 65945 -842
rect 65887 -1230 65945 -1218
rect 66005 -842 66063 -830
rect 66005 -1218 66017 -842
rect 66051 -1218 66063 -842
rect 66005 -1230 66063 -1218
rect 66123 -842 66181 -830
rect 66123 -1218 66135 -842
rect 66169 -1218 66181 -842
rect 66123 -1230 66181 -1218
rect 66241 -842 66299 -830
rect 66241 -1218 66253 -842
rect 66287 -1218 66299 -842
rect 66241 -1230 66299 -1218
rect 66359 -842 66417 -830
rect 66359 -1218 66371 -842
rect 66405 -1218 66417 -842
rect 66359 -1230 66417 -1218
rect 70509 -540 70909 -528
rect 70509 -574 70521 -540
rect 70897 -574 70909 -540
rect 70509 -586 70909 -574
rect 70509 -658 70909 -646
rect 70509 -692 70521 -658
rect 70897 -692 70909 -658
rect 70509 -704 70909 -692
rect 70509 -776 70909 -764
rect 70509 -810 70521 -776
rect 70897 -810 70909 -776
rect 70509 -822 70909 -810
rect 70509 -889 70909 -877
rect 70509 -923 70521 -889
rect 70897 -923 70909 -889
rect 70509 -935 70909 -923
rect 70509 -1007 70909 -995
rect 70509 -1041 70521 -1007
rect 70897 -1041 70909 -1007
rect 70509 -1053 70909 -1041
rect 70509 -1125 70909 -1113
rect 70509 -1159 70521 -1125
rect 70897 -1159 70909 -1125
rect 70509 -1171 70909 -1159
rect 70509 -1243 70909 -1231
rect 70509 -1277 70521 -1243
rect 70897 -1277 70909 -1243
rect 70509 -1289 70909 -1277
rect 70509 -1361 70909 -1349
rect 70509 -1395 70521 -1361
rect 70897 -1395 70909 -1361
rect 70509 -1407 70909 -1395
rect 70509 -1479 70909 -1467
rect 70509 -1513 70521 -1479
rect 70897 -1513 70909 -1479
rect 70509 -1525 70909 -1513
rect 64546 -1637 64604 -1625
rect 55858 -1762 55916 -1750
rect 24411 -2148 24469 -2136
rect 24530 -1960 24588 -1948
rect 24530 -2136 24542 -1960
rect 24576 -2136 24588 -1960
rect 24530 -2148 24588 -2136
rect 24648 -1960 24706 -1948
rect 24648 -2136 24660 -1960
rect 24694 -2136 24706 -1960
rect 24648 -2148 24706 -2136
rect 24766 -1960 24824 -1948
rect 24766 -2136 24778 -1960
rect 24812 -2136 24824 -1960
rect 24766 -2148 24824 -2136
rect 24884 -1960 24942 -1948
rect 24884 -2136 24896 -1960
rect 24930 -2136 24942 -1960
rect 29950 -1913 30350 -1901
rect 29950 -1947 29962 -1913
rect 30338 -1947 30350 -1913
rect 29950 -1959 30350 -1947
rect 30643 -1856 31043 -1844
rect 30643 -1890 30655 -1856
rect 31031 -1890 31043 -1856
rect 30643 -1902 31043 -1890
rect 24884 -2148 24942 -2136
rect 29950 -2031 30350 -2019
rect 29950 -2065 29962 -2031
rect 30338 -2065 30350 -2031
rect 29950 -2077 30350 -2065
rect 30643 -1974 31043 -1962
rect 30643 -2008 30655 -1974
rect 31031 -2008 31043 -1974
rect 30643 -2020 31043 -2008
rect 30643 -2092 31043 -2080
rect 30643 -2126 30655 -2092
rect 31031 -2126 31043 -2092
rect 29950 -2149 30350 -2137
rect 30643 -2138 31043 -2126
rect 29950 -2183 29962 -2149
rect 30338 -2183 30350 -2149
rect 29950 -2195 30350 -2183
rect 29950 -2267 30350 -2255
rect 29950 -2301 29962 -2267
rect 30338 -2301 30350 -2267
rect 29950 -2313 30350 -2301
rect 29950 -2385 30350 -2373
rect 29950 -2419 29962 -2385
rect 30338 -2419 30350 -2385
rect 29950 -2431 30350 -2419
rect 30643 -2210 31043 -2198
rect 30643 -2244 30655 -2210
rect 31031 -2244 31043 -2210
rect 30643 -2256 31043 -2244
rect 70509 -1597 70909 -1585
rect 70509 -1631 70521 -1597
rect 70897 -1631 70909 -1597
rect 70509 -1643 70909 -1631
rect 70509 -1716 70909 -1704
rect 70509 -1750 70521 -1716
rect 70897 -1750 70909 -1716
rect 70509 -1762 70909 -1750
rect 70509 -1834 70909 -1822
rect 70509 -1868 70521 -1834
rect 70897 -1868 70909 -1834
rect 70509 -1880 70909 -1868
rect 70509 -1952 70909 -1940
rect 70509 -1986 70521 -1952
rect 70897 -1986 70909 -1952
rect 70509 -1998 70909 -1986
rect 70509 -2070 70909 -2058
rect 70509 -2104 70521 -2070
rect 70897 -2104 70909 -2070
rect 70509 -2116 70909 -2104
rect 70709 -2189 70909 -2177
rect 70709 -2223 70721 -2189
rect 70897 -2223 70909 -2189
rect 70709 -2235 70909 -2223
rect 30643 -2328 31043 -2316
rect 30643 -2362 30655 -2328
rect 31031 -2362 31043 -2328
rect 30643 -2374 31043 -2362
rect 70709 -2307 70909 -2295
rect 70709 -2341 70721 -2307
rect 70897 -2341 70909 -2307
rect 70709 -2353 70909 -2341
rect 29950 -2503 30350 -2491
rect 29950 -2537 29962 -2503
rect 30338 -2537 30350 -2503
rect 29950 -2549 30350 -2537
rect 30150 -2632 30350 -2620
rect 30150 -2666 30162 -2632
rect 30338 -2666 30350 -2632
rect 30150 -2678 30350 -2666
rect 30643 -2446 31043 -2434
rect 30643 -2480 30655 -2446
rect 31031 -2480 31043 -2446
rect 30643 -2492 31043 -2480
rect 70709 -2425 70909 -2413
rect 70709 -2459 70721 -2425
rect 70897 -2459 70909 -2425
rect 70709 -2471 70909 -2459
rect 70709 -2543 70909 -2531
rect 70709 -2577 70721 -2543
rect 70897 -2577 70909 -2543
rect 70709 -2589 70909 -2577
rect 30150 -2750 30350 -2738
rect 30150 -2784 30162 -2750
rect 30338 -2784 30350 -2750
rect 30150 -2796 30350 -2784
rect 30150 -2868 30350 -2856
rect 30150 -2902 30162 -2868
rect 30338 -2902 30350 -2868
rect 30150 -2914 30350 -2902
rect 30150 -2986 30350 -2974
rect 30150 -3020 30162 -2986
rect 30338 -3020 30350 -2986
rect 30150 -3032 30350 -3020
<< ndiffc >>
rect 39837 23708 39871 24084
rect 39955 23708 39989 24084
rect 40073 23708 40107 24084
rect 40190 23908 40224 24084
rect 40308 23908 40342 24084
rect 41835 23634 41869 23810
rect 41953 23634 41987 23810
rect 42071 23634 42105 23810
rect 42189 23634 42223 23810
rect 42977 23638 43011 23814
rect 43095 23638 43129 23814
rect 43213 23638 43247 23814
rect 43331 23638 43365 23814
rect 46350 23705 46384 24081
rect 46468 23705 46502 24081
rect 46586 23705 46620 24081
rect 46703 23905 46737 24081
rect 46821 23905 46855 24081
rect 48348 23631 48382 23807
rect 48466 23631 48500 23807
rect 48584 23631 48618 23807
rect 48702 23631 48736 23807
rect 49490 23635 49524 23811
rect 49608 23635 49642 23811
rect 49726 23635 49760 23811
rect 49844 23635 49878 23811
rect 52884 23700 52918 24076
rect 53002 23700 53036 24076
rect 53120 23700 53154 24076
rect 53237 23900 53271 24076
rect 53355 23900 53389 24076
rect 54882 23626 54916 23802
rect 55000 23626 55034 23802
rect 55118 23626 55152 23802
rect 55236 23626 55270 23802
rect 56024 23630 56058 23806
rect 56142 23630 56176 23806
rect 56260 23630 56294 23806
rect 56378 23630 56412 23806
rect 59442 23704 59476 24080
rect 59560 23704 59594 24080
rect 59678 23704 59712 24080
rect 59795 23904 59829 24080
rect 59913 23904 59947 24080
rect 61440 23630 61474 23806
rect 61558 23630 61592 23806
rect 61676 23630 61710 23806
rect 61794 23630 61828 23806
rect 62582 23634 62616 23810
rect 62700 23634 62734 23810
rect 62818 23634 62852 23810
rect 62936 23634 62970 23810
rect 39851 22058 39885 22434
rect 39969 22058 40003 22434
rect 40087 22058 40121 22434
rect 40204 22258 40238 22434
rect 40322 22258 40356 22434
rect 3880 20475 3914 20651
rect 3998 20475 4032 20651
rect 4076 20275 4110 20651
rect 4194 20275 4228 20651
rect 4312 20275 4346 20651
rect 4430 20275 4464 20651
rect 4548 20275 4582 20651
rect 4622 20475 4656 20651
rect 4740 20475 4774 20651
rect 7024 20475 7058 20651
rect 7142 20475 7176 20651
rect 7220 20275 7254 20651
rect 7338 20275 7372 20651
rect 7456 20275 7490 20651
rect 7574 20275 7608 20651
rect 7692 20275 7726 20651
rect 7766 20475 7800 20651
rect 7884 20475 7918 20651
rect 10156 20471 10190 20647
rect 10274 20471 10308 20647
rect 10352 20271 10386 20647
rect 10470 20271 10504 20647
rect 10588 20271 10622 20647
rect 10706 20271 10740 20647
rect 10824 20271 10858 20647
rect 10898 20471 10932 20647
rect 11016 20471 11050 20647
rect 13300 20471 13334 20647
rect 13418 20471 13452 20647
rect 13496 20271 13530 20647
rect 13614 20271 13648 20647
rect 13732 20271 13766 20647
rect 13850 20271 13884 20647
rect 13968 20271 14002 20647
rect 14042 20471 14076 20647
rect 14160 20471 14194 20647
rect 16502 20475 16536 20651
rect 16620 20475 16654 20651
rect 16698 20275 16732 20651
rect 16816 20275 16850 20651
rect 16934 20275 16968 20651
rect 17052 20275 17086 20651
rect 17170 20275 17204 20651
rect 17244 20475 17278 20651
rect 17362 20475 17396 20651
rect 19646 20475 19680 20651
rect 19764 20475 19798 20651
rect 19842 20275 19876 20651
rect 19960 20275 19994 20651
rect 20078 20275 20112 20651
rect 20196 20275 20230 20651
rect 20314 20275 20348 20651
rect 20388 20475 20422 20651
rect 46364 22055 46398 22431
rect 46482 22055 46516 22431
rect 46600 22055 46634 22431
rect 46717 22255 46751 22431
rect 46835 22255 46869 22431
rect 41203 20853 41237 21029
rect 20506 20475 20540 20651
rect 22778 20471 22812 20647
rect 22896 20471 22930 20647
rect 22974 20271 23008 20647
rect 23092 20271 23126 20647
rect 23210 20271 23244 20647
rect 23328 20271 23362 20647
rect 23446 20271 23480 20647
rect 23520 20471 23554 20647
rect 23638 20471 23672 20647
rect 25922 20471 25956 20647
rect 26040 20471 26074 20647
rect 26118 20271 26152 20647
rect 26236 20271 26270 20647
rect 26354 20271 26388 20647
rect 26472 20271 26506 20647
rect 26590 20271 26624 20647
rect 26664 20471 26698 20647
rect 26782 20471 26816 20647
rect 39846 20454 39880 20830
rect 39964 20454 39998 20830
rect 40082 20454 40116 20830
rect 40199 20654 40233 20830
rect 41321 20853 41355 21029
rect 40317 20654 40351 20830
rect 41623 20653 41657 21029
rect 41741 20653 41775 21029
rect 41859 20653 41893 21029
rect 41977 20653 42011 21029
rect 42095 20653 42129 21029
rect 42501 20853 42535 21029
rect 42619 20853 42653 21029
rect 43101 20853 43135 21029
rect 43219 20853 43253 21029
rect 43521 20653 43555 21029
rect 43639 20653 43673 21029
rect 43757 20653 43791 21029
rect 43875 20653 43909 21029
rect 43993 20653 44027 21029
rect 44399 20853 44433 21029
rect 44517 20853 44551 21029
rect 52898 22050 52932 22426
rect 53016 22050 53050 22426
rect 53134 22050 53168 22426
rect 53251 22250 53285 22426
rect 53369 22250 53403 22426
rect 47716 20850 47750 21026
rect 46359 20451 46393 20827
rect 46477 20451 46511 20827
rect 46595 20451 46629 20827
rect 46712 20651 46746 20827
rect 47834 20850 47868 21026
rect 46830 20651 46864 20827
rect 48136 20650 48170 21026
rect 48254 20650 48288 21026
rect 48372 20650 48406 21026
rect 48490 20650 48524 21026
rect 48608 20650 48642 21026
rect 49014 20850 49048 21026
rect 49132 20850 49166 21026
rect 49614 20850 49648 21026
rect 49732 20850 49766 21026
rect 50034 20650 50068 21026
rect 50152 20650 50186 21026
rect 50270 20650 50304 21026
rect 50388 20650 50422 21026
rect 50506 20650 50540 21026
rect 50912 20850 50946 21026
rect 51030 20850 51064 21026
rect 59456 22054 59490 22430
rect 59574 22054 59608 22430
rect 59692 22054 59726 22430
rect 59809 22254 59843 22430
rect 59927 22254 59961 22430
rect 54250 20845 54284 21021
rect 52893 20446 52927 20822
rect 53011 20446 53045 20822
rect 53129 20446 53163 20822
rect 53246 20646 53280 20822
rect 54368 20845 54402 21021
rect 53364 20646 53398 20822
rect 54670 20645 54704 21021
rect 54788 20645 54822 21021
rect 54906 20645 54940 21021
rect 55024 20645 55058 21021
rect 55142 20645 55176 21021
rect 55548 20845 55582 21021
rect 55666 20845 55700 21021
rect 56148 20845 56182 21021
rect 56266 20845 56300 21021
rect 56568 20645 56602 21021
rect 56686 20645 56720 21021
rect 56804 20645 56838 21021
rect 56922 20645 56956 21021
rect 57040 20645 57074 21021
rect 57446 20845 57480 21021
rect 57564 20845 57598 21021
rect 60808 20849 60842 21025
rect 59451 20450 59485 20826
rect 59569 20450 59603 20826
rect 59687 20450 59721 20826
rect 59804 20650 59838 20826
rect 60926 20849 60960 21025
rect 59922 20650 59956 20826
rect 61228 20649 61262 21025
rect 61346 20649 61380 21025
rect 61464 20649 61498 21025
rect 61582 20649 61616 21025
rect 61700 20649 61734 21025
rect 62106 20849 62140 21025
rect 62224 20849 62258 21025
rect 62706 20849 62740 21025
rect 62824 20849 62858 21025
rect 63126 20649 63160 21025
rect 63244 20649 63278 21025
rect 63362 20649 63396 21025
rect 63480 20649 63514 21025
rect 63598 20649 63632 21025
rect 64004 20849 64038 21025
rect 64122 20849 64156 21025
rect 71858 21193 72034 21227
rect 71858 21075 72034 21109
rect 71858 21001 72234 21035
rect 71858 20883 72234 20917
rect 71858 20765 72234 20799
rect 71858 20647 72234 20681
rect 71858 20529 72234 20563
rect 71858 20451 72034 20485
rect 71858 20333 72034 20367
rect 40055 18030 40089 18206
rect 40173 18030 40207 18206
rect 40291 18030 40325 18206
rect 43078 18300 43112 18476
rect 43196 18300 43230 18476
rect 40409 18030 40443 18206
rect 41197 18026 41231 18202
rect 41315 18026 41349 18202
rect 41433 18026 41467 18202
rect 41551 18026 41585 18202
rect 43313 18100 43347 18476
rect 43431 18100 43465 18476
rect 43549 18100 43583 18476
rect 46613 18026 46647 18202
rect 46731 18026 46765 18202
rect 46849 18026 46883 18202
rect 49636 18296 49670 18472
rect 49754 18296 49788 18472
rect 46967 18026 47001 18202
rect 47755 18022 47789 18198
rect 47873 18022 47907 18198
rect 47991 18022 48025 18198
rect 48109 18022 48143 18198
rect 49871 18096 49905 18472
rect 49989 18096 50023 18472
rect 50107 18096 50141 18472
rect 53147 18031 53181 18207
rect 53265 18031 53299 18207
rect 53383 18031 53417 18207
rect 56170 18301 56204 18477
rect 56288 18301 56322 18477
rect 53501 18031 53535 18207
rect 54289 18027 54323 18203
rect 54407 18027 54441 18203
rect 54525 18027 54559 18203
rect 54643 18027 54677 18203
rect 56405 18101 56439 18477
rect 56523 18101 56557 18477
rect 56641 18101 56675 18477
rect 59660 18034 59694 18210
rect 59778 18034 59812 18210
rect 59896 18034 59930 18210
rect 62683 18304 62717 18480
rect 62801 18304 62835 18480
rect 60014 18034 60048 18210
rect 60802 18030 60836 18206
rect 60920 18030 60954 18206
rect 61038 18030 61072 18206
rect 61156 18030 61190 18206
rect 62918 18104 62952 18480
rect 63036 18104 63070 18480
rect 63154 18104 63188 18480
rect 71858 18049 72034 18083
rect 71858 17931 72034 17965
rect 71858 17857 72234 17891
rect 71858 17739 72234 17773
rect 71858 17621 72234 17655
rect 71858 17503 72234 17537
rect 4964 15838 4998 16014
rect 5082 15838 5116 16014
rect 5200 15838 5234 16014
rect 5318 15838 5352 16014
rect 6132 15838 6166 16014
rect 6250 15838 6284 16014
rect 6368 15838 6402 16014
rect 6486 15838 6520 16014
rect 7300 15836 7334 16012
rect 7418 15836 7452 16012
rect 7536 15836 7570 16012
rect 7654 15836 7688 16012
rect 8468 15836 8502 16012
rect 8586 15836 8620 16012
rect 8704 15836 8738 16012
rect 8822 15836 8856 16012
rect 9642 15836 9676 16012
rect 9760 15836 9794 16012
rect 9878 15836 9912 16012
rect 9996 15836 10030 16012
rect 10810 15836 10844 16012
rect 10928 15836 10962 16012
rect 11046 15836 11080 16012
rect 11164 15836 11198 16012
rect 11978 15836 12012 16012
rect 12096 15836 12130 16012
rect 12214 15836 12248 16012
rect 12332 15836 12366 16012
rect 13146 15834 13180 16010
rect 13264 15834 13298 16010
rect 13382 15834 13416 16010
rect 13500 15834 13534 16010
rect 14157 15988 14191 16164
rect 14275 15988 14309 16164
rect 14392 15788 14426 16164
rect 14510 15788 14544 16164
rect 14628 15788 14662 16164
rect 15605 15988 15639 16164
rect 15723 15988 15757 16164
rect 15840 15788 15874 16164
rect 15958 15788 15992 16164
rect 43064 16650 43098 16826
rect 43182 16650 43216 16826
rect 16076 15788 16110 16164
rect 17103 15986 17137 16162
rect 17221 15986 17255 16162
rect 17338 15786 17372 16162
rect 17456 15786 17490 16162
rect 17574 15786 17608 16162
rect 18551 15986 18585 16162
rect 18669 15986 18703 16162
rect 18786 15786 18820 16162
rect 18904 15786 18938 16162
rect 19022 15786 19056 16162
rect 20071 15988 20105 16164
rect 20189 15988 20223 16164
rect 20306 15788 20340 16164
rect 20424 15788 20458 16164
rect 20542 15788 20576 16164
rect 21519 15988 21553 16164
rect 21637 15988 21671 16164
rect 21754 15788 21788 16164
rect 21872 15788 21906 16164
rect 21990 15788 22024 16164
rect 23017 15986 23051 16162
rect 23135 15986 23169 16162
rect 23252 15786 23286 16162
rect 23370 15786 23404 16162
rect 23488 15786 23522 16162
rect 24465 15986 24499 16162
rect 24583 15986 24617 16162
rect 24700 15786 24734 16162
rect 24818 15786 24852 16162
rect 24936 15786 24970 16162
rect 43299 16450 43333 16826
rect 43417 16450 43451 16826
rect 43535 16450 43569 16826
rect 49622 16646 49656 16822
rect 49740 16646 49774 16822
rect 38869 15245 38903 15421
rect 38987 15245 39021 15421
rect 39393 15045 39427 15421
rect 39511 15045 39545 15421
rect 39629 15045 39663 15421
rect 39747 15045 39781 15421
rect 39865 15045 39899 15421
rect 40167 15245 40201 15421
rect 40285 15245 40319 15421
rect 40767 15245 40801 15421
rect 40885 15245 40919 15421
rect 41291 15045 41325 15421
rect 41409 15045 41443 15421
rect 41527 15045 41561 15421
rect 41645 15045 41679 15421
rect 41763 15045 41797 15421
rect 42065 15245 42099 15421
rect 42183 15245 42217 15421
rect 49857 16446 49891 16822
rect 49975 16446 50009 16822
rect 50093 16446 50127 16822
rect 56156 16651 56190 16827
rect 56274 16651 56308 16827
rect 45427 15241 45461 15417
rect 43069 15046 43103 15222
rect 43187 15046 43221 15222
rect 1378 13337 1412 13513
rect 1496 13337 1530 13513
rect 1574 13137 1608 13513
rect 1692 13137 1726 13513
rect 1810 13137 1844 13513
rect 1928 13137 1962 13513
rect 2046 13137 2080 13513
rect 2120 13337 2154 13513
rect 2238 13337 2272 13513
rect 4522 13337 4556 13513
rect 4640 13337 4674 13513
rect 4718 13137 4752 13513
rect 4836 13137 4870 13513
rect 4954 13137 4988 13513
rect 5072 13137 5106 13513
rect 5190 13137 5224 13513
rect 5264 13337 5298 13513
rect 43304 14846 43338 15222
rect 43422 14846 43456 15222
rect 45545 15241 45579 15417
rect 43540 14846 43574 15222
rect 45951 15041 45985 15417
rect 46069 15041 46103 15417
rect 46187 15041 46221 15417
rect 46305 15041 46339 15417
rect 46423 15041 46457 15417
rect 46725 15241 46759 15417
rect 46843 15241 46877 15417
rect 47325 15241 47359 15417
rect 47443 15241 47477 15417
rect 47849 15041 47883 15417
rect 47967 15041 48001 15417
rect 48085 15041 48119 15417
rect 48203 15041 48237 15417
rect 48321 15041 48355 15417
rect 48623 15241 48657 15417
rect 48741 15241 48775 15417
rect 56391 16451 56425 16827
rect 56509 16451 56543 16827
rect 56627 16451 56661 16827
rect 71858 17385 72234 17419
rect 71858 17307 72034 17341
rect 62669 16654 62703 16830
rect 62787 16654 62821 16830
rect 51961 15246 51995 15422
rect 52079 15246 52113 15422
rect 49627 15042 49661 15218
rect 49745 15042 49779 15218
rect 49862 14842 49896 15218
rect 49980 14842 50014 15218
rect 50098 14842 50132 15218
rect 52485 15046 52519 15422
rect 52603 15046 52637 15422
rect 52721 15046 52755 15422
rect 52839 15046 52873 15422
rect 52957 15046 52991 15422
rect 53259 15246 53293 15422
rect 53377 15246 53411 15422
rect 53859 15246 53893 15422
rect 53977 15246 54011 15422
rect 54383 15046 54417 15422
rect 54501 15046 54535 15422
rect 54619 15046 54653 15422
rect 54737 15046 54771 15422
rect 54855 15046 54889 15422
rect 55157 15246 55191 15422
rect 55275 15246 55309 15422
rect 62904 16454 62938 16830
rect 63022 16454 63056 16830
rect 63140 16454 63174 16830
rect 71858 17189 72034 17223
rect 58474 15249 58508 15425
rect 58592 15249 58626 15425
rect 56161 15047 56195 15223
rect 56279 15047 56313 15223
rect 56396 14847 56430 15223
rect 56514 14847 56548 15223
rect 56632 14847 56666 15223
rect 58998 15049 59032 15425
rect 59116 15049 59150 15425
rect 59234 15049 59268 15425
rect 59352 15049 59386 15425
rect 59470 15049 59504 15425
rect 59772 15249 59806 15425
rect 59890 15249 59924 15425
rect 60372 15249 60406 15425
rect 60490 15249 60524 15425
rect 60896 15049 60930 15425
rect 61014 15049 61048 15425
rect 61132 15049 61166 15425
rect 61250 15049 61284 15425
rect 61368 15049 61402 15425
rect 61670 15249 61704 15425
rect 61788 15249 61822 15425
rect 62674 15050 62708 15226
rect 62792 15050 62826 15226
rect 62909 14850 62943 15226
rect 63027 14850 63061 15226
rect 63145 14850 63179 15226
rect 71854 14917 72030 14951
rect 71854 14799 72030 14833
rect 71854 14725 72230 14759
rect 5382 13337 5416 13513
rect 7654 13333 7688 13509
rect 7772 13333 7806 13509
rect 7850 13133 7884 13509
rect 7968 13133 8002 13509
rect 8086 13133 8120 13509
rect 8204 13133 8238 13509
rect 8322 13133 8356 13509
rect 8396 13333 8430 13509
rect 8514 13333 8548 13509
rect 10798 13333 10832 13509
rect 10916 13333 10950 13509
rect 10994 13133 11028 13509
rect 11112 13133 11146 13509
rect 11230 13133 11264 13509
rect 11348 13133 11382 13509
rect 11466 13133 11500 13509
rect 11540 13333 11574 13509
rect 11658 13333 11692 13509
rect 14000 13337 14034 13513
rect 14118 13337 14152 13513
rect 14196 13137 14230 13513
rect 14314 13137 14348 13513
rect 14432 13137 14466 13513
rect 14550 13137 14584 13513
rect 14668 13137 14702 13513
rect 14742 13337 14776 13513
rect 14860 13337 14894 13513
rect 17144 13337 17178 13513
rect 17262 13337 17296 13513
rect 17340 13137 17374 13513
rect 17458 13137 17492 13513
rect 17576 13137 17610 13513
rect 17694 13137 17728 13513
rect 17812 13137 17846 13513
rect 17886 13337 17920 13513
rect 71854 14607 72230 14641
rect 71854 14489 72230 14523
rect 71854 14371 72230 14405
rect 71854 14253 72230 14287
rect 71854 14175 72030 14209
rect 18004 13337 18038 13513
rect 20276 13333 20310 13509
rect 20394 13333 20428 13509
rect 20472 13133 20506 13509
rect 20590 13133 20624 13509
rect 20708 13133 20742 13509
rect 20826 13133 20860 13509
rect 20944 13133 20978 13509
rect 21018 13333 21052 13509
rect 21136 13333 21170 13509
rect 23420 13333 23454 13509
rect 23538 13333 23572 13509
rect 23616 13133 23650 13509
rect 23734 13133 23768 13509
rect 23852 13133 23886 13509
rect 23970 13133 24004 13509
rect 24088 13133 24122 13509
rect 24162 13333 24196 13509
rect 24280 13333 24314 13509
rect 71854 14057 72030 14091
rect 31391 13009 31567 13043
rect 31391 12891 31567 12925
rect 31391 12589 31767 12623
rect 31391 12471 31767 12505
rect 31391 12353 31767 12387
rect 1378 10603 1412 10779
rect 1496 10603 1530 10779
rect 1574 10403 1608 10779
rect 1692 10403 1726 10779
rect 1810 10403 1844 10779
rect 1928 10403 1962 10779
rect 2046 10403 2080 10779
rect 2120 10603 2154 10779
rect 2238 10603 2272 10779
rect 4522 10603 4556 10779
rect 4640 10603 4674 10779
rect 4718 10403 4752 10779
rect 4836 10403 4870 10779
rect 4954 10403 4988 10779
rect 5072 10403 5106 10779
rect 5190 10403 5224 10779
rect 5264 10603 5298 10779
rect 31391 12235 31767 12269
rect 31391 12117 31767 12151
rect 5382 10603 5416 10779
rect 7654 10599 7688 10775
rect 7772 10599 7806 10775
rect 7850 10399 7884 10775
rect 7968 10399 8002 10775
rect 8086 10399 8120 10775
rect 8204 10399 8238 10775
rect 8322 10399 8356 10775
rect 8396 10599 8430 10775
rect 8514 10599 8548 10775
rect 10798 10599 10832 10775
rect 10916 10599 10950 10775
rect 10994 10399 11028 10775
rect 11112 10399 11146 10775
rect 11230 10399 11264 10775
rect 11348 10399 11382 10775
rect 11466 10399 11500 10775
rect 11540 10599 11574 10775
rect 11658 10599 11692 10775
rect 14000 10603 14034 10779
rect 14118 10603 14152 10779
rect 14196 10403 14230 10779
rect 14314 10403 14348 10779
rect 14432 10403 14466 10779
rect 14550 10403 14584 10779
rect 14668 10403 14702 10779
rect 14742 10603 14776 10779
rect 14860 10603 14894 10779
rect 17144 10603 17178 10779
rect 17262 10603 17296 10779
rect 17340 10403 17374 10779
rect 17458 10403 17492 10779
rect 17576 10403 17610 10779
rect 17694 10403 17728 10779
rect 17812 10403 17846 10779
rect 17886 10603 17920 10779
rect 31391 11711 31567 11745
rect 31391 11593 31567 11627
rect 41807 11324 41841 11700
rect 41925 11324 41959 11700
rect 42043 11324 42077 11700
rect 42160 11524 42194 11700
rect 42278 11524 42312 11700
rect 48356 11323 48390 11699
rect 48474 11323 48508 11699
rect 48592 11323 48626 11699
rect 48709 11523 48743 11699
rect 48827 11523 48861 11699
rect 55010 11344 55044 11720
rect 55128 11344 55162 11720
rect 55246 11344 55280 11720
rect 55363 11544 55397 11720
rect 55481 11544 55515 11720
rect 63663 11177 63697 11553
rect 63781 11177 63815 11553
rect 63899 11177 63933 11553
rect 64016 11377 64050 11553
rect 64134 11377 64168 11553
rect 71854 11773 72030 11807
rect 71854 11655 72030 11689
rect 71854 11581 72230 11615
rect 31389 10941 31565 10975
rect 18004 10603 18038 10779
rect 20276 10599 20310 10775
rect 20394 10599 20428 10775
rect 20472 10399 20506 10775
rect 20590 10399 20624 10775
rect 20708 10399 20742 10775
rect 20826 10399 20860 10775
rect 20944 10399 20978 10775
rect 21018 10599 21052 10775
rect 21136 10599 21170 10775
rect 23420 10599 23454 10775
rect 23538 10599 23572 10775
rect 23616 10399 23650 10775
rect 23734 10399 23768 10775
rect 23852 10399 23886 10775
rect 23970 10399 24004 10775
rect 24088 10399 24122 10775
rect 24162 10599 24196 10775
rect 24280 10599 24314 10775
rect 31389 10823 31565 10857
rect 31389 10521 31765 10555
rect 31389 10403 31765 10437
rect 31389 10285 31765 10319
rect 31389 10167 31765 10201
rect 31389 10049 31765 10083
rect 71854 11463 72230 11497
rect 71854 11345 72230 11379
rect 71854 11227 72230 11261
rect 67264 10769 67298 11145
rect 67382 10769 67416 11145
rect 67500 10769 67534 11145
rect 67617 10969 67651 11145
rect 67735 10969 67769 11145
rect 71854 11109 72230 11143
rect 71854 11031 72030 11065
rect 31389 9643 31565 9677
rect 31389 9525 31565 9559
rect 35143 9424 35177 9800
rect 35261 9424 35295 9800
rect 35379 9424 35413 9800
rect 35496 9624 35530 9800
rect 35614 9624 35648 9800
rect 1388 7871 1422 8047
rect 1506 7871 1540 8047
rect 1584 7671 1618 8047
rect 1702 7671 1736 8047
rect 1820 7671 1854 8047
rect 1938 7671 1972 8047
rect 2056 7671 2090 8047
rect 2130 7871 2164 8047
rect 2248 7871 2282 8047
rect 4532 7871 4566 8047
rect 4650 7871 4684 8047
rect 4728 7671 4762 8047
rect 4846 7671 4880 8047
rect 4964 7671 4998 8047
rect 5082 7671 5116 8047
rect 5200 7671 5234 8047
rect 5274 7871 5308 8047
rect 38033 9157 38067 9533
rect 38151 9157 38185 9533
rect 38269 9157 38303 9533
rect 38386 9357 38420 9533
rect 38504 9357 38538 9533
rect 65359 10184 65393 10360
rect 65477 10184 65511 10360
rect 40031 9083 40065 9259
rect 40149 9083 40183 9259
rect 40267 9083 40301 9259
rect 40385 9083 40419 9259
rect 41173 9087 41207 9263
rect 41291 9087 41325 9263
rect 41409 9087 41443 9263
rect 41527 9087 41561 9263
rect 44582 9245 44616 9621
rect 44700 9245 44734 9621
rect 44818 9245 44852 9621
rect 44935 9445 44969 9621
rect 45053 9445 45087 9621
rect 46580 9171 46614 9347
rect 46698 9171 46732 9347
rect 46816 9171 46850 9347
rect 46934 9171 46968 9347
rect 47722 9175 47756 9351
rect 47840 9175 47874 9351
rect 47958 9175 47992 9351
rect 48076 9175 48110 9351
rect 51236 9177 51270 9553
rect 51354 9177 51388 9553
rect 51472 9177 51506 9553
rect 51589 9377 51623 9553
rect 51707 9377 51741 9553
rect 65779 9984 65813 10360
rect 65897 9984 65931 10360
rect 66015 9984 66049 10360
rect 66133 9984 66167 10360
rect 66251 9984 66285 10360
rect 66657 10184 66691 10360
rect 66775 10184 66809 10360
rect 71854 10913 72030 10947
rect 53234 9103 53268 9279
rect 53352 9103 53386 9279
rect 53470 9103 53504 9279
rect 53588 9103 53622 9279
rect 54376 9107 54410 9283
rect 54494 9107 54528 9283
rect 54612 9107 54646 9283
rect 54730 9107 54764 9283
rect 57861 9245 57895 9621
rect 57979 9245 58013 9621
rect 58097 9245 58131 9621
rect 58214 9445 58248 9621
rect 58332 9445 58366 9621
rect 59859 9171 59893 9347
rect 59977 9171 60011 9347
rect 60095 9171 60129 9347
rect 60213 9171 60247 9347
rect 61001 9175 61035 9351
rect 61119 9175 61153 9351
rect 61237 9175 61271 9351
rect 61355 9175 61389 9351
rect 5392 7871 5426 8047
rect 7664 7867 7698 8043
rect 7782 7867 7816 8043
rect 7860 7667 7894 8043
rect 7978 7667 8012 8043
rect 8096 7667 8130 8043
rect 8214 7667 8248 8043
rect 8332 7667 8366 8043
rect 8406 7867 8440 8043
rect 8524 7867 8558 8043
rect 10808 7867 10842 8043
rect 10926 7867 10960 8043
rect 11004 7667 11038 8043
rect 11122 7667 11156 8043
rect 11240 7667 11274 8043
rect 11358 7667 11392 8043
rect 11476 7667 11510 8043
rect 11550 7867 11584 8043
rect 11668 7867 11702 8043
rect 14010 7871 14044 8047
rect 14128 7871 14162 8047
rect 14206 7671 14240 8047
rect 14324 7671 14358 8047
rect 14442 7671 14476 8047
rect 14560 7671 14594 8047
rect 14678 7671 14712 8047
rect 14752 7871 14786 8047
rect 14870 7871 14904 8047
rect 17154 7871 17188 8047
rect 17272 7871 17306 8047
rect 17350 7671 17384 8047
rect 17468 7671 17502 8047
rect 17586 7671 17620 8047
rect 17704 7671 17738 8047
rect 17822 7671 17856 8047
rect 17896 7871 17930 8047
rect 31391 8872 31567 8906
rect 31391 8754 31567 8788
rect 63658 8606 63692 8982
rect 63776 8606 63810 8982
rect 63894 8606 63928 8982
rect 64011 8806 64045 8982
rect 64129 8806 64163 8982
rect 31391 8452 31767 8486
rect 31391 8334 31767 8368
rect 31391 8216 31767 8250
rect 18014 7871 18048 8047
rect 20286 7867 20320 8043
rect 20404 7867 20438 8043
rect 20482 7667 20516 8043
rect 20600 7667 20634 8043
rect 20718 7667 20752 8043
rect 20836 7667 20870 8043
rect 20954 7667 20988 8043
rect 21028 7867 21062 8043
rect 21146 7867 21180 8043
rect 23430 7867 23464 8043
rect 23548 7867 23582 8043
rect 23626 7667 23660 8043
rect 23744 7667 23778 8043
rect 23862 7667 23896 8043
rect 23980 7667 24014 8043
rect 24098 7667 24132 8043
rect 24172 7867 24206 8043
rect 24290 7867 24324 8043
rect 31391 8098 31767 8132
rect 31391 7980 31767 8014
rect 71858 8571 72034 8605
rect 71858 8453 72034 8487
rect 71858 8379 72234 8413
rect 31391 7574 31567 7608
rect 31391 7456 31567 7490
rect 38047 7507 38081 7883
rect 38165 7507 38199 7883
rect 38283 7507 38317 7883
rect 38400 7707 38434 7883
rect 38518 7707 38552 7883
rect 44596 7595 44630 7971
rect 44714 7595 44748 7971
rect 44832 7595 44866 7971
rect 44949 7795 44983 7971
rect 45067 7795 45101 7971
rect 31389 6804 31565 6838
rect 35135 6839 35169 7215
rect 35253 6839 35287 7215
rect 35371 6839 35405 7215
rect 35488 7039 35522 7215
rect 35606 7039 35640 7215
rect 31389 6686 31565 6720
rect 3247 5987 3281 6163
rect 3365 5987 3399 6163
rect 3985 5987 4019 6163
rect 4103 5987 4137 6163
rect 4723 5983 4757 6159
rect 4841 5983 4875 6159
rect 5461 5983 5495 6159
rect 5579 5983 5613 6159
rect 6201 5983 6235 6159
rect 6319 5983 6353 6159
rect 6943 5983 6977 6159
rect 7061 5983 7095 6159
rect 7681 5987 7715 6163
rect 7799 5987 7833 6163
rect 8419 5985 8453 6161
rect 8537 5985 8571 6161
rect 9367 4834 9401 5010
rect 9485 4834 9519 5010
rect 9891 4634 9925 5010
rect 10009 4634 10043 5010
rect 10127 4634 10161 5010
rect 10245 4634 10279 5010
rect 10363 4634 10397 5010
rect 10665 4834 10699 5010
rect 10783 4834 10817 5010
rect 11435 4832 11469 5008
rect 11553 4832 11587 5008
rect 11959 4632 11993 5008
rect 12077 4632 12111 5008
rect 12195 4632 12229 5008
rect 12313 4632 12347 5008
rect 12431 4632 12465 5008
rect 12733 4832 12767 5008
rect 12851 4832 12885 5008
rect 13504 4834 13538 5010
rect 13622 4834 13656 5010
rect 14028 4634 14062 5010
rect 14146 4634 14180 5010
rect 14264 4634 14298 5010
rect 14382 4634 14416 5010
rect 14500 4634 14534 5010
rect 14802 4834 14836 5010
rect 31389 6384 31765 6418
rect 31389 6266 31765 6300
rect 71858 8261 72234 8295
rect 71858 8143 72234 8177
rect 71858 8025 72234 8059
rect 39399 6302 39433 6478
rect 31389 6148 31765 6182
rect 14920 4834 14954 5010
rect 15572 4832 15606 5008
rect 15690 4832 15724 5008
rect 16096 4632 16130 5008
rect 16214 4632 16248 5008
rect 16332 4632 16366 5008
rect 16450 4632 16484 5008
rect 16568 4632 16602 5008
rect 16870 4832 16904 5008
rect 16988 4832 17022 5008
rect 17641 4832 17675 5008
rect 17759 4832 17793 5008
rect 18165 4632 18199 5008
rect 18283 4632 18317 5008
rect 18401 4632 18435 5008
rect 18519 4632 18553 5008
rect 18637 4632 18671 5008
rect 18939 4832 18973 5008
rect 31389 6030 31765 6064
rect 31389 5912 31765 5946
rect 38042 5903 38076 6279
rect 38160 5903 38194 6279
rect 38278 5903 38312 6279
rect 38395 6103 38429 6279
rect 39517 6302 39551 6478
rect 38513 6103 38547 6279
rect 39819 6102 39853 6478
rect 39937 6102 39971 6478
rect 40055 6102 40089 6478
rect 40173 6102 40207 6478
rect 40291 6102 40325 6478
rect 40697 6302 40731 6478
rect 40815 6302 40849 6478
rect 41297 6302 41331 6478
rect 41415 6302 41449 6478
rect 41717 6102 41751 6478
rect 41835 6102 41869 6478
rect 41953 6102 41987 6478
rect 42071 6102 42105 6478
rect 42189 6102 42223 6478
rect 42595 6302 42629 6478
rect 42713 6302 42747 6478
rect 51250 7527 51284 7903
rect 51368 7527 51402 7903
rect 51486 7527 51520 7903
rect 51603 7727 51637 7903
rect 51721 7727 51755 7903
rect 57875 7595 57909 7971
rect 57993 7595 58027 7971
rect 58111 7595 58145 7971
rect 58228 7795 58262 7971
rect 58346 7795 58380 7971
rect 45948 6390 45982 6566
rect 44591 5991 44625 6367
rect 44709 5991 44743 6367
rect 44827 5991 44861 6367
rect 44944 6191 44978 6367
rect 46066 6390 46100 6566
rect 45062 6191 45096 6367
rect 46368 6190 46402 6566
rect 46486 6190 46520 6566
rect 46604 6190 46638 6566
rect 46722 6190 46756 6566
rect 46840 6190 46874 6566
rect 47246 6390 47280 6566
rect 47364 6390 47398 6566
rect 47846 6390 47880 6566
rect 47964 6390 47998 6566
rect 48266 6190 48300 6566
rect 48384 6190 48418 6566
rect 48502 6190 48536 6566
rect 48620 6190 48654 6566
rect 48738 6190 48772 6566
rect 49144 6390 49178 6566
rect 49262 6390 49296 6566
rect 52602 6322 52636 6498
rect 19057 4832 19091 5008
rect 19709 4830 19743 5006
rect 19827 4830 19861 5006
rect 20233 4630 20267 5006
rect 20351 4630 20385 5006
rect 20469 4630 20503 5006
rect 20587 4630 20621 5006
rect 20705 4630 20739 5006
rect 21007 4830 21041 5006
rect 21125 4830 21159 5006
rect 21778 4832 21812 5008
rect 21896 4832 21930 5008
rect 22302 4632 22336 5008
rect 22420 4632 22454 5008
rect 22538 4632 22572 5008
rect 22656 4632 22690 5008
rect 22774 4632 22808 5008
rect 23076 4832 23110 5008
rect 51245 5923 51279 6299
rect 51363 5923 51397 6299
rect 51481 5923 51515 6299
rect 51598 6123 51632 6299
rect 52720 6322 52754 6498
rect 51716 6123 51750 6299
rect 53022 6122 53056 6498
rect 53140 6122 53174 6498
rect 53258 6122 53292 6498
rect 53376 6122 53410 6498
rect 53494 6122 53528 6498
rect 53900 6322 53934 6498
rect 54018 6322 54052 6498
rect 54500 6322 54534 6498
rect 54618 6322 54652 6498
rect 54920 6122 54954 6498
rect 55038 6122 55072 6498
rect 55156 6122 55190 6498
rect 55274 6122 55308 6498
rect 55392 6122 55426 6498
rect 55798 6322 55832 6498
rect 55916 6322 55950 6498
rect 71858 7907 72234 7941
rect 71858 7829 72034 7863
rect 59227 6390 59261 6566
rect 57870 5991 57904 6367
rect 57988 5991 58022 6367
rect 58106 5991 58140 6367
rect 58223 6191 58257 6367
rect 59345 6390 59379 6566
rect 58341 6191 58375 6367
rect 59647 6190 59681 6566
rect 59765 6190 59799 6566
rect 59883 6190 59917 6566
rect 60001 6190 60035 6566
rect 60119 6190 60153 6566
rect 60525 6390 60559 6566
rect 60643 6390 60677 6566
rect 61125 6390 61159 6566
rect 61243 6390 61277 6566
rect 61545 6190 61579 6566
rect 61663 6190 61697 6566
rect 61781 6190 61815 6566
rect 61899 6190 61933 6566
rect 62017 6190 62051 6566
rect 62423 6390 62457 6566
rect 62541 6390 62575 6566
rect 67266 6678 67300 7054
rect 67384 6678 67418 7054
rect 67502 6678 67536 7054
rect 67619 6878 67653 7054
rect 67737 6878 67771 7054
rect 71858 7711 72034 7745
rect 65361 6093 65395 6269
rect 65479 6093 65513 6269
rect 63658 5573 63692 5949
rect 63776 5573 63810 5949
rect 63894 5573 63928 5949
rect 64011 5773 64045 5949
rect 64129 5773 64163 5949
rect 65781 5893 65815 6269
rect 65899 5893 65933 6269
rect 66017 5893 66051 6269
rect 66135 5893 66169 6269
rect 66253 5893 66287 6269
rect 66659 6093 66693 6269
rect 66777 6093 66811 6269
rect 31389 5506 31565 5540
rect 31389 5388 31565 5422
rect 71858 5427 72034 5461
rect 71858 5309 72034 5343
rect 71858 5235 72234 5269
rect 23194 4832 23228 5008
rect 23846 4830 23880 5006
rect 23964 4830 23998 5006
rect 24370 4630 24404 5006
rect 24488 4630 24522 5006
rect 24606 4630 24640 5006
rect 24724 4630 24758 5006
rect 24842 4630 24876 5006
rect 25144 4830 25178 5006
rect 25262 4830 25296 5006
rect 71858 5117 72234 5151
rect 71858 4999 72234 5033
rect 71858 4881 72234 4915
rect 31389 4735 31565 4769
rect 31389 4617 31565 4651
rect 31389 4315 31765 4349
rect 31389 4197 31765 4231
rect 31389 4079 31765 4113
rect 31389 3961 31765 3995
rect 31389 3843 31765 3877
rect 35116 3561 35150 3937
rect 35234 3561 35268 3937
rect 35352 3561 35386 3937
rect 35469 3761 35503 3937
rect 35587 3761 35621 3937
rect 31389 3437 31565 3471
rect 31389 3319 31565 3353
rect 38025 3377 38059 3753
rect 38143 3377 38177 3753
rect 38261 3377 38295 3753
rect 38378 3577 38412 3753
rect 38496 3577 38530 3753
rect 40023 3303 40057 3479
rect 40141 3303 40175 3479
rect 40259 3303 40293 3479
rect 40377 3303 40411 3479
rect 41165 3307 41199 3483
rect 41283 3307 41317 3483
rect 41401 3307 41435 3483
rect 41519 3307 41553 3483
rect 44576 3375 44610 3751
rect 44694 3375 44728 3751
rect 44812 3375 44846 3751
rect 44929 3575 44963 3751
rect 45047 3575 45081 3751
rect 71858 4763 72234 4797
rect 71858 4685 72034 4719
rect 46574 3301 46608 3477
rect 46692 3301 46726 3477
rect 46810 3301 46844 3477
rect 46928 3301 46962 3477
rect 47716 3305 47750 3481
rect 47834 3305 47868 3481
rect 47952 3305 47986 3481
rect 48070 3305 48104 3481
rect 51231 3376 51265 3752
rect 51349 3376 51383 3752
rect 51467 3376 51501 3752
rect 51584 3576 51618 3752
rect 51702 3576 51736 3752
rect 53229 3302 53263 3478
rect 53347 3302 53381 3478
rect 53465 3302 53499 3478
rect 53583 3302 53617 3478
rect 54371 3306 54405 3482
rect 54489 3306 54523 3482
rect 54607 3306 54641 3482
rect 54725 3306 54759 3482
rect 57853 3377 57887 3753
rect 57971 3377 58005 3753
rect 58089 3377 58123 3753
rect 58206 3577 58240 3753
rect 58324 3577 58358 3753
rect 63729 3653 63763 4029
rect 63847 3653 63881 4029
rect 63965 3653 63999 4029
rect 64082 3853 64116 4029
rect 64200 3853 64234 4029
rect 59851 3303 59885 3479
rect 59969 3303 60003 3479
rect 60087 3303 60121 3479
rect 60205 3303 60239 3479
rect 60993 3307 61027 3483
rect 61111 3307 61145 3483
rect 61229 3307 61263 3483
rect 61347 3307 61381 3483
rect 71858 4567 72034 4601
rect 67266 3183 67300 3559
rect 67384 3183 67418 3559
rect 67502 3183 67536 3559
rect 67619 3383 67653 3559
rect 67737 3383 67771 3559
rect 31387 2667 31563 2701
rect 31387 2549 31563 2583
rect 31387 2247 31763 2281
rect 31387 2129 31763 2163
rect 65361 2598 65395 2774
rect 65479 2598 65513 2774
rect 65781 2398 65815 2774
rect 65899 2398 65933 2774
rect 66017 2398 66051 2774
rect 66135 2398 66169 2774
rect 66253 2398 66287 2774
rect 66659 2598 66693 2774
rect 66777 2598 66811 2774
rect 31387 2011 31763 2045
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 31387 1893 31763 1927
rect 31387 1775 31763 1809
rect 38039 1727 38073 2103
rect 38157 1727 38191 2103
rect 38275 1727 38309 2103
rect 38392 1927 38426 2103
rect 38510 1927 38544 2103
rect 31387 1369 31563 1403
rect 31387 1251 31563 1285
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 35132 801 35166 1177
rect 35250 801 35284 1177
rect 35368 801 35402 1177
rect 35485 1001 35519 1177
rect 35603 1001 35637 1177
rect 31389 598 31565 632
rect 31389 480 31565 514
rect 44590 1725 44624 2101
rect 44708 1725 44742 2101
rect 44826 1725 44860 2101
rect 44943 1925 44977 2101
rect 45061 1925 45095 2101
rect 39391 522 39425 698
rect 31389 178 31765 212
rect 38034 123 38068 499
rect 38152 123 38186 499
rect 38270 123 38304 499
rect 38387 323 38421 499
rect 39509 522 39543 698
rect 38505 323 38539 499
rect 39811 322 39845 698
rect 39929 322 39963 698
rect 40047 322 40081 698
rect 40165 322 40199 698
rect 40283 322 40317 698
rect 40689 522 40723 698
rect 40807 522 40841 698
rect 41289 522 41323 698
rect 41407 522 41441 698
rect 41709 322 41743 698
rect 41827 322 41861 698
rect 41945 322 41979 698
rect 42063 322 42097 698
rect 42181 322 42215 698
rect 42587 522 42621 698
rect 42705 522 42739 698
rect 51245 1726 51279 2102
rect 51363 1726 51397 2102
rect 51481 1726 51515 2102
rect 51598 1926 51632 2102
rect 51716 1926 51750 2102
rect 45942 520 45976 696
rect 31389 60 31765 94
rect 44585 121 44619 497
rect 44703 121 44737 497
rect 44821 121 44855 497
rect 44938 321 44972 497
rect 46060 520 46094 696
rect 45056 321 45090 497
rect 46362 320 46396 696
rect 46480 320 46514 696
rect 46598 320 46632 696
rect 46716 320 46750 696
rect 46834 320 46868 696
rect 47240 520 47274 696
rect 47358 520 47392 696
rect 47840 520 47874 696
rect 47958 520 47992 696
rect 48260 320 48294 696
rect 48378 320 48412 696
rect 48496 320 48530 696
rect 48614 320 48648 696
rect 48732 320 48766 696
rect 49138 520 49172 696
rect 49256 520 49290 696
rect 57867 1727 57901 2103
rect 57985 1727 58019 2103
rect 58103 1727 58137 2103
rect 58220 1927 58254 2103
rect 58338 1927 58372 2103
rect 71854 2295 72030 2329
rect 71854 2177 72030 2211
rect 71854 2103 72230 2137
rect 71854 1985 72230 2019
rect 52597 521 52631 697
rect 31389 -58 31765 -24
rect 31389 -176 31765 -142
rect 51240 122 51274 498
rect 51358 122 51392 498
rect 51476 122 51510 498
rect 51593 322 51627 498
rect 52715 521 52749 697
rect 51711 322 51745 498
rect 53017 321 53051 697
rect 53135 321 53169 697
rect 53253 321 53287 697
rect 53371 321 53405 697
rect 53489 321 53523 697
rect 53895 521 53929 697
rect 54013 521 54047 697
rect 54495 521 54529 697
rect 54613 521 54647 697
rect 54915 321 54949 697
rect 55033 321 55067 697
rect 55151 321 55185 697
rect 55269 321 55303 697
rect 55387 321 55421 697
rect 55793 521 55827 697
rect 55911 521 55945 697
rect 71854 1867 72230 1901
rect 71854 1749 72230 1783
rect 71854 1631 72230 1665
rect 71854 1553 72030 1587
rect 59219 522 59253 698
rect 57862 123 57896 499
rect 57980 123 58014 499
rect 58098 123 58132 499
rect 58215 323 58249 499
rect 59337 522 59371 698
rect 58333 323 58367 499
rect 59639 322 59673 698
rect 59757 322 59791 698
rect 59875 322 59909 698
rect 59993 322 60027 698
rect 60111 322 60145 698
rect 60517 522 60551 698
rect 60635 522 60669 698
rect 61117 522 61151 698
rect 61235 522 61269 698
rect 61537 322 61571 698
rect 61655 322 61689 698
rect 61773 322 61807 698
rect 61891 322 61925 698
rect 62009 322 62043 698
rect 62415 522 62449 698
rect 62533 522 62567 698
rect 63726 583 63760 959
rect 63844 583 63878 959
rect 63962 583 63996 959
rect 64079 783 64113 959
rect 64197 783 64231 959
rect 71854 1435 72030 1469
rect 31389 -294 31765 -260
rect 31389 -700 31565 -666
rect 31389 -818 31565 -784
rect 41842 -1306 41876 -930
rect 41960 -1306 41994 -930
rect 42078 -1306 42112 -930
rect 42195 -1306 42229 -1130
rect 42313 -1306 42347 -1130
rect 48396 -1301 48430 -925
rect 48514 -1301 48548 -925
rect 48632 -1301 48666 -925
rect 48749 -1301 48783 -1125
rect 48867 -1301 48901 -1125
rect 55045 -1313 55079 -937
rect 31387 -1470 31563 -1436
rect 31387 -1588 31563 -1554
rect 55163 -1313 55197 -937
rect 55281 -1313 55315 -937
rect 55398 -1313 55432 -1137
rect 55516 -1313 55550 -1137
rect 67266 -1165 67300 -789
rect 67384 -1165 67418 -789
rect 67502 -1165 67536 -789
rect 67619 -965 67653 -789
rect 67737 -965 67771 -789
rect 71854 -849 72030 -815
rect 71854 -967 72030 -933
rect 71854 -1041 72230 -1007
rect 71854 -1159 72230 -1125
rect 71854 -1277 72230 -1243
rect 71854 -1395 72230 -1361
rect 31387 -1890 31763 -1856
rect 65361 -1750 65395 -1574
rect 65479 -1750 65513 -1574
rect 1126 -3273 1160 -3097
rect 1244 -3273 1278 -3097
rect 1318 -3473 1352 -3097
rect 1436 -3473 1470 -3097
rect 1554 -3473 1588 -3097
rect 1672 -3473 1706 -3097
rect 1790 -3473 1824 -3097
rect 1868 -3273 1902 -3097
rect 1986 -3273 2020 -3097
rect 4270 -3273 4304 -3097
rect 4388 -3273 4422 -3097
rect 4462 -3473 4496 -3097
rect 4580 -3473 4614 -3097
rect 4698 -3473 4732 -3097
rect 4816 -3473 4850 -3097
rect 4934 -3473 4968 -3097
rect 5012 -3273 5046 -3097
rect 5130 -3273 5164 -3097
rect 7402 -3269 7436 -3093
rect 7520 -3269 7554 -3093
rect 7594 -3469 7628 -3093
rect 7712 -3469 7746 -3093
rect 7830 -3469 7864 -3093
rect 7948 -3469 7982 -3093
rect 8066 -3469 8100 -3093
rect 8144 -3269 8178 -3093
rect 8262 -3269 8296 -3093
rect 10546 -3269 10580 -3093
rect 10664 -3269 10698 -3093
rect 10738 -3469 10772 -3093
rect 10856 -3469 10890 -3093
rect 10974 -3469 11008 -3093
rect 11092 -3469 11126 -3093
rect 11210 -3469 11244 -3093
rect 11288 -3269 11322 -3093
rect 31387 -2008 31763 -1974
rect 31387 -2126 31763 -2092
rect 31387 -2244 31763 -2210
rect 63733 -2262 63767 -1886
rect 63851 -2262 63885 -1886
rect 63969 -2262 64003 -1886
rect 64086 -2062 64120 -1886
rect 64204 -2062 64238 -1886
rect 65781 -1950 65815 -1574
rect 65899 -1950 65933 -1574
rect 66017 -1950 66051 -1574
rect 66135 -1950 66169 -1574
rect 66253 -1950 66287 -1574
rect 66659 -1750 66693 -1574
rect 66777 -1750 66811 -1574
rect 71854 -1513 72230 -1479
rect 71854 -1591 72030 -1557
rect 31387 -2362 31763 -2328
rect 71854 -1709 72030 -1675
rect 31387 -2768 31563 -2734
rect 31387 -2886 31563 -2852
rect 11406 -3269 11440 -3093
rect 13748 -3273 13782 -3097
rect 13866 -3273 13900 -3097
rect 13940 -3473 13974 -3097
rect 14058 -3473 14092 -3097
rect 14176 -3473 14210 -3097
rect 14294 -3473 14328 -3097
rect 14412 -3473 14446 -3097
rect 14490 -3273 14524 -3097
rect 14608 -3273 14642 -3097
rect 16892 -3273 16926 -3097
rect 17010 -3273 17044 -3097
rect 17084 -3473 17118 -3097
rect 17202 -3473 17236 -3097
rect 17320 -3473 17354 -3097
rect 17438 -3473 17472 -3097
rect 17556 -3473 17590 -3097
rect 17634 -3273 17668 -3097
rect 17752 -3273 17786 -3097
rect 20024 -3269 20058 -3093
rect 20142 -3269 20176 -3093
rect 20216 -3469 20250 -3093
rect 20334 -3469 20368 -3093
rect 20452 -3469 20486 -3093
rect 20570 -3469 20604 -3093
rect 20688 -3469 20722 -3093
rect 20766 -3269 20800 -3093
rect 20884 -3269 20918 -3093
rect 23168 -3269 23202 -3093
rect 23286 -3269 23320 -3093
rect 23360 -3469 23394 -3093
rect 23478 -3469 23512 -3093
rect 23596 -3469 23630 -3093
rect 23714 -3469 23748 -3093
rect 23832 -3469 23866 -3093
rect 23910 -3269 23944 -3093
rect 24028 -3269 24062 -3093
<< pdiffc >>
rect 39600 24345 39634 24521
rect 39718 24345 39752 24521
rect 39836 24345 39870 24521
rect 39954 24345 39988 24521
rect 40072 24345 40106 24521
rect 40190 24345 40224 24521
rect 40308 24345 40342 24521
rect 40426 24345 40460 24521
rect 40544 24345 40578 24521
rect 40662 24345 40696 24521
rect 41925 24217 41959 24593
rect 42043 24217 42077 24593
rect 42161 24217 42195 24593
rect 42279 24217 42313 24593
rect 42397 24217 42431 24593
rect 42515 24217 42549 24593
rect 42633 24217 42667 24593
rect 43067 24221 43101 24597
rect 43185 24221 43219 24597
rect 43303 24221 43337 24597
rect 43421 24221 43455 24597
rect 43539 24221 43573 24597
rect 43657 24221 43691 24597
rect 43775 24221 43809 24597
rect 46113 24342 46147 24518
rect 46231 24342 46265 24518
rect 46349 24342 46383 24518
rect 46467 24342 46501 24518
rect 46585 24342 46619 24518
rect 46703 24342 46737 24518
rect 46821 24342 46855 24518
rect 46939 24342 46973 24518
rect 47057 24342 47091 24518
rect 47175 24342 47209 24518
rect 48438 24214 48472 24590
rect 48556 24214 48590 24590
rect 48674 24214 48708 24590
rect 48792 24214 48826 24590
rect 48910 24214 48944 24590
rect 49028 24214 49062 24590
rect 49146 24214 49180 24590
rect 49580 24218 49614 24594
rect 49698 24218 49732 24594
rect 49816 24218 49850 24594
rect 49934 24218 49968 24594
rect 50052 24218 50086 24594
rect 50170 24218 50204 24594
rect 50288 24218 50322 24594
rect 52647 24337 52681 24513
rect 52765 24337 52799 24513
rect 52883 24337 52917 24513
rect 53001 24337 53035 24513
rect 53119 24337 53153 24513
rect 53237 24337 53271 24513
rect 53355 24337 53389 24513
rect 53473 24337 53507 24513
rect 53591 24337 53625 24513
rect 53709 24337 53743 24513
rect 42354 23634 42388 23810
rect 42472 23634 42506 23810
rect 42590 23634 42624 23810
rect 42708 23634 42742 23810
rect 43496 23638 43530 23814
rect 43614 23638 43648 23814
rect 43732 23638 43766 23814
rect 43850 23638 43884 23814
rect 54972 24209 55006 24585
rect 55090 24209 55124 24585
rect 55208 24209 55242 24585
rect 55326 24209 55360 24585
rect 55444 24209 55478 24585
rect 55562 24209 55596 24585
rect 55680 24209 55714 24585
rect 56114 24213 56148 24589
rect 56232 24213 56266 24589
rect 56350 24213 56384 24589
rect 56468 24213 56502 24589
rect 56586 24213 56620 24589
rect 56704 24213 56738 24589
rect 56822 24213 56856 24589
rect 59205 24341 59239 24517
rect 59323 24341 59357 24517
rect 59441 24341 59475 24517
rect 59559 24341 59593 24517
rect 59677 24341 59711 24517
rect 59795 24341 59829 24517
rect 59913 24341 59947 24517
rect 60031 24341 60065 24517
rect 60149 24341 60183 24517
rect 60267 24341 60301 24517
rect 48867 23631 48901 23807
rect 48985 23631 49019 23807
rect 49103 23631 49137 23807
rect 49221 23631 49255 23807
rect 50009 23635 50043 23811
rect 50127 23635 50161 23811
rect 50245 23635 50279 23811
rect 50363 23635 50397 23811
rect 61530 24213 61564 24589
rect 61648 24213 61682 24589
rect 61766 24213 61800 24589
rect 61884 24213 61918 24589
rect 62002 24213 62036 24589
rect 62120 24213 62154 24589
rect 62238 24213 62272 24589
rect 62672 24217 62706 24593
rect 62790 24217 62824 24593
rect 62908 24217 62942 24593
rect 63026 24217 63060 24593
rect 63144 24217 63178 24593
rect 63262 24217 63296 24593
rect 63380 24217 63414 24593
rect 55401 23626 55435 23802
rect 55519 23626 55553 23802
rect 55637 23626 55671 23802
rect 55755 23626 55789 23802
rect 56543 23630 56577 23806
rect 56661 23630 56695 23806
rect 56779 23630 56813 23806
rect 56897 23630 56931 23806
rect 61959 23630 61993 23806
rect 62077 23630 62111 23806
rect 62195 23630 62229 23806
rect 62313 23630 62347 23806
rect 63101 23634 63135 23810
rect 63219 23634 63253 23810
rect 63337 23634 63371 23810
rect 63455 23634 63489 23810
rect 39614 22695 39648 22871
rect 39732 22695 39766 22871
rect 39850 22695 39884 22871
rect 39968 22695 40002 22871
rect 40086 22695 40120 22871
rect 40204 22695 40238 22871
rect 40322 22695 40356 22871
rect 40440 22695 40474 22871
rect 40558 22695 40592 22871
rect 40676 22695 40710 22871
rect 46127 22692 46161 22868
rect 46245 22692 46279 22868
rect 46363 22692 46397 22868
rect 46481 22692 46515 22868
rect 46599 22692 46633 22868
rect 46717 22692 46751 22868
rect 46835 22692 46869 22868
rect 46953 22692 46987 22868
rect 47071 22692 47105 22868
rect 47189 22692 47223 22868
rect 52661 22687 52695 22863
rect 3012 21608 3046 21784
rect 3130 21608 3164 21784
rect 3248 21608 3282 21784
rect 3366 21608 3400 21784
rect 3485 21608 3519 21984
rect 3603 21608 3637 21984
rect 3721 21608 3755 21984
rect 3839 21608 3873 21984
rect 3958 21608 3992 21984
rect 4076 21608 4110 21984
rect 4194 21608 4228 21984
rect 4312 21608 4346 21984
rect 4430 21608 4464 21984
rect 4548 21608 4582 21984
rect 4666 21608 4700 21984
rect 4779 21608 4813 21984
rect 4897 21608 4931 21984
rect 5015 21608 5049 21984
rect 5133 21608 5167 21984
rect 5220 21608 5254 21784
rect 5338 21608 5372 21784
rect 5456 21608 5490 21784
rect 5574 21608 5608 21784
rect 6156 21608 6190 21784
rect 6274 21608 6308 21784
rect 6392 21608 6426 21784
rect 6510 21608 6544 21784
rect 6629 21608 6663 21984
rect 6747 21608 6781 21984
rect 6865 21608 6899 21984
rect 6983 21608 7017 21984
rect 7102 21608 7136 21984
rect 7220 21608 7254 21984
rect 7338 21608 7372 21984
rect 7456 21608 7490 21984
rect 7574 21608 7608 21984
rect 7692 21608 7726 21984
rect 7810 21608 7844 21984
rect 7923 21608 7957 21984
rect 8041 21608 8075 21984
rect 8159 21608 8193 21984
rect 8277 21608 8311 21984
rect 8364 21608 8398 21784
rect 8482 21608 8516 21784
rect 8600 21608 8634 21784
rect 8718 21608 8752 21784
rect 9288 21604 9322 21780
rect 9406 21604 9440 21780
rect 9524 21604 9558 21780
rect 9642 21604 9676 21780
rect 9761 21604 9795 21980
rect 9879 21604 9913 21980
rect 9997 21604 10031 21980
rect 10115 21604 10149 21980
rect 10234 21604 10268 21980
rect 10352 21604 10386 21980
rect 10470 21604 10504 21980
rect 10588 21604 10622 21980
rect 10706 21604 10740 21980
rect 10824 21604 10858 21980
rect 10942 21604 10976 21980
rect 11055 21604 11089 21980
rect 11173 21604 11207 21980
rect 11291 21604 11325 21980
rect 11409 21604 11443 21980
rect 11496 21604 11530 21780
rect 11614 21604 11648 21780
rect 11732 21604 11766 21780
rect 11850 21604 11884 21780
rect 12432 21604 12466 21780
rect 12550 21604 12584 21780
rect 12668 21604 12702 21780
rect 12786 21604 12820 21780
rect 12905 21604 12939 21980
rect 13023 21604 13057 21980
rect 13141 21604 13175 21980
rect 13259 21604 13293 21980
rect 13378 21604 13412 21980
rect 13496 21604 13530 21980
rect 13614 21604 13648 21980
rect 13732 21604 13766 21980
rect 13850 21604 13884 21980
rect 13968 21604 14002 21980
rect 14086 21604 14120 21980
rect 14199 21604 14233 21980
rect 14317 21604 14351 21980
rect 14435 21604 14469 21980
rect 14553 21604 14587 21980
rect 14640 21604 14674 21780
rect 14758 21604 14792 21780
rect 14876 21604 14910 21780
rect 14994 21604 15028 21780
rect 15634 21608 15668 21784
rect 15752 21608 15786 21784
rect 15870 21608 15904 21784
rect 15988 21608 16022 21784
rect 16107 21608 16141 21984
rect 16225 21608 16259 21984
rect 16343 21608 16377 21984
rect 16461 21608 16495 21984
rect 16580 21608 16614 21984
rect 16698 21608 16732 21984
rect 16816 21608 16850 21984
rect 16934 21608 16968 21984
rect 17052 21608 17086 21984
rect 17170 21608 17204 21984
rect 17288 21608 17322 21984
rect 17401 21608 17435 21984
rect 17519 21608 17553 21984
rect 17637 21608 17671 21984
rect 17755 21608 17789 21984
rect 17842 21608 17876 21784
rect 17960 21608 17994 21784
rect 18078 21608 18112 21784
rect 18196 21608 18230 21784
rect 18778 21608 18812 21784
rect 18896 21608 18930 21784
rect 19014 21608 19048 21784
rect 19132 21608 19166 21784
rect 19251 21608 19285 21984
rect 19369 21608 19403 21984
rect 19487 21608 19521 21984
rect 19605 21608 19639 21984
rect 19724 21608 19758 21984
rect 19842 21608 19876 21984
rect 19960 21608 19994 21984
rect 20078 21608 20112 21984
rect 20196 21608 20230 21984
rect 20314 21608 20348 21984
rect 20432 21608 20466 21984
rect 20545 21608 20579 21984
rect 20663 21608 20697 21984
rect 20781 21608 20815 21984
rect 20899 21608 20933 21984
rect 20986 21608 21020 21784
rect 21104 21608 21138 21784
rect 21222 21608 21256 21784
rect 21340 21608 21374 21784
rect 21910 21604 21944 21780
rect 22028 21604 22062 21780
rect 22146 21604 22180 21780
rect 22264 21604 22298 21780
rect 22383 21604 22417 21980
rect 22501 21604 22535 21980
rect 22619 21604 22653 21980
rect 22737 21604 22771 21980
rect 22856 21604 22890 21980
rect 22974 21604 23008 21980
rect 23092 21604 23126 21980
rect 23210 21604 23244 21980
rect 23328 21604 23362 21980
rect 23446 21604 23480 21980
rect 23564 21604 23598 21980
rect 23677 21604 23711 21980
rect 23795 21604 23829 21980
rect 23913 21604 23947 21980
rect 24031 21604 24065 21980
rect 24118 21604 24152 21780
rect 24236 21604 24270 21780
rect 24354 21604 24388 21780
rect 24472 21604 24506 21780
rect 25054 21604 25088 21780
rect 25172 21604 25206 21780
rect 25290 21604 25324 21780
rect 25408 21604 25442 21780
rect 25527 21604 25561 21980
rect 25645 21604 25679 21980
rect 25763 21604 25797 21980
rect 25881 21604 25915 21980
rect 26000 21604 26034 21980
rect 26118 21604 26152 21980
rect 26236 21604 26270 21980
rect 26354 21604 26388 21980
rect 26472 21604 26506 21980
rect 26590 21604 26624 21980
rect 26708 21604 26742 21980
rect 26821 21604 26855 21980
rect 26939 21604 26973 21980
rect 27057 21604 27091 21980
rect 27175 21604 27209 21980
rect 41078 22078 41112 22254
rect 41196 22078 41230 22254
rect 41314 22078 41348 22254
rect 41432 22078 41466 22254
rect 41562 22078 41596 22454
rect 41680 22078 41714 22454
rect 41798 22078 41832 22454
rect 41916 22078 41950 22454
rect 42034 22078 42068 22454
rect 42152 22078 42186 22454
rect 42270 22078 42304 22454
rect 42399 22078 42433 22254
rect 42517 22078 42551 22254
rect 42635 22078 42669 22254
rect 42753 22078 42787 22254
rect 42976 22078 43010 22254
rect 43094 22078 43128 22254
rect 43212 22078 43246 22254
rect 43330 22078 43364 22254
rect 43460 22078 43494 22454
rect 43578 22078 43612 22454
rect 43696 22078 43730 22454
rect 43814 22078 43848 22454
rect 43932 22078 43966 22454
rect 44050 22078 44084 22454
rect 44168 22078 44202 22454
rect 52779 22687 52813 22863
rect 52897 22687 52931 22863
rect 53015 22687 53049 22863
rect 53133 22687 53167 22863
rect 53251 22687 53285 22863
rect 53369 22687 53403 22863
rect 53487 22687 53521 22863
rect 53605 22687 53639 22863
rect 53723 22687 53757 22863
rect 59219 22691 59253 22867
rect 59337 22691 59371 22867
rect 59455 22691 59489 22867
rect 59573 22691 59607 22867
rect 59691 22691 59725 22867
rect 59809 22691 59843 22867
rect 59927 22691 59961 22867
rect 60045 22691 60079 22867
rect 60163 22691 60197 22867
rect 60281 22691 60315 22867
rect 44297 22078 44331 22254
rect 44415 22078 44449 22254
rect 44533 22078 44567 22254
rect 44651 22078 44685 22254
rect 27262 21604 27296 21780
rect 27380 21604 27414 21780
rect 27498 21604 27532 21780
rect 27616 21604 27650 21780
rect 39609 21091 39643 21267
rect 39727 21091 39761 21267
rect 39845 21091 39879 21267
rect 39963 21091 39997 21267
rect 40081 21091 40115 21267
rect 40199 21091 40233 21267
rect 40317 21091 40351 21267
rect 40435 21091 40469 21267
rect 40553 21091 40587 21267
rect 40671 21091 40705 21267
rect 41505 21385 41539 21761
rect 41623 21385 41657 21761
rect 41741 21385 41775 21761
rect 41859 21385 41893 21761
rect 41977 21385 42011 21761
rect 42095 21385 42129 21761
rect 42213 21385 42247 21761
rect 47591 22075 47625 22251
rect 47709 22075 47743 22251
rect 47827 22075 47861 22251
rect 47945 22075 47979 22251
rect 48075 22075 48109 22451
rect 48193 22075 48227 22451
rect 48311 22075 48345 22451
rect 48429 22075 48463 22451
rect 48547 22075 48581 22451
rect 48665 22075 48699 22451
rect 48783 22075 48817 22451
rect 48912 22075 48946 22251
rect 49030 22075 49064 22251
rect 49148 22075 49182 22251
rect 49266 22075 49300 22251
rect 49489 22075 49523 22251
rect 49607 22075 49641 22251
rect 49725 22075 49759 22251
rect 49843 22075 49877 22251
rect 49973 22075 50007 22451
rect 50091 22075 50125 22451
rect 50209 22075 50243 22451
rect 50327 22075 50361 22451
rect 50445 22075 50479 22451
rect 50563 22075 50597 22451
rect 50681 22075 50715 22451
rect 50810 22075 50844 22251
rect 50928 22075 50962 22251
rect 51046 22075 51080 22251
rect 51164 22075 51198 22251
rect 43403 21385 43437 21761
rect 43521 21385 43555 21761
rect 43639 21385 43673 21761
rect 43757 21385 43791 21761
rect 43875 21385 43909 21761
rect 43993 21385 44027 21761
rect 44111 21385 44145 21761
rect 46122 21088 46156 21264
rect 46240 21088 46274 21264
rect 46358 21088 46392 21264
rect 46476 21088 46510 21264
rect 46594 21088 46628 21264
rect 46712 21088 46746 21264
rect 46830 21088 46864 21264
rect 46948 21088 46982 21264
rect 47066 21088 47100 21264
rect 47184 21088 47218 21264
rect 48018 21382 48052 21758
rect 48136 21382 48170 21758
rect 48254 21382 48288 21758
rect 48372 21382 48406 21758
rect 48490 21382 48524 21758
rect 48608 21382 48642 21758
rect 48726 21382 48760 21758
rect 54125 22070 54159 22246
rect 54243 22070 54277 22246
rect 54361 22070 54395 22246
rect 54479 22070 54513 22246
rect 54609 22070 54643 22446
rect 54727 22070 54761 22446
rect 54845 22070 54879 22446
rect 54963 22070 54997 22446
rect 55081 22070 55115 22446
rect 55199 22070 55233 22446
rect 55317 22070 55351 22446
rect 55446 22070 55480 22246
rect 55564 22070 55598 22246
rect 55682 22070 55716 22246
rect 55800 22070 55834 22246
rect 56023 22070 56057 22246
rect 56141 22070 56175 22246
rect 56259 22070 56293 22246
rect 56377 22070 56411 22246
rect 56507 22070 56541 22446
rect 56625 22070 56659 22446
rect 56743 22070 56777 22446
rect 56861 22070 56895 22446
rect 56979 22070 57013 22446
rect 57097 22070 57131 22446
rect 57215 22070 57249 22446
rect 57344 22070 57378 22246
rect 57462 22070 57496 22246
rect 57580 22070 57614 22246
rect 57698 22070 57732 22246
rect 49916 21382 49950 21758
rect 50034 21382 50068 21758
rect 50152 21382 50186 21758
rect 50270 21382 50304 21758
rect 50388 21382 50422 21758
rect 50506 21382 50540 21758
rect 50624 21382 50658 21758
rect 52656 21083 52690 21259
rect 52774 21083 52808 21259
rect 52892 21083 52926 21259
rect 53010 21083 53044 21259
rect 53128 21083 53162 21259
rect 53246 21083 53280 21259
rect 53364 21083 53398 21259
rect 53482 21083 53516 21259
rect 53600 21083 53634 21259
rect 53718 21083 53752 21259
rect 54552 21377 54586 21753
rect 54670 21377 54704 21753
rect 54788 21377 54822 21753
rect 54906 21377 54940 21753
rect 55024 21377 55058 21753
rect 55142 21377 55176 21753
rect 55260 21377 55294 21753
rect 60683 22074 60717 22250
rect 60801 22074 60835 22250
rect 60919 22074 60953 22250
rect 61037 22074 61071 22250
rect 61167 22074 61201 22450
rect 61285 22074 61319 22450
rect 61403 22074 61437 22450
rect 61521 22074 61555 22450
rect 61639 22074 61673 22450
rect 61757 22074 61791 22450
rect 61875 22074 61909 22450
rect 62004 22074 62038 22250
rect 62122 22074 62156 22250
rect 62240 22074 62274 22250
rect 62358 22074 62392 22250
rect 62581 22074 62615 22250
rect 62699 22074 62733 22250
rect 62817 22074 62851 22250
rect 62935 22074 62969 22250
rect 63065 22074 63099 22450
rect 63183 22074 63217 22450
rect 63301 22074 63335 22450
rect 63419 22074 63453 22450
rect 63537 22074 63571 22450
rect 63655 22074 63689 22450
rect 63773 22074 63807 22450
rect 63902 22074 63936 22250
rect 64020 22074 64054 22250
rect 64138 22074 64172 22250
rect 64256 22074 64290 22250
rect 56450 21377 56484 21753
rect 56568 21377 56602 21753
rect 56686 21377 56720 21753
rect 56804 21377 56838 21753
rect 56922 21377 56956 21753
rect 57040 21377 57074 21753
rect 57158 21377 57192 21753
rect 59214 21087 59248 21263
rect 59332 21087 59366 21263
rect 59450 21087 59484 21263
rect 59568 21087 59602 21263
rect 59686 21087 59720 21263
rect 59804 21087 59838 21263
rect 59922 21087 59956 21263
rect 60040 21087 60074 21263
rect 60158 21087 60192 21263
rect 60276 21087 60310 21263
rect 61110 21381 61144 21757
rect 61228 21381 61262 21757
rect 61346 21381 61380 21757
rect 61464 21381 61498 21757
rect 61582 21381 61616 21757
rect 61700 21381 61734 21757
rect 61818 21381 61852 21757
rect 70725 22027 70901 22061
rect 70725 21909 70901 21943
rect 63008 21381 63042 21757
rect 63126 21381 63160 21757
rect 63244 21381 63278 21757
rect 63362 21381 63396 21757
rect 63480 21381 63514 21757
rect 63598 21381 63632 21757
rect 63716 21381 63750 21757
rect 70725 21791 70901 21825
rect 70725 21673 70901 21707
rect 70525 21586 70901 21620
rect 70525 21468 70901 21502
rect 70525 21350 70901 21384
rect 70525 21232 70901 21266
rect 70525 21119 70901 21153
rect 70525 21001 70901 21035
rect 70525 20883 70901 20917
rect 70525 20765 70901 20799
rect 70525 20647 70901 20681
rect 70525 20529 70901 20563
rect 70525 20411 70901 20445
rect 70525 20292 70901 20326
rect 70525 20174 70901 20208
rect 70525 20056 70901 20090
rect 70525 19938 70901 19972
rect 70725 19819 70901 19853
rect 70725 19701 70901 19735
rect 70725 19583 70901 19617
rect 70725 19465 70901 19499
rect 39611 18613 39645 18989
rect 39729 18613 39763 18989
rect 39847 18613 39881 18989
rect 39965 18613 39999 18989
rect 40083 18613 40117 18989
rect 40201 18613 40235 18989
rect 40319 18613 40353 18989
rect 40753 18609 40787 18985
rect 40871 18609 40905 18985
rect 40989 18609 41023 18985
rect 41107 18609 41141 18985
rect 41225 18609 41259 18985
rect 41343 18609 41377 18985
rect 41461 18609 41495 18985
rect 42724 18737 42758 18913
rect 42842 18737 42876 18913
rect 42960 18737 42994 18913
rect 43078 18737 43112 18913
rect 43196 18737 43230 18913
rect 43314 18737 43348 18913
rect 43432 18737 43466 18913
rect 43550 18737 43584 18913
rect 43668 18737 43702 18913
rect 43786 18737 43820 18913
rect 46169 18609 46203 18985
rect 46287 18609 46321 18985
rect 46405 18609 46439 18985
rect 46523 18609 46557 18985
rect 46641 18609 46675 18985
rect 46759 18609 46793 18985
rect 46877 18609 46911 18985
rect 47311 18605 47345 18981
rect 39536 18030 39570 18206
rect 39654 18030 39688 18206
rect 39772 18030 39806 18206
rect 39890 18030 39924 18206
rect 40678 18026 40712 18202
rect 40796 18026 40830 18202
rect 40914 18026 40948 18202
rect 41032 18026 41066 18202
rect 47429 18605 47463 18981
rect 47547 18605 47581 18981
rect 47665 18605 47699 18981
rect 47783 18605 47817 18981
rect 47901 18605 47935 18981
rect 48019 18605 48053 18981
rect 49282 18733 49316 18909
rect 49400 18733 49434 18909
rect 49518 18733 49552 18909
rect 49636 18733 49670 18909
rect 49754 18733 49788 18909
rect 49872 18733 49906 18909
rect 49990 18733 50024 18909
rect 50108 18733 50142 18909
rect 50226 18733 50260 18909
rect 50344 18733 50378 18909
rect 52703 18614 52737 18990
rect 52821 18614 52855 18990
rect 52939 18614 52973 18990
rect 53057 18614 53091 18990
rect 53175 18614 53209 18990
rect 53293 18614 53327 18990
rect 53411 18614 53445 18990
rect 53845 18610 53879 18986
rect 46094 18026 46128 18202
rect 46212 18026 46246 18202
rect 46330 18026 46364 18202
rect 46448 18026 46482 18202
rect 47236 18022 47270 18198
rect 47354 18022 47388 18198
rect 47472 18022 47506 18198
rect 47590 18022 47624 18198
rect 53963 18610 53997 18986
rect 54081 18610 54115 18986
rect 54199 18610 54233 18986
rect 54317 18610 54351 18986
rect 54435 18610 54469 18986
rect 54553 18610 54587 18986
rect 55816 18738 55850 18914
rect 55934 18738 55968 18914
rect 56052 18738 56086 18914
rect 56170 18738 56204 18914
rect 56288 18738 56322 18914
rect 56406 18738 56440 18914
rect 56524 18738 56558 18914
rect 56642 18738 56676 18914
rect 56760 18738 56794 18914
rect 56878 18738 56912 18914
rect 59216 18617 59250 18993
rect 59334 18617 59368 18993
rect 59452 18617 59486 18993
rect 59570 18617 59604 18993
rect 59688 18617 59722 18993
rect 59806 18617 59840 18993
rect 59924 18617 59958 18993
rect 60358 18613 60392 18989
rect 52628 18031 52662 18207
rect 52746 18031 52780 18207
rect 52864 18031 52898 18207
rect 52982 18031 53016 18207
rect 53770 18027 53804 18203
rect 53888 18027 53922 18203
rect 54006 18027 54040 18203
rect 54124 18027 54158 18203
rect 60476 18613 60510 18989
rect 60594 18613 60628 18989
rect 60712 18613 60746 18989
rect 60830 18613 60864 18989
rect 60948 18613 60982 18989
rect 61066 18613 61100 18989
rect 62329 18741 62363 18917
rect 62447 18741 62481 18917
rect 62565 18741 62599 18917
rect 62683 18741 62717 18917
rect 62801 18741 62835 18917
rect 62919 18741 62953 18917
rect 63037 18741 63071 18917
rect 63155 18741 63189 18917
rect 63273 18741 63307 18917
rect 63391 18741 63425 18917
rect 70725 18883 70901 18917
rect 70725 18765 70901 18799
rect 70725 18647 70901 18681
rect 70725 18529 70901 18563
rect 59141 18034 59175 18210
rect 59259 18034 59293 18210
rect 59377 18034 59411 18210
rect 59495 18034 59529 18210
rect 60283 18030 60317 18206
rect 60401 18030 60435 18206
rect 60519 18030 60553 18206
rect 60637 18030 60671 18206
rect 70525 18442 70901 18476
rect 70525 18324 70901 18358
rect 70525 18206 70901 18240
rect 70525 18088 70901 18122
rect 70525 17975 70901 18009
rect 70525 17857 70901 17891
rect 70525 17739 70901 17773
rect 70525 17621 70901 17655
rect 70525 17503 70901 17537
rect 42710 17087 42744 17263
rect 4520 16420 4554 16796
rect 4638 16420 4672 16796
rect 4756 16420 4790 16796
rect 4874 16420 4908 16796
rect 4992 16420 5026 16796
rect 5110 16420 5144 16796
rect 5228 16420 5262 16796
rect 5688 16422 5722 16798
rect 5806 16422 5840 16798
rect 5924 16422 5958 16798
rect 6042 16422 6076 16798
rect 6160 16422 6194 16798
rect 6278 16422 6312 16798
rect 42828 17087 42862 17263
rect 42946 17087 42980 17263
rect 43064 17087 43098 17263
rect 43182 17087 43216 17263
rect 43300 17087 43334 17263
rect 43418 17087 43452 17263
rect 43536 17087 43570 17263
rect 43654 17087 43688 17263
rect 43772 17087 43806 17263
rect 49268 17083 49302 17259
rect 49386 17083 49420 17259
rect 49504 17083 49538 17259
rect 49622 17083 49656 17259
rect 49740 17083 49774 17259
rect 49858 17083 49892 17259
rect 49976 17083 50010 17259
rect 50094 17083 50128 17259
rect 50212 17083 50246 17259
rect 50330 17083 50364 17259
rect 55802 17088 55836 17264
rect 55920 17088 55954 17264
rect 56038 17088 56072 17264
rect 56156 17088 56190 17264
rect 56274 17088 56308 17264
rect 56392 17088 56426 17264
rect 56510 17088 56544 17264
rect 56628 17088 56662 17264
rect 56746 17088 56780 17264
rect 56864 17088 56898 17264
rect 70525 17385 70901 17419
rect 62315 17091 62349 17267
rect 62433 17091 62467 17267
rect 62551 17091 62585 17267
rect 62669 17091 62703 17267
rect 62787 17091 62821 17267
rect 62905 17091 62939 17267
rect 63023 17091 63057 17267
rect 63141 17091 63175 17267
rect 63259 17091 63293 17267
rect 63377 17091 63411 17267
rect 70525 17267 70901 17301
rect 70525 17148 70901 17182
rect 6396 16422 6430 16798
rect 6856 16420 6890 16796
rect 6974 16420 7008 16796
rect 7092 16420 7126 16796
rect 7210 16420 7244 16796
rect 7328 16420 7362 16796
rect 7446 16420 7480 16796
rect 7564 16420 7598 16796
rect 8024 16422 8058 16798
rect 8142 16422 8176 16798
rect 8260 16422 8294 16798
rect 8378 16422 8412 16798
rect 8496 16422 8530 16798
rect 8614 16422 8648 16798
rect 8732 16422 8766 16798
rect 9198 16420 9232 16796
rect 4445 15832 4479 16008
rect 4563 15832 4597 16008
rect 4681 15832 4715 16008
rect 4799 15832 4833 16008
rect 5613 15831 5647 16007
rect 5731 15831 5765 16007
rect 5849 15831 5883 16007
rect 5967 15831 6001 16007
rect 9316 16420 9350 16796
rect 9434 16420 9468 16796
rect 9552 16420 9586 16796
rect 9670 16420 9704 16796
rect 9788 16420 9822 16796
rect 9906 16420 9940 16796
rect 10366 16418 10400 16794
rect 6781 15831 6815 16007
rect 6899 15831 6933 16007
rect 7017 15831 7051 16007
rect 7135 15831 7169 16007
rect 10484 16418 10518 16794
rect 10602 16418 10636 16794
rect 10720 16418 10754 16794
rect 10838 16418 10872 16794
rect 10956 16418 10990 16794
rect 11074 16418 11108 16794
rect 11534 16420 11568 16796
rect 11652 16420 11686 16796
rect 11770 16420 11804 16796
rect 11888 16420 11922 16796
rect 12006 16420 12040 16796
rect 12124 16420 12158 16796
rect 12242 16420 12276 16796
rect 12702 16420 12736 16796
rect 12820 16420 12854 16796
rect 12938 16420 12972 16796
rect 13056 16420 13090 16796
rect 13174 16420 13208 16796
rect 13292 16420 13326 16796
rect 13410 16420 13444 16796
rect 13803 16425 13837 16601
rect 13921 16425 13955 16601
rect 14039 16425 14073 16601
rect 14157 16425 14191 16601
rect 14275 16425 14309 16601
rect 14393 16425 14427 16601
rect 14511 16425 14545 16601
rect 14629 16425 14663 16601
rect 14747 16425 14781 16601
rect 14865 16425 14899 16601
rect 15251 16425 15285 16601
rect 15369 16425 15403 16601
rect 15487 16425 15521 16601
rect 15605 16425 15639 16601
rect 15723 16425 15757 16601
rect 15841 16425 15875 16601
rect 15959 16425 15993 16601
rect 16077 16425 16111 16601
rect 16195 16425 16229 16601
rect 16313 16425 16347 16601
rect 16749 16423 16783 16599
rect 7950 15832 7984 16008
rect 8068 15832 8102 16008
rect 8186 15832 8220 16008
rect 8304 15832 8338 16008
rect 9122 15836 9156 16012
rect 9240 15836 9274 16012
rect 9358 15836 9392 16012
rect 9476 15836 9510 16012
rect 10291 15836 10325 16012
rect 10409 15836 10443 16012
rect 10527 15836 10561 16012
rect 10645 15836 10679 16012
rect 11459 15836 11493 16012
rect 11577 15836 11611 16012
rect 11695 15836 11729 16012
rect 11813 15836 11847 16012
rect 16867 16423 16901 16599
rect 16985 16423 17019 16599
rect 17103 16423 17137 16599
rect 17221 16423 17255 16599
rect 17339 16423 17373 16599
rect 17457 16423 17491 16599
rect 17575 16423 17609 16599
rect 17693 16423 17727 16599
rect 17811 16423 17845 16599
rect 18197 16423 18231 16599
rect 18315 16423 18349 16599
rect 18433 16423 18467 16599
rect 18551 16423 18585 16599
rect 18669 16423 18703 16599
rect 18787 16423 18821 16599
rect 18905 16423 18939 16599
rect 19023 16423 19057 16599
rect 19141 16423 19175 16599
rect 19259 16423 19293 16599
rect 19717 16425 19751 16601
rect 19835 16425 19869 16601
rect 19953 16425 19987 16601
rect 20071 16425 20105 16601
rect 20189 16425 20223 16601
rect 20307 16425 20341 16601
rect 20425 16425 20459 16601
rect 20543 16425 20577 16601
rect 20661 16425 20695 16601
rect 20779 16425 20813 16601
rect 21165 16425 21199 16601
rect 21283 16425 21317 16601
rect 21401 16425 21435 16601
rect 21519 16425 21553 16601
rect 21637 16425 21671 16601
rect 21755 16425 21789 16601
rect 21873 16425 21907 16601
rect 21991 16425 22025 16601
rect 22109 16425 22143 16601
rect 22227 16425 22261 16601
rect 22663 16423 22697 16599
rect 12626 15830 12660 16006
rect 12744 15830 12778 16006
rect 12862 15830 12896 16006
rect 12980 15830 13014 16006
rect 22781 16423 22815 16599
rect 22899 16423 22933 16599
rect 23017 16423 23051 16599
rect 23135 16423 23169 16599
rect 23253 16423 23287 16599
rect 23371 16423 23405 16599
rect 23489 16423 23523 16599
rect 23607 16423 23641 16599
rect 23725 16423 23759 16599
rect 24111 16423 24145 16599
rect 24229 16423 24263 16599
rect 24347 16423 24381 16599
rect 24465 16423 24499 16599
rect 24583 16423 24617 16599
rect 24701 16423 24735 16599
rect 24819 16423 24853 16599
rect 24937 16423 24971 16599
rect 25055 16423 25089 16599
rect 25173 16423 25207 16599
rect 38735 16470 38769 16646
rect 38853 16470 38887 16646
rect 38971 16470 39005 16646
rect 39089 16470 39123 16646
rect 39218 16470 39252 16846
rect 39336 16470 39370 16846
rect 39454 16470 39488 16846
rect 39572 16470 39606 16846
rect 39690 16470 39724 16846
rect 39808 16470 39842 16846
rect 39926 16470 39960 16846
rect 40056 16470 40090 16646
rect 40174 16470 40208 16646
rect 40292 16470 40326 16646
rect 40410 16470 40444 16646
rect 40633 16470 40667 16646
rect 40751 16470 40785 16646
rect 40869 16470 40903 16646
rect 40987 16470 41021 16646
rect 41116 16470 41150 16846
rect 41234 16470 41268 16846
rect 41352 16470 41386 16846
rect 41470 16470 41504 16846
rect 41588 16470 41622 16846
rect 41706 16470 41740 16846
rect 41824 16470 41858 16846
rect 41954 16470 41988 16646
rect 42072 16470 42106 16646
rect 42190 16470 42224 16646
rect 42308 16470 42342 16646
rect 39275 15777 39309 16153
rect 39393 15777 39427 16153
rect 39511 15777 39545 16153
rect 39629 15777 39663 16153
rect 39747 15777 39781 16153
rect 39865 15777 39899 16153
rect 39983 15777 40017 16153
rect 45293 16466 45327 16642
rect 45411 16466 45445 16642
rect 45529 16466 45563 16642
rect 45647 16466 45681 16642
rect 45776 16466 45810 16842
rect 45894 16466 45928 16842
rect 46012 16466 46046 16842
rect 46130 16466 46164 16842
rect 46248 16466 46282 16842
rect 46366 16466 46400 16842
rect 46484 16466 46518 16842
rect 46614 16466 46648 16642
rect 46732 16466 46766 16642
rect 46850 16466 46884 16642
rect 46968 16466 47002 16642
rect 47191 16466 47225 16642
rect 47309 16466 47343 16642
rect 47427 16466 47461 16642
rect 47545 16466 47579 16642
rect 47674 16466 47708 16842
rect 47792 16466 47826 16842
rect 47910 16466 47944 16842
rect 48028 16466 48062 16842
rect 48146 16466 48180 16842
rect 48264 16466 48298 16842
rect 48382 16466 48416 16842
rect 48512 16466 48546 16642
rect 48630 16466 48664 16642
rect 48748 16466 48782 16642
rect 48866 16466 48900 16642
rect 41173 15777 41207 16153
rect 41291 15777 41325 16153
rect 41409 15777 41443 16153
rect 41527 15777 41561 16153
rect 41645 15777 41679 16153
rect 41763 15777 41797 16153
rect 41881 15777 41915 16153
rect 42715 15483 42749 15659
rect 42833 15483 42867 15659
rect 42951 15483 42985 15659
rect 43069 15483 43103 15659
rect 43187 15483 43221 15659
rect 43305 15483 43339 15659
rect 43423 15483 43457 15659
rect 43541 15483 43575 15659
rect 43659 15483 43693 15659
rect 43777 15483 43811 15659
rect 45833 15773 45867 16149
rect 45951 15773 45985 16149
rect 46069 15773 46103 16149
rect 46187 15773 46221 16149
rect 46305 15773 46339 16149
rect 46423 15773 46457 16149
rect 46541 15773 46575 16149
rect 51827 16471 51861 16647
rect 51945 16471 51979 16647
rect 52063 16471 52097 16647
rect 52181 16471 52215 16647
rect 52310 16471 52344 16847
rect 52428 16471 52462 16847
rect 52546 16471 52580 16847
rect 52664 16471 52698 16847
rect 52782 16471 52816 16847
rect 52900 16471 52934 16847
rect 53018 16471 53052 16847
rect 53148 16471 53182 16647
rect 53266 16471 53300 16647
rect 53384 16471 53418 16647
rect 53502 16471 53536 16647
rect 53725 16471 53759 16647
rect 53843 16471 53877 16647
rect 53961 16471 53995 16647
rect 54079 16471 54113 16647
rect 54208 16471 54242 16847
rect 54326 16471 54360 16847
rect 54444 16471 54478 16847
rect 54562 16471 54596 16847
rect 54680 16471 54714 16847
rect 54798 16471 54832 16847
rect 54916 16471 54950 16847
rect 55046 16471 55080 16647
rect 55164 16471 55198 16647
rect 55282 16471 55316 16647
rect 55400 16471 55434 16647
rect 47731 15773 47765 16149
rect 47849 15773 47883 16149
rect 47967 15773 48001 16149
rect 48085 15773 48119 16149
rect 48203 15773 48237 16149
rect 48321 15773 48355 16149
rect 48439 15773 48473 16149
rect 49273 15479 49307 15655
rect 49391 15479 49425 15655
rect 49509 15479 49543 15655
rect 49627 15479 49661 15655
rect 49745 15479 49779 15655
rect 49863 15479 49897 15655
rect 49981 15479 50015 15655
rect 50099 15479 50133 15655
rect 50217 15479 50251 15655
rect 50335 15479 50369 15655
rect 52367 15778 52401 16154
rect 52485 15778 52519 16154
rect 52603 15778 52637 16154
rect 52721 15778 52755 16154
rect 52839 15778 52873 16154
rect 52957 15778 52991 16154
rect 53075 15778 53109 16154
rect 510 14470 544 14646
rect 628 14470 662 14646
rect 746 14470 780 14646
rect 864 14470 898 14646
rect 983 14470 1017 14846
rect 1101 14470 1135 14846
rect 1219 14470 1253 14846
rect 1337 14470 1371 14846
rect 1456 14470 1490 14846
rect 1574 14470 1608 14846
rect 1692 14470 1726 14846
rect 1810 14470 1844 14846
rect 1928 14470 1962 14846
rect 2046 14470 2080 14846
rect 2164 14470 2198 14846
rect 2277 14470 2311 14846
rect 2395 14470 2429 14846
rect 2513 14470 2547 14846
rect 2631 14470 2665 14846
rect 2718 14470 2752 14646
rect 2836 14470 2870 14646
rect 2954 14470 2988 14646
rect 3072 14470 3106 14646
rect 3654 14470 3688 14646
rect 3772 14470 3806 14646
rect 3890 14470 3924 14646
rect 4008 14470 4042 14646
rect 4127 14470 4161 14846
rect 4245 14470 4279 14846
rect 4363 14470 4397 14846
rect 4481 14470 4515 14846
rect 4600 14470 4634 14846
rect 4718 14470 4752 14846
rect 4836 14470 4870 14846
rect 4954 14470 4988 14846
rect 5072 14470 5106 14846
rect 5190 14470 5224 14846
rect 5308 14470 5342 14846
rect 5421 14470 5455 14846
rect 5539 14470 5573 14846
rect 5657 14470 5691 14846
rect 5775 14470 5809 14846
rect 5862 14470 5896 14646
rect 5980 14470 6014 14646
rect 6098 14470 6132 14646
rect 6216 14470 6250 14646
rect 6786 14466 6820 14642
rect 6904 14466 6938 14642
rect 7022 14466 7056 14642
rect 7140 14466 7174 14642
rect 7259 14466 7293 14842
rect 7377 14466 7411 14842
rect 7495 14466 7529 14842
rect 7613 14466 7647 14842
rect 7732 14466 7766 14842
rect 7850 14466 7884 14842
rect 7968 14466 8002 14842
rect 8086 14466 8120 14842
rect 8204 14466 8238 14842
rect 8322 14466 8356 14842
rect 8440 14466 8474 14842
rect 8553 14466 8587 14842
rect 8671 14466 8705 14842
rect 8789 14466 8823 14842
rect 8907 14466 8941 14842
rect 8994 14466 9028 14642
rect 9112 14466 9146 14642
rect 9230 14466 9264 14642
rect 9348 14466 9382 14642
rect 9930 14466 9964 14642
rect 10048 14466 10082 14642
rect 10166 14466 10200 14642
rect 10284 14466 10318 14642
rect 10403 14466 10437 14842
rect 10521 14466 10555 14842
rect 10639 14466 10673 14842
rect 10757 14466 10791 14842
rect 10876 14466 10910 14842
rect 10994 14466 11028 14842
rect 11112 14466 11146 14842
rect 11230 14466 11264 14842
rect 11348 14466 11382 14842
rect 11466 14466 11500 14842
rect 11584 14466 11618 14842
rect 11697 14466 11731 14842
rect 11815 14466 11849 14842
rect 11933 14466 11967 14842
rect 12051 14466 12085 14842
rect 12138 14466 12172 14642
rect 12256 14466 12290 14642
rect 12374 14466 12408 14642
rect 12492 14466 12526 14642
rect 13132 14470 13166 14646
rect 13250 14470 13284 14646
rect 13368 14470 13402 14646
rect 13486 14470 13520 14646
rect 13605 14470 13639 14846
rect 13723 14470 13757 14846
rect 13841 14470 13875 14846
rect 13959 14470 13993 14846
rect 14078 14470 14112 14846
rect 14196 14470 14230 14846
rect 14314 14470 14348 14846
rect 14432 14470 14466 14846
rect 14550 14470 14584 14846
rect 14668 14470 14702 14846
rect 14786 14470 14820 14846
rect 14899 14470 14933 14846
rect 15017 14470 15051 14846
rect 15135 14470 15169 14846
rect 15253 14470 15287 14846
rect 15340 14470 15374 14646
rect 15458 14470 15492 14646
rect 15576 14470 15610 14646
rect 15694 14470 15728 14646
rect 16276 14470 16310 14646
rect 16394 14470 16428 14646
rect 16512 14470 16546 14646
rect 16630 14470 16664 14646
rect 16749 14470 16783 14846
rect 16867 14470 16901 14846
rect 16985 14470 17019 14846
rect 17103 14470 17137 14846
rect 17222 14470 17256 14846
rect 17340 14470 17374 14846
rect 17458 14470 17492 14846
rect 17576 14470 17610 14846
rect 17694 14470 17728 14846
rect 17812 14470 17846 14846
rect 17930 14470 17964 14846
rect 18043 14470 18077 14846
rect 18161 14470 18195 14846
rect 18279 14470 18313 14846
rect 18397 14470 18431 14846
rect 18484 14470 18518 14646
rect 18602 14470 18636 14646
rect 18720 14470 18754 14646
rect 18838 14470 18872 14646
rect 19408 14466 19442 14642
rect 19526 14466 19560 14642
rect 19644 14466 19678 14642
rect 19762 14466 19796 14642
rect 19881 14466 19915 14842
rect 19999 14466 20033 14842
rect 20117 14466 20151 14842
rect 20235 14466 20269 14842
rect 20354 14466 20388 14842
rect 20472 14466 20506 14842
rect 20590 14466 20624 14842
rect 20708 14466 20742 14842
rect 20826 14466 20860 14842
rect 20944 14466 20978 14842
rect 21062 14466 21096 14842
rect 21175 14466 21209 14842
rect 21293 14466 21327 14842
rect 21411 14466 21445 14842
rect 21529 14466 21563 14842
rect 21616 14466 21650 14642
rect 21734 14466 21768 14642
rect 21852 14466 21886 14642
rect 21970 14466 22004 14642
rect 22552 14466 22586 14642
rect 22670 14466 22704 14642
rect 22788 14466 22822 14642
rect 22906 14466 22940 14642
rect 23025 14466 23059 14842
rect 23143 14466 23177 14842
rect 23261 14466 23295 14842
rect 23379 14466 23413 14842
rect 23498 14466 23532 14842
rect 23616 14466 23650 14842
rect 23734 14466 23768 14842
rect 23852 14466 23886 14842
rect 23970 14466 24004 14842
rect 24088 14466 24122 14842
rect 24206 14466 24240 14842
rect 24319 14466 24353 14842
rect 24437 14466 24471 14842
rect 24555 14466 24589 14842
rect 24673 14466 24707 14842
rect 58340 16474 58374 16650
rect 58458 16474 58492 16650
rect 58576 16474 58610 16650
rect 58694 16474 58728 16650
rect 58823 16474 58857 16850
rect 58941 16474 58975 16850
rect 59059 16474 59093 16850
rect 59177 16474 59211 16850
rect 59295 16474 59329 16850
rect 59413 16474 59447 16850
rect 59531 16474 59565 16850
rect 59661 16474 59695 16650
rect 59779 16474 59813 16650
rect 59897 16474 59931 16650
rect 60015 16474 60049 16650
rect 60238 16474 60272 16650
rect 60356 16474 60390 16650
rect 60474 16474 60508 16650
rect 60592 16474 60626 16650
rect 60721 16474 60755 16850
rect 60839 16474 60873 16850
rect 60957 16474 60991 16850
rect 61075 16474 61109 16850
rect 61193 16474 61227 16850
rect 61311 16474 61345 16850
rect 61429 16474 61463 16850
rect 70525 17030 70901 17064
rect 70525 16912 70901 16946
rect 61559 16474 61593 16650
rect 61677 16474 61711 16650
rect 61795 16474 61829 16650
rect 61913 16474 61947 16650
rect 54265 15778 54299 16154
rect 54383 15778 54417 16154
rect 54501 15778 54535 16154
rect 54619 15778 54653 16154
rect 54737 15778 54771 16154
rect 54855 15778 54889 16154
rect 54973 15778 55007 16154
rect 55807 15484 55841 15660
rect 55925 15484 55959 15660
rect 56043 15484 56077 15660
rect 56161 15484 56195 15660
rect 56279 15484 56313 15660
rect 56397 15484 56431 15660
rect 56515 15484 56549 15660
rect 56633 15484 56667 15660
rect 56751 15484 56785 15660
rect 56869 15484 56903 15660
rect 58880 15781 58914 16157
rect 58998 15781 59032 16157
rect 59116 15781 59150 16157
rect 59234 15781 59268 16157
rect 59352 15781 59386 16157
rect 59470 15781 59504 16157
rect 59588 15781 59622 16157
rect 70525 16794 70901 16828
rect 70725 16675 70901 16709
rect 70725 16557 70901 16591
rect 70725 16439 70901 16473
rect 70725 16321 70901 16355
rect 60778 15781 60812 16157
rect 60896 15781 60930 16157
rect 61014 15781 61048 16157
rect 61132 15781 61166 16157
rect 61250 15781 61284 16157
rect 61368 15781 61402 16157
rect 61486 15781 61520 16157
rect 70721 15751 70897 15785
rect 62320 15487 62354 15663
rect 62438 15487 62472 15663
rect 62556 15487 62590 15663
rect 62674 15487 62708 15663
rect 62792 15487 62826 15663
rect 62910 15487 62944 15663
rect 63028 15487 63062 15663
rect 63146 15487 63180 15663
rect 63264 15487 63298 15663
rect 63382 15487 63416 15663
rect 70721 15633 70897 15667
rect 70721 15515 70897 15549
rect 24760 14466 24794 14642
rect 24878 14466 24912 14642
rect 24996 14466 25030 14642
rect 25114 14466 25148 14642
rect 70721 15397 70897 15431
rect 70521 15310 70897 15344
rect 70521 15192 70897 15226
rect 70521 15074 70897 15108
rect 70521 14956 70897 14990
rect 70521 14843 70897 14877
rect 70521 14725 70897 14759
rect 70521 14607 70897 14641
rect 70521 14489 70897 14523
rect 70521 14371 70897 14405
rect 70521 14253 70897 14287
rect 70521 14135 70897 14169
rect 70521 14016 70897 14050
rect 70521 13898 70897 13932
rect 70521 13780 70897 13814
rect 70521 13662 70897 13696
rect 70721 13543 70897 13577
rect 70721 13425 70897 13459
rect 70721 13307 70897 13341
rect 70721 13189 70897 13223
rect 30166 13134 30342 13168
rect 30166 13016 30342 13050
rect 30166 12898 30342 12932
rect 30166 12780 30342 12814
rect 29966 12650 30342 12684
rect 30659 12707 31035 12741
rect 29966 12532 30342 12566
rect 30659 12589 31035 12623
rect 70721 12607 70897 12641
rect 29966 12414 30342 12448
rect 30659 12471 31035 12505
rect 70721 12489 70897 12523
rect 30659 12353 31035 12387
rect 29966 12296 30342 12330
rect 510 11736 544 11912
rect 628 11736 662 11912
rect 746 11736 780 11912
rect 864 11736 898 11912
rect 983 11736 1017 12112
rect 1101 11736 1135 12112
rect 1219 11736 1253 12112
rect 1337 11736 1371 12112
rect 1456 11736 1490 12112
rect 1574 11736 1608 12112
rect 1692 11736 1726 12112
rect 1810 11736 1844 12112
rect 1928 11736 1962 12112
rect 2046 11736 2080 12112
rect 2164 11736 2198 12112
rect 2277 11736 2311 12112
rect 2395 11736 2429 12112
rect 2513 11736 2547 12112
rect 2631 11736 2665 12112
rect 2718 11736 2752 11912
rect 2836 11736 2870 11912
rect 2954 11736 2988 11912
rect 3072 11736 3106 11912
rect 3654 11736 3688 11912
rect 3772 11736 3806 11912
rect 3890 11736 3924 11912
rect 4008 11736 4042 11912
rect 4127 11736 4161 12112
rect 4245 11736 4279 12112
rect 4363 11736 4397 12112
rect 4481 11736 4515 12112
rect 4600 11736 4634 12112
rect 4718 11736 4752 12112
rect 4836 11736 4870 12112
rect 4954 11736 4988 12112
rect 5072 11736 5106 12112
rect 5190 11736 5224 12112
rect 5308 11736 5342 12112
rect 5421 11736 5455 12112
rect 5539 11736 5573 12112
rect 5657 11736 5691 12112
rect 5775 11736 5809 12112
rect 5862 11736 5896 11912
rect 5980 11736 6014 11912
rect 6098 11736 6132 11912
rect 6216 11736 6250 11912
rect 6786 11732 6820 11908
rect 6904 11732 6938 11908
rect 7022 11732 7056 11908
rect 7140 11732 7174 11908
rect 7259 11732 7293 12108
rect 7377 11732 7411 12108
rect 7495 11732 7529 12108
rect 7613 11732 7647 12108
rect 7732 11732 7766 12108
rect 7850 11732 7884 12108
rect 7968 11732 8002 12108
rect 8086 11732 8120 12108
rect 8204 11732 8238 12108
rect 8322 11732 8356 12108
rect 8440 11732 8474 12108
rect 8553 11732 8587 12108
rect 8671 11732 8705 12108
rect 8789 11732 8823 12108
rect 8907 11732 8941 12108
rect 8994 11732 9028 11908
rect 9112 11732 9146 11908
rect 9230 11732 9264 11908
rect 9348 11732 9382 11908
rect 9930 11732 9964 11908
rect 10048 11732 10082 11908
rect 10166 11732 10200 11908
rect 10284 11732 10318 11908
rect 10403 11732 10437 12108
rect 10521 11732 10555 12108
rect 10639 11732 10673 12108
rect 10757 11732 10791 12108
rect 10876 11732 10910 12108
rect 10994 11732 11028 12108
rect 11112 11732 11146 12108
rect 11230 11732 11264 12108
rect 11348 11732 11382 12108
rect 11466 11732 11500 12108
rect 11584 11732 11618 12108
rect 11697 11732 11731 12108
rect 11815 11732 11849 12108
rect 11933 11732 11967 12108
rect 12051 11732 12085 12108
rect 12138 11732 12172 11908
rect 12256 11732 12290 11908
rect 12374 11732 12408 11908
rect 12492 11732 12526 11908
rect 13132 11736 13166 11912
rect 13250 11736 13284 11912
rect 13368 11736 13402 11912
rect 13486 11736 13520 11912
rect 13605 11736 13639 12112
rect 13723 11736 13757 12112
rect 13841 11736 13875 12112
rect 13959 11736 13993 12112
rect 14078 11736 14112 12112
rect 14196 11736 14230 12112
rect 14314 11736 14348 12112
rect 14432 11736 14466 12112
rect 14550 11736 14584 12112
rect 14668 11736 14702 12112
rect 14786 11736 14820 12112
rect 14899 11736 14933 12112
rect 15017 11736 15051 12112
rect 15135 11736 15169 12112
rect 15253 11736 15287 12112
rect 15340 11736 15374 11912
rect 15458 11736 15492 11912
rect 15576 11736 15610 11912
rect 15694 11736 15728 11912
rect 16276 11736 16310 11912
rect 16394 11736 16428 11912
rect 16512 11736 16546 11912
rect 16630 11736 16664 11912
rect 16749 11736 16783 12112
rect 16867 11736 16901 12112
rect 16985 11736 17019 12112
rect 17103 11736 17137 12112
rect 17222 11736 17256 12112
rect 17340 11736 17374 12112
rect 17458 11736 17492 12112
rect 17576 11736 17610 12112
rect 17694 11736 17728 12112
rect 17812 11736 17846 12112
rect 17930 11736 17964 12112
rect 18043 11736 18077 12112
rect 18161 11736 18195 12112
rect 18279 11736 18313 12112
rect 18397 11736 18431 12112
rect 18484 11736 18518 11912
rect 18602 11736 18636 11912
rect 18720 11736 18754 11912
rect 18838 11736 18872 11912
rect 19408 11732 19442 11908
rect 19526 11732 19560 11908
rect 19644 11732 19678 11908
rect 19762 11732 19796 11908
rect 19881 11732 19915 12108
rect 19999 11732 20033 12108
rect 20117 11732 20151 12108
rect 20235 11732 20269 12108
rect 20354 11732 20388 12108
rect 20472 11732 20506 12108
rect 20590 11732 20624 12108
rect 20708 11732 20742 12108
rect 20826 11732 20860 12108
rect 20944 11732 20978 12108
rect 21062 11732 21096 12108
rect 21175 11732 21209 12108
rect 21293 11732 21327 12108
rect 21411 11732 21445 12108
rect 21529 11732 21563 12108
rect 21616 11732 21650 11908
rect 21734 11732 21768 11908
rect 21852 11732 21886 11908
rect 21970 11732 22004 11908
rect 22552 11732 22586 11908
rect 22670 11732 22704 11908
rect 22788 11732 22822 11908
rect 22906 11732 22940 11908
rect 23025 11732 23059 12108
rect 23143 11732 23177 12108
rect 23261 11732 23295 12108
rect 23379 11732 23413 12108
rect 23498 11732 23532 12108
rect 23616 11732 23650 12108
rect 23734 11732 23768 12108
rect 23852 11732 23886 12108
rect 23970 11732 24004 12108
rect 24088 11732 24122 12108
rect 24206 11732 24240 12108
rect 24319 11732 24353 12108
rect 24437 11732 24471 12108
rect 24555 11732 24589 12108
rect 24673 11732 24707 12108
rect 29966 12178 30342 12212
rect 29966 12060 30342 12094
rect 30659 12235 31035 12269
rect 70721 12371 70897 12405
rect 30659 12117 31035 12151
rect 29966 11942 30342 11976
rect 24760 11732 24794 11908
rect 24878 11732 24912 11908
rect 24996 11732 25030 11908
rect 25114 11732 25148 11908
rect 30166 11813 30342 11847
rect 30659 11999 31035 12033
rect 41570 11961 41604 12137
rect 41688 11961 41722 12137
rect 41806 11961 41840 12137
rect 41924 11961 41958 12137
rect 42042 11961 42076 12137
rect 42160 11961 42194 12137
rect 42278 11961 42312 12137
rect 42396 11961 42430 12137
rect 42514 11961 42548 12137
rect 42632 11961 42666 12137
rect 48119 11960 48153 12136
rect 30166 11695 30342 11729
rect 48237 11960 48271 12136
rect 48355 11960 48389 12136
rect 48473 11960 48507 12136
rect 48591 11960 48625 12136
rect 48709 11960 48743 12136
rect 48827 11960 48861 12136
rect 48945 11960 48979 12136
rect 49063 11960 49097 12136
rect 49181 11960 49215 12136
rect 54773 11981 54807 12157
rect 54891 11981 54925 12157
rect 55009 11981 55043 12157
rect 55127 11981 55161 12157
rect 55245 11981 55279 12157
rect 55363 11981 55397 12157
rect 55481 11981 55515 12157
rect 55599 11981 55633 12157
rect 55717 11981 55751 12157
rect 55835 11981 55869 12157
rect 70721 12253 70897 12287
rect 70521 12166 70897 12200
rect 70521 12048 70897 12082
rect 30166 11577 30342 11611
rect 30166 11459 30342 11493
rect 63426 11814 63460 11990
rect 63544 11814 63578 11990
rect 63662 11814 63696 11990
rect 63780 11814 63814 11990
rect 63898 11814 63932 11990
rect 64016 11814 64050 11990
rect 64134 11814 64168 11990
rect 64252 11814 64286 11990
rect 64370 11814 64404 11990
rect 64488 11814 64522 11990
rect 70521 11930 70897 11964
rect 30164 11066 30340 11100
rect 65234 11409 65268 11585
rect 65352 11409 65386 11585
rect 65470 11409 65504 11585
rect 65588 11409 65622 11585
rect 65718 11409 65752 11785
rect 65836 11409 65870 11785
rect 65954 11409 65988 11785
rect 66072 11409 66106 11785
rect 66190 11409 66224 11785
rect 66308 11409 66342 11785
rect 66426 11409 66460 11785
rect 70521 11812 70897 11846
rect 70521 11699 70897 11733
rect 66555 11409 66589 11585
rect 66673 11409 66707 11585
rect 66791 11409 66825 11585
rect 66909 11409 66943 11585
rect 67027 11406 67061 11582
rect 67145 11406 67179 11582
rect 67263 11406 67297 11582
rect 67381 11406 67415 11582
rect 67499 11406 67533 11582
rect 67617 11406 67651 11582
rect 67735 11406 67769 11582
rect 67853 11406 67887 11582
rect 67971 11406 68005 11582
rect 68089 11406 68123 11582
rect 70521 11581 70897 11615
rect 30164 10948 30340 10982
rect 30164 10830 30340 10864
rect 30164 10712 30340 10746
rect 29964 10582 30340 10616
rect 30657 10639 31033 10673
rect 29964 10464 30340 10498
rect 30657 10521 31033 10555
rect 29964 10346 30340 10380
rect 30657 10403 31033 10437
rect 30657 10285 31033 10319
rect 29964 10228 30340 10262
rect 29964 10110 30340 10144
rect 29964 9992 30340 10026
rect 30657 10167 31033 10201
rect 30657 10049 31033 10083
rect 34906 10061 34940 10237
rect 35024 10061 35058 10237
rect 35142 10061 35176 10237
rect 35260 10061 35294 10237
rect 35378 10061 35412 10237
rect 35496 10061 35530 10237
rect 35614 10061 35648 10237
rect 35732 10061 35766 10237
rect 35850 10061 35884 10237
rect 35968 10061 36002 10237
rect 65661 10716 65695 11092
rect 65779 10716 65813 11092
rect 65897 10716 65931 11092
rect 66015 10716 66049 11092
rect 66133 10716 66167 11092
rect 66251 10716 66285 11092
rect 66369 10716 66403 11092
rect 70521 11463 70897 11497
rect 70521 11345 70897 11379
rect 70521 11227 70897 11261
rect 70521 11109 70897 11143
rect 70521 10991 70897 11025
rect 70521 10872 70897 10906
rect 70521 10754 70897 10788
rect 70521 10636 70897 10670
rect 70521 10518 70897 10552
rect 70721 10399 70897 10433
rect 29964 9874 30340 9908
rect 30164 9745 30340 9779
rect 30657 9931 31033 9965
rect 30164 9627 30340 9661
rect 30164 9509 30340 9543
rect 520 9004 554 9180
rect 638 9004 672 9180
rect 756 9004 790 9180
rect 874 9004 908 9180
rect 993 9004 1027 9380
rect 1111 9004 1145 9380
rect 1229 9004 1263 9380
rect 1347 9004 1381 9380
rect 1466 9004 1500 9380
rect 1584 9004 1618 9380
rect 1702 9004 1736 9380
rect 1820 9004 1854 9380
rect 1938 9004 1972 9380
rect 2056 9004 2090 9380
rect 2174 9004 2208 9380
rect 2287 9004 2321 9380
rect 2405 9004 2439 9380
rect 2523 9004 2557 9380
rect 2641 9004 2675 9380
rect 2728 9004 2762 9180
rect 2846 9004 2880 9180
rect 2964 9004 2998 9180
rect 3082 9004 3116 9180
rect 3664 9004 3698 9180
rect 3782 9004 3816 9180
rect 3900 9004 3934 9180
rect 4018 9004 4052 9180
rect 4137 9004 4171 9380
rect 4255 9004 4289 9380
rect 4373 9004 4407 9380
rect 4491 9004 4525 9380
rect 4610 9004 4644 9380
rect 4728 9004 4762 9380
rect 4846 9004 4880 9380
rect 4964 9004 4998 9380
rect 5082 9004 5116 9380
rect 5200 9004 5234 9380
rect 5318 9004 5352 9380
rect 5431 9004 5465 9380
rect 5549 9004 5583 9380
rect 5667 9004 5701 9380
rect 5785 9004 5819 9380
rect 5872 9004 5906 9180
rect 5990 9004 6024 9180
rect 6108 9004 6142 9180
rect 6226 9004 6260 9180
rect 6796 9000 6830 9176
rect 6914 9000 6948 9176
rect 7032 9000 7066 9176
rect 7150 9000 7184 9176
rect 7269 9000 7303 9376
rect 7387 9000 7421 9376
rect 7505 9000 7539 9376
rect 7623 9000 7657 9376
rect 7742 9000 7776 9376
rect 7860 9000 7894 9376
rect 7978 9000 8012 9376
rect 8096 9000 8130 9376
rect 8214 9000 8248 9376
rect 8332 9000 8366 9376
rect 8450 9000 8484 9376
rect 8563 9000 8597 9376
rect 8681 9000 8715 9376
rect 8799 9000 8833 9376
rect 8917 9000 8951 9376
rect 9004 9000 9038 9176
rect 9122 9000 9156 9176
rect 9240 9000 9274 9176
rect 9358 9000 9392 9176
rect 9940 9000 9974 9176
rect 10058 9000 10092 9176
rect 10176 9000 10210 9176
rect 10294 9000 10328 9176
rect 10413 9000 10447 9376
rect 10531 9000 10565 9376
rect 10649 9000 10683 9376
rect 10767 9000 10801 9376
rect 10886 9000 10920 9376
rect 11004 9000 11038 9376
rect 11122 9000 11156 9376
rect 11240 9000 11274 9376
rect 11358 9000 11392 9376
rect 11476 9000 11510 9376
rect 11594 9000 11628 9376
rect 11707 9000 11741 9376
rect 11825 9000 11859 9376
rect 11943 9000 11977 9376
rect 12061 9000 12095 9376
rect 12148 9000 12182 9176
rect 12266 9000 12300 9176
rect 12384 9000 12418 9176
rect 12502 9000 12536 9176
rect 13142 9004 13176 9180
rect 13260 9004 13294 9180
rect 13378 9004 13412 9180
rect 13496 9004 13530 9180
rect 13615 9004 13649 9380
rect 13733 9004 13767 9380
rect 13851 9004 13885 9380
rect 13969 9004 14003 9380
rect 14088 9004 14122 9380
rect 14206 9004 14240 9380
rect 14324 9004 14358 9380
rect 14442 9004 14476 9380
rect 14560 9004 14594 9380
rect 14678 9004 14712 9380
rect 14796 9004 14830 9380
rect 14909 9004 14943 9380
rect 15027 9004 15061 9380
rect 15145 9004 15179 9380
rect 15263 9004 15297 9380
rect 15350 9004 15384 9180
rect 15468 9004 15502 9180
rect 15586 9004 15620 9180
rect 15704 9004 15738 9180
rect 16286 9004 16320 9180
rect 16404 9004 16438 9180
rect 16522 9004 16556 9180
rect 16640 9004 16674 9180
rect 16759 9004 16793 9380
rect 16877 9004 16911 9380
rect 16995 9004 17029 9380
rect 17113 9004 17147 9380
rect 17232 9004 17266 9380
rect 17350 9004 17384 9380
rect 17468 9004 17502 9380
rect 17586 9004 17620 9380
rect 17704 9004 17738 9380
rect 17822 9004 17856 9380
rect 17940 9004 17974 9380
rect 18053 9004 18087 9380
rect 18171 9004 18205 9380
rect 18289 9004 18323 9380
rect 30164 9391 30340 9425
rect 37796 9794 37830 9970
rect 37914 9794 37948 9970
rect 38032 9794 38066 9970
rect 38150 9794 38184 9970
rect 38268 9794 38302 9970
rect 38386 9794 38420 9970
rect 38504 9794 38538 9970
rect 38622 9794 38656 9970
rect 38740 9794 38774 9970
rect 38858 9794 38892 9970
rect 40121 9666 40155 10042
rect 40239 9666 40273 10042
rect 40357 9666 40391 10042
rect 40475 9666 40509 10042
rect 40593 9666 40627 10042
rect 40711 9666 40745 10042
rect 40829 9666 40863 10042
rect 41263 9670 41297 10046
rect 41381 9670 41415 10046
rect 41499 9670 41533 10046
rect 41617 9670 41651 10046
rect 41735 9670 41769 10046
rect 41853 9670 41887 10046
rect 41971 9670 42005 10046
rect 44345 9882 44379 10058
rect 44463 9882 44497 10058
rect 44581 9882 44615 10058
rect 44699 9882 44733 10058
rect 44817 9882 44851 10058
rect 44935 9882 44969 10058
rect 45053 9882 45087 10058
rect 45171 9882 45205 10058
rect 45289 9882 45323 10058
rect 45407 9882 45441 10058
rect 18407 9004 18441 9380
rect 18494 9004 18528 9180
rect 18612 9004 18646 9180
rect 18730 9004 18764 9180
rect 18848 9004 18882 9180
rect 19418 9000 19452 9176
rect 19536 9000 19570 9176
rect 19654 9000 19688 9176
rect 19772 9000 19806 9176
rect 19891 9000 19925 9376
rect 20009 9000 20043 9376
rect 20127 9000 20161 9376
rect 20245 9000 20279 9376
rect 20364 9000 20398 9376
rect 20482 9000 20516 9376
rect 20600 9000 20634 9376
rect 20718 9000 20752 9376
rect 20836 9000 20870 9376
rect 20954 9000 20988 9376
rect 21072 9000 21106 9376
rect 21185 9000 21219 9376
rect 21303 9000 21337 9376
rect 21421 9000 21455 9376
rect 21539 9000 21573 9376
rect 21626 9000 21660 9176
rect 21744 9000 21778 9176
rect 21862 9000 21896 9176
rect 21980 9000 22014 9176
rect 22562 9000 22596 9176
rect 22680 9000 22714 9176
rect 22798 9000 22832 9176
rect 22916 9000 22950 9176
rect 23035 9000 23069 9376
rect 23153 9000 23187 9376
rect 23271 9000 23305 9376
rect 23389 9000 23423 9376
rect 23508 9000 23542 9376
rect 23626 9000 23660 9376
rect 23744 9000 23778 9376
rect 23862 9000 23896 9376
rect 23980 9000 24014 9376
rect 24098 9000 24132 9376
rect 24216 9000 24250 9376
rect 24329 9000 24363 9376
rect 24447 9000 24481 9376
rect 24565 9000 24599 9376
rect 24683 9000 24717 9376
rect 24770 9000 24804 9176
rect 24888 9000 24922 9176
rect 25006 9000 25040 9176
rect 25124 9000 25158 9176
rect 46670 9754 46704 10130
rect 46788 9754 46822 10130
rect 46906 9754 46940 10130
rect 47024 9754 47058 10130
rect 47142 9754 47176 10130
rect 47260 9754 47294 10130
rect 47378 9754 47412 10130
rect 47812 9758 47846 10134
rect 47930 9758 47964 10134
rect 48048 9758 48082 10134
rect 48166 9758 48200 10134
rect 48284 9758 48318 10134
rect 48402 9758 48436 10134
rect 48520 9758 48554 10134
rect 50999 9814 51033 9990
rect 51117 9814 51151 9990
rect 51235 9814 51269 9990
rect 51353 9814 51387 9990
rect 51471 9814 51505 9990
rect 51589 9814 51623 9990
rect 51707 9814 51741 9990
rect 51825 9814 51859 9990
rect 51943 9814 51977 9990
rect 52061 9814 52095 9990
rect 40550 9083 40584 9259
rect 40668 9083 40702 9259
rect 40786 9083 40820 9259
rect 40904 9083 40938 9259
rect 41692 9087 41726 9263
rect 41810 9087 41844 9263
rect 41928 9087 41962 9263
rect 42046 9087 42080 9263
rect 53324 9686 53358 10062
rect 53442 9686 53476 10062
rect 53560 9686 53594 10062
rect 53678 9686 53712 10062
rect 53796 9686 53830 10062
rect 53914 9686 53948 10062
rect 54032 9686 54066 10062
rect 54466 9690 54500 10066
rect 54584 9690 54618 10066
rect 54702 9690 54736 10066
rect 54820 9690 54854 10066
rect 54938 9690 54972 10066
rect 55056 9690 55090 10066
rect 55174 9690 55208 10066
rect 57624 9882 57658 10058
rect 57742 9882 57776 10058
rect 57860 9882 57894 10058
rect 57978 9882 58012 10058
rect 58096 9882 58130 10058
rect 58214 9882 58248 10058
rect 58332 9882 58366 10058
rect 58450 9882 58484 10058
rect 58568 9882 58602 10058
rect 58686 9882 58720 10058
rect 47099 9171 47133 9347
rect 47217 9171 47251 9347
rect 47335 9171 47369 9347
rect 47453 9171 47487 9347
rect 48241 9175 48275 9351
rect 48359 9175 48393 9351
rect 48477 9175 48511 9351
rect 48595 9175 48629 9351
rect 59949 9754 59983 10130
rect 60067 9754 60101 10130
rect 60185 9754 60219 10130
rect 60303 9754 60337 10130
rect 60421 9754 60455 10130
rect 60539 9754 60573 10130
rect 60657 9754 60691 10130
rect 61091 9758 61125 10134
rect 61209 9758 61243 10134
rect 61327 9758 61361 10134
rect 61445 9758 61479 10134
rect 61563 9758 61597 10134
rect 61681 9758 61715 10134
rect 61799 9758 61833 10134
rect 70721 10281 70897 10315
rect 70721 10163 70897 10197
rect 70721 10045 70897 10079
rect 53753 9103 53787 9279
rect 53871 9103 53905 9279
rect 53989 9103 54023 9279
rect 54107 9103 54141 9279
rect 54895 9107 54929 9283
rect 55013 9107 55047 9283
rect 55131 9107 55165 9283
rect 55249 9107 55283 9283
rect 60378 9171 60412 9347
rect 60496 9171 60530 9347
rect 60614 9171 60648 9347
rect 60732 9171 60766 9347
rect 61520 9175 61554 9351
rect 61638 9175 61672 9351
rect 61756 9175 61790 9351
rect 61874 9175 61908 9351
rect 63421 9243 63455 9419
rect 63539 9243 63573 9419
rect 63657 9243 63691 9419
rect 63775 9243 63809 9419
rect 63893 9243 63927 9419
rect 64011 9243 64045 9419
rect 64129 9243 64163 9419
rect 64247 9243 64281 9419
rect 64365 9243 64399 9419
rect 64483 9243 64517 9419
rect 70725 9405 70901 9439
rect 70725 9287 70901 9321
rect 30166 8997 30342 9031
rect 30166 8879 30342 8913
rect 70725 9169 70901 9203
rect 70725 9051 70901 9085
rect 30166 8761 30342 8795
rect 30166 8643 30342 8677
rect 29966 8513 30342 8547
rect 30659 8570 31035 8604
rect 29966 8395 30342 8429
rect 30659 8452 31035 8486
rect 70525 8964 70901 8998
rect 70525 8846 70901 8880
rect 70525 8728 70901 8762
rect 70525 8610 70901 8644
rect 29966 8277 30342 8311
rect 30659 8334 31035 8368
rect 30659 8216 31035 8250
rect 29966 8159 30342 8193
rect 29966 8041 30342 8075
rect 29966 7923 30342 7957
rect 30659 8098 31035 8132
rect 37810 8144 37844 8320
rect 37928 8144 37962 8320
rect 38046 8144 38080 8320
rect 38164 8144 38198 8320
rect 38282 8144 38316 8320
rect 38400 8144 38434 8320
rect 38518 8144 38552 8320
rect 38636 8144 38670 8320
rect 38754 8144 38788 8320
rect 38872 8144 38906 8320
rect 44359 8232 44393 8408
rect 44477 8232 44511 8408
rect 44595 8232 44629 8408
rect 44713 8232 44747 8408
rect 44831 8232 44865 8408
rect 44949 8232 44983 8408
rect 45067 8232 45101 8408
rect 45185 8232 45219 8408
rect 45303 8232 45337 8408
rect 45421 8232 45455 8408
rect 70525 8497 70901 8531
rect 30659 7980 31035 8014
rect 29966 7805 30342 7839
rect 30166 7676 30342 7710
rect 30659 7862 31035 7896
rect 51013 8164 51047 8340
rect 51131 8164 51165 8340
rect 51249 8164 51283 8340
rect 51367 8164 51401 8340
rect 51485 8164 51519 8340
rect 51603 8164 51637 8340
rect 51721 8164 51755 8340
rect 51839 8164 51873 8340
rect 51957 8164 51991 8340
rect 52075 8164 52109 8340
rect 57638 8232 57672 8408
rect 57756 8232 57790 8408
rect 57874 8232 57908 8408
rect 57992 8232 58026 8408
rect 58110 8232 58144 8408
rect 58228 8232 58262 8408
rect 58346 8232 58380 8408
rect 58464 8232 58498 8408
rect 58582 8232 58616 8408
rect 58700 8232 58734 8408
rect 70525 8379 70901 8413
rect 30166 7558 30342 7592
rect 30166 7440 30342 7474
rect 34898 7476 34932 7652
rect 35016 7476 35050 7652
rect 35134 7476 35168 7652
rect 35252 7476 35286 7652
rect 35370 7476 35404 7652
rect 35488 7476 35522 7652
rect 35606 7476 35640 7652
rect 35724 7476 35758 7652
rect 35842 7476 35876 7652
rect 35960 7476 35994 7652
rect 30166 7322 30342 7356
rect 39274 7527 39308 7703
rect 39392 7527 39426 7703
rect 39510 7527 39544 7703
rect 39628 7527 39662 7703
rect 39758 7527 39792 7903
rect 39876 7527 39910 7903
rect 39994 7527 40028 7903
rect 40112 7527 40146 7903
rect 40230 7527 40264 7903
rect 40348 7527 40382 7903
rect 40466 7527 40500 7903
rect 40595 7527 40629 7703
rect 40713 7527 40747 7703
rect 40831 7527 40865 7703
rect 40949 7527 40983 7703
rect 41172 7527 41206 7703
rect 41290 7527 41324 7703
rect 41408 7527 41442 7703
rect 41526 7527 41560 7703
rect 41656 7527 41690 7903
rect 41774 7527 41808 7903
rect 41892 7527 41926 7903
rect 42010 7527 42044 7903
rect 42128 7527 42162 7903
rect 42246 7527 42280 7903
rect 42364 7527 42398 7903
rect 42493 7527 42527 7703
rect 42611 7527 42645 7703
rect 42729 7527 42763 7703
rect 42847 7527 42881 7703
rect 30164 6929 30340 6963
rect 30164 6811 30340 6845
rect 30164 6693 30340 6727
rect 3129 6369 3163 6545
rect 3247 6369 3281 6545
rect 3365 6369 3399 6545
rect 3483 6369 3517 6545
rect 3867 6369 3901 6545
rect 3985 6369 4019 6545
rect 4103 6369 4137 6545
rect 4221 6369 4255 6545
rect 4605 6369 4639 6545
rect 4723 6369 4757 6545
rect 4841 6369 4875 6545
rect 4959 6369 4993 6545
rect 5343 6369 5377 6545
rect 5461 6369 5495 6545
rect 5579 6369 5613 6545
rect 5697 6369 5731 6545
rect 6083 6369 6117 6545
rect 6201 6369 6235 6545
rect 6319 6369 6353 6545
rect 6437 6369 6471 6545
rect 6825 6371 6859 6547
rect 6943 6371 6977 6547
rect 7061 6371 7095 6547
rect 7179 6371 7213 6547
rect 7563 6375 7597 6551
rect 7681 6375 7715 6551
rect 7799 6375 7833 6551
rect 30164 6575 30340 6609
rect 7917 6375 7951 6551
rect 8301 6371 8335 6547
rect 8419 6371 8453 6547
rect 8537 6371 8571 6547
rect 8655 6371 8689 6547
rect 9233 6059 9267 6235
rect 9351 6059 9385 6235
rect 9469 6059 9503 6235
rect 9587 6059 9621 6235
rect 9716 6059 9750 6435
rect 9834 6059 9868 6435
rect 9952 6059 9986 6435
rect 10070 6059 10104 6435
rect 10188 6059 10222 6435
rect 10306 6059 10340 6435
rect 10424 6059 10458 6435
rect 10554 6059 10588 6235
rect 10672 6059 10706 6235
rect 10790 6059 10824 6235
rect 10908 6059 10942 6235
rect 11301 6057 11335 6233
rect 11419 6057 11453 6233
rect 11537 6057 11571 6233
rect 11655 6057 11689 6233
rect 11784 6057 11818 6433
rect 11902 6057 11936 6433
rect 12020 6057 12054 6433
rect 12138 6057 12172 6433
rect 12256 6057 12290 6433
rect 12374 6057 12408 6433
rect 12492 6057 12526 6433
rect 12622 6057 12656 6233
rect 12740 6057 12774 6233
rect 12858 6057 12892 6233
rect 12976 6057 13010 6233
rect 13370 6059 13404 6235
rect 13488 6059 13522 6235
rect 13606 6059 13640 6235
rect 13724 6059 13758 6235
rect 13853 6059 13887 6435
rect 13971 6059 14005 6435
rect 14089 6059 14123 6435
rect 14207 6059 14241 6435
rect 14325 6059 14359 6435
rect 14443 6059 14477 6435
rect 14561 6059 14595 6435
rect 14691 6059 14725 6235
rect 14809 6059 14843 6235
rect 14927 6059 14961 6235
rect 15045 6059 15079 6235
rect 15438 6057 15472 6233
rect 9773 5366 9807 5742
rect 9891 5366 9925 5742
rect 10009 5366 10043 5742
rect 10127 5366 10161 5742
rect 10245 5366 10279 5742
rect 10363 5366 10397 5742
rect 10481 5366 10515 5742
rect 15556 6057 15590 6233
rect 15674 6057 15708 6233
rect 15792 6057 15826 6233
rect 15921 6057 15955 6433
rect 16039 6057 16073 6433
rect 16157 6057 16191 6433
rect 16275 6057 16309 6433
rect 16393 6057 16427 6433
rect 16511 6057 16545 6433
rect 16629 6057 16663 6433
rect 16759 6057 16793 6233
rect 16877 6057 16911 6233
rect 16995 6057 17029 6233
rect 17113 6057 17147 6233
rect 17507 6057 17541 6233
rect 17625 6057 17659 6233
rect 17743 6057 17777 6233
rect 17861 6057 17895 6233
rect 17990 6057 18024 6433
rect 18108 6057 18142 6433
rect 18226 6057 18260 6433
rect 18344 6057 18378 6433
rect 18462 6057 18496 6433
rect 18580 6057 18614 6433
rect 18698 6057 18732 6433
rect 18828 6057 18862 6233
rect 18946 6057 18980 6233
rect 19064 6057 19098 6233
rect 19182 6057 19216 6233
rect 19575 6055 19609 6231
rect 11841 5364 11875 5740
rect 11959 5364 11993 5740
rect 12077 5364 12111 5740
rect 12195 5364 12229 5740
rect 12313 5364 12347 5740
rect 12431 5364 12465 5740
rect 12549 5364 12583 5740
rect 13910 5366 13944 5742
rect 14028 5366 14062 5742
rect 14146 5366 14180 5742
rect 14264 5366 14298 5742
rect 14382 5366 14416 5742
rect 14500 5366 14534 5742
rect 14618 5366 14652 5742
rect 15978 5364 16012 5740
rect 16096 5364 16130 5740
rect 16214 5364 16248 5740
rect 16332 5364 16366 5740
rect 16450 5364 16484 5740
rect 16568 5364 16602 5740
rect 16686 5364 16720 5740
rect 19693 6055 19727 6231
rect 19811 6055 19845 6231
rect 19929 6055 19963 6231
rect 20058 6055 20092 6431
rect 20176 6055 20210 6431
rect 20294 6055 20328 6431
rect 20412 6055 20446 6431
rect 20530 6055 20564 6431
rect 20648 6055 20682 6431
rect 20766 6055 20800 6431
rect 20896 6055 20930 6231
rect 21014 6055 21048 6231
rect 21132 6055 21166 6231
rect 21250 6055 21284 6231
rect 21644 6057 21678 6233
rect 21762 6057 21796 6233
rect 21880 6057 21914 6233
rect 21998 6057 22032 6233
rect 22127 6057 22161 6433
rect 22245 6057 22279 6433
rect 22363 6057 22397 6433
rect 22481 6057 22515 6433
rect 22599 6057 22633 6433
rect 22717 6057 22751 6433
rect 29964 6445 30340 6479
rect 22835 6057 22869 6433
rect 22965 6057 22999 6233
rect 23083 6057 23117 6233
rect 23201 6057 23235 6233
rect 23319 6057 23353 6233
rect 23712 6055 23746 6231
rect 18047 5364 18081 5740
rect 18165 5364 18199 5740
rect 18283 5364 18317 5740
rect 18401 5364 18435 5740
rect 18519 5364 18553 5740
rect 18637 5364 18671 5740
rect 18755 5364 18789 5740
rect 23830 6055 23864 6231
rect 23948 6055 23982 6231
rect 24066 6055 24100 6231
rect 24195 6055 24229 6431
rect 24313 6055 24347 6431
rect 24431 6055 24465 6431
rect 24549 6055 24583 6431
rect 24667 6055 24701 6431
rect 24785 6055 24819 6431
rect 30657 6502 31033 6536
rect 37805 6540 37839 6716
rect 37923 6540 37957 6716
rect 38041 6540 38075 6716
rect 38159 6540 38193 6716
rect 38277 6540 38311 6716
rect 38395 6540 38429 6716
rect 38513 6540 38547 6716
rect 38631 6540 38665 6716
rect 38749 6540 38783 6716
rect 38867 6540 38901 6716
rect 39701 6834 39735 7210
rect 39819 6834 39853 7210
rect 39937 6834 39971 7210
rect 40055 6834 40089 7210
rect 40173 6834 40207 7210
rect 40291 6834 40325 7210
rect 40409 6834 40443 7210
rect 24903 6055 24937 6431
rect 29964 6327 30340 6361
rect 30657 6384 31033 6418
rect 25033 6055 25067 6231
rect 25151 6055 25185 6231
rect 25269 6055 25303 6231
rect 25387 6055 25421 6231
rect 29964 6209 30340 6243
rect 30657 6266 31033 6300
rect 45823 7615 45857 7791
rect 45941 7615 45975 7791
rect 46059 7615 46093 7791
rect 46177 7615 46211 7791
rect 46307 7615 46341 7991
rect 46425 7615 46459 7991
rect 46543 7615 46577 7991
rect 46661 7615 46695 7991
rect 46779 7615 46813 7991
rect 46897 7615 46931 7991
rect 47015 7615 47049 7991
rect 47144 7615 47178 7791
rect 47262 7615 47296 7791
rect 47380 7615 47414 7791
rect 47498 7615 47532 7791
rect 47721 7615 47755 7791
rect 47839 7615 47873 7791
rect 47957 7615 47991 7791
rect 48075 7615 48109 7791
rect 48205 7615 48239 7991
rect 48323 7615 48357 7991
rect 48441 7615 48475 7991
rect 48559 7615 48593 7991
rect 48677 7615 48711 7991
rect 48795 7615 48829 7991
rect 48913 7615 48947 7991
rect 70525 8261 70901 8295
rect 70525 8143 70901 8177
rect 70525 8025 70901 8059
rect 49042 7615 49076 7791
rect 49160 7615 49194 7791
rect 49278 7615 49312 7791
rect 49396 7615 49430 7791
rect 41599 6834 41633 7210
rect 41717 6834 41751 7210
rect 41835 6834 41869 7210
rect 41953 6834 41987 7210
rect 42071 6834 42105 7210
rect 42189 6834 42223 7210
rect 42307 6834 42341 7210
rect 44354 6628 44388 6804
rect 44472 6628 44506 6804
rect 44590 6628 44624 6804
rect 44708 6628 44742 6804
rect 44826 6628 44860 6804
rect 44944 6628 44978 6804
rect 45062 6628 45096 6804
rect 45180 6628 45214 6804
rect 45298 6628 45332 6804
rect 45416 6628 45450 6804
rect 46250 6922 46284 7298
rect 46368 6922 46402 7298
rect 46486 6922 46520 7298
rect 46604 6922 46638 7298
rect 46722 6922 46756 7298
rect 46840 6922 46874 7298
rect 46958 6922 46992 7298
rect 30657 6148 31033 6182
rect 29964 6091 30340 6125
rect 20115 5362 20149 5738
rect 20233 5362 20267 5738
rect 20351 5362 20385 5738
rect 20469 5362 20503 5738
rect 20587 5362 20621 5738
rect 20705 5362 20739 5738
rect 20823 5362 20857 5738
rect 22184 5364 22218 5740
rect 22302 5364 22336 5740
rect 22420 5364 22454 5740
rect 22538 5364 22572 5740
rect 22656 5364 22690 5740
rect 22774 5364 22808 5740
rect 22892 5364 22926 5740
rect 24252 5362 24286 5738
rect 24370 5362 24404 5738
rect 24488 5362 24522 5738
rect 24606 5362 24640 5738
rect 24724 5362 24758 5738
rect 24842 5362 24876 5738
rect 24960 5362 24994 5738
rect 29964 5973 30340 6007
rect 29964 5855 30340 5889
rect 30657 6030 31033 6064
rect 30657 5912 31033 5946
rect 52477 7547 52511 7723
rect 52595 7547 52629 7723
rect 52713 7547 52747 7723
rect 52831 7547 52865 7723
rect 52961 7547 52995 7923
rect 53079 7547 53113 7923
rect 53197 7547 53231 7923
rect 53315 7547 53349 7923
rect 53433 7547 53467 7923
rect 53551 7547 53585 7923
rect 53669 7547 53703 7923
rect 53798 7547 53832 7723
rect 53916 7547 53950 7723
rect 54034 7547 54068 7723
rect 54152 7547 54186 7723
rect 54375 7547 54409 7723
rect 54493 7547 54527 7723
rect 54611 7547 54645 7723
rect 54729 7547 54763 7723
rect 54859 7547 54893 7923
rect 54977 7547 55011 7923
rect 55095 7547 55129 7923
rect 55213 7547 55247 7923
rect 55331 7547 55365 7923
rect 55449 7547 55483 7923
rect 55567 7547 55601 7923
rect 55696 7547 55730 7723
rect 55814 7547 55848 7723
rect 55932 7547 55966 7723
rect 56050 7547 56084 7723
rect 48148 6922 48182 7298
rect 48266 6922 48300 7298
rect 48384 6922 48418 7298
rect 48502 6922 48536 7298
rect 48620 6922 48654 7298
rect 48738 6922 48772 7298
rect 48856 6922 48890 7298
rect 51008 6560 51042 6736
rect 51126 6560 51160 6736
rect 51244 6560 51278 6736
rect 51362 6560 51396 6736
rect 51480 6560 51514 6736
rect 51598 6560 51632 6736
rect 51716 6560 51750 6736
rect 51834 6560 51868 6736
rect 51952 6560 51986 6736
rect 52070 6560 52104 6736
rect 52904 6854 52938 7230
rect 53022 6854 53056 7230
rect 53140 6854 53174 7230
rect 53258 6854 53292 7230
rect 53376 6854 53410 7230
rect 53494 6854 53528 7230
rect 53612 6854 53646 7230
rect 59102 7615 59136 7791
rect 59220 7615 59254 7791
rect 59338 7615 59372 7791
rect 59456 7615 59490 7791
rect 59586 7615 59620 7991
rect 59704 7615 59738 7991
rect 59822 7615 59856 7991
rect 59940 7615 59974 7991
rect 60058 7615 60092 7991
rect 60176 7615 60210 7991
rect 60294 7615 60328 7991
rect 60423 7615 60457 7791
rect 60541 7615 60575 7791
rect 60659 7615 60693 7791
rect 60777 7615 60811 7791
rect 61000 7615 61034 7791
rect 61118 7615 61152 7791
rect 61236 7615 61270 7791
rect 61354 7615 61388 7791
rect 61484 7615 61518 7991
rect 61602 7615 61636 7991
rect 61720 7615 61754 7991
rect 61838 7615 61872 7991
rect 61956 7615 61990 7991
rect 62074 7615 62108 7991
rect 62192 7615 62226 7991
rect 70525 7907 70901 7941
rect 62321 7615 62355 7791
rect 62439 7615 62473 7791
rect 62557 7615 62591 7791
rect 62675 7615 62709 7791
rect 70525 7789 70901 7823
rect 54802 6854 54836 7230
rect 54920 6854 54954 7230
rect 55038 6854 55072 7230
rect 55156 6854 55190 7230
rect 55274 6854 55308 7230
rect 55392 6854 55426 7230
rect 55510 6854 55544 7230
rect 57633 6628 57667 6804
rect 57751 6628 57785 6804
rect 57869 6628 57903 6804
rect 57987 6628 58021 6804
rect 58105 6628 58139 6804
rect 58223 6628 58257 6804
rect 58341 6628 58375 6804
rect 58459 6628 58493 6804
rect 58577 6628 58611 6804
rect 58695 6628 58729 6804
rect 59529 6922 59563 7298
rect 59647 6922 59681 7298
rect 59765 6922 59799 7298
rect 59883 6922 59917 7298
rect 60001 6922 60035 7298
rect 60119 6922 60153 7298
rect 60237 6922 60271 7298
rect 29964 5737 30340 5771
rect 30164 5608 30340 5642
rect 30657 5794 31033 5828
rect 61427 6922 61461 7298
rect 61545 6922 61579 7298
rect 61663 6922 61697 7298
rect 61781 6922 61815 7298
rect 61899 6922 61933 7298
rect 62017 6922 62051 7298
rect 62135 6922 62169 7298
rect 65236 7318 65270 7494
rect 65354 7318 65388 7494
rect 65472 7318 65506 7494
rect 65590 7318 65624 7494
rect 65720 7318 65754 7694
rect 65838 7318 65872 7694
rect 65956 7318 65990 7694
rect 66074 7318 66108 7694
rect 66192 7318 66226 7694
rect 66310 7318 66344 7694
rect 66428 7318 66462 7694
rect 70525 7670 70901 7704
rect 66557 7318 66591 7494
rect 66675 7318 66709 7494
rect 66793 7318 66827 7494
rect 70525 7552 70901 7586
rect 66911 7318 66945 7494
rect 67029 7315 67063 7491
rect 67147 7315 67181 7491
rect 67265 7315 67299 7491
rect 67383 7315 67417 7491
rect 67501 7315 67535 7491
rect 67619 7315 67653 7491
rect 67737 7315 67771 7491
rect 67855 7315 67889 7491
rect 67973 7315 68007 7491
rect 68091 7315 68125 7491
rect 70525 7434 70901 7468
rect 70525 7316 70901 7350
rect 63421 6210 63455 6386
rect 63539 6210 63573 6386
rect 63657 6210 63691 6386
rect 63775 6210 63809 6386
rect 63893 6210 63927 6386
rect 64011 6210 64045 6386
rect 64129 6210 64163 6386
rect 64247 6210 64281 6386
rect 64365 6210 64399 6386
rect 64483 6210 64517 6386
rect 65663 6625 65697 7001
rect 65781 6625 65815 7001
rect 65899 6625 65933 7001
rect 66017 6625 66051 7001
rect 66135 6625 66169 7001
rect 66253 6625 66287 7001
rect 66371 6625 66405 7001
rect 70725 7197 70901 7231
rect 70725 7079 70901 7113
rect 70725 6961 70901 6995
rect 70725 6843 70901 6877
rect 30164 5490 30340 5524
rect 70725 6261 70901 6295
rect 70725 6143 70901 6177
rect 70725 6025 70901 6059
rect 70725 5907 70901 5941
rect 70525 5820 70901 5854
rect 70525 5702 70901 5736
rect 70525 5584 70901 5618
rect 70525 5466 70901 5500
rect 30164 5372 30340 5406
rect 70525 5353 70901 5387
rect 30164 5254 30340 5288
rect 70525 5235 70901 5269
rect 70525 5117 70901 5151
rect 70525 4999 70901 5033
rect 30164 4860 30340 4894
rect 30164 4742 30340 4776
rect 70525 4881 70901 4915
rect 70525 4763 70901 4797
rect 30164 4624 30340 4658
rect 30164 4506 30340 4540
rect 29964 4376 30340 4410
rect 30657 4433 31033 4467
rect 29964 4258 30340 4292
rect 30657 4315 31033 4349
rect 29964 4140 30340 4174
rect 30657 4197 31033 4231
rect 34879 4198 34913 4374
rect 34997 4198 35031 4374
rect 35115 4198 35149 4374
rect 35233 4198 35267 4374
rect 35351 4198 35385 4374
rect 35469 4198 35503 4374
rect 35587 4198 35621 4374
rect 35705 4198 35739 4374
rect 35823 4198 35857 4374
rect 35941 4198 35975 4374
rect 30657 4079 31033 4113
rect 29964 4022 30340 4056
rect 29964 3904 30340 3938
rect 29964 3786 30340 3820
rect 30657 3961 31033 3995
rect 37788 4014 37822 4190
rect 37906 4014 37940 4190
rect 38024 4014 38058 4190
rect 38142 4014 38176 4190
rect 38260 4014 38294 4190
rect 38378 4014 38412 4190
rect 38496 4014 38530 4190
rect 38614 4014 38648 4190
rect 38732 4014 38766 4190
rect 38850 4014 38884 4190
rect 30657 3843 31033 3877
rect 29964 3668 30340 3702
rect 30164 3539 30340 3573
rect 30657 3725 31033 3759
rect 40113 3886 40147 4262
rect 40231 3886 40265 4262
rect 40349 3886 40383 4262
rect 40467 3886 40501 4262
rect 40585 3886 40619 4262
rect 40703 3886 40737 4262
rect 40821 3886 40855 4262
rect 41255 3890 41289 4266
rect 41373 3890 41407 4266
rect 41491 3890 41525 4266
rect 41609 3890 41643 4266
rect 41727 3890 41761 4266
rect 41845 3890 41879 4266
rect 70525 4645 70901 4679
rect 70525 4526 70901 4560
rect 41963 3890 41997 4266
rect 44339 4012 44373 4188
rect 44457 4012 44491 4188
rect 44575 4012 44609 4188
rect 44693 4012 44727 4188
rect 44811 4012 44845 4188
rect 44929 4012 44963 4188
rect 45047 4012 45081 4188
rect 45165 4012 45199 4188
rect 45283 4012 45317 4188
rect 45401 4012 45435 4188
rect 30164 3421 30340 3455
rect 30164 3303 30340 3337
rect 46664 3884 46698 4260
rect 46782 3884 46816 4260
rect 46900 3884 46934 4260
rect 47018 3884 47052 4260
rect 47136 3884 47170 4260
rect 47254 3884 47288 4260
rect 47372 3884 47406 4260
rect 47806 3888 47840 4264
rect 47924 3888 47958 4264
rect 48042 3888 48076 4264
rect 48160 3888 48194 4264
rect 48278 3888 48312 4264
rect 48396 3888 48430 4264
rect 48514 3888 48548 4264
rect 50994 4013 51028 4189
rect 51112 4013 51146 4189
rect 51230 4013 51264 4189
rect 51348 4013 51382 4189
rect 51466 4013 51500 4189
rect 51584 4013 51618 4189
rect 51702 4013 51736 4189
rect 51820 4013 51854 4189
rect 51938 4013 51972 4189
rect 52056 4013 52090 4189
rect 40542 3303 40576 3479
rect 40660 3303 40694 3479
rect 40778 3303 40812 3479
rect 40896 3303 40930 3479
rect 41684 3307 41718 3483
rect 41802 3307 41836 3483
rect 41920 3307 41954 3483
rect 42038 3307 42072 3483
rect 53319 3885 53353 4261
rect 53437 3885 53471 4261
rect 53555 3885 53589 4261
rect 53673 3885 53707 4261
rect 53791 3885 53825 4261
rect 53909 3885 53943 4261
rect 54027 3885 54061 4261
rect 54461 3889 54495 4265
rect 54579 3889 54613 4265
rect 54697 3889 54731 4265
rect 54815 3889 54849 4265
rect 54933 3889 54967 4265
rect 55051 3889 55085 4265
rect 63492 4290 63526 4466
rect 63610 4290 63644 4466
rect 63728 4290 63762 4466
rect 63846 4290 63880 4466
rect 63964 4290 63998 4466
rect 64082 4290 64116 4466
rect 64200 4290 64234 4466
rect 64318 4290 64352 4466
rect 64436 4290 64470 4466
rect 64554 4290 64588 4466
rect 70525 4408 70901 4442
rect 70525 4290 70901 4324
rect 55169 3889 55203 4265
rect 57616 4014 57650 4190
rect 57734 4014 57768 4190
rect 57852 4014 57886 4190
rect 57970 4014 58004 4190
rect 58088 4014 58122 4190
rect 58206 4014 58240 4190
rect 58324 4014 58358 4190
rect 58442 4014 58476 4190
rect 58560 4014 58594 4190
rect 58678 4014 58712 4190
rect 30164 3185 30340 3219
rect 47093 3301 47127 3477
rect 47211 3301 47245 3477
rect 47329 3301 47363 3477
rect 47447 3301 47481 3477
rect 48235 3305 48269 3481
rect 48353 3305 48387 3481
rect 48471 3305 48505 3481
rect 48589 3305 48623 3481
rect 59941 3886 59975 4262
rect 60059 3886 60093 4262
rect 60177 3886 60211 4262
rect 60295 3886 60329 4262
rect 60413 3886 60447 4262
rect 60531 3886 60565 4262
rect 60649 3886 60683 4262
rect 61083 3890 61117 4266
rect 61201 3890 61235 4266
rect 61319 3890 61353 4266
rect 61437 3890 61471 4266
rect 61555 3890 61589 4266
rect 61673 3890 61707 4266
rect 61791 3890 61825 4266
rect 53748 3302 53782 3478
rect 53866 3302 53900 3478
rect 53984 3302 54018 3478
rect 54102 3302 54136 3478
rect 54890 3306 54924 3482
rect 55008 3306 55042 3482
rect 55126 3306 55160 3482
rect 55244 3306 55278 3482
rect 65236 3823 65270 3999
rect 65354 3823 65388 3999
rect 65472 3823 65506 3999
rect 65590 3823 65624 3999
rect 65720 3823 65754 4199
rect 65838 3823 65872 4199
rect 65956 3823 65990 4199
rect 66074 3823 66108 4199
rect 66192 3823 66226 4199
rect 66310 3823 66344 4199
rect 66428 3823 66462 4199
rect 70525 4172 70901 4206
rect 66557 3823 66591 3999
rect 66675 3823 66709 3999
rect 66793 3823 66827 3999
rect 70725 4053 70901 4087
rect 66911 3823 66945 3999
rect 67029 3820 67063 3996
rect 67147 3820 67181 3996
rect 67265 3820 67299 3996
rect 67383 3820 67417 3996
rect 67501 3820 67535 3996
rect 67619 3820 67653 3996
rect 67737 3820 67771 3996
rect 67855 3820 67889 3996
rect 67973 3820 68007 3996
rect 68091 3820 68125 3996
rect 70725 3935 70901 3969
rect 60370 3303 60404 3479
rect 60488 3303 60522 3479
rect 60606 3303 60640 3479
rect 60724 3303 60758 3479
rect 61512 3307 61546 3483
rect 61630 3307 61664 3483
rect 61748 3307 61782 3483
rect 61866 3307 61900 3483
rect 30162 2792 30338 2826
rect 30162 2674 30338 2708
rect 65663 3130 65697 3506
rect 65781 3130 65815 3506
rect 65899 3130 65933 3506
rect 66017 3130 66051 3506
rect 66135 3130 66169 3506
rect 66253 3130 66287 3506
rect 66371 3130 66405 3506
rect 70725 3817 70901 3851
rect 70725 3699 70901 3733
rect 70721 3129 70897 3163
rect 70721 3011 70897 3045
rect 70721 2893 70897 2927
rect 30162 2556 30338 2590
rect 30162 2438 30338 2472
rect 29962 2308 30338 2342
rect 30655 2365 31031 2399
rect 37802 2364 37836 2540
rect 37920 2364 37954 2540
rect 38038 2364 38072 2540
rect 38156 2364 38190 2540
rect 38274 2364 38308 2540
rect 38392 2364 38426 2540
rect 38510 2364 38544 2540
rect 38628 2364 38662 2540
rect 38746 2364 38780 2540
rect 38864 2364 38898 2540
rect 44353 2362 44387 2538
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 29962 2190 30338 2224
rect 30655 2247 31031 2281
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 29962 2072 30338 2106
rect 30655 2129 31031 2163
rect 44471 2362 44505 2538
rect 44589 2362 44623 2538
rect 44707 2362 44741 2538
rect 44825 2362 44859 2538
rect 44943 2362 44977 2538
rect 45061 2362 45095 2538
rect 45179 2362 45213 2538
rect 45297 2362 45331 2538
rect 45415 2362 45449 2538
rect 51008 2363 51042 2539
rect 51126 2363 51160 2539
rect 51244 2363 51278 2539
rect 51362 2363 51396 2539
rect 51480 2363 51514 2539
rect 51598 2363 51632 2539
rect 51716 2363 51750 2539
rect 51834 2363 51868 2539
rect 51952 2363 51986 2539
rect 52070 2363 52104 2539
rect 57630 2364 57664 2540
rect 57748 2364 57782 2540
rect 57866 2364 57900 2540
rect 57984 2364 58018 2540
rect 58102 2364 58136 2540
rect 58220 2364 58254 2540
rect 58338 2364 58372 2540
rect 58456 2364 58490 2540
rect 58574 2364 58608 2540
rect 58692 2364 58726 2540
rect 70721 2775 70897 2809
rect 70521 2688 70897 2722
rect 70521 2570 70897 2604
rect 70521 2452 70897 2486
rect 30655 2011 31031 2045
rect 29962 1954 30338 1988
rect 29962 1836 30338 1870
rect 29962 1718 30338 1752
rect 30655 1893 31031 1927
rect 30655 1775 31031 1809
rect 29962 1600 30338 1634
rect 30162 1471 30338 1505
rect 30655 1657 31031 1691
rect 39266 1747 39300 1923
rect 39384 1747 39418 1923
rect 39502 1747 39536 1923
rect 39620 1747 39654 1923
rect 39750 1747 39784 2123
rect 39868 1747 39902 2123
rect 39986 1747 40020 2123
rect 40104 1747 40138 2123
rect 40222 1747 40256 2123
rect 40340 1747 40374 2123
rect 40458 1747 40492 2123
rect 40587 1747 40621 1923
rect 40705 1747 40739 1923
rect 40823 1747 40857 1923
rect 40941 1747 40975 1923
rect 41164 1747 41198 1923
rect 41282 1747 41316 1923
rect 41400 1747 41434 1923
rect 41518 1747 41552 1923
rect 41648 1747 41682 2123
rect 41766 1747 41800 2123
rect 41884 1747 41918 2123
rect 42002 1747 42036 2123
rect 42120 1747 42154 2123
rect 42238 1747 42272 2123
rect 42356 1747 42390 2123
rect 42485 1747 42519 1923
rect 42603 1747 42637 1923
rect 42721 1747 42755 1923
rect 42839 1747 42873 1923
rect 30162 1353 30338 1387
rect 34895 1438 34929 1614
rect 35013 1438 35047 1614
rect 35131 1438 35165 1614
rect 35249 1438 35283 1614
rect 35367 1438 35401 1614
rect 35485 1438 35519 1614
rect 35603 1438 35637 1614
rect 35721 1438 35755 1614
rect 35839 1438 35873 1614
rect 35957 1438 35991 1614
rect 30162 1235 30338 1269
rect 30162 1117 30338 1151
rect 30164 723 30340 757
rect 30164 605 30340 639
rect 37797 760 37831 936
rect 37915 760 37949 936
rect 38033 760 38067 936
rect 38151 760 38185 936
rect 38269 760 38303 936
rect 38387 760 38421 936
rect 38505 760 38539 936
rect 38623 760 38657 936
rect 38741 760 38775 936
rect 38859 760 38893 936
rect 39693 1054 39727 1430
rect 39811 1054 39845 1430
rect 39929 1054 39963 1430
rect 40047 1054 40081 1430
rect 40165 1054 40199 1430
rect 40283 1054 40317 1430
rect 40401 1054 40435 1430
rect 30164 487 30340 521
rect 45817 1745 45851 1921
rect 45935 1745 45969 1921
rect 46053 1745 46087 1921
rect 46171 1745 46205 1921
rect 46301 1745 46335 2121
rect 46419 1745 46453 2121
rect 46537 1745 46571 2121
rect 46655 1745 46689 2121
rect 46773 1745 46807 2121
rect 46891 1745 46925 2121
rect 47009 1745 47043 2121
rect 47138 1745 47172 1921
rect 47256 1745 47290 1921
rect 47374 1745 47408 1921
rect 47492 1745 47526 1921
rect 47715 1745 47749 1921
rect 47833 1745 47867 1921
rect 47951 1745 47985 1921
rect 48069 1745 48103 1921
rect 48199 1745 48233 2121
rect 48317 1745 48351 2121
rect 48435 1745 48469 2121
rect 48553 1745 48587 2121
rect 48671 1745 48705 2121
rect 48789 1745 48823 2121
rect 48907 1745 48941 2121
rect 49036 1745 49070 1921
rect 49154 1745 49188 1921
rect 49272 1745 49306 1921
rect 49390 1745 49424 1921
rect 41591 1054 41625 1430
rect 41709 1054 41743 1430
rect 41827 1054 41861 1430
rect 41945 1054 41979 1430
rect 42063 1054 42097 1430
rect 42181 1054 42215 1430
rect 42299 1054 42333 1430
rect 44348 758 44382 934
rect 44466 758 44500 934
rect 44584 758 44618 934
rect 44702 758 44736 934
rect 44820 758 44854 934
rect 44938 758 44972 934
rect 45056 758 45090 934
rect 45174 758 45208 934
rect 45292 758 45326 934
rect 45410 758 45444 934
rect 46244 1052 46278 1428
rect 46362 1052 46396 1428
rect 46480 1052 46514 1428
rect 46598 1052 46632 1428
rect 46716 1052 46750 1428
rect 46834 1052 46868 1428
rect 46952 1052 46986 1428
rect 30164 369 30340 403
rect 29964 239 30340 273
rect 30657 296 31033 330
rect 29964 121 30340 155
rect 30657 178 31033 212
rect 52472 1746 52506 1922
rect 52590 1746 52624 1922
rect 52708 1746 52742 1922
rect 52826 1746 52860 1922
rect 52956 1746 52990 2122
rect 53074 1746 53108 2122
rect 53192 1746 53226 2122
rect 53310 1746 53344 2122
rect 53428 1746 53462 2122
rect 53546 1746 53580 2122
rect 53664 1746 53698 2122
rect 53793 1746 53827 1922
rect 53911 1746 53945 1922
rect 54029 1746 54063 1922
rect 54147 1746 54181 1922
rect 54370 1746 54404 1922
rect 54488 1746 54522 1922
rect 54606 1746 54640 1922
rect 54724 1746 54758 1922
rect 54854 1746 54888 2122
rect 54972 1746 55006 2122
rect 55090 1746 55124 2122
rect 55208 1746 55242 2122
rect 55326 1746 55360 2122
rect 55444 1746 55478 2122
rect 55562 1746 55596 2122
rect 70521 2334 70897 2368
rect 55691 1746 55725 1922
rect 55809 1746 55843 1922
rect 55927 1746 55961 1922
rect 56045 1746 56079 1922
rect 48142 1052 48176 1428
rect 48260 1052 48294 1428
rect 48378 1052 48412 1428
rect 48496 1052 48530 1428
rect 48614 1052 48648 1428
rect 48732 1052 48766 1428
rect 48850 1052 48884 1428
rect 51003 759 51037 935
rect 51121 759 51155 935
rect 51239 759 51273 935
rect 51357 759 51391 935
rect 51475 759 51509 935
rect 51593 759 51627 935
rect 51711 759 51745 935
rect 51829 759 51863 935
rect 51947 759 51981 935
rect 52065 759 52099 935
rect 52899 1053 52933 1429
rect 53017 1053 53051 1429
rect 53135 1053 53169 1429
rect 53253 1053 53287 1429
rect 53371 1053 53405 1429
rect 53489 1053 53523 1429
rect 53607 1053 53641 1429
rect 29964 3 30340 37
rect 30657 60 31033 94
rect 59094 1747 59128 1923
rect 59212 1747 59246 1923
rect 59330 1747 59364 1923
rect 59448 1747 59482 1923
rect 59578 1747 59612 2123
rect 59696 1747 59730 2123
rect 59814 1747 59848 2123
rect 59932 1747 59966 2123
rect 60050 1747 60084 2123
rect 60168 1747 60202 2123
rect 60286 1747 60320 2123
rect 60415 1747 60449 1923
rect 60533 1747 60567 1923
rect 60651 1747 60685 1923
rect 60769 1747 60803 1923
rect 60992 1747 61026 1923
rect 61110 1747 61144 1923
rect 61228 1747 61262 1923
rect 61346 1747 61380 1923
rect 61476 1747 61510 2123
rect 61594 1747 61628 2123
rect 61712 1747 61746 2123
rect 61830 1747 61864 2123
rect 61948 1747 61982 2123
rect 62066 1747 62100 2123
rect 62184 1747 62218 2123
rect 70521 2221 70897 2255
rect 70521 2103 70897 2137
rect 62313 1747 62347 1923
rect 62431 1747 62465 1923
rect 62549 1747 62583 1923
rect 62667 1747 62701 1923
rect 70521 1985 70897 2019
rect 70521 1867 70897 1901
rect 54797 1053 54831 1429
rect 54915 1053 54949 1429
rect 55033 1053 55067 1429
rect 55151 1053 55185 1429
rect 55269 1053 55303 1429
rect 55387 1053 55421 1429
rect 55505 1053 55539 1429
rect 57625 760 57659 936
rect 57743 760 57777 936
rect 57861 760 57895 936
rect 57979 760 58013 936
rect 58097 760 58131 936
rect 58215 760 58249 936
rect 58333 760 58367 936
rect 58451 760 58485 936
rect 58569 760 58603 936
rect 58687 760 58721 936
rect 59521 1054 59555 1430
rect 59639 1054 59673 1430
rect 59757 1054 59791 1430
rect 59875 1054 59909 1430
rect 59993 1054 60027 1430
rect 60111 1054 60145 1430
rect 60229 1054 60263 1430
rect 30657 -58 31033 -24
rect 29964 -115 30340 -81
rect 29964 -233 30340 -199
rect 29964 -351 30340 -317
rect 30657 -176 31033 -142
rect 70521 1749 70897 1783
rect 70521 1631 70897 1665
rect 70521 1513 70897 1547
rect 61419 1054 61453 1430
rect 61537 1054 61571 1430
rect 61655 1054 61689 1430
rect 61773 1054 61807 1430
rect 61891 1054 61925 1430
rect 62009 1054 62043 1430
rect 62127 1054 62161 1430
rect 63489 1220 63523 1396
rect 63607 1220 63641 1396
rect 63725 1220 63759 1396
rect 63843 1220 63877 1396
rect 63961 1220 63995 1396
rect 64079 1220 64113 1396
rect 64197 1220 64231 1396
rect 64315 1220 64349 1396
rect 64433 1220 64467 1396
rect 64551 1220 64585 1396
rect 70521 1394 70897 1428
rect 70521 1276 70897 1310
rect 70521 1158 70897 1192
rect 70521 1040 70897 1074
rect 70721 921 70897 955
rect 70721 803 70897 837
rect 70721 685 70897 719
rect 70721 567 70897 601
rect 70721 -15 70897 19
rect 30657 -294 31033 -260
rect 29964 -469 30340 -435
rect 30164 -598 30340 -564
rect 30657 -412 31033 -378
rect 65236 -525 65270 -349
rect 65354 -525 65388 -349
rect 65472 -525 65506 -349
rect 65590 -525 65624 -349
rect 65720 -525 65754 -149
rect 65838 -525 65872 -149
rect 65956 -525 65990 -149
rect 66074 -525 66108 -149
rect 66192 -525 66226 -149
rect 66310 -525 66344 -149
rect 66428 -525 66462 -149
rect 70721 -133 70897 -99
rect 70721 -251 70897 -217
rect 66557 -525 66591 -349
rect 66675 -525 66709 -349
rect 66793 -525 66827 -349
rect 66911 -525 66945 -349
rect 67029 -528 67063 -352
rect 30164 -716 30340 -682
rect 30164 -834 30340 -800
rect 67147 -528 67181 -352
rect 67265 -528 67299 -352
rect 67383 -528 67417 -352
rect 67501 -528 67535 -352
rect 67619 -528 67653 -352
rect 67737 -528 67771 -352
rect 67855 -528 67889 -352
rect 67973 -528 68007 -352
rect 68091 -528 68125 -352
rect 70721 -369 70897 -335
rect 70521 -456 70897 -422
rect 30164 -952 30340 -918
rect 30162 -1345 30338 -1311
rect 30162 -1463 30338 -1429
rect 30162 -1581 30338 -1547
rect 292 -2140 326 -1964
rect 410 -2140 444 -1964
rect 528 -2140 562 -1964
rect 646 -2140 680 -1964
rect 733 -2140 767 -1764
rect 851 -2140 885 -1764
rect 969 -2140 1003 -1764
rect 1087 -2140 1121 -1764
rect 1200 -2140 1234 -1764
rect 1318 -2140 1352 -1764
rect 1436 -2140 1470 -1764
rect 1554 -2140 1588 -1764
rect 1672 -2140 1706 -1764
rect 1790 -2140 1824 -1764
rect 1908 -2140 1942 -1764
rect 2027 -2140 2061 -1764
rect 2145 -2140 2179 -1764
rect 2263 -2140 2297 -1764
rect 2381 -2140 2415 -1764
rect 2500 -2140 2534 -1964
rect 2618 -2140 2652 -1964
rect 2736 -2140 2770 -1964
rect 2854 -2140 2888 -1964
rect 3436 -2140 3470 -1964
rect 3554 -2140 3588 -1964
rect 3672 -2140 3706 -1964
rect 3790 -2140 3824 -1964
rect 3877 -2140 3911 -1764
rect 3995 -2140 4029 -1764
rect 4113 -2140 4147 -1764
rect 4231 -2140 4265 -1764
rect 4344 -2140 4378 -1764
rect 4462 -2140 4496 -1764
rect 4580 -2140 4614 -1764
rect 4698 -2140 4732 -1764
rect 4816 -2140 4850 -1764
rect 4934 -2140 4968 -1764
rect 5052 -2140 5086 -1764
rect 5171 -2140 5205 -1764
rect 5289 -2140 5323 -1764
rect 5407 -2140 5441 -1764
rect 5525 -2140 5559 -1764
rect 5644 -2140 5678 -1964
rect 5762 -2140 5796 -1964
rect 5880 -2140 5914 -1964
rect 5998 -2140 6032 -1964
rect 6568 -2136 6602 -1960
rect 6686 -2136 6720 -1960
rect 6804 -2136 6838 -1960
rect 6922 -2136 6956 -1960
rect 7009 -2136 7043 -1760
rect 7127 -2136 7161 -1760
rect 7245 -2136 7279 -1760
rect 7363 -2136 7397 -1760
rect 7476 -2136 7510 -1760
rect 7594 -2136 7628 -1760
rect 7712 -2136 7746 -1760
rect 7830 -2136 7864 -1760
rect 7948 -2136 7982 -1760
rect 8066 -2136 8100 -1760
rect 8184 -2136 8218 -1760
rect 8303 -2136 8337 -1760
rect 8421 -2136 8455 -1760
rect 8539 -2136 8573 -1760
rect 8657 -2136 8691 -1760
rect 8776 -2136 8810 -1960
rect 8894 -2136 8928 -1960
rect 9012 -2136 9046 -1960
rect 9130 -2136 9164 -1960
rect 9712 -2136 9746 -1960
rect 9830 -2136 9864 -1960
rect 9948 -2136 9982 -1960
rect 10066 -2136 10100 -1960
rect 10153 -2136 10187 -1760
rect 10271 -2136 10305 -1760
rect 10389 -2136 10423 -1760
rect 10507 -2136 10541 -1760
rect 10620 -2136 10654 -1760
rect 10738 -2136 10772 -1760
rect 10856 -2136 10890 -1760
rect 10974 -2136 11008 -1760
rect 11092 -2136 11126 -1760
rect 11210 -2136 11244 -1760
rect 11328 -2136 11362 -1760
rect 11447 -2136 11481 -1760
rect 11565 -2136 11599 -1760
rect 11683 -2136 11717 -1760
rect 30162 -1699 30338 -1665
rect 11801 -2136 11835 -1760
rect 11920 -2136 11954 -1960
rect 12038 -2136 12072 -1960
rect 12156 -2136 12190 -1960
rect 12274 -2136 12308 -1960
rect 12914 -2140 12948 -1964
rect 13032 -2140 13066 -1964
rect 13150 -2140 13184 -1964
rect 13268 -2140 13302 -1964
rect 13355 -2140 13389 -1764
rect 13473 -2140 13507 -1764
rect 13591 -2140 13625 -1764
rect 13709 -2140 13743 -1764
rect 13822 -2140 13856 -1764
rect 13940 -2140 13974 -1764
rect 14058 -2140 14092 -1764
rect 14176 -2140 14210 -1764
rect 14294 -2140 14328 -1764
rect 14412 -2140 14446 -1764
rect 14530 -2140 14564 -1764
rect 14649 -2140 14683 -1764
rect 14767 -2140 14801 -1764
rect 14885 -2140 14919 -1764
rect 15003 -2140 15037 -1764
rect 15122 -2140 15156 -1964
rect 15240 -2140 15274 -1964
rect 15358 -2140 15392 -1964
rect 15476 -2140 15510 -1964
rect 16058 -2140 16092 -1964
rect 16176 -2140 16210 -1964
rect 16294 -2140 16328 -1964
rect 16412 -2140 16446 -1964
rect 16499 -2140 16533 -1764
rect 16617 -2140 16651 -1764
rect 16735 -2140 16769 -1764
rect 16853 -2140 16887 -1764
rect 16966 -2140 17000 -1764
rect 17084 -2140 17118 -1764
rect 17202 -2140 17236 -1764
rect 17320 -2140 17354 -1764
rect 17438 -2140 17472 -1764
rect 17556 -2140 17590 -1764
rect 17674 -2140 17708 -1764
rect 17793 -2140 17827 -1764
rect 17911 -2140 17945 -1764
rect 18029 -2140 18063 -1764
rect 18147 -2140 18181 -1764
rect 18266 -2140 18300 -1964
rect 18384 -2140 18418 -1964
rect 18502 -2140 18536 -1964
rect 18620 -2140 18654 -1964
rect 19190 -2136 19224 -1960
rect 19308 -2136 19342 -1960
rect 19426 -2136 19460 -1960
rect 19544 -2136 19578 -1960
rect 19631 -2136 19665 -1760
rect 19749 -2136 19783 -1760
rect 19867 -2136 19901 -1760
rect 19985 -2136 20019 -1760
rect 20098 -2136 20132 -1760
rect 20216 -2136 20250 -1760
rect 20334 -2136 20368 -1760
rect 20452 -2136 20486 -1760
rect 20570 -2136 20604 -1760
rect 20688 -2136 20722 -1760
rect 20806 -2136 20840 -1760
rect 20925 -2136 20959 -1760
rect 21043 -2136 21077 -1760
rect 21161 -2136 21195 -1760
rect 21279 -2136 21313 -1760
rect 21398 -2136 21432 -1960
rect 21516 -2136 21550 -1960
rect 21634 -2136 21668 -1960
rect 21752 -2136 21786 -1960
rect 22334 -2136 22368 -1960
rect 22452 -2136 22486 -1960
rect 22570 -2136 22604 -1960
rect 22688 -2136 22722 -1960
rect 22775 -2136 22809 -1760
rect 22893 -2136 22927 -1760
rect 23011 -2136 23045 -1760
rect 23129 -2136 23163 -1760
rect 23242 -2136 23276 -1760
rect 23360 -2136 23394 -1760
rect 23478 -2136 23512 -1760
rect 23596 -2136 23630 -1760
rect 23714 -2136 23748 -1760
rect 23832 -2136 23866 -1760
rect 23950 -2136 23984 -1760
rect 24069 -2136 24103 -1760
rect 24187 -2136 24221 -1760
rect 24305 -2136 24339 -1760
rect 24423 -2136 24457 -1760
rect 29962 -1829 30338 -1795
rect 30655 -1772 31031 -1738
rect 41605 -1743 41639 -1567
rect 41723 -1743 41757 -1567
rect 41841 -1743 41875 -1567
rect 41959 -1743 41993 -1567
rect 42077 -1743 42111 -1567
rect 42195 -1743 42229 -1567
rect 42313 -1743 42347 -1567
rect 42431 -1743 42465 -1567
rect 42549 -1743 42583 -1567
rect 42667 -1743 42701 -1567
rect 48159 -1738 48193 -1562
rect 48277 -1738 48311 -1562
rect 48395 -1738 48429 -1562
rect 48513 -1738 48547 -1562
rect 48631 -1738 48665 -1562
rect 48749 -1738 48783 -1562
rect 48867 -1738 48901 -1562
rect 48985 -1738 49019 -1562
rect 49103 -1738 49137 -1562
rect 49221 -1738 49255 -1562
rect 54808 -1750 54842 -1574
rect 54926 -1750 54960 -1574
rect 55044 -1750 55078 -1574
rect 55162 -1750 55196 -1574
rect 55280 -1750 55314 -1574
rect 55398 -1750 55432 -1574
rect 55516 -1750 55550 -1574
rect 55634 -1750 55668 -1574
rect 55752 -1750 55786 -1574
rect 55870 -1750 55904 -1574
rect 63496 -1625 63530 -1449
rect 63614 -1625 63648 -1449
rect 63732 -1625 63766 -1449
rect 63850 -1625 63884 -1449
rect 63968 -1625 64002 -1449
rect 64086 -1625 64120 -1449
rect 64204 -1625 64238 -1449
rect 64322 -1625 64356 -1449
rect 64440 -1625 64474 -1449
rect 64558 -1625 64592 -1449
rect 65663 -1218 65697 -842
rect 65781 -1218 65815 -842
rect 65899 -1218 65933 -842
rect 66017 -1218 66051 -842
rect 66135 -1218 66169 -842
rect 66253 -1218 66287 -842
rect 66371 -1218 66405 -842
rect 70521 -574 70897 -540
rect 70521 -692 70897 -658
rect 70521 -810 70897 -776
rect 70521 -923 70897 -889
rect 70521 -1041 70897 -1007
rect 70521 -1159 70897 -1125
rect 70521 -1277 70897 -1243
rect 70521 -1395 70897 -1361
rect 70521 -1513 70897 -1479
rect 24542 -2136 24576 -1960
rect 24660 -2136 24694 -1960
rect 24778 -2136 24812 -1960
rect 24896 -2136 24930 -1960
rect 29962 -1947 30338 -1913
rect 30655 -1890 31031 -1856
rect 29962 -2065 30338 -2031
rect 30655 -2008 31031 -1974
rect 30655 -2126 31031 -2092
rect 29962 -2183 30338 -2149
rect 29962 -2301 30338 -2267
rect 29962 -2419 30338 -2385
rect 30655 -2244 31031 -2210
rect 70521 -1631 70897 -1597
rect 70521 -1750 70897 -1716
rect 70521 -1868 70897 -1834
rect 70521 -1986 70897 -1952
rect 70521 -2104 70897 -2070
rect 70721 -2223 70897 -2189
rect 30655 -2362 31031 -2328
rect 70721 -2341 70897 -2307
rect 29962 -2537 30338 -2503
rect 30162 -2666 30338 -2632
rect 30655 -2480 31031 -2446
rect 70721 -2459 70897 -2425
rect 70721 -2577 70897 -2543
rect 30162 -2784 30338 -2750
rect 30162 -2902 30338 -2868
rect 30162 -3020 30338 -2986
<< psubdiff >>
rect 40361 23758 40595 23792
rect 40361 23668 40407 23758
rect 40570 23668 40595 23758
rect 40361 23637 40595 23668
rect 46874 23755 47108 23789
rect 46874 23665 46920 23755
rect 47083 23665 47108 23755
rect 46874 23634 47108 23665
rect 53408 23750 53642 23784
rect 53408 23660 53454 23750
rect 53617 23660 53642 23750
rect 53408 23629 53642 23660
rect 59966 23754 60200 23788
rect 59966 23664 60012 23754
rect 60175 23664 60200 23754
rect 59966 23633 60200 23664
rect 41858 23387 42013 23433
rect 41858 23224 41889 23387
rect 41979 23224 42013 23387
rect 41858 23199 42013 23224
rect 43000 23385 43155 23431
rect 43000 23222 43031 23385
rect 43121 23222 43155 23385
rect 48371 23384 48526 23430
rect 43000 23197 43155 23222
rect 48371 23221 48402 23384
rect 48492 23221 48526 23384
rect 48371 23196 48526 23221
rect 49513 23382 49668 23428
rect 49513 23219 49544 23382
rect 49634 23219 49668 23382
rect 54905 23379 55060 23425
rect 49513 23194 49668 23219
rect 54905 23216 54936 23379
rect 55026 23216 55060 23379
rect 54905 23191 55060 23216
rect 56047 23377 56202 23423
rect 56047 23214 56078 23377
rect 56168 23214 56202 23377
rect 61463 23383 61618 23429
rect 56047 23189 56202 23214
rect 61463 23220 61494 23383
rect 61584 23220 61618 23383
rect 61463 23195 61618 23220
rect 62605 23381 62760 23427
rect 62605 23218 62636 23381
rect 62726 23218 62760 23381
rect 62605 23193 62760 23218
rect 40375 22108 40609 22142
rect 40375 22018 40421 22108
rect 40584 22018 40609 22108
rect 40375 21987 40609 22018
rect 46888 22105 47122 22139
rect 46888 22015 46934 22105
rect 47097 22015 47122 22105
rect 46888 21984 47122 22015
rect 53422 22100 53656 22134
rect 53422 22010 53468 22100
rect 53631 22010 53656 22100
rect 53422 21979 53656 22010
rect 40370 20504 40604 20538
rect 40370 20414 40416 20504
rect 40579 20414 40604 20504
rect 59980 22104 60214 22138
rect 59980 22014 60026 22104
rect 60189 22014 60214 22104
rect 59980 21983 60214 22014
rect 46883 20501 47117 20535
rect 40370 20383 40604 20414
rect 41802 20344 41957 20390
rect 46883 20411 46929 20501
rect 47092 20411 47117 20501
rect 53417 20496 53651 20530
rect 46883 20380 47117 20411
rect 41802 20181 41833 20344
rect 41923 20181 41957 20344
rect 41802 20156 41957 20181
rect 48315 20341 48470 20387
rect 53417 20406 53463 20496
rect 53626 20406 53651 20496
rect 72477 20817 72583 20859
rect 59975 20500 60209 20534
rect 53417 20375 53651 20406
rect 48315 20178 48346 20341
rect 48436 20178 48470 20341
rect 48315 20153 48470 20178
rect 54849 20336 55004 20382
rect 59975 20410 60021 20500
rect 60184 20410 60209 20500
rect 59975 20379 60209 20410
rect 54849 20173 54880 20336
rect 54970 20173 55004 20336
rect 54849 20148 55004 20173
rect 61407 20340 61562 20386
rect 61407 20177 61438 20340
rect 61528 20177 61562 20340
rect 61407 20152 61562 20177
rect 72477 20713 72501 20817
rect 72547 20713 72583 20817
rect 72477 20673 72583 20713
rect 4220 20008 4406 20032
rect 4220 19962 4260 20008
rect 4364 19962 4406 20008
rect 4220 19926 4406 19962
rect 7364 20008 7550 20032
rect 7364 19962 7404 20008
rect 7508 19962 7550 20008
rect 7364 19926 7550 19962
rect 10496 20004 10682 20028
rect 10496 19958 10536 20004
rect 10640 19958 10682 20004
rect 10496 19922 10682 19958
rect 13640 20004 13826 20028
rect 13640 19958 13680 20004
rect 13784 19958 13826 20004
rect 13640 19922 13826 19958
rect 16842 20008 17028 20032
rect 16842 19962 16882 20008
rect 16986 19962 17028 20008
rect 16842 19926 17028 19962
rect 19986 20008 20172 20032
rect 19986 19962 20026 20008
rect 20130 19962 20172 20008
rect 19986 19926 20172 19962
rect 23118 20004 23304 20028
rect 23118 19958 23158 20004
rect 23262 19958 23304 20004
rect 23118 19922 23304 19958
rect 26262 20004 26448 20028
rect 26262 19958 26302 20004
rect 26406 19958 26448 20004
rect 26262 19922 26448 19958
rect 42825 18150 43059 18184
rect 42825 18060 42850 18150
rect 43013 18060 43059 18150
rect 42825 18029 43059 18060
rect 49383 18146 49617 18180
rect 49383 18056 49408 18146
rect 49571 18056 49617 18146
rect 49383 18025 49617 18056
rect 55917 18151 56151 18185
rect 55917 18061 55942 18151
rect 56105 18061 56151 18151
rect 55917 18030 56151 18061
rect 62430 18154 62664 18188
rect 62430 18064 62455 18154
rect 62618 18064 62664 18154
rect 62430 18033 62664 18064
rect 40265 17777 40420 17823
rect 40265 17614 40299 17777
rect 40389 17614 40420 17777
rect 40265 17589 40420 17614
rect 41407 17779 41562 17825
rect 41407 17616 41441 17779
rect 41531 17616 41562 17779
rect 46823 17773 46978 17819
rect 41407 17591 41562 17616
rect 46823 17610 46857 17773
rect 46947 17610 46978 17773
rect 46823 17585 46978 17610
rect 47965 17775 48120 17821
rect 47965 17612 47999 17775
rect 48089 17612 48120 17775
rect 53357 17778 53512 17824
rect 47965 17587 48120 17612
rect 53357 17615 53391 17778
rect 53481 17615 53512 17778
rect 53357 17590 53512 17615
rect 54499 17780 54654 17826
rect 54499 17617 54533 17780
rect 54623 17617 54654 17780
rect 59870 17781 60025 17827
rect 54499 17592 54654 17617
rect 59870 17618 59904 17781
rect 59994 17618 60025 17781
rect 59870 17593 60025 17618
rect 61012 17783 61167 17829
rect 61012 17620 61046 17783
rect 61136 17620 61167 17783
rect 61012 17595 61167 17620
rect 72477 17673 72583 17715
rect 42811 16500 43045 16534
rect 5034 15704 5230 15734
rect 5034 15638 5072 15704
rect 5190 15638 5230 15704
rect 5034 15590 5230 15638
rect 6202 15704 6398 15734
rect 6202 15638 6240 15704
rect 6358 15638 6398 15704
rect 6202 15590 6398 15638
rect 7370 15704 7566 15734
rect 7370 15638 7408 15704
rect 7526 15638 7566 15704
rect 7370 15590 7566 15638
rect 8538 15704 8734 15734
rect 8538 15638 8576 15704
rect 8694 15638 8734 15704
rect 8538 15590 8734 15638
rect 9712 15702 9908 15732
rect 9712 15636 9750 15702
rect 9868 15636 9908 15702
rect 9712 15588 9908 15636
rect 10880 15702 11076 15732
rect 10880 15636 10918 15702
rect 11036 15636 11076 15702
rect 10880 15588 11076 15636
rect 12048 15702 12244 15732
rect 12048 15636 12086 15702
rect 12204 15636 12244 15702
rect 12048 15588 12244 15636
rect 13216 15702 13412 15732
rect 13216 15636 13254 15702
rect 13372 15636 13412 15702
rect 13216 15588 13412 15636
rect 14198 15633 14410 15663
rect 14198 15577 14236 15633
rect 14370 15577 14410 15633
rect 14198 15555 14410 15577
rect 15646 15633 15858 15663
rect 15646 15577 15684 15633
rect 15818 15577 15858 15633
rect 15646 15555 15858 15577
rect 17144 15631 17356 15661
rect 17144 15575 17182 15631
rect 17316 15575 17356 15631
rect 17144 15553 17356 15575
rect 18592 15631 18804 15661
rect 18592 15575 18630 15631
rect 18764 15575 18804 15631
rect 18592 15553 18804 15575
rect 20112 15633 20324 15663
rect 20112 15577 20150 15633
rect 20284 15577 20324 15633
rect 20112 15555 20324 15577
rect 21560 15633 21772 15663
rect 21560 15577 21598 15633
rect 21732 15577 21772 15633
rect 21560 15555 21772 15577
rect 23058 15631 23270 15661
rect 23058 15575 23096 15631
rect 23230 15575 23270 15631
rect 23058 15553 23270 15575
rect 24506 15631 24718 15661
rect 24506 15575 24544 15631
rect 24678 15575 24718 15631
rect 24506 15553 24718 15575
rect 42811 16410 42836 16500
rect 42999 16410 43045 16500
rect 49369 16496 49603 16530
rect 42811 16379 43045 16410
rect 49369 16406 49394 16496
rect 49557 16406 49603 16496
rect 55903 16501 56137 16535
rect 49369 16375 49603 16406
rect 42816 14896 43050 14930
rect 42816 14806 42841 14896
rect 43004 14806 43050 14896
rect 55903 16411 55928 16501
rect 56091 16411 56137 16501
rect 72477 17569 72501 17673
rect 72547 17569 72583 17673
rect 72477 17529 72583 17569
rect 62416 16504 62650 16538
rect 55903 16380 56137 16411
rect 49374 14892 49608 14926
rect 41463 14736 41618 14782
rect 42816 14775 43050 14806
rect 49374 14802 49399 14892
rect 49562 14802 49608 14892
rect 62416 16414 62441 16504
rect 62604 16414 62650 16504
rect 62416 16383 62650 16414
rect 55908 14897 56142 14931
rect 41463 14573 41497 14736
rect 41587 14573 41618 14736
rect 41463 14548 41618 14573
rect 48021 14732 48176 14778
rect 49374 14771 49608 14802
rect 55908 14807 55933 14897
rect 56096 14807 56142 14897
rect 62421 14900 62655 14934
rect 48021 14569 48055 14732
rect 48145 14569 48176 14732
rect 48021 14544 48176 14569
rect 54555 14737 54710 14783
rect 55908 14776 56142 14807
rect 62421 14810 62446 14900
rect 62609 14810 62655 14900
rect 54555 14574 54589 14737
rect 54679 14574 54710 14737
rect 54555 14549 54710 14574
rect 61068 14740 61223 14786
rect 62421 14779 62655 14810
rect 61068 14577 61102 14740
rect 61192 14577 61223 14740
rect 61068 14552 61223 14577
rect 72473 14541 72579 14583
rect 72473 14437 72497 14541
rect 72543 14437 72579 14541
rect 72473 14397 72579 14437
rect 1718 12870 1904 12894
rect 1718 12824 1758 12870
rect 1862 12824 1904 12870
rect 1718 12788 1904 12824
rect 4862 12870 5048 12894
rect 4862 12824 4902 12870
rect 5006 12824 5048 12870
rect 4862 12788 5048 12824
rect 7994 12866 8180 12890
rect 7994 12820 8034 12866
rect 8138 12820 8180 12866
rect 7994 12784 8180 12820
rect 11138 12866 11324 12890
rect 11138 12820 11178 12866
rect 11282 12820 11324 12866
rect 11138 12784 11324 12820
rect 14340 12870 14526 12894
rect 14340 12824 14380 12870
rect 14484 12824 14526 12870
rect 14340 12788 14526 12824
rect 17484 12870 17670 12894
rect 17484 12824 17524 12870
rect 17628 12824 17670 12870
rect 17484 12788 17670 12824
rect 20616 12866 20802 12890
rect 20616 12820 20656 12866
rect 20760 12820 20802 12866
rect 20616 12784 20802 12820
rect 23760 12866 23946 12890
rect 23760 12820 23800 12866
rect 23904 12820 23946 12866
rect 23760 12784 23946 12820
rect 31935 12433 32033 12491
rect 31935 12301 31955 12433
rect 32011 12301 32033 12433
rect 31935 12239 32033 12301
rect 42059 11169 42271 11199
rect 42059 11113 42099 11169
rect 42233 11113 42271 11169
rect 42059 11091 42271 11113
rect 48608 11168 48820 11198
rect 48608 11112 48648 11168
rect 48782 11112 48820 11168
rect 48608 11090 48820 11112
rect 55262 11189 55474 11219
rect 55262 11133 55302 11189
rect 55436 11133 55474 11189
rect 55262 11111 55474 11133
rect 63915 11022 64127 11052
rect 63915 10966 63955 11022
rect 64089 10966 64127 11022
rect 63915 10944 64127 10966
rect 31933 10365 32031 10423
rect 1718 10136 1904 10160
rect 1718 10090 1758 10136
rect 1862 10090 1904 10136
rect 1718 10054 1904 10090
rect 4862 10136 5048 10160
rect 4862 10090 4902 10136
rect 5006 10090 5048 10136
rect 4862 10054 5048 10090
rect 7994 10132 8180 10156
rect 7994 10086 8034 10132
rect 8138 10086 8180 10132
rect 7994 10050 8180 10086
rect 11138 10132 11324 10156
rect 11138 10086 11178 10132
rect 11282 10086 11324 10132
rect 11138 10050 11324 10086
rect 14340 10136 14526 10160
rect 14340 10090 14380 10136
rect 14484 10090 14526 10136
rect 14340 10054 14526 10090
rect 17484 10136 17670 10160
rect 17484 10090 17524 10136
rect 17628 10090 17670 10136
rect 17484 10054 17670 10090
rect 20616 10132 20802 10156
rect 20616 10086 20656 10132
rect 20760 10086 20802 10132
rect 20616 10050 20802 10086
rect 23760 10132 23946 10156
rect 23760 10086 23800 10132
rect 23904 10086 23946 10132
rect 23760 10050 23946 10086
rect 31933 10233 31953 10365
rect 32009 10233 32031 10365
rect 31933 10171 32031 10233
rect 72473 11397 72579 11439
rect 72473 11293 72497 11397
rect 72543 11293 72579 11397
rect 72473 11253 72579 11293
rect 67516 10614 67728 10644
rect 67516 10558 67556 10614
rect 67690 10558 67728 10614
rect 67516 10536 67728 10558
rect 35395 9269 35607 9299
rect 35395 9213 35435 9269
rect 35569 9213 35607 9269
rect 35395 9191 35607 9213
rect 38557 9207 38791 9241
rect 38557 9117 38603 9207
rect 38766 9117 38791 9207
rect 38557 9086 38791 9117
rect 45106 9295 45340 9329
rect 45106 9205 45152 9295
rect 45315 9205 45340 9295
rect 45106 9174 45340 9205
rect 65926 9813 66168 9825
rect 51760 9227 51994 9261
rect 51760 9137 51806 9227
rect 51969 9137 51994 9227
rect 51760 9106 51994 9137
rect 65926 9711 65973 9813
rect 66108 9711 66168 9813
rect 65926 9694 66168 9711
rect 58385 9295 58619 9329
rect 58385 9205 58431 9295
rect 58594 9205 58619 9295
rect 58385 9174 58619 9205
rect 46603 8924 46758 8970
rect 40054 8836 40209 8882
rect 40054 8673 40085 8836
rect 40175 8673 40209 8836
rect 40054 8648 40209 8673
rect 41196 8834 41351 8880
rect 41196 8671 41227 8834
rect 41317 8671 41351 8834
rect 41196 8646 41351 8671
rect 46603 8761 46634 8924
rect 46724 8761 46758 8924
rect 46603 8736 46758 8761
rect 47745 8922 47900 8968
rect 47745 8759 47776 8922
rect 47866 8759 47900 8922
rect 59882 8924 60037 8970
rect 53257 8856 53412 8902
rect 47745 8734 47900 8759
rect 53257 8693 53288 8856
rect 53378 8693 53412 8856
rect 53257 8668 53412 8693
rect 54399 8854 54554 8900
rect 54399 8691 54430 8854
rect 54520 8691 54554 8854
rect 54399 8666 54554 8691
rect 59882 8761 59913 8924
rect 60003 8761 60037 8924
rect 59882 8736 60037 8761
rect 61024 8922 61179 8968
rect 61024 8759 61055 8922
rect 61145 8759 61179 8922
rect 61024 8734 61179 8759
rect 31935 8296 32033 8354
rect 31935 8164 31955 8296
rect 32011 8164 32033 8296
rect 31935 8102 32033 8164
rect 63910 8451 64122 8481
rect 63910 8395 63950 8451
rect 64084 8395 64122 8451
rect 63910 8373 64122 8395
rect 38571 7557 38805 7591
rect 1728 7404 1914 7428
rect 1728 7358 1768 7404
rect 1872 7358 1914 7404
rect 1728 7322 1914 7358
rect 4872 7404 5058 7428
rect 4872 7358 4912 7404
rect 5016 7358 5058 7404
rect 4872 7322 5058 7358
rect 8004 7400 8190 7424
rect 8004 7354 8044 7400
rect 8148 7354 8190 7400
rect 8004 7318 8190 7354
rect 11148 7400 11334 7424
rect 11148 7354 11188 7400
rect 11292 7354 11334 7400
rect 11148 7318 11334 7354
rect 14350 7404 14536 7428
rect 14350 7358 14390 7404
rect 14494 7358 14536 7404
rect 14350 7322 14536 7358
rect 17494 7404 17680 7428
rect 17494 7358 17534 7404
rect 17638 7358 17680 7404
rect 17494 7322 17680 7358
rect 20626 7400 20812 7424
rect 20626 7354 20666 7400
rect 20770 7354 20812 7400
rect 20626 7318 20812 7354
rect 23770 7400 23956 7424
rect 23770 7354 23810 7400
rect 23914 7354 23956 7400
rect 23770 7318 23956 7354
rect 38571 7467 38617 7557
rect 38780 7467 38805 7557
rect 45120 7645 45354 7679
rect 38571 7436 38805 7467
rect 35387 6684 35599 6714
rect 3261 5871 3521 5917
rect 3261 5801 3315 5871
rect 3459 5801 3521 5871
rect 3261 5767 3521 5801
rect 3999 5871 4259 5917
rect 3999 5801 4053 5871
rect 4197 5801 4259 5871
rect 3999 5767 4259 5801
rect 4737 5871 4997 5917
rect 4737 5801 4791 5871
rect 4935 5801 4997 5871
rect 4737 5767 4997 5801
rect 5475 5871 5735 5917
rect 5475 5801 5529 5871
rect 5673 5801 5735 5871
rect 5475 5767 5735 5801
rect 6215 5871 6475 5917
rect 6215 5801 6269 5871
rect 6413 5801 6475 5871
rect 6215 5767 6475 5801
rect 6957 5871 7217 5917
rect 6957 5801 7011 5871
rect 7155 5801 7217 5871
rect 6957 5767 7217 5801
rect 7695 5871 7955 5917
rect 7695 5801 7749 5871
rect 7893 5801 7955 5871
rect 7695 5767 7955 5801
rect 8433 5873 8693 5919
rect 8433 5803 8487 5873
rect 8631 5803 8693 5873
rect 8433 5769 8693 5803
rect 35387 6628 35427 6684
rect 35561 6628 35599 6684
rect 35387 6606 35599 6628
rect 45120 7555 45166 7645
rect 45329 7555 45354 7645
rect 72477 8195 72583 8237
rect 45120 7524 45354 7555
rect 31933 6228 32031 6286
rect 31933 6096 31953 6228
rect 32009 6096 32031 6228
rect 31933 6034 32031 6096
rect 51774 7577 52008 7611
rect 51774 7487 51820 7577
rect 51983 7487 52008 7577
rect 58399 7645 58633 7679
rect 51774 7456 52008 7487
rect 38566 5953 38800 5987
rect 58399 7555 58445 7645
rect 58608 7555 58633 7645
rect 58399 7524 58633 7555
rect 45115 6041 45349 6075
rect 38566 5863 38612 5953
rect 38775 5863 38800 5953
rect 45115 5951 45161 6041
rect 45324 5951 45349 6041
rect 45115 5920 45349 5951
rect 38566 5832 38800 5863
rect 46547 5881 46702 5927
rect 72477 8091 72501 8195
rect 72547 8091 72583 8195
rect 72477 8051 72583 8091
rect 51769 5973 52003 6007
rect 67518 6523 67730 6553
rect 67518 6467 67558 6523
rect 67692 6467 67730 6523
rect 67518 6445 67730 6467
rect 58394 6041 58628 6075
rect 39998 5793 40153 5839
rect 39998 5630 40029 5793
rect 40119 5630 40153 5793
rect 46547 5718 46578 5881
rect 46668 5718 46702 5881
rect 51769 5883 51815 5973
rect 51978 5883 52003 5973
rect 58394 5951 58440 6041
rect 58603 5951 58628 6041
rect 58394 5920 58628 5951
rect 51769 5852 52003 5883
rect 59826 5881 59981 5927
rect 46547 5693 46702 5718
rect 53201 5813 53356 5859
rect 39998 5605 40153 5630
rect 53201 5650 53232 5813
rect 53322 5650 53356 5813
rect 59826 5718 59857 5881
rect 59947 5718 59981 5881
rect 59826 5693 59981 5718
rect 53201 5625 53356 5650
rect 65928 5722 66170 5734
rect 65928 5620 65975 5722
rect 66110 5620 66170 5722
rect 65928 5603 66170 5620
rect 63910 5418 64122 5448
rect 63910 5362 63950 5418
rect 64084 5362 64122 5418
rect 63910 5340 64122 5362
rect 72477 5051 72583 5093
rect 10013 4446 10265 4466
rect 10013 4390 10075 4446
rect 10207 4390 10265 4446
rect 10013 4368 10265 4390
rect 12081 4444 12333 4464
rect 12081 4388 12143 4444
rect 12275 4388 12333 4444
rect 12081 4366 12333 4388
rect 14150 4446 14402 4466
rect 14150 4390 14212 4446
rect 14344 4390 14402 4446
rect 14150 4368 14402 4390
rect 16218 4444 16470 4464
rect 16218 4388 16280 4444
rect 16412 4388 16470 4444
rect 16218 4366 16470 4388
rect 18287 4444 18539 4464
rect 18287 4388 18349 4444
rect 18481 4388 18539 4444
rect 18287 4366 18539 4388
rect 20355 4442 20607 4462
rect 20355 4386 20417 4442
rect 20549 4386 20607 4442
rect 20355 4364 20607 4386
rect 22424 4444 22676 4464
rect 22424 4388 22486 4444
rect 22618 4388 22676 4444
rect 22424 4366 22676 4388
rect 24492 4442 24744 4462
rect 24492 4386 24554 4442
rect 24686 4386 24744 4442
rect 24492 4364 24744 4386
rect 31933 4159 32031 4217
rect 31933 4027 31953 4159
rect 32009 4027 32031 4159
rect 31933 3965 32031 4027
rect 35368 3406 35580 3436
rect 35368 3350 35408 3406
rect 35542 3350 35580 3406
rect 38549 3427 38783 3461
rect 35368 3328 35580 3350
rect 38549 3337 38595 3427
rect 38758 3337 38783 3427
rect 38549 3306 38783 3337
rect 72477 4947 72501 5051
rect 72547 4947 72583 5051
rect 72477 4907 72583 4947
rect 45100 3425 45334 3459
rect 45100 3335 45146 3425
rect 45309 3335 45334 3425
rect 45100 3304 45334 3335
rect 51755 3426 51989 3460
rect 51755 3336 51801 3426
rect 51964 3336 51989 3426
rect 51755 3305 51989 3336
rect 63981 3498 64193 3528
rect 58377 3427 58611 3461
rect 58377 3337 58423 3427
rect 58586 3337 58611 3427
rect 58377 3306 58611 3337
rect 63981 3442 64021 3498
rect 64155 3442 64193 3498
rect 63981 3420 64193 3442
rect 40046 3056 40201 3102
rect 40046 2893 40077 3056
rect 40167 2893 40201 3056
rect 40046 2868 40201 2893
rect 41188 3054 41343 3100
rect 41188 2891 41219 3054
rect 41309 2891 41343 3054
rect 46597 3054 46752 3100
rect 41188 2866 41343 2891
rect 46597 2891 46628 3054
rect 46718 2891 46752 3054
rect 46597 2866 46752 2891
rect 47739 3052 47894 3098
rect 47739 2889 47770 3052
rect 47860 2889 47894 3052
rect 53252 3055 53407 3101
rect 47739 2864 47894 2889
rect 53252 2892 53283 3055
rect 53373 2892 53407 3055
rect 53252 2867 53407 2892
rect 54394 3053 54549 3099
rect 54394 2890 54425 3053
rect 54515 2890 54549 3053
rect 59874 3056 60029 3102
rect 54394 2865 54549 2890
rect 59874 2893 59905 3056
rect 59995 2893 60029 3056
rect 59874 2868 60029 2893
rect 61016 3054 61171 3100
rect 61016 2891 61047 3054
rect 61137 2891 61171 3054
rect 61016 2866 61171 2891
rect 67518 3028 67730 3058
rect 67518 2972 67558 3028
rect 67692 2972 67730 3028
rect 67518 2950 67730 2972
rect 31931 2091 32029 2149
rect 31931 1959 31951 2091
rect 32007 1959 32029 2091
rect 31931 1897 32029 1959
rect 38563 1777 38797 1811
rect 38563 1687 38609 1777
rect 38772 1687 38797 1777
rect 38563 1656 38797 1687
rect 35384 646 35596 676
rect 35384 590 35424 646
rect 35558 590 35596 646
rect 35384 568 35596 590
rect 45114 1775 45348 1809
rect 45114 1685 45160 1775
rect 45323 1685 45348 1775
rect 45114 1654 45348 1685
rect 1462 152 1648 176
rect 1462 106 1504 152
rect 1608 106 1648 152
rect 1462 70 1648 106
rect 4606 152 4792 176
rect 4606 106 4648 152
rect 4752 106 4792 152
rect 4606 70 4792 106
rect 7738 156 7924 180
rect 7738 110 7780 156
rect 7884 110 7924 156
rect 7738 74 7924 110
rect 10882 156 11068 180
rect 10882 110 10924 156
rect 11028 110 11068 156
rect 10882 74 11068 110
rect 14084 152 14270 176
rect 14084 106 14126 152
rect 14230 106 14270 152
rect 14084 70 14270 106
rect 17228 152 17414 176
rect 17228 106 17270 152
rect 17374 106 17414 152
rect 17228 70 17414 106
rect 20360 156 20546 180
rect 20360 110 20402 156
rect 20506 110 20546 156
rect 20360 74 20546 110
rect 23504 156 23690 180
rect 23504 110 23546 156
rect 23650 110 23690 156
rect 23504 74 23690 110
rect 51769 1776 52003 1810
rect 51769 1686 51815 1776
rect 51978 1686 52003 1776
rect 65928 2227 66170 2239
rect 51769 1655 52003 1686
rect 38558 173 38792 207
rect 31933 22 32031 80
rect 38558 83 38604 173
rect 38767 83 38792 173
rect 58391 1777 58625 1811
rect 58391 1687 58437 1777
rect 58600 1687 58625 1777
rect 65928 2125 65975 2227
rect 66110 2125 66170 2227
rect 65928 2108 66170 2125
rect 72473 1919 72579 1961
rect 58391 1656 58625 1687
rect 45109 171 45343 205
rect 38558 52 38792 83
rect 31933 -110 31953 22
rect 32009 -110 32031 22
rect 31933 -172 32031 -110
rect 39990 13 40145 59
rect 45109 81 45155 171
rect 45318 81 45343 171
rect 72473 1815 72497 1919
rect 72543 1815 72579 1919
rect 72473 1775 72579 1815
rect 51764 172 51998 206
rect 45109 50 45343 81
rect 39990 -150 40021 13
rect 40111 -150 40145 13
rect 39990 -175 40145 -150
rect 46541 11 46696 57
rect 51764 82 51810 172
rect 51973 82 51998 172
rect 63978 428 64190 458
rect 63978 372 64018 428
rect 64152 372 64190 428
rect 63978 350 64190 372
rect 58386 173 58620 207
rect 51764 51 51998 82
rect 46541 -152 46572 11
rect 46662 -152 46696 11
rect 46541 -177 46696 -152
rect 53196 12 53351 58
rect 58386 83 58432 173
rect 58595 83 58620 173
rect 58386 52 58620 83
rect 53196 -151 53227 12
rect 53317 -151 53351 12
rect 53196 -176 53351 -151
rect 59818 13 59973 59
rect 59818 -150 59849 13
rect 59939 -150 59973 13
rect 59818 -175 59973 -150
rect 42094 -719 42306 -697
rect 42094 -775 42134 -719
rect 42268 -775 42306 -719
rect 42094 -805 42306 -775
rect 48648 -714 48860 -692
rect 48648 -770 48688 -714
rect 48822 -770 48860 -714
rect 48648 -800 48860 -770
rect 55297 -726 55509 -704
rect 55297 -782 55337 -726
rect 55471 -782 55509 -726
rect 55297 -812 55509 -782
rect 67518 -1320 67730 -1290
rect 67518 -1376 67558 -1320
rect 67692 -1376 67730 -1320
rect 67518 -1398 67730 -1376
rect 72473 -1225 72579 -1183
rect 31931 -2046 32029 -1988
rect 31931 -2178 31951 -2046
rect 32007 -2178 32029 -2046
rect 31931 -2240 32029 -2178
rect 72473 -1329 72497 -1225
rect 72543 -1329 72579 -1225
rect 72473 -1369 72579 -1329
rect 65928 -2121 66170 -2109
rect 65928 -2223 65975 -2121
rect 66110 -2223 66170 -2121
rect 65928 -2240 66170 -2223
rect 63985 -2417 64197 -2387
rect 63985 -2473 64025 -2417
rect 64159 -2473 64197 -2417
rect 63985 -2495 64197 -2473
rect 1494 -3740 1680 -3716
rect 1494 -3786 1536 -3740
rect 1640 -3786 1680 -3740
rect 1494 -3822 1680 -3786
rect 4638 -3740 4824 -3716
rect 4638 -3786 4680 -3740
rect 4784 -3786 4824 -3740
rect 4638 -3822 4824 -3786
rect 7770 -3736 7956 -3712
rect 7770 -3782 7812 -3736
rect 7916 -3782 7956 -3736
rect 7770 -3818 7956 -3782
rect 10914 -3736 11100 -3712
rect 10914 -3782 10956 -3736
rect 11060 -3782 11100 -3736
rect 10914 -3818 11100 -3782
rect 14116 -3740 14302 -3716
rect 14116 -3786 14158 -3740
rect 14262 -3786 14302 -3740
rect 14116 -3822 14302 -3786
rect 17260 -3740 17446 -3716
rect 17260 -3786 17302 -3740
rect 17406 -3786 17446 -3740
rect 17260 -3822 17446 -3786
rect 20392 -3736 20578 -3712
rect 20392 -3782 20434 -3736
rect 20538 -3782 20578 -3736
rect 20392 -3818 20578 -3782
rect 23536 -3736 23722 -3712
rect 23536 -3782 23578 -3736
rect 23682 -3782 23722 -3736
rect 23536 -3818 23722 -3782
<< nsubdiff >>
rect 42513 24989 42666 25029
rect 40031 24935 40184 24975
rect 40031 24786 40074 24935
rect 40141 24786 40184 24935
rect 40031 24717 40184 24786
rect 42513 24840 42556 24989
rect 42623 24840 42666 24989
rect 42513 24771 42666 24840
rect 43660 24989 43813 25029
rect 43660 24840 43703 24989
rect 43770 24840 43813 24989
rect 49026 24986 49179 25026
rect 43660 24771 43813 24840
rect 46544 24932 46697 24972
rect 46544 24783 46587 24932
rect 46654 24783 46697 24932
rect 46544 24714 46697 24783
rect 49026 24837 49069 24986
rect 49136 24837 49179 24986
rect 49026 24768 49179 24837
rect 50173 24986 50326 25026
rect 50173 24837 50216 24986
rect 50283 24837 50326 24986
rect 55560 24981 55713 25021
rect 50173 24768 50326 24837
rect 53078 24927 53231 24967
rect 53078 24778 53121 24927
rect 53188 24778 53231 24927
rect 53078 24709 53231 24778
rect 55560 24832 55603 24981
rect 55670 24832 55713 24981
rect 55560 24763 55713 24832
rect 56707 24981 56860 25021
rect 56707 24832 56750 24981
rect 56817 24832 56860 24981
rect 62118 24985 62271 25025
rect 56707 24763 56860 24832
rect 59636 24931 59789 24971
rect 59636 24782 59679 24931
rect 59746 24782 59789 24931
rect 59636 24713 59789 24782
rect 62118 24836 62161 24985
rect 62228 24836 62271 24985
rect 62118 24767 62271 24836
rect 63265 24985 63418 25025
rect 63265 24836 63308 24985
rect 63375 24836 63418 24985
rect 63265 24767 63418 24836
rect 40045 23285 40198 23325
rect 40045 23136 40088 23285
rect 40155 23136 40198 23285
rect 46558 23282 46711 23322
rect 40045 23067 40198 23136
rect 46558 23133 46601 23282
rect 46668 23133 46711 23282
rect 53092 23277 53245 23317
rect 46558 23064 46711 23133
rect 53092 23128 53135 23277
rect 53202 23128 53245 23277
rect 59650 23281 59803 23321
rect 53092 23059 53245 23128
rect 59650 23132 59693 23281
rect 59760 23132 59803 23281
rect 59650 23063 59803 23132
rect 43756 22942 43909 22982
rect 43756 22793 43799 22942
rect 43866 22793 43909 22942
rect 50269 22939 50422 22979
rect 43756 22724 43909 22793
rect 50269 22790 50312 22939
rect 50379 22790 50422 22939
rect 56803 22934 56956 22974
rect 63361 22938 63514 22978
rect 50269 22721 50422 22790
rect 4172 22254 4476 22310
rect 4172 22178 4226 22254
rect 4422 22178 4476 22254
rect 4172 22164 4476 22178
rect 7316 22254 7620 22310
rect 7316 22178 7370 22254
rect 7566 22178 7620 22254
rect 7316 22164 7620 22178
rect 10448 22250 10752 22306
rect 10448 22174 10502 22250
rect 10698 22174 10752 22250
rect 10448 22160 10752 22174
rect 13592 22250 13896 22306
rect 13592 22174 13646 22250
rect 13842 22174 13896 22250
rect 13592 22160 13896 22174
rect 16794 22254 17098 22310
rect 16794 22178 16848 22254
rect 17044 22178 17098 22254
rect 16794 22164 17098 22178
rect 19938 22254 20242 22310
rect 19938 22178 19992 22254
rect 20188 22178 20242 22254
rect 19938 22164 20242 22178
rect 23070 22250 23374 22306
rect 23070 22174 23124 22250
rect 23320 22174 23374 22250
rect 23070 22160 23374 22174
rect 26214 22250 26518 22306
rect 26214 22174 26268 22250
rect 26464 22174 26518 22250
rect 26214 22160 26518 22174
rect 56803 22785 56846 22934
rect 56913 22785 56956 22934
rect 56803 22716 56956 22785
rect 63361 22789 63404 22938
rect 63471 22789 63514 22938
rect 63361 22720 63514 22789
rect 40040 21681 40193 21721
rect 40040 21532 40083 21681
rect 40150 21532 40193 21681
rect 40040 21463 40193 21532
rect 46553 21678 46706 21718
rect 46553 21529 46596 21678
rect 46663 21529 46706 21678
rect 46553 21460 46706 21529
rect 53087 21673 53240 21713
rect 53087 21524 53130 21673
rect 53197 21524 53240 21673
rect 53087 21455 53240 21524
rect 59645 21677 59798 21717
rect 59645 21528 59688 21677
rect 59755 21528 59798 21677
rect 59645 21459 59798 21528
rect 70199 20875 70345 20929
rect 70199 20679 70255 20875
rect 70331 20679 70345 20875
rect 70199 20625 70345 20679
rect 39607 19381 39760 19421
rect 39607 19232 39650 19381
rect 39717 19232 39760 19381
rect 39607 19163 39760 19232
rect 40754 19381 40907 19421
rect 40754 19232 40797 19381
rect 40864 19232 40907 19381
rect 46165 19377 46318 19417
rect 40754 19163 40907 19232
rect 43236 19327 43389 19367
rect 43236 19178 43279 19327
rect 43346 19178 43389 19327
rect 43236 19109 43389 19178
rect 46165 19228 46208 19377
rect 46275 19228 46318 19377
rect 46165 19159 46318 19228
rect 47312 19377 47465 19417
rect 47312 19228 47355 19377
rect 47422 19228 47465 19377
rect 52699 19382 52852 19422
rect 47312 19159 47465 19228
rect 49794 19323 49947 19363
rect 49794 19174 49837 19323
rect 49904 19174 49947 19323
rect 49794 19105 49947 19174
rect 52699 19233 52742 19382
rect 52809 19233 52852 19382
rect 52699 19164 52852 19233
rect 53846 19382 53999 19422
rect 53846 19233 53889 19382
rect 53956 19233 53999 19382
rect 59212 19385 59365 19425
rect 53846 19164 53999 19233
rect 56328 19328 56481 19368
rect 56328 19179 56371 19328
rect 56438 19179 56481 19328
rect 56328 19110 56481 19179
rect 59212 19236 59255 19385
rect 59322 19236 59365 19385
rect 59212 19167 59365 19236
rect 60359 19385 60512 19425
rect 60359 19236 60402 19385
rect 60469 19236 60512 19385
rect 60359 19167 60512 19236
rect 62841 19331 62994 19371
rect 62841 19182 62884 19331
rect 62951 19182 62994 19331
rect 62841 19113 62994 19182
rect 43222 17677 43375 17717
rect 43222 17528 43265 17677
rect 43332 17528 43375 17677
rect 49780 17673 49933 17713
rect 43222 17459 43375 17528
rect 49780 17524 49823 17673
rect 49890 17524 49933 17673
rect 56314 17678 56467 17718
rect 49780 17455 49933 17524
rect 56314 17529 56357 17678
rect 56424 17529 56467 17678
rect 70199 17731 70345 17785
rect 62827 17681 62980 17721
rect 56314 17460 56467 17529
rect 62827 17532 62870 17681
rect 62937 17532 62980 17681
rect 62827 17463 62980 17532
rect 70199 17535 70255 17731
rect 70331 17535 70345 17731
rect 70199 17481 70345 17535
rect 39511 17334 39664 17374
rect 39511 17185 39554 17334
rect 39621 17185 39664 17334
rect 46069 17330 46222 17370
rect 39511 17116 39664 17185
rect 4524 17048 4790 17086
rect 4524 16976 4590 17048
rect 4734 16976 4790 17048
rect 5692 17048 5958 17086
rect 4524 16946 4790 16976
rect 5692 16976 5758 17048
rect 5902 16976 5958 17048
rect 6860 17048 7126 17086
rect 5692 16946 5958 16976
rect 6860 16976 6926 17048
rect 7070 16976 7126 17048
rect 8028 17048 8294 17086
rect 6860 16946 7126 16976
rect 8028 16976 8094 17048
rect 8238 16976 8294 17048
rect 9202 17046 9468 17084
rect 8028 16946 8294 16976
rect 9202 16974 9268 17046
rect 9412 16974 9468 17046
rect 10370 17046 10636 17084
rect 9202 16944 9468 16974
rect 10370 16974 10436 17046
rect 10580 16974 10636 17046
rect 11538 17046 11804 17084
rect 10370 16944 10636 16974
rect 11538 16974 11604 17046
rect 11748 16974 11804 17046
rect 12706 17046 12972 17084
rect 46069 17181 46112 17330
rect 46179 17181 46222 17330
rect 52603 17335 52756 17375
rect 46069 17112 46222 17181
rect 11538 16944 11804 16974
rect 12706 16974 12772 17046
rect 12916 16974 12972 17046
rect 52603 17186 52646 17335
rect 52713 17186 52756 17335
rect 59116 17338 59269 17378
rect 52603 17117 52756 17186
rect 59116 17189 59159 17338
rect 59226 17189 59269 17338
rect 59116 17120 59269 17189
rect 12706 16944 12972 16974
rect 14406 16841 14650 16879
rect 14406 16771 14458 16841
rect 14594 16771 14650 16841
rect 14406 16749 14650 16771
rect 15854 16841 16098 16879
rect 15854 16771 15906 16841
rect 16042 16771 16098 16841
rect 15854 16749 16098 16771
rect 17352 16839 17596 16877
rect 17352 16769 17404 16839
rect 17540 16769 17596 16839
rect 17352 16747 17596 16769
rect 18800 16839 19044 16877
rect 18800 16769 18852 16839
rect 18988 16769 19044 16839
rect 18800 16747 19044 16769
rect 20320 16841 20564 16879
rect 20320 16771 20372 16841
rect 20508 16771 20564 16841
rect 20320 16749 20564 16771
rect 21768 16841 22012 16879
rect 21768 16771 21820 16841
rect 21956 16771 22012 16841
rect 21768 16749 22012 16771
rect 23266 16839 23510 16877
rect 23266 16769 23318 16839
rect 23454 16769 23510 16839
rect 23266 16747 23510 16769
rect 24714 16839 24958 16877
rect 24714 16769 24766 16839
rect 24902 16769 24958 16839
rect 24714 16747 24958 16769
rect 43227 16073 43380 16113
rect 43227 15924 43270 16073
rect 43337 15924 43380 16073
rect 43227 15855 43380 15924
rect 1670 15116 1974 15172
rect 1670 15040 1724 15116
rect 1920 15040 1974 15116
rect 1670 15026 1974 15040
rect 4814 15116 5118 15172
rect 4814 15040 4868 15116
rect 5064 15040 5118 15116
rect 4814 15026 5118 15040
rect 7946 15112 8250 15168
rect 7946 15036 8000 15112
rect 8196 15036 8250 15112
rect 7946 15022 8250 15036
rect 11090 15112 11394 15168
rect 11090 15036 11144 15112
rect 11340 15036 11394 15112
rect 11090 15022 11394 15036
rect 14292 15116 14596 15172
rect 14292 15040 14346 15116
rect 14542 15040 14596 15116
rect 14292 15026 14596 15040
rect 17436 15116 17740 15172
rect 17436 15040 17490 15116
rect 17686 15040 17740 15116
rect 17436 15026 17740 15040
rect 20568 15112 20872 15168
rect 20568 15036 20622 15112
rect 20818 15036 20872 15112
rect 20568 15022 20872 15036
rect 23712 15112 24016 15168
rect 23712 15036 23766 15112
rect 23962 15036 24016 15112
rect 23712 15022 24016 15036
rect 49785 16069 49938 16109
rect 49785 15920 49828 16069
rect 49895 15920 49938 16069
rect 49785 15851 49938 15920
rect 56319 16074 56472 16114
rect 56319 15925 56362 16074
rect 56429 15925 56472 16074
rect 56319 15856 56472 15925
rect 62832 16077 62985 16117
rect 62832 15928 62875 16077
rect 62942 15928 62985 16077
rect 62832 15859 62985 15928
rect 70195 14599 70341 14653
rect 70195 14403 70251 14599
rect 70327 14403 70341 14599
rect 70195 14349 70341 14403
rect 1670 12382 1974 12438
rect 1670 12306 1724 12382
rect 1920 12306 1974 12382
rect 1670 12292 1974 12306
rect 4814 12382 5118 12438
rect 4814 12306 4868 12382
rect 5064 12306 5118 12382
rect 4814 12292 5118 12306
rect 7946 12378 8250 12434
rect 7946 12302 8000 12378
rect 8196 12302 8250 12378
rect 7946 12288 8250 12302
rect 11090 12378 11394 12434
rect 11090 12302 11144 12378
rect 11340 12302 11394 12378
rect 11090 12288 11394 12302
rect 14292 12382 14596 12438
rect 14292 12306 14346 12382
rect 14542 12306 14596 12382
rect 14292 12292 14596 12306
rect 17436 12382 17740 12438
rect 17436 12306 17490 12382
rect 17686 12306 17740 12382
rect 17436 12292 17740 12306
rect 20568 12378 20872 12434
rect 20568 12302 20622 12378
rect 20818 12302 20872 12378
rect 20568 12288 20872 12302
rect 23712 12378 24016 12434
rect 23712 12302 23766 12378
rect 23962 12302 24016 12378
rect 23712 12288 24016 12302
rect 29643 12383 29787 12507
rect 29643 12261 29695 12383
rect 29739 12261 29787 12383
rect 29643 12107 29787 12261
rect 41819 12377 42063 12415
rect 41819 12307 41875 12377
rect 42011 12307 42063 12377
rect 41819 12285 42063 12307
rect 48368 12376 48612 12414
rect 48368 12306 48424 12376
rect 48560 12306 48612 12376
rect 48368 12284 48612 12306
rect 55022 12397 55266 12435
rect 55022 12327 55078 12397
rect 55214 12327 55266 12397
rect 55022 12305 55266 12327
rect 65868 12289 66289 12323
rect 63675 12230 63919 12268
rect 63675 12160 63731 12230
rect 63867 12160 63919 12230
rect 63675 12138 63919 12160
rect 65868 12144 65931 12289
rect 66240 12144 66289 12289
rect 65868 12123 66289 12144
rect 67276 11822 67520 11860
rect 67276 11752 67332 11822
rect 67468 11752 67520 11822
rect 67276 11730 67520 11752
rect 70195 11455 70341 11509
rect 47258 10526 47411 10566
rect 29641 10315 29785 10439
rect 29641 10193 29693 10315
rect 29737 10193 29785 10315
rect 35155 10477 35399 10515
rect 35155 10407 35211 10477
rect 35347 10407 35399 10477
rect 40709 10438 40862 10478
rect 35155 10385 35399 10407
rect 29641 10039 29785 10193
rect 38227 10384 38380 10424
rect 38227 10235 38270 10384
rect 38337 10235 38380 10384
rect 38227 10166 38380 10235
rect 40709 10289 40752 10438
rect 40819 10289 40862 10438
rect 40709 10220 40862 10289
rect 41856 10438 42009 10478
rect 41856 10289 41899 10438
rect 41966 10289 42009 10438
rect 41856 10220 42009 10289
rect 44776 10472 44929 10512
rect 44776 10323 44819 10472
rect 44886 10323 44929 10472
rect 44776 10254 44929 10323
rect 47258 10377 47301 10526
rect 47368 10377 47411 10526
rect 47258 10308 47411 10377
rect 48405 10526 48558 10566
rect 48405 10377 48448 10526
rect 48515 10377 48558 10526
rect 60537 10526 60690 10566
rect 53912 10458 54065 10498
rect 48405 10308 48558 10377
rect 51430 10404 51583 10444
rect 51430 10255 51473 10404
rect 51540 10255 51583 10404
rect 51430 10186 51583 10255
rect 53912 10309 53955 10458
rect 54022 10309 54065 10458
rect 53912 10240 54065 10309
rect 55059 10458 55212 10498
rect 55059 10309 55102 10458
rect 55169 10309 55212 10458
rect 55059 10240 55212 10309
rect 58055 10472 58208 10512
rect 58055 10323 58098 10472
rect 58165 10323 58208 10472
rect 58055 10254 58208 10323
rect 60537 10377 60580 10526
rect 60647 10377 60690 10526
rect 60537 10308 60690 10377
rect 61684 10526 61837 10566
rect 61684 10377 61727 10526
rect 61794 10377 61837 10526
rect 61684 10308 61837 10377
rect 70195 11259 70251 11455
rect 70327 11259 70341 11455
rect 70195 11205 70341 11259
rect 1680 9650 1984 9706
rect 1680 9574 1734 9650
rect 1930 9574 1984 9650
rect 1680 9560 1984 9574
rect 4824 9650 5128 9706
rect 4824 9574 4878 9650
rect 5074 9574 5128 9650
rect 4824 9560 5128 9574
rect 7956 9646 8260 9702
rect 7956 9570 8010 9646
rect 8206 9570 8260 9646
rect 7956 9556 8260 9570
rect 11100 9646 11404 9702
rect 11100 9570 11154 9646
rect 11350 9570 11404 9646
rect 11100 9556 11404 9570
rect 14302 9650 14606 9706
rect 14302 9574 14356 9650
rect 14552 9574 14606 9650
rect 14302 9560 14606 9574
rect 17446 9650 17750 9706
rect 17446 9574 17500 9650
rect 17696 9574 17750 9650
rect 17446 9560 17750 9574
rect 20578 9646 20882 9702
rect 20578 9570 20632 9646
rect 20828 9570 20882 9646
rect 20578 9556 20882 9570
rect 23722 9646 24026 9702
rect 23722 9570 23776 9646
rect 23972 9570 24026 9646
rect 23722 9556 24026 9570
rect 63670 9659 63914 9697
rect 63670 9589 63726 9659
rect 63862 9589 63914 9659
rect 63670 9567 63914 9589
rect 38241 8734 38394 8774
rect 38241 8585 38284 8734
rect 38351 8585 38394 8734
rect 44790 8822 44943 8862
rect 44790 8673 44833 8822
rect 44900 8673 44943 8822
rect 51444 8754 51597 8794
rect 44790 8604 44943 8673
rect 51444 8605 51487 8754
rect 51554 8605 51597 8754
rect 58069 8822 58222 8862
rect 58069 8673 58112 8822
rect 58179 8673 58222 8822
rect 38241 8516 38394 8585
rect 51444 8536 51597 8605
rect 58069 8604 58222 8673
rect 48501 8479 48654 8519
rect 29643 8246 29787 8370
rect 29643 8124 29695 8246
rect 29739 8124 29787 8246
rect 41952 8391 42105 8431
rect 29643 7970 29787 8124
rect 41952 8242 41995 8391
rect 42062 8242 42105 8391
rect 41952 8173 42105 8242
rect 48501 8330 48544 8479
rect 48611 8330 48654 8479
rect 61780 8479 61933 8519
rect 55155 8411 55308 8451
rect 48501 8261 48654 8330
rect 35147 7892 35391 7930
rect 55155 8262 55198 8411
rect 55265 8262 55308 8411
rect 55155 8193 55308 8262
rect 61780 8330 61823 8479
rect 61890 8330 61933 8479
rect 61780 8261 61933 8330
rect 70199 8253 70345 8307
rect 35147 7822 35203 7892
rect 35339 7822 35391 7892
rect 35147 7800 35391 7822
rect 3175 6751 3471 6765
rect 3175 6689 3253 6751
rect 3393 6689 3471 6751
rect 3175 6633 3471 6689
rect 3913 6751 4209 6765
rect 3913 6689 3991 6751
rect 4131 6689 4209 6751
rect 3913 6633 4209 6689
rect 4651 6751 4947 6765
rect 4651 6689 4729 6751
rect 4869 6689 4947 6751
rect 4651 6633 4947 6689
rect 5389 6751 5685 6765
rect 5389 6689 5467 6751
rect 5607 6689 5685 6751
rect 5389 6633 5685 6689
rect 6129 6751 6425 6765
rect 6129 6689 6207 6751
rect 6347 6689 6425 6751
rect 6129 6633 6425 6689
rect 6871 6751 7167 6765
rect 6871 6689 6949 6751
rect 7089 6689 7167 6751
rect 6871 6633 7167 6689
rect 7609 6751 7905 6765
rect 7609 6689 7687 6751
rect 7827 6689 7905 6751
rect 7609 6633 7905 6689
rect 8347 6753 8643 6767
rect 8347 6691 8425 6753
rect 8565 6691 8643 6753
rect 8347 6635 8643 6691
rect 9881 6706 10281 6758
rect 9881 6662 10035 6706
rect 10157 6662 10281 6706
rect 9881 6614 10281 6662
rect 11949 6704 12349 6756
rect 11949 6660 12103 6704
rect 12225 6660 12349 6704
rect 11949 6612 12349 6660
rect 14018 6706 14418 6758
rect 14018 6662 14172 6706
rect 14294 6662 14418 6706
rect 14018 6614 14418 6662
rect 16086 6704 16486 6756
rect 16086 6660 16240 6704
rect 16362 6660 16486 6704
rect 16086 6612 16486 6660
rect 18155 6704 18555 6756
rect 18155 6660 18309 6704
rect 18431 6660 18555 6704
rect 18155 6612 18555 6660
rect 20223 6702 20623 6754
rect 20223 6658 20377 6702
rect 20499 6658 20623 6702
rect 20223 6610 20623 6658
rect 22292 6704 22692 6756
rect 22292 6660 22446 6704
rect 22568 6660 22692 6704
rect 22292 6612 22692 6660
rect 24360 6702 24760 6754
rect 38236 7130 38389 7170
rect 38236 6981 38279 7130
rect 38346 6981 38389 7130
rect 38236 6912 38389 6981
rect 24360 6658 24514 6702
rect 24636 6658 24760 6702
rect 24360 6610 24760 6658
rect 29641 6178 29785 6302
rect 29641 6056 29693 6178
rect 29737 6056 29785 6178
rect 65870 8198 66291 8232
rect 65870 8053 65933 8198
rect 66242 8053 66291 8198
rect 65870 8032 66291 8053
rect 70199 8057 70255 8253
rect 70331 8057 70345 8253
rect 70199 8003 70345 8057
rect 44785 7218 44938 7258
rect 44785 7069 44828 7218
rect 44895 7069 44938 7218
rect 44785 7000 44938 7069
rect 29641 5902 29785 6056
rect 51439 7150 51592 7190
rect 51439 7001 51482 7150
rect 51549 7001 51592 7150
rect 51439 6932 51592 7001
rect 67278 7731 67522 7769
rect 58064 7218 58217 7258
rect 58064 7069 58107 7218
rect 58174 7069 58217 7218
rect 58064 7000 58217 7069
rect 67278 7661 67334 7731
rect 67470 7661 67522 7731
rect 67278 7639 67522 7661
rect 63670 6626 63914 6664
rect 63670 6556 63726 6626
rect 63862 6556 63914 6626
rect 63670 6534 63914 6556
rect 70199 5109 70345 5163
rect 70199 4913 70255 5109
rect 70331 4913 70345 5109
rect 70199 4859 70345 4913
rect 63741 4706 63985 4744
rect 40701 4658 40854 4698
rect 35128 4614 35372 4652
rect 35128 4544 35184 4614
rect 35320 4544 35372 4614
rect 35128 4522 35372 4544
rect 38219 4604 38372 4644
rect 38219 4455 38262 4604
rect 38329 4455 38372 4604
rect 38219 4386 38372 4455
rect 40701 4509 40744 4658
rect 40811 4509 40854 4658
rect 40701 4440 40854 4509
rect 41848 4658 42001 4698
rect 41848 4509 41891 4658
rect 41958 4509 42001 4658
rect 47252 4656 47405 4696
rect 41848 4440 42001 4509
rect 44770 4602 44923 4642
rect 44770 4453 44813 4602
rect 44880 4453 44923 4602
rect 29641 4109 29785 4233
rect 29641 3987 29693 4109
rect 29737 3987 29785 4109
rect 44770 4384 44923 4453
rect 47252 4507 47295 4656
rect 47362 4507 47405 4656
rect 47252 4438 47405 4507
rect 48399 4656 48552 4696
rect 48399 4507 48442 4656
rect 48509 4507 48552 4656
rect 53907 4657 54060 4697
rect 48399 4438 48552 4507
rect 51425 4603 51578 4643
rect 51425 4454 51468 4603
rect 51535 4454 51578 4603
rect 51425 4385 51578 4454
rect 53907 4508 53950 4657
rect 54017 4508 54060 4657
rect 53907 4439 54060 4508
rect 55054 4657 55207 4697
rect 55054 4508 55097 4657
rect 55164 4508 55207 4657
rect 60529 4658 60682 4698
rect 55054 4439 55207 4508
rect 58047 4604 58200 4644
rect 58047 4455 58090 4604
rect 58157 4455 58200 4604
rect 29641 3833 29785 3987
rect 58047 4386 58200 4455
rect 60529 4509 60572 4658
rect 60639 4509 60682 4658
rect 60529 4440 60682 4509
rect 61676 4658 61829 4698
rect 61676 4509 61719 4658
rect 61786 4509 61829 4658
rect 63741 4636 63797 4706
rect 63933 4636 63985 4706
rect 63741 4614 63985 4636
rect 65870 4703 66291 4737
rect 65870 4558 65933 4703
rect 66242 4558 66291 4703
rect 65870 4537 66291 4558
rect 61676 4440 61829 4509
rect 67278 4236 67522 4274
rect 67278 4166 67334 4236
rect 67470 4166 67522 4236
rect 67278 4144 67522 4166
rect 38233 2954 38386 2994
rect 38233 2805 38276 2954
rect 38343 2805 38386 2954
rect 44784 2952 44937 2992
rect 38233 2736 38386 2805
rect 44784 2803 44827 2952
rect 44894 2803 44937 2952
rect 51439 2953 51592 2993
rect 44784 2734 44937 2803
rect 51439 2804 51482 2953
rect 51549 2804 51592 2953
rect 58061 2954 58214 2994
rect 51439 2735 51592 2804
rect 58061 2805 58104 2954
rect 58171 2805 58214 2954
rect 58061 2736 58214 2805
rect 41944 2611 42097 2651
rect 1392 2398 1696 2454
rect 1392 2322 1446 2398
rect 1642 2322 1696 2398
rect 1392 2308 1696 2322
rect 4536 2398 4840 2454
rect 4536 2322 4590 2398
rect 4786 2322 4840 2398
rect 4536 2308 4840 2322
rect 7668 2402 7972 2458
rect 7668 2326 7722 2402
rect 7918 2326 7972 2402
rect 7668 2312 7972 2326
rect 10812 2402 11116 2458
rect 10812 2326 10866 2402
rect 11062 2326 11116 2402
rect 10812 2312 11116 2326
rect 14014 2398 14318 2454
rect 14014 2322 14068 2398
rect 14264 2322 14318 2398
rect 14014 2308 14318 2322
rect 17158 2398 17462 2454
rect 17158 2322 17212 2398
rect 17408 2322 17462 2398
rect 17158 2308 17462 2322
rect 20290 2402 20594 2458
rect 20290 2326 20344 2402
rect 20540 2326 20594 2402
rect 20290 2312 20594 2326
rect 23434 2402 23738 2458
rect 23434 2326 23488 2402
rect 23684 2326 23738 2402
rect 23434 2312 23738 2326
rect 41944 2462 41987 2611
rect 42054 2462 42097 2611
rect 48495 2609 48648 2649
rect 41944 2393 42097 2462
rect 29639 2041 29783 2165
rect 29639 1919 29691 2041
rect 29735 1919 29783 2041
rect 48495 2460 48538 2609
rect 48605 2460 48648 2609
rect 55150 2610 55303 2650
rect 48495 2391 48648 2460
rect 55150 2461 55193 2610
rect 55260 2461 55303 2610
rect 61772 2611 61925 2651
rect 55150 2392 55303 2461
rect 61772 2462 61815 2611
rect 61882 2462 61925 2611
rect 61772 2393 61925 2462
rect 29639 1765 29783 1919
rect 35144 1854 35388 1892
rect 35144 1784 35200 1854
rect 35336 1784 35388 1854
rect 35144 1762 35388 1784
rect 38228 1350 38381 1390
rect 38228 1201 38271 1350
rect 38338 1201 38381 1350
rect 38228 1132 38381 1201
rect 44779 1348 44932 1388
rect 44779 1199 44822 1348
rect 44889 1199 44932 1348
rect 44779 1130 44932 1199
rect 29641 -28 29785 96
rect 29641 -150 29693 -28
rect 29737 -150 29785 -28
rect 51434 1349 51587 1389
rect 51434 1200 51477 1349
rect 51544 1200 51587 1349
rect 51434 1131 51587 1200
rect 70195 1977 70341 2031
rect 70195 1781 70251 1977
rect 70327 1781 70341 1977
rect 58056 1350 58209 1390
rect 58056 1201 58099 1350
rect 58166 1201 58209 1350
rect 58056 1132 58209 1201
rect 29641 -304 29785 -150
rect 70195 1727 70341 1781
rect 63738 1636 63982 1674
rect 63738 1566 63794 1636
rect 63930 1566 63982 1636
rect 63738 1544 63982 1566
rect 65870 355 66291 389
rect 65870 210 65933 355
rect 66242 210 66291 355
rect 65870 189 66291 210
rect 67278 -112 67522 -74
rect 67278 -182 67334 -112
rect 67470 -182 67522 -112
rect 67278 -204 67522 -182
rect 1424 -1494 1728 -1438
rect 1424 -1570 1478 -1494
rect 1674 -1570 1728 -1494
rect 1424 -1584 1728 -1570
rect 4568 -1494 4872 -1438
rect 4568 -1570 4622 -1494
rect 4818 -1570 4872 -1494
rect 4568 -1584 4872 -1570
rect 7700 -1490 8004 -1434
rect 7700 -1566 7754 -1490
rect 7950 -1566 8004 -1490
rect 7700 -1580 8004 -1566
rect 10844 -1490 11148 -1434
rect 10844 -1566 10898 -1490
rect 11094 -1566 11148 -1490
rect 10844 -1580 11148 -1566
rect 14046 -1494 14350 -1438
rect 14046 -1570 14100 -1494
rect 14296 -1570 14350 -1494
rect 14046 -1584 14350 -1570
rect 17190 -1494 17494 -1438
rect 17190 -1570 17244 -1494
rect 17440 -1570 17494 -1494
rect 17190 -1584 17494 -1570
rect 20322 -1490 20626 -1434
rect 20322 -1566 20376 -1490
rect 20572 -1566 20626 -1490
rect 20322 -1580 20626 -1566
rect 23466 -1490 23770 -1434
rect 23466 -1566 23520 -1490
rect 23716 -1566 23770 -1490
rect 23466 -1580 23770 -1566
rect 63745 -1209 63989 -1171
rect 63745 -1279 63801 -1209
rect 63937 -1279 63989 -1209
rect 63745 -1301 63989 -1279
rect 70195 -1167 70341 -1113
rect 70195 -1363 70251 -1167
rect 70327 -1363 70341 -1167
rect 70195 -1417 70341 -1363
rect 29639 -2096 29783 -1972
rect 29639 -2218 29691 -2096
rect 29735 -2218 29783 -2096
rect 41854 -1913 42098 -1891
rect 41854 -1983 41910 -1913
rect 42046 -1983 42098 -1913
rect 41854 -2021 42098 -1983
rect 48408 -1908 48652 -1886
rect 48408 -1978 48464 -1908
rect 48600 -1978 48652 -1908
rect 48408 -2016 48652 -1978
rect 55057 -1920 55301 -1898
rect 55057 -1990 55113 -1920
rect 55249 -1990 55301 -1920
rect 55057 -2028 55301 -1990
rect 29639 -2372 29783 -2218
<< psubdiffcont >>
rect 40407 23668 40570 23758
rect 46920 23665 47083 23755
rect 53454 23660 53617 23750
rect 60012 23664 60175 23754
rect 41889 23224 41979 23387
rect 43031 23222 43121 23385
rect 48402 23221 48492 23384
rect 49544 23219 49634 23382
rect 54936 23216 55026 23379
rect 56078 23214 56168 23377
rect 61494 23220 61584 23383
rect 62636 23218 62726 23381
rect 40421 22018 40584 22108
rect 46934 22015 47097 22105
rect 53468 22010 53631 22100
rect 40416 20414 40579 20504
rect 60026 22014 60189 22104
rect 46929 20411 47092 20501
rect 41833 20181 41923 20344
rect 53463 20406 53626 20496
rect 48346 20178 48436 20341
rect 60021 20410 60184 20500
rect 54880 20173 54970 20336
rect 61438 20177 61528 20340
rect 72501 20713 72547 20817
rect 4260 19962 4364 20008
rect 7404 19962 7508 20008
rect 10536 19958 10640 20004
rect 13680 19958 13784 20004
rect 16882 19962 16986 20008
rect 20026 19962 20130 20008
rect 23158 19958 23262 20004
rect 26302 19958 26406 20004
rect 42850 18060 43013 18150
rect 49408 18056 49571 18146
rect 55942 18061 56105 18151
rect 62455 18064 62618 18154
rect 40299 17614 40389 17777
rect 41441 17616 41531 17779
rect 46857 17610 46947 17773
rect 47999 17612 48089 17775
rect 53391 17615 53481 17778
rect 54533 17617 54623 17780
rect 59904 17618 59994 17781
rect 61046 17620 61136 17783
rect 5072 15638 5190 15704
rect 6240 15638 6358 15704
rect 7408 15638 7526 15704
rect 8576 15638 8694 15704
rect 9750 15636 9868 15702
rect 10918 15636 11036 15702
rect 12086 15636 12204 15702
rect 13254 15636 13372 15702
rect 14236 15577 14370 15633
rect 15684 15577 15818 15633
rect 17182 15575 17316 15631
rect 18630 15575 18764 15631
rect 20150 15577 20284 15633
rect 21598 15577 21732 15633
rect 23096 15575 23230 15631
rect 24544 15575 24678 15631
rect 42836 16410 42999 16500
rect 49394 16406 49557 16496
rect 42841 14806 43004 14896
rect 55928 16411 56091 16501
rect 72501 17569 72547 17673
rect 49399 14802 49562 14892
rect 62441 16414 62604 16504
rect 41497 14573 41587 14736
rect 55933 14807 56096 14897
rect 48055 14569 48145 14732
rect 62446 14810 62609 14900
rect 54589 14574 54679 14737
rect 61102 14577 61192 14740
rect 72497 14437 72543 14541
rect 1758 12824 1862 12870
rect 4902 12824 5006 12870
rect 8034 12820 8138 12866
rect 11178 12820 11282 12866
rect 14380 12824 14484 12870
rect 17524 12824 17628 12870
rect 20656 12820 20760 12866
rect 23800 12820 23904 12866
rect 31955 12301 32011 12433
rect 42099 11113 42233 11169
rect 48648 11112 48782 11168
rect 55302 11133 55436 11189
rect 63955 10966 64089 11022
rect 1758 10090 1862 10136
rect 4902 10090 5006 10136
rect 8034 10086 8138 10132
rect 11178 10086 11282 10132
rect 14380 10090 14484 10136
rect 17524 10090 17628 10136
rect 20656 10086 20760 10132
rect 23800 10086 23904 10132
rect 31953 10233 32009 10365
rect 72497 11293 72543 11397
rect 67556 10558 67690 10614
rect 35435 9213 35569 9269
rect 38603 9117 38766 9207
rect 45152 9205 45315 9295
rect 51806 9137 51969 9227
rect 65973 9711 66108 9813
rect 58431 9205 58594 9295
rect 40085 8673 40175 8836
rect 41227 8671 41317 8834
rect 46634 8761 46724 8924
rect 47776 8759 47866 8922
rect 53288 8693 53378 8856
rect 54430 8691 54520 8854
rect 59913 8761 60003 8924
rect 61055 8759 61145 8922
rect 31955 8164 32011 8296
rect 63950 8395 64084 8451
rect 1768 7358 1872 7404
rect 4912 7358 5016 7404
rect 8044 7354 8148 7400
rect 11188 7354 11292 7400
rect 14390 7358 14494 7404
rect 17534 7358 17638 7404
rect 20666 7354 20770 7400
rect 23810 7354 23914 7400
rect 38617 7467 38780 7557
rect 3315 5801 3459 5871
rect 4053 5801 4197 5871
rect 4791 5801 4935 5871
rect 5529 5801 5673 5871
rect 6269 5801 6413 5871
rect 7011 5801 7155 5871
rect 7749 5801 7893 5871
rect 8487 5803 8631 5873
rect 35427 6628 35561 6684
rect 45166 7555 45329 7645
rect 31953 6096 32009 6228
rect 51820 7487 51983 7577
rect 58445 7555 58608 7645
rect 38612 5863 38775 5953
rect 45161 5951 45324 6041
rect 72501 8091 72547 8195
rect 67558 6467 67692 6523
rect 40029 5630 40119 5793
rect 46578 5718 46668 5881
rect 51815 5883 51978 5973
rect 58440 5951 58603 6041
rect 53232 5650 53322 5813
rect 59857 5718 59947 5881
rect 65975 5620 66110 5722
rect 63950 5362 64084 5418
rect 10075 4390 10207 4446
rect 12143 4388 12275 4444
rect 14212 4390 14344 4446
rect 16280 4388 16412 4444
rect 18349 4388 18481 4444
rect 20417 4386 20549 4442
rect 22486 4388 22618 4444
rect 24554 4386 24686 4442
rect 31953 4027 32009 4159
rect 35408 3350 35542 3406
rect 38595 3337 38758 3427
rect 72501 4947 72547 5051
rect 45146 3335 45309 3425
rect 51801 3336 51964 3426
rect 58423 3337 58586 3427
rect 64021 3442 64155 3498
rect 40077 2893 40167 3056
rect 41219 2891 41309 3054
rect 46628 2891 46718 3054
rect 47770 2889 47860 3052
rect 53283 2892 53373 3055
rect 54425 2890 54515 3053
rect 59905 2893 59995 3056
rect 61047 2891 61137 3054
rect 67558 2972 67692 3028
rect 31951 1959 32007 2091
rect 38609 1687 38772 1777
rect 35424 590 35558 646
rect 45160 1685 45323 1775
rect 1504 106 1608 152
rect 4648 106 4752 152
rect 7780 110 7884 156
rect 10924 110 11028 156
rect 14126 106 14230 152
rect 17270 106 17374 152
rect 20402 110 20506 156
rect 23546 110 23650 156
rect 51815 1686 51978 1776
rect 38604 83 38767 173
rect 58437 1687 58600 1777
rect 65975 2125 66110 2227
rect 31953 -110 32009 22
rect 45155 81 45318 171
rect 72497 1815 72543 1919
rect 40021 -150 40111 13
rect 51810 82 51973 172
rect 64018 372 64152 428
rect 46572 -152 46662 11
rect 58432 83 58595 173
rect 53227 -151 53317 12
rect 59849 -150 59939 13
rect 42134 -775 42268 -719
rect 48688 -770 48822 -714
rect 55337 -782 55471 -726
rect 67558 -1376 67692 -1320
rect 31951 -2178 32007 -2046
rect 72497 -1329 72543 -1225
rect 65975 -2223 66110 -2121
rect 64025 -2473 64159 -2417
rect 1536 -3786 1640 -3740
rect 4680 -3786 4784 -3740
rect 7812 -3782 7916 -3736
rect 10956 -3782 11060 -3736
rect 14158 -3786 14262 -3740
rect 17302 -3786 17406 -3740
rect 20434 -3782 20538 -3736
rect 23578 -3782 23682 -3736
<< nsubdiffcont >>
rect 40074 24786 40141 24935
rect 42556 24840 42623 24989
rect 43703 24840 43770 24989
rect 46587 24783 46654 24932
rect 49069 24837 49136 24986
rect 50216 24837 50283 24986
rect 53121 24778 53188 24927
rect 55603 24832 55670 24981
rect 56750 24832 56817 24981
rect 59679 24782 59746 24931
rect 62161 24836 62228 24985
rect 63308 24836 63375 24985
rect 40088 23136 40155 23285
rect 46601 23133 46668 23282
rect 53135 23128 53202 23277
rect 59693 23132 59760 23281
rect 43799 22793 43866 22942
rect 50312 22790 50379 22939
rect 4226 22178 4422 22254
rect 7370 22178 7566 22254
rect 10502 22174 10698 22250
rect 13646 22174 13842 22250
rect 16848 22178 17044 22254
rect 19992 22178 20188 22254
rect 23124 22174 23320 22250
rect 26268 22174 26464 22250
rect 56846 22785 56913 22934
rect 63404 22789 63471 22938
rect 40083 21532 40150 21681
rect 46596 21529 46663 21678
rect 53130 21524 53197 21673
rect 59688 21528 59755 21677
rect 70255 20679 70331 20875
rect 39650 19232 39717 19381
rect 40797 19232 40864 19381
rect 43279 19178 43346 19327
rect 46208 19228 46275 19377
rect 47355 19228 47422 19377
rect 49837 19174 49904 19323
rect 52742 19233 52809 19382
rect 53889 19233 53956 19382
rect 56371 19179 56438 19328
rect 59255 19236 59322 19385
rect 60402 19236 60469 19385
rect 62884 19182 62951 19331
rect 43265 17528 43332 17677
rect 49823 17524 49890 17673
rect 56357 17529 56424 17678
rect 62870 17532 62937 17681
rect 70255 17535 70331 17731
rect 39554 17185 39621 17334
rect 4590 16976 4734 17048
rect 5758 16976 5902 17048
rect 6926 16976 7070 17048
rect 8094 16976 8238 17048
rect 9268 16974 9412 17046
rect 10436 16974 10580 17046
rect 11604 16974 11748 17046
rect 46112 17181 46179 17330
rect 12772 16974 12916 17046
rect 52646 17186 52713 17335
rect 59159 17189 59226 17338
rect 14458 16771 14594 16841
rect 15906 16771 16042 16841
rect 17404 16769 17540 16839
rect 18852 16769 18988 16839
rect 20372 16771 20508 16841
rect 21820 16771 21956 16841
rect 23318 16769 23454 16839
rect 24766 16769 24902 16839
rect 43270 15924 43337 16073
rect 1724 15040 1920 15116
rect 4868 15040 5064 15116
rect 8000 15036 8196 15112
rect 11144 15036 11340 15112
rect 14346 15040 14542 15116
rect 17490 15040 17686 15116
rect 20622 15036 20818 15112
rect 23766 15036 23962 15112
rect 49828 15920 49895 16069
rect 56362 15925 56429 16074
rect 62875 15928 62942 16077
rect 70251 14403 70327 14599
rect 1724 12306 1920 12382
rect 4868 12306 5064 12382
rect 8000 12302 8196 12378
rect 11144 12302 11340 12378
rect 14346 12306 14542 12382
rect 17490 12306 17686 12382
rect 20622 12302 20818 12378
rect 23766 12302 23962 12378
rect 29695 12261 29739 12383
rect 41875 12307 42011 12377
rect 48424 12306 48560 12376
rect 55078 12327 55214 12397
rect 63731 12160 63867 12230
rect 65931 12144 66240 12289
rect 67332 11752 67468 11822
rect 29693 10193 29737 10315
rect 35211 10407 35347 10477
rect 38270 10235 38337 10384
rect 40752 10289 40819 10438
rect 41899 10289 41966 10438
rect 44819 10323 44886 10472
rect 47301 10377 47368 10526
rect 48448 10377 48515 10526
rect 51473 10255 51540 10404
rect 53955 10309 54022 10458
rect 55102 10309 55169 10458
rect 58098 10323 58165 10472
rect 60580 10377 60647 10526
rect 61727 10377 61794 10526
rect 70251 11259 70327 11455
rect 1734 9574 1930 9650
rect 4878 9574 5074 9650
rect 8010 9570 8206 9646
rect 11154 9570 11350 9646
rect 14356 9574 14552 9650
rect 17500 9574 17696 9650
rect 20632 9570 20828 9646
rect 23776 9570 23972 9646
rect 63726 9589 63862 9659
rect 38284 8585 38351 8734
rect 44833 8673 44900 8822
rect 51487 8605 51554 8754
rect 58112 8673 58179 8822
rect 29695 8124 29739 8246
rect 41995 8242 42062 8391
rect 48544 8330 48611 8479
rect 55198 8262 55265 8411
rect 61823 8330 61890 8479
rect 35203 7822 35339 7892
rect 3253 6689 3393 6751
rect 3991 6689 4131 6751
rect 4729 6689 4869 6751
rect 5467 6689 5607 6751
rect 6207 6689 6347 6751
rect 6949 6689 7089 6751
rect 7687 6689 7827 6751
rect 8425 6691 8565 6753
rect 10035 6662 10157 6706
rect 12103 6660 12225 6704
rect 14172 6662 14294 6706
rect 16240 6660 16362 6704
rect 18309 6660 18431 6704
rect 20377 6658 20499 6702
rect 22446 6660 22568 6704
rect 38279 6981 38346 7130
rect 24514 6658 24636 6702
rect 29693 6056 29737 6178
rect 65933 8053 66242 8198
rect 70255 8057 70331 8253
rect 44828 7069 44895 7218
rect 51482 7001 51549 7150
rect 58107 7069 58174 7218
rect 67334 7661 67470 7731
rect 63726 6556 63862 6626
rect 70255 4913 70331 5109
rect 35184 4544 35320 4614
rect 38262 4455 38329 4604
rect 40744 4509 40811 4658
rect 41891 4509 41958 4658
rect 44813 4453 44880 4602
rect 29693 3987 29737 4109
rect 47295 4507 47362 4656
rect 48442 4507 48509 4656
rect 51468 4454 51535 4603
rect 53950 4508 54017 4657
rect 55097 4508 55164 4657
rect 58090 4455 58157 4604
rect 60572 4509 60639 4658
rect 61719 4509 61786 4658
rect 63797 4636 63933 4706
rect 65933 4558 66242 4703
rect 67334 4166 67470 4236
rect 38276 2805 38343 2954
rect 44827 2803 44894 2952
rect 51482 2804 51549 2953
rect 58104 2805 58171 2954
rect 1446 2322 1642 2398
rect 4590 2322 4786 2398
rect 7722 2326 7918 2402
rect 10866 2326 11062 2402
rect 14068 2322 14264 2398
rect 17212 2322 17408 2398
rect 20344 2326 20540 2402
rect 23488 2326 23684 2402
rect 41987 2462 42054 2611
rect 29691 1919 29735 2041
rect 48538 2460 48605 2609
rect 55193 2461 55260 2610
rect 61815 2462 61882 2611
rect 35200 1784 35336 1854
rect 38271 1201 38338 1350
rect 44822 1199 44889 1348
rect 29693 -150 29737 -28
rect 51477 1200 51544 1349
rect 70251 1781 70327 1977
rect 58099 1201 58166 1350
rect 63794 1566 63930 1636
rect 65933 210 66242 355
rect 67334 -182 67470 -112
rect 1478 -1570 1674 -1494
rect 4622 -1570 4818 -1494
rect 7754 -1566 7950 -1490
rect 10898 -1566 11094 -1490
rect 14100 -1570 14296 -1494
rect 17244 -1570 17440 -1494
rect 20376 -1566 20572 -1490
rect 23520 -1566 23716 -1490
rect 63801 -1279 63937 -1209
rect 70251 -1363 70327 -1167
rect 29691 -2218 29735 -2096
rect 41910 -1983 42046 -1913
rect 48464 -1978 48600 -1908
rect 55113 -1990 55249 -1920
<< poly >>
rect 41794 24769 41860 24785
rect 42924 24775 42990 24791
rect 41794 24735 41810 24769
rect 41844 24762 41860 24769
rect 41844 24735 42369 24762
rect 41794 24719 42369 24735
rect 42924 24741 42940 24775
rect 42974 24766 42990 24775
rect 42974 24741 43511 24766
rect 42924 24723 43511 24741
rect 42325 24667 42369 24719
rect 43467 24671 43511 24723
rect 48307 24766 48373 24782
rect 49437 24772 49503 24788
rect 48307 24732 48323 24766
rect 48357 24759 48373 24766
rect 48357 24732 48882 24759
rect 48307 24716 48882 24732
rect 49437 24738 49453 24772
rect 49487 24763 49503 24772
rect 49487 24738 50024 24763
rect 49437 24720 50024 24738
rect 41794 24651 42267 24667
rect 41794 24617 41810 24651
rect 41844 24626 42267 24651
rect 41844 24625 42031 24626
rect 41844 24617 41860 24625
rect 41794 24601 41860 24617
rect 41971 24605 42031 24625
rect 42089 24605 42149 24626
rect 42207 24605 42267 24626
rect 42325 24626 42621 24667
rect 42325 24605 42385 24626
rect 42443 24605 42503 24626
rect 42561 24605 42621 24626
rect 42924 24655 43409 24671
rect 42924 24621 42940 24655
rect 42974 24630 43409 24655
rect 42974 24629 43173 24630
rect 42974 24621 42990 24629
rect 42924 24605 42990 24621
rect 43113 24609 43173 24629
rect 43231 24609 43291 24630
rect 43349 24609 43409 24630
rect 43467 24630 43763 24671
rect 48838 24664 48882 24716
rect 49980 24668 50024 24720
rect 54841 24761 54907 24777
rect 55971 24767 56037 24783
rect 54841 24727 54857 24761
rect 54891 24754 54907 24761
rect 54891 24727 55416 24754
rect 54841 24711 55416 24727
rect 55971 24733 55987 24767
rect 56021 24758 56037 24767
rect 56021 24733 56558 24758
rect 55971 24715 56558 24733
rect 43467 24609 43527 24630
rect 43585 24609 43645 24630
rect 43703 24609 43763 24630
rect 48307 24648 48780 24664
rect 48307 24614 48323 24648
rect 48357 24623 48780 24648
rect 48357 24622 48544 24623
rect 48357 24614 48373 24622
rect 39646 24554 39942 24590
rect 39646 24533 39706 24554
rect 39764 24533 39824 24554
rect 39882 24533 39942 24554
rect 40000 24553 40296 24589
rect 40000 24533 40060 24553
rect 40118 24533 40178 24553
rect 40236 24533 40296 24553
rect 40354 24553 40650 24589
rect 40354 24533 40414 24553
rect 40472 24533 40532 24553
rect 40590 24533 40650 24553
rect 39646 24307 39706 24333
rect 39764 24307 39824 24333
rect 39882 24307 39942 24333
rect 40000 24313 40060 24333
rect 40000 24307 40061 24313
rect 40118 24307 40178 24333
rect 40236 24307 40296 24333
rect 39883 24122 39941 24307
rect 39883 24096 39943 24122
rect 40001 24096 40061 24307
rect 40354 24301 40414 24333
rect 40472 24307 40532 24333
rect 40590 24307 40650 24333
rect 40351 24285 40417 24301
rect 40351 24251 40367 24285
rect 40401 24251 40417 24285
rect 40351 24235 40417 24251
rect 48307 24598 48373 24614
rect 48484 24602 48544 24622
rect 48602 24602 48662 24623
rect 48720 24602 48780 24623
rect 48838 24623 49134 24664
rect 48838 24602 48898 24623
rect 48956 24602 49016 24623
rect 49074 24602 49134 24623
rect 49437 24652 49922 24668
rect 49437 24618 49453 24652
rect 49487 24627 49922 24652
rect 49487 24626 49686 24627
rect 49487 24618 49503 24626
rect 49437 24602 49503 24618
rect 49626 24606 49686 24626
rect 49744 24606 49804 24627
rect 49862 24606 49922 24627
rect 49980 24627 50276 24668
rect 55372 24659 55416 24711
rect 56514 24663 56558 24715
rect 61399 24765 61465 24781
rect 62529 24771 62595 24787
rect 61399 24731 61415 24765
rect 61449 24758 61465 24765
rect 61449 24731 61974 24758
rect 61399 24715 61974 24731
rect 62529 24737 62545 24771
rect 62579 24762 62595 24771
rect 62579 24737 63116 24762
rect 62529 24719 63116 24737
rect 61930 24663 61974 24715
rect 63072 24667 63116 24719
rect 49980 24606 50040 24627
rect 50098 24606 50158 24627
rect 50216 24606 50276 24627
rect 54841 24643 55314 24659
rect 54841 24609 54857 24643
rect 54891 24618 55314 24643
rect 54891 24617 55078 24618
rect 54891 24609 54907 24617
rect 46159 24551 46455 24587
rect 46159 24530 46219 24551
rect 46277 24530 46337 24551
rect 46395 24530 46455 24551
rect 46513 24550 46809 24586
rect 46513 24530 46573 24550
rect 46631 24530 46691 24550
rect 46749 24530 46809 24550
rect 46867 24550 47163 24586
rect 46867 24530 46927 24550
rect 46985 24530 47045 24550
rect 47103 24530 47163 24550
rect 46159 24304 46219 24330
rect 46277 24304 46337 24330
rect 46395 24304 46455 24330
rect 46513 24310 46573 24330
rect 46513 24304 46574 24310
rect 46631 24304 46691 24330
rect 46749 24304 46809 24330
rect 41971 24188 42031 24205
rect 40233 24168 40299 24184
rect 40233 24134 40249 24168
rect 40283 24134 40299 24168
rect 40233 24118 40299 24134
rect 40236 24096 40296 24118
rect 41971 24099 42032 24188
rect 42089 24179 42149 24205
rect 42207 24179 42267 24205
rect 41881 24046 42032 24099
rect 40236 23870 40296 23896
rect 41881 23822 41941 24046
rect 42325 24004 42385 24205
rect 42443 24179 42503 24205
rect 42561 24179 42621 24205
rect 43113 24192 43173 24209
rect 43113 24103 43174 24192
rect 43231 24183 43291 24209
rect 43349 24183 43409 24209
rect 41999 23953 42385 24004
rect 43023 24050 43174 24103
rect 41999 23822 42059 23953
rect 42114 23895 42180 23911
rect 42114 23861 42130 23895
rect 42164 23861 42180 23895
rect 42114 23845 42180 23861
rect 42117 23822 42177 23845
rect 42400 23822 42460 23848
rect 42518 23822 42578 23848
rect 42636 23822 42696 23848
rect 43023 23826 43083 24050
rect 43467 24008 43527 24209
rect 43585 24183 43645 24209
rect 43703 24183 43763 24209
rect 46396 24119 46454 24304
rect 46396 24093 46456 24119
rect 46514 24093 46574 24304
rect 46867 24298 46927 24330
rect 46985 24304 47045 24330
rect 47103 24304 47163 24330
rect 46864 24282 46930 24298
rect 46864 24248 46880 24282
rect 46914 24248 46930 24282
rect 46864 24232 46930 24248
rect 54841 24593 54907 24609
rect 55018 24597 55078 24617
rect 55136 24597 55196 24618
rect 55254 24597 55314 24618
rect 55372 24618 55668 24659
rect 55372 24597 55432 24618
rect 55490 24597 55550 24618
rect 55608 24597 55668 24618
rect 55971 24647 56456 24663
rect 55971 24613 55987 24647
rect 56021 24622 56456 24647
rect 56021 24621 56220 24622
rect 56021 24613 56037 24621
rect 55971 24597 56037 24613
rect 56160 24601 56220 24621
rect 56278 24601 56338 24622
rect 56396 24601 56456 24622
rect 56514 24622 56810 24663
rect 56514 24601 56574 24622
rect 56632 24601 56692 24622
rect 56750 24601 56810 24622
rect 61399 24647 61872 24663
rect 61399 24613 61415 24647
rect 61449 24622 61872 24647
rect 61449 24621 61636 24622
rect 61449 24613 61465 24621
rect 52693 24546 52989 24582
rect 52693 24525 52753 24546
rect 52811 24525 52871 24546
rect 52929 24525 52989 24546
rect 53047 24545 53343 24581
rect 53047 24525 53107 24545
rect 53165 24525 53225 24545
rect 53283 24525 53343 24545
rect 53401 24545 53697 24581
rect 53401 24525 53461 24545
rect 53519 24525 53579 24545
rect 53637 24525 53697 24545
rect 52693 24299 52753 24325
rect 52811 24299 52871 24325
rect 52929 24299 52989 24325
rect 53047 24305 53107 24325
rect 53047 24299 53108 24305
rect 53165 24299 53225 24325
rect 53283 24299 53343 24325
rect 48484 24185 48544 24202
rect 46746 24165 46812 24181
rect 46746 24131 46762 24165
rect 46796 24131 46812 24165
rect 46746 24115 46812 24131
rect 46749 24093 46809 24115
rect 48484 24096 48545 24185
rect 48602 24176 48662 24202
rect 48720 24176 48780 24202
rect 43141 23957 43527 24008
rect 43141 23826 43201 23957
rect 43256 23899 43322 23915
rect 43256 23865 43272 23899
rect 43306 23865 43322 23899
rect 43256 23849 43322 23865
rect 43259 23826 43319 23849
rect 43542 23826 43602 23852
rect 43660 23826 43720 23852
rect 43778 23826 43838 23852
rect 39883 23674 39943 23696
rect 40001 23674 40061 23696
rect 39880 23658 39946 23674
rect 39880 23624 39896 23658
rect 39930 23624 39946 23658
rect 39880 23608 39946 23624
rect 39998 23658 40064 23674
rect 39998 23624 40014 23658
rect 40048 23624 40064 23658
rect 39998 23608 40064 23624
rect 48394 24043 48545 24096
rect 46749 23867 46809 23893
rect 48394 23819 48454 24043
rect 48838 24001 48898 24202
rect 48956 24176 49016 24202
rect 49074 24176 49134 24202
rect 49626 24189 49686 24206
rect 49626 24100 49687 24189
rect 49744 24180 49804 24206
rect 49862 24180 49922 24206
rect 48512 23950 48898 24001
rect 49536 24047 49687 24100
rect 48512 23819 48572 23950
rect 48627 23892 48693 23908
rect 48627 23858 48643 23892
rect 48677 23858 48693 23892
rect 48627 23842 48693 23858
rect 48630 23819 48690 23842
rect 48913 23819 48973 23845
rect 49031 23819 49091 23845
rect 49149 23819 49209 23845
rect 49536 23823 49596 24047
rect 49980 24005 50040 24206
rect 50098 24180 50158 24206
rect 50216 24180 50276 24206
rect 52930 24114 52988 24299
rect 52930 24088 52990 24114
rect 53048 24088 53108 24299
rect 53401 24293 53461 24325
rect 53519 24299 53579 24325
rect 53637 24299 53697 24325
rect 53398 24277 53464 24293
rect 53398 24243 53414 24277
rect 53448 24243 53464 24277
rect 53398 24227 53464 24243
rect 61399 24597 61465 24613
rect 61576 24601 61636 24621
rect 61694 24601 61754 24622
rect 61812 24601 61872 24622
rect 61930 24622 62226 24663
rect 61930 24601 61990 24622
rect 62048 24601 62108 24622
rect 62166 24601 62226 24622
rect 62529 24651 63014 24667
rect 62529 24617 62545 24651
rect 62579 24626 63014 24651
rect 62579 24625 62778 24626
rect 62579 24617 62595 24625
rect 62529 24601 62595 24617
rect 62718 24605 62778 24625
rect 62836 24605 62896 24626
rect 62954 24605 63014 24626
rect 63072 24626 63368 24667
rect 63072 24605 63132 24626
rect 63190 24605 63250 24626
rect 63308 24605 63368 24626
rect 59251 24550 59547 24586
rect 59251 24529 59311 24550
rect 59369 24529 59429 24550
rect 59487 24529 59547 24550
rect 59605 24549 59901 24585
rect 59605 24529 59665 24549
rect 59723 24529 59783 24549
rect 59841 24529 59901 24549
rect 59959 24549 60255 24585
rect 59959 24529 60019 24549
rect 60077 24529 60137 24549
rect 60195 24529 60255 24549
rect 59251 24303 59311 24329
rect 59369 24303 59429 24329
rect 59487 24303 59547 24329
rect 59605 24309 59665 24329
rect 59605 24303 59666 24309
rect 59723 24303 59783 24329
rect 59841 24303 59901 24329
rect 55018 24180 55078 24197
rect 53280 24160 53346 24176
rect 53280 24126 53296 24160
rect 53330 24126 53346 24160
rect 53280 24110 53346 24126
rect 53283 24088 53343 24110
rect 55018 24091 55079 24180
rect 55136 24171 55196 24197
rect 55254 24171 55314 24197
rect 49654 23954 50040 24005
rect 49654 23823 49714 23954
rect 49769 23896 49835 23912
rect 49769 23862 49785 23896
rect 49819 23862 49835 23896
rect 49769 23846 49835 23862
rect 49772 23823 49832 23846
rect 50055 23823 50115 23849
rect 50173 23823 50233 23849
rect 50291 23823 50351 23849
rect 46396 23671 46456 23693
rect 46514 23671 46574 23693
rect 46393 23655 46459 23671
rect 41881 23596 41941 23622
rect 41999 23596 42059 23622
rect 42117 23590 42177 23622
rect 42400 23590 42460 23622
rect 42518 23590 42578 23622
rect 42636 23590 42696 23622
rect 43023 23600 43083 23626
rect 43141 23600 43201 23626
rect 42117 23549 42696 23590
rect 43259 23594 43319 23626
rect 43542 23594 43602 23626
rect 43660 23594 43720 23626
rect 43778 23594 43838 23626
rect 46393 23621 46409 23655
rect 46443 23621 46459 23655
rect 46393 23605 46459 23621
rect 46511 23655 46577 23671
rect 46511 23621 46527 23655
rect 46561 23621 46577 23655
rect 46511 23605 46577 23621
rect 54928 24038 55079 24091
rect 53283 23862 53343 23888
rect 54928 23814 54988 24038
rect 55372 23996 55432 24197
rect 55490 24171 55550 24197
rect 55608 24171 55668 24197
rect 56160 24184 56220 24201
rect 56160 24095 56221 24184
rect 56278 24175 56338 24201
rect 56396 24175 56456 24201
rect 55046 23945 55432 23996
rect 56070 24042 56221 24095
rect 55046 23814 55106 23945
rect 55161 23887 55227 23903
rect 55161 23853 55177 23887
rect 55211 23853 55227 23887
rect 55161 23837 55227 23853
rect 55164 23814 55224 23837
rect 55447 23814 55507 23840
rect 55565 23814 55625 23840
rect 55683 23814 55743 23840
rect 56070 23818 56130 24042
rect 56514 24000 56574 24201
rect 56632 24175 56692 24201
rect 56750 24175 56810 24201
rect 59488 24118 59546 24303
rect 59488 24092 59548 24118
rect 59606 24092 59666 24303
rect 59959 24297 60019 24329
rect 60077 24303 60137 24329
rect 60195 24303 60255 24329
rect 59956 24281 60022 24297
rect 59956 24247 59972 24281
rect 60006 24247 60022 24281
rect 59956 24231 60022 24247
rect 61576 24184 61636 24201
rect 59838 24164 59904 24180
rect 59838 24130 59854 24164
rect 59888 24130 59904 24164
rect 59838 24114 59904 24130
rect 59841 24092 59901 24114
rect 61576 24095 61637 24184
rect 61694 24175 61754 24201
rect 61812 24175 61872 24201
rect 56188 23949 56574 24000
rect 56188 23818 56248 23949
rect 56303 23891 56369 23907
rect 56303 23857 56319 23891
rect 56353 23857 56369 23891
rect 56303 23841 56369 23857
rect 56306 23818 56366 23841
rect 56589 23818 56649 23844
rect 56707 23818 56767 23844
rect 56825 23818 56885 23844
rect 52930 23666 52990 23688
rect 53048 23666 53108 23688
rect 52927 23650 52993 23666
rect 43259 23553 43838 23594
rect 48394 23593 48454 23619
rect 48512 23593 48572 23619
rect 48630 23587 48690 23619
rect 48913 23587 48973 23619
rect 49031 23587 49091 23619
rect 49149 23587 49209 23619
rect 49536 23597 49596 23623
rect 49654 23597 49714 23623
rect 48630 23546 49209 23587
rect 49772 23591 49832 23623
rect 50055 23591 50115 23623
rect 50173 23591 50233 23623
rect 50291 23591 50351 23623
rect 52927 23616 52943 23650
rect 52977 23616 52993 23650
rect 52927 23600 52993 23616
rect 53045 23650 53111 23666
rect 53045 23616 53061 23650
rect 53095 23616 53111 23650
rect 53045 23600 53111 23616
rect 61486 24042 61637 24095
rect 59841 23866 59901 23892
rect 61486 23818 61546 24042
rect 61930 24000 61990 24201
rect 62048 24175 62108 24201
rect 62166 24175 62226 24201
rect 62718 24188 62778 24205
rect 62718 24099 62779 24188
rect 62836 24179 62896 24205
rect 62954 24179 63014 24205
rect 61604 23949 61990 24000
rect 62628 24046 62779 24099
rect 61604 23818 61664 23949
rect 61719 23891 61785 23907
rect 61719 23857 61735 23891
rect 61769 23857 61785 23891
rect 61719 23841 61785 23857
rect 61722 23818 61782 23841
rect 62005 23818 62065 23844
rect 62123 23818 62183 23844
rect 62241 23818 62301 23844
rect 62628 23822 62688 24046
rect 63072 24004 63132 24205
rect 63190 24179 63250 24205
rect 63308 24179 63368 24205
rect 62746 23953 63132 24004
rect 62746 23822 62806 23953
rect 62861 23895 62927 23911
rect 62861 23861 62877 23895
rect 62911 23861 62927 23895
rect 62861 23845 62927 23861
rect 62864 23822 62924 23845
rect 63147 23822 63207 23848
rect 63265 23822 63325 23848
rect 63383 23822 63443 23848
rect 59488 23670 59548 23692
rect 59606 23670 59666 23692
rect 59485 23654 59551 23670
rect 59485 23620 59501 23654
rect 59535 23620 59551 23654
rect 49772 23550 50351 23591
rect 54928 23588 54988 23614
rect 55046 23588 55106 23614
rect 55164 23582 55224 23614
rect 55447 23582 55507 23614
rect 55565 23582 55625 23614
rect 55683 23582 55743 23614
rect 56070 23592 56130 23618
rect 56188 23592 56248 23618
rect 55164 23541 55743 23582
rect 56306 23586 56366 23618
rect 56589 23586 56649 23618
rect 56707 23586 56767 23618
rect 56825 23586 56885 23618
rect 59485 23604 59551 23620
rect 59603 23654 59669 23670
rect 59603 23620 59619 23654
rect 59653 23620 59669 23654
rect 59603 23604 59669 23620
rect 61486 23592 61546 23618
rect 61604 23592 61664 23618
rect 56306 23545 56885 23586
rect 61722 23586 61782 23618
rect 62005 23586 62065 23618
rect 62123 23586 62183 23618
rect 62241 23586 62301 23618
rect 62628 23596 62688 23622
rect 62746 23596 62806 23622
rect 61722 23545 62301 23586
rect 62864 23590 62924 23622
rect 63147 23590 63207 23622
rect 63265 23590 63325 23622
rect 63383 23590 63443 23622
rect 62864 23549 63443 23590
rect 39660 22904 39956 22940
rect 39660 22883 39720 22904
rect 39778 22883 39838 22904
rect 39896 22883 39956 22904
rect 40014 22903 40310 22939
rect 40014 22883 40074 22903
rect 40132 22883 40192 22903
rect 40250 22883 40310 22903
rect 40368 22903 40664 22939
rect 40368 22883 40428 22903
rect 40486 22883 40546 22903
rect 40604 22883 40664 22903
rect 46173 22901 46469 22937
rect 46173 22880 46233 22901
rect 46291 22880 46351 22901
rect 46409 22880 46469 22901
rect 46527 22900 46823 22936
rect 46527 22880 46587 22900
rect 46645 22880 46705 22900
rect 46763 22880 46823 22900
rect 46881 22900 47177 22936
rect 46881 22880 46941 22900
rect 46999 22880 47059 22900
rect 47117 22880 47177 22900
rect 39660 22657 39720 22683
rect 39778 22657 39838 22683
rect 39896 22657 39956 22683
rect 40014 22663 40074 22683
rect 40014 22657 40075 22663
rect 40132 22657 40192 22683
rect 40250 22657 40310 22683
rect 39897 22472 39955 22657
rect 39897 22446 39957 22472
rect 40015 22446 40075 22657
rect 40368 22651 40428 22683
rect 40486 22657 40546 22683
rect 40604 22657 40664 22683
rect 52707 22896 53003 22932
rect 52707 22875 52767 22896
rect 52825 22875 52885 22896
rect 52943 22875 53003 22896
rect 53061 22895 53357 22931
rect 53061 22875 53121 22895
rect 53179 22875 53239 22895
rect 53297 22875 53357 22895
rect 53415 22895 53711 22931
rect 53415 22875 53475 22895
rect 53533 22875 53593 22895
rect 53651 22875 53711 22895
rect 46173 22654 46233 22680
rect 46291 22654 46351 22680
rect 46409 22654 46469 22680
rect 46527 22660 46587 22680
rect 46527 22654 46588 22660
rect 46645 22654 46705 22680
rect 46763 22654 46823 22680
rect 40365 22635 40431 22651
rect 40365 22601 40381 22635
rect 40415 22601 40431 22635
rect 40365 22585 40431 22601
rect 40247 22518 40313 22534
rect 40247 22484 40263 22518
rect 40297 22484 40313 22518
rect 40247 22468 40313 22484
rect 41608 22481 41904 22532
rect 40250 22446 40310 22468
rect 41608 22466 41668 22481
rect 41726 22466 41786 22481
rect 41844 22466 41904 22481
rect 41962 22466 42022 22492
rect 42080 22466 42140 22492
rect 42198 22466 42258 22492
rect 43506 22481 43802 22532
rect 43506 22466 43566 22481
rect 43624 22466 43684 22481
rect 43742 22466 43802 22481
rect 43860 22466 43920 22492
rect 43978 22466 44038 22492
rect 44096 22466 44156 22492
rect 46410 22469 46468 22654
rect 3531 22011 3827 22050
rect 3531 21996 3591 22011
rect 3649 21996 3709 22011
rect 3767 21996 3827 22011
rect 4004 22011 4300 22050
rect 4004 21996 4064 22011
rect 4122 21996 4182 22011
rect 4240 21996 4300 22011
rect 4358 22011 4654 22050
rect 4358 21996 4418 22011
rect 4476 21996 4536 22011
rect 4594 21996 4654 22011
rect 4825 22011 5121 22050
rect 4825 21996 4885 22011
rect 4943 21996 5003 22011
rect 5061 21996 5121 22011
rect 6675 22011 6971 22050
rect 6675 21996 6735 22011
rect 6793 21996 6853 22011
rect 6911 21996 6971 22011
rect 7148 22011 7444 22050
rect 7148 21996 7208 22011
rect 7266 21996 7326 22011
rect 7384 21996 7444 22011
rect 7502 22011 7798 22050
rect 7502 21996 7562 22011
rect 7620 21996 7680 22011
rect 7738 21996 7798 22011
rect 7969 22011 8265 22050
rect 7969 21996 8029 22011
rect 8087 21996 8147 22011
rect 8205 21996 8265 22011
rect 9807 22007 10103 22046
rect 3058 21812 3354 21851
rect 3058 21796 3118 21812
rect 3176 21796 3236 21812
rect 3294 21796 3354 21812
rect 5266 21812 5562 21851
rect 5266 21796 5326 21812
rect 5384 21796 5444 21812
rect 5502 21796 5562 21812
rect 6202 21812 6498 21851
rect 6202 21796 6262 21812
rect 6320 21796 6380 21812
rect 6438 21796 6498 21812
rect 9807 21992 9867 22007
rect 9925 21992 9985 22007
rect 10043 21992 10103 22007
rect 10280 22007 10576 22046
rect 10280 21992 10340 22007
rect 10398 21992 10458 22007
rect 10516 21992 10576 22007
rect 10634 22007 10930 22046
rect 10634 21992 10694 22007
rect 10752 21992 10812 22007
rect 10870 21992 10930 22007
rect 11101 22007 11397 22046
rect 11101 21992 11161 22007
rect 11219 21992 11279 22007
rect 11337 21992 11397 22007
rect 12951 22007 13247 22046
rect 12951 21992 13011 22007
rect 13069 21992 13129 22007
rect 13187 21992 13247 22007
rect 13424 22007 13720 22046
rect 13424 21992 13484 22007
rect 13542 21992 13602 22007
rect 13660 21992 13720 22007
rect 13778 22007 14074 22046
rect 13778 21992 13838 22007
rect 13896 21992 13956 22007
rect 14014 21992 14074 22007
rect 14245 22007 14541 22046
rect 14245 21992 14305 22007
rect 14363 21992 14423 22007
rect 14481 21992 14541 22007
rect 16153 22011 16449 22050
rect 16153 21996 16213 22011
rect 16271 21996 16331 22011
rect 16389 21996 16449 22011
rect 16626 22011 16922 22050
rect 16626 21996 16686 22011
rect 16744 21996 16804 22011
rect 16862 21996 16922 22011
rect 16980 22011 17276 22050
rect 16980 21996 17040 22011
rect 17098 21996 17158 22011
rect 17216 21996 17276 22011
rect 17447 22011 17743 22050
rect 17447 21996 17507 22011
rect 17565 21996 17625 22011
rect 17683 21996 17743 22011
rect 19297 22011 19593 22050
rect 19297 21996 19357 22011
rect 19415 21996 19475 22011
rect 19533 21996 19593 22011
rect 19770 22011 20066 22050
rect 19770 21996 19830 22011
rect 19888 21996 19948 22011
rect 20006 21996 20066 22011
rect 20124 22011 20420 22050
rect 20124 21996 20184 22011
rect 20242 21996 20302 22011
rect 20360 21996 20420 22011
rect 20591 22011 20887 22050
rect 41124 22266 41184 22292
rect 41242 22266 41302 22292
rect 41360 22266 41420 22292
rect 40250 22220 40310 22246
rect 20591 21996 20651 22011
rect 20709 21996 20769 22011
rect 20827 21996 20887 22011
rect 22429 22007 22725 22046
rect 8410 21812 8706 21851
rect 8410 21796 8470 21812
rect 8528 21796 8588 21812
rect 8646 21796 8706 21812
rect 9334 21808 9630 21847
rect 9334 21792 9394 21808
rect 9452 21792 9512 21808
rect 9570 21792 9630 21808
rect 3058 21447 3118 21596
rect 3176 21570 3236 21596
rect 3294 21570 3354 21596
rect 3531 21570 3591 21596
rect 3162 21447 3228 21450
rect 3058 21434 3228 21447
rect 3058 21400 3178 21434
rect 3212 21400 3228 21434
rect 3058 21387 3228 21400
rect 3058 20911 3118 21387
rect 3162 21384 3228 21387
rect 3649 21180 3709 21596
rect 3767 21570 3827 21596
rect 4004 21570 4064 21596
rect 4122 21271 4182 21596
rect 4240 21570 4300 21596
rect 4358 21570 4418 21596
rect 4476 21570 4536 21596
rect 4594 21570 4654 21596
rect 4825 21570 4885 21596
rect 4476 21410 4535 21570
rect 4472 21409 4535 21410
rect 4472 21393 4538 21409
rect 4472 21359 4488 21393
rect 4522 21359 4538 21393
rect 4472 21343 4538 21359
rect 4340 21294 4435 21309
rect 4340 21271 4358 21294
rect 4122 21239 4358 21271
rect 4416 21239 4435 21294
rect 4122 21222 4435 21239
rect 3649 21163 4187 21180
rect 3649 21129 4134 21163
rect 4168 21129 4187 21163
rect 3649 21123 4187 21129
rect 4118 21113 4187 21123
rect 4122 21111 4187 21113
rect 3058 20866 3986 20911
rect 3926 20663 3986 20866
rect 4122 20663 4182 21111
rect 4237 20773 4303 20789
rect 4237 20739 4253 20773
rect 4287 20739 4303 20773
rect 4237 20723 4303 20739
rect 4240 20663 4300 20723
rect 4358 20663 4418 21222
rect 4943 21178 5003 21596
rect 5061 21570 5121 21596
rect 5266 21570 5326 21596
rect 5384 21570 5444 21596
rect 5502 21310 5562 21596
rect 5426 21293 5562 21310
rect 5426 21238 5445 21293
rect 5503 21238 5562 21293
rect 5426 21223 5562 21238
rect 4476 21121 5003 21178
rect 4476 21022 4536 21121
rect 4466 21009 4547 21022
rect 4466 20954 4476 21009
rect 4534 20954 4547 21009
rect 4466 20943 4547 20954
rect 4476 20663 4536 20943
rect 5502 20911 5562 21223
rect 4668 20866 5562 20911
rect 6202 21447 6262 21596
rect 6320 21570 6380 21596
rect 6438 21570 6498 21596
rect 6675 21570 6735 21596
rect 6306 21447 6372 21450
rect 6202 21434 6372 21447
rect 6202 21400 6322 21434
rect 6356 21400 6372 21434
rect 6202 21387 6372 21400
rect 6202 20911 6262 21387
rect 6306 21384 6372 21387
rect 6793 21180 6853 21596
rect 6911 21570 6971 21596
rect 7148 21570 7208 21596
rect 7266 21271 7326 21596
rect 7384 21570 7444 21596
rect 7502 21570 7562 21596
rect 7620 21570 7680 21596
rect 7738 21570 7798 21596
rect 7969 21570 8029 21596
rect 7620 21410 7679 21570
rect 7616 21409 7679 21410
rect 7616 21393 7682 21409
rect 7616 21359 7632 21393
rect 7666 21359 7682 21393
rect 7616 21343 7682 21359
rect 7484 21294 7579 21309
rect 7484 21271 7502 21294
rect 7266 21239 7502 21271
rect 7560 21239 7579 21294
rect 7266 21222 7579 21239
rect 6793 21163 7331 21180
rect 6793 21129 7278 21163
rect 7312 21129 7331 21163
rect 6793 21123 7331 21129
rect 7262 21113 7331 21123
rect 7266 21111 7331 21113
rect 6202 20866 7130 20911
rect 4668 20663 4728 20866
rect 7070 20663 7130 20866
rect 7266 20663 7326 21111
rect 7381 20773 7447 20789
rect 7381 20739 7397 20773
rect 7431 20739 7447 20773
rect 7381 20723 7447 20739
rect 7384 20663 7444 20723
rect 7502 20663 7562 21222
rect 8087 21178 8147 21596
rect 8205 21570 8265 21596
rect 8410 21570 8470 21596
rect 8528 21570 8588 21596
rect 8646 21310 8706 21596
rect 11542 21808 11838 21847
rect 11542 21792 11602 21808
rect 11660 21792 11720 21808
rect 11778 21792 11838 21808
rect 12478 21808 12774 21847
rect 12478 21792 12538 21808
rect 12596 21792 12656 21808
rect 12714 21792 12774 21808
rect 14686 21808 14982 21847
rect 14686 21792 14746 21808
rect 14804 21792 14864 21808
rect 14922 21792 14982 21808
rect 15680 21812 15976 21851
rect 15680 21796 15740 21812
rect 15798 21796 15858 21812
rect 15916 21796 15976 21812
rect 17888 21812 18184 21851
rect 17888 21796 17948 21812
rect 18006 21796 18066 21812
rect 18124 21796 18184 21812
rect 18824 21812 19120 21851
rect 18824 21796 18884 21812
rect 18942 21796 19002 21812
rect 19060 21796 19120 21812
rect 22429 21992 22489 22007
rect 22547 21992 22607 22007
rect 22665 21992 22725 22007
rect 22902 22007 23198 22046
rect 22902 21992 22962 22007
rect 23020 21992 23080 22007
rect 23138 21992 23198 22007
rect 23256 22007 23552 22046
rect 23256 21992 23316 22007
rect 23374 21992 23434 22007
rect 23492 21992 23552 22007
rect 23723 22007 24019 22046
rect 23723 21992 23783 22007
rect 23841 21992 23901 22007
rect 23959 21992 24019 22007
rect 25573 22007 25869 22046
rect 25573 21992 25633 22007
rect 25691 21992 25751 22007
rect 25809 21992 25869 22007
rect 26046 22007 26342 22046
rect 26046 21992 26106 22007
rect 26164 21992 26224 22007
rect 26282 21992 26342 22007
rect 26400 22007 26696 22046
rect 26400 21992 26460 22007
rect 26518 21992 26578 22007
rect 26636 21992 26696 22007
rect 26867 22007 27163 22046
rect 39897 22024 39957 22046
rect 40015 22030 40075 22046
rect 26867 21992 26927 22007
rect 26985 21992 27045 22007
rect 27103 21992 27163 22007
rect 39894 22008 39960 22024
rect 21032 21812 21328 21851
rect 21032 21796 21092 21812
rect 21150 21796 21210 21812
rect 21268 21796 21328 21812
rect 21956 21808 22252 21847
rect 21956 21792 22016 21808
rect 22074 21792 22134 21808
rect 22192 21792 22252 21808
rect 8570 21293 8706 21310
rect 8570 21238 8589 21293
rect 8647 21238 8706 21293
rect 8570 21223 8706 21238
rect 7620 21121 8147 21178
rect 7620 21022 7680 21121
rect 7610 21009 7691 21022
rect 7610 20954 7620 21009
rect 7678 20954 7691 21009
rect 7610 20943 7691 20954
rect 7620 20663 7680 20943
rect 8646 20911 8706 21223
rect 7812 20866 8706 20911
rect 9334 21443 9394 21592
rect 9452 21566 9512 21592
rect 9570 21566 9630 21592
rect 9807 21566 9867 21592
rect 9438 21443 9504 21446
rect 9334 21430 9504 21443
rect 9334 21396 9454 21430
rect 9488 21396 9504 21430
rect 9334 21383 9504 21396
rect 9334 20907 9394 21383
rect 9438 21380 9504 21383
rect 9925 21176 9985 21592
rect 10043 21566 10103 21592
rect 10280 21566 10340 21592
rect 10398 21267 10458 21592
rect 10516 21566 10576 21592
rect 10634 21566 10694 21592
rect 10752 21566 10812 21592
rect 10870 21566 10930 21592
rect 11101 21566 11161 21592
rect 10752 21406 10811 21566
rect 10748 21405 10811 21406
rect 10748 21389 10814 21405
rect 10748 21355 10764 21389
rect 10798 21355 10814 21389
rect 10748 21339 10814 21355
rect 10616 21290 10711 21305
rect 10616 21267 10634 21290
rect 10398 21235 10634 21267
rect 10692 21235 10711 21290
rect 10398 21218 10711 21235
rect 9925 21159 10463 21176
rect 9925 21125 10410 21159
rect 10444 21125 10463 21159
rect 9925 21119 10463 21125
rect 10394 21109 10463 21119
rect 10398 21107 10463 21109
rect 7812 20663 7872 20866
rect 9334 20862 10262 20907
rect 3926 20182 3986 20463
rect 4668 20437 4728 20463
rect 4122 20237 4182 20263
rect 4240 20237 4300 20263
rect 4358 20237 4418 20263
rect 4476 20237 4536 20263
rect 4295 20182 4361 20190
rect 3926 20174 4361 20182
rect 3926 20140 4311 20174
rect 4345 20140 4361 20174
rect 3926 20131 4361 20140
rect 7070 20182 7130 20463
rect 10202 20659 10262 20862
rect 10398 20659 10458 21107
rect 10513 20769 10579 20785
rect 10513 20735 10529 20769
rect 10563 20735 10579 20769
rect 10513 20719 10579 20735
rect 10516 20659 10576 20719
rect 10634 20659 10694 21218
rect 11219 21174 11279 21592
rect 11337 21566 11397 21592
rect 11542 21566 11602 21592
rect 11660 21566 11720 21592
rect 11778 21306 11838 21592
rect 11702 21289 11838 21306
rect 11702 21234 11721 21289
rect 11779 21234 11838 21289
rect 11702 21219 11838 21234
rect 10752 21117 11279 21174
rect 10752 21018 10812 21117
rect 10742 21005 10823 21018
rect 10742 20950 10752 21005
rect 10810 20950 10823 21005
rect 10742 20939 10823 20950
rect 10752 20659 10812 20939
rect 11778 20907 11838 21219
rect 10944 20862 11838 20907
rect 12478 21443 12538 21592
rect 12596 21566 12656 21592
rect 12714 21566 12774 21592
rect 12951 21566 13011 21592
rect 12582 21443 12648 21446
rect 12478 21430 12648 21443
rect 12478 21396 12598 21430
rect 12632 21396 12648 21430
rect 12478 21383 12648 21396
rect 12478 20907 12538 21383
rect 12582 21380 12648 21383
rect 13069 21176 13129 21592
rect 13187 21566 13247 21592
rect 13424 21566 13484 21592
rect 13542 21267 13602 21592
rect 13660 21566 13720 21592
rect 13778 21566 13838 21592
rect 13896 21566 13956 21592
rect 14014 21566 14074 21592
rect 14245 21566 14305 21592
rect 13896 21406 13955 21566
rect 13892 21405 13955 21406
rect 13892 21389 13958 21405
rect 13892 21355 13908 21389
rect 13942 21355 13958 21389
rect 13892 21339 13958 21355
rect 13760 21290 13855 21305
rect 13760 21267 13778 21290
rect 13542 21235 13778 21267
rect 13836 21235 13855 21290
rect 13542 21218 13855 21235
rect 13069 21159 13607 21176
rect 13069 21125 13554 21159
rect 13588 21125 13607 21159
rect 13069 21119 13607 21125
rect 13538 21109 13607 21119
rect 13542 21107 13607 21109
rect 12478 20862 13406 20907
rect 10944 20659 11004 20862
rect 13346 20659 13406 20862
rect 13542 20659 13602 21107
rect 13657 20769 13723 20785
rect 13657 20735 13673 20769
rect 13707 20735 13723 20769
rect 13657 20719 13723 20735
rect 13660 20659 13720 20719
rect 13778 20659 13838 21218
rect 14363 21174 14423 21592
rect 14481 21566 14541 21592
rect 14686 21566 14746 21592
rect 14804 21566 14864 21592
rect 14922 21306 14982 21592
rect 14846 21289 14982 21306
rect 14846 21234 14865 21289
rect 14923 21234 14982 21289
rect 14846 21219 14982 21234
rect 13896 21117 14423 21174
rect 13896 21018 13956 21117
rect 13886 21005 13967 21018
rect 13886 20950 13896 21005
rect 13954 20950 13967 21005
rect 13886 20939 13967 20950
rect 13896 20659 13956 20939
rect 14922 20907 14982 21219
rect 14088 20862 14982 20907
rect 15680 21447 15740 21596
rect 15798 21570 15858 21596
rect 15916 21570 15976 21596
rect 16153 21570 16213 21596
rect 15784 21447 15850 21450
rect 15680 21434 15850 21447
rect 15680 21400 15800 21434
rect 15834 21400 15850 21434
rect 15680 21387 15850 21400
rect 15680 20911 15740 21387
rect 15784 21384 15850 21387
rect 16271 21180 16331 21596
rect 16389 21570 16449 21596
rect 16626 21570 16686 21596
rect 16744 21271 16804 21596
rect 16862 21570 16922 21596
rect 16980 21570 17040 21596
rect 17098 21570 17158 21596
rect 17216 21570 17276 21596
rect 17447 21570 17507 21596
rect 17098 21410 17157 21570
rect 17094 21409 17157 21410
rect 17094 21393 17160 21409
rect 17094 21359 17110 21393
rect 17144 21359 17160 21393
rect 17094 21343 17160 21359
rect 16962 21294 17057 21309
rect 16962 21271 16980 21294
rect 16744 21239 16980 21271
rect 17038 21239 17057 21294
rect 16744 21222 17057 21239
rect 16271 21163 16809 21180
rect 16271 21129 16756 21163
rect 16790 21129 16809 21163
rect 16271 21123 16809 21129
rect 16740 21113 16809 21123
rect 16744 21111 16809 21113
rect 15680 20866 16608 20911
rect 14088 20659 14148 20862
rect 16548 20663 16608 20866
rect 16744 20663 16804 21111
rect 16859 20773 16925 20789
rect 16859 20739 16875 20773
rect 16909 20739 16925 20773
rect 16859 20723 16925 20739
rect 16862 20663 16922 20723
rect 16980 20663 17040 21222
rect 17565 21178 17625 21596
rect 17683 21570 17743 21596
rect 17888 21570 17948 21596
rect 18006 21570 18066 21596
rect 18124 21310 18184 21596
rect 18048 21293 18184 21310
rect 18048 21238 18067 21293
rect 18125 21238 18184 21293
rect 18048 21223 18184 21238
rect 17098 21121 17625 21178
rect 17098 21022 17158 21121
rect 17088 21009 17169 21022
rect 17088 20954 17098 21009
rect 17156 20954 17169 21009
rect 17088 20943 17169 20954
rect 17098 20663 17158 20943
rect 18124 20911 18184 21223
rect 17290 20866 18184 20911
rect 18824 21447 18884 21596
rect 18942 21570 19002 21596
rect 19060 21570 19120 21596
rect 19297 21570 19357 21596
rect 18928 21447 18994 21450
rect 18824 21434 18994 21447
rect 18824 21400 18944 21434
rect 18978 21400 18994 21434
rect 18824 21387 18994 21400
rect 18824 20911 18884 21387
rect 18928 21384 18994 21387
rect 19415 21180 19475 21596
rect 19533 21570 19593 21596
rect 19770 21570 19830 21596
rect 19888 21271 19948 21596
rect 20006 21570 20066 21596
rect 20124 21570 20184 21596
rect 20242 21570 20302 21596
rect 20360 21570 20420 21596
rect 20591 21570 20651 21596
rect 20242 21410 20301 21570
rect 20238 21409 20301 21410
rect 20238 21393 20304 21409
rect 20238 21359 20254 21393
rect 20288 21359 20304 21393
rect 20238 21343 20304 21359
rect 20106 21294 20201 21309
rect 20106 21271 20124 21294
rect 19888 21239 20124 21271
rect 20182 21239 20201 21294
rect 19888 21222 20201 21239
rect 19415 21163 19953 21180
rect 19415 21129 19900 21163
rect 19934 21129 19953 21163
rect 19415 21123 19953 21129
rect 19884 21113 19953 21123
rect 19888 21111 19953 21113
rect 18824 20866 19752 20911
rect 17290 20663 17350 20866
rect 19692 20663 19752 20866
rect 19888 20663 19948 21111
rect 20003 20773 20069 20789
rect 20003 20739 20019 20773
rect 20053 20739 20069 20773
rect 20003 20723 20069 20739
rect 20006 20663 20066 20723
rect 20124 20663 20184 21222
rect 20709 21178 20769 21596
rect 20827 21570 20887 21596
rect 21032 21570 21092 21596
rect 21150 21570 21210 21596
rect 21268 21310 21328 21596
rect 24164 21808 24460 21847
rect 24164 21792 24224 21808
rect 24282 21792 24342 21808
rect 24400 21792 24460 21808
rect 25100 21808 25396 21847
rect 25100 21792 25160 21808
rect 25218 21792 25278 21808
rect 25336 21792 25396 21808
rect 39894 21974 39910 22008
rect 39944 21974 39960 22008
rect 39894 21958 39960 21974
rect 40009 22008 40083 22030
rect 40009 21974 40028 22008
rect 40062 21974 40083 22008
rect 42445 22283 42741 22334
rect 42445 22266 42505 22283
rect 42563 22266 42623 22283
rect 42681 22266 42741 22283
rect 43022 22266 43082 22292
rect 43140 22266 43200 22292
rect 43258 22266 43318 22292
rect 46410 22443 46470 22469
rect 46528 22443 46588 22654
rect 46881 22648 46941 22680
rect 46999 22654 47059 22680
rect 47117 22654 47177 22680
rect 59265 22900 59561 22936
rect 59265 22879 59325 22900
rect 59383 22879 59443 22900
rect 59501 22879 59561 22900
rect 59619 22899 59915 22935
rect 59619 22879 59679 22899
rect 59737 22879 59797 22899
rect 59855 22879 59915 22899
rect 59973 22899 60269 22935
rect 59973 22879 60033 22899
rect 60091 22879 60151 22899
rect 60209 22879 60269 22899
rect 52707 22649 52767 22675
rect 52825 22649 52885 22675
rect 52943 22649 53003 22675
rect 53061 22655 53121 22675
rect 53061 22649 53122 22655
rect 53179 22649 53239 22675
rect 53297 22649 53357 22675
rect 46878 22632 46944 22648
rect 46878 22598 46894 22632
rect 46928 22598 46944 22632
rect 46878 22582 46944 22598
rect 46760 22515 46826 22531
rect 46760 22481 46776 22515
rect 46810 22481 46826 22515
rect 46760 22465 46826 22481
rect 48121 22478 48417 22529
rect 46763 22443 46823 22465
rect 48121 22463 48181 22478
rect 48239 22463 48299 22478
rect 48357 22463 48417 22478
rect 48475 22463 48535 22489
rect 48593 22463 48653 22489
rect 48711 22463 48771 22489
rect 50019 22478 50315 22529
rect 50019 22463 50079 22478
rect 50137 22463 50197 22478
rect 50255 22463 50315 22478
rect 50373 22463 50433 22489
rect 50491 22463 50551 22489
rect 50609 22463 50669 22489
rect 52944 22464 53002 22649
rect 44343 22283 44639 22334
rect 44343 22266 44403 22283
rect 44461 22266 44521 22283
rect 44579 22266 44639 22283
rect 41124 22049 41184 22066
rect 41242 22049 41302 22066
rect 41360 22049 41420 22066
rect 41608 22049 41668 22066
rect 41124 21998 41668 22049
rect 41726 22040 41786 22066
rect 41844 22040 41904 22066
rect 41962 22047 42022 22066
rect 42080 22047 42140 22066
rect 42198 22047 42258 22066
rect 42445 22047 42505 22066
rect 42563 22047 42623 22066
rect 40009 21917 40083 21974
rect 41249 21917 41309 21998
rect 41962 21996 42505 22047
rect 42547 22040 42623 22047
rect 42681 22040 42741 22066
rect 43022 22049 43082 22066
rect 43140 22049 43200 22066
rect 43258 22049 43318 22066
rect 43506 22049 43566 22066
rect 42547 21996 42622 22040
rect 43022 21998 43566 22049
rect 43624 22040 43684 22066
rect 43742 22040 43802 22066
rect 43860 22047 43920 22066
rect 43978 22047 44038 22066
rect 44096 22047 44156 22066
rect 44343 22047 44403 22066
rect 44461 22047 44521 22066
rect 40009 21892 41309 21917
rect 27308 21808 27604 21847
rect 40008 21844 41309 21892
rect 42547 21876 42607 21996
rect 27308 21792 27368 21808
rect 27426 21792 27486 21808
rect 27544 21792 27604 21808
rect 21192 21293 21328 21310
rect 21192 21238 21211 21293
rect 21269 21238 21328 21293
rect 21192 21223 21328 21238
rect 20242 21121 20769 21178
rect 20242 21022 20302 21121
rect 20232 21009 20313 21022
rect 20232 20954 20242 21009
rect 20300 20954 20313 21009
rect 20232 20943 20313 20954
rect 20242 20663 20302 20943
rect 21268 20911 21328 21223
rect 20434 20866 21328 20911
rect 21956 21443 22016 21592
rect 22074 21566 22134 21592
rect 22192 21566 22252 21592
rect 22429 21566 22489 21592
rect 22060 21443 22126 21446
rect 21956 21430 22126 21443
rect 21956 21396 22076 21430
rect 22110 21396 22126 21430
rect 21956 21383 22126 21396
rect 21956 20907 22016 21383
rect 22060 21380 22126 21383
rect 22547 21176 22607 21592
rect 22665 21566 22725 21592
rect 22902 21566 22962 21592
rect 23020 21267 23080 21592
rect 23138 21566 23198 21592
rect 23256 21566 23316 21592
rect 23374 21566 23434 21592
rect 23492 21566 23552 21592
rect 23723 21566 23783 21592
rect 23374 21406 23433 21566
rect 23370 21405 23433 21406
rect 23370 21389 23436 21405
rect 23370 21355 23386 21389
rect 23420 21355 23436 21389
rect 23370 21339 23436 21355
rect 23238 21290 23333 21305
rect 23238 21267 23256 21290
rect 23020 21235 23256 21267
rect 23314 21235 23333 21290
rect 23020 21218 23333 21235
rect 22547 21159 23085 21176
rect 22547 21125 23032 21159
rect 23066 21125 23085 21159
rect 22547 21119 23085 21125
rect 23016 21109 23085 21119
rect 23020 21107 23085 21109
rect 20434 20663 20494 20866
rect 21956 20862 22884 20907
rect 7812 20437 7872 20463
rect 7266 20237 7326 20263
rect 7384 20237 7444 20263
rect 7502 20237 7562 20263
rect 7620 20237 7680 20263
rect 7439 20182 7505 20190
rect 7070 20174 7505 20182
rect 7070 20140 7455 20174
rect 7489 20140 7505 20174
rect 7070 20131 7505 20140
rect 4295 20124 4361 20131
rect 7439 20124 7505 20131
rect 10202 20178 10262 20459
rect 10944 20433 11004 20459
rect 10398 20233 10458 20259
rect 10516 20233 10576 20259
rect 10634 20233 10694 20259
rect 10752 20233 10812 20259
rect 10571 20178 10637 20186
rect 10202 20170 10637 20178
rect 10202 20136 10587 20170
rect 10621 20136 10637 20170
rect 10202 20127 10637 20136
rect 13346 20178 13406 20459
rect 14088 20433 14148 20459
rect 13542 20233 13602 20259
rect 13660 20233 13720 20259
rect 13778 20233 13838 20259
rect 13896 20233 13956 20259
rect 13715 20178 13781 20186
rect 13346 20170 13781 20178
rect 13346 20136 13731 20170
rect 13765 20136 13781 20170
rect 13346 20127 13781 20136
rect 16548 20182 16608 20463
rect 17290 20437 17350 20463
rect 16744 20237 16804 20263
rect 16862 20237 16922 20263
rect 16980 20237 17040 20263
rect 17098 20237 17158 20263
rect 16917 20182 16983 20190
rect 16548 20174 16983 20182
rect 16548 20140 16933 20174
rect 16967 20140 16983 20174
rect 16548 20131 16983 20140
rect 19692 20182 19752 20463
rect 22824 20659 22884 20862
rect 23020 20659 23080 21107
rect 23135 20769 23201 20785
rect 23135 20735 23151 20769
rect 23185 20735 23201 20769
rect 23135 20719 23201 20735
rect 23138 20659 23198 20719
rect 23256 20659 23316 21218
rect 23841 21174 23901 21592
rect 23959 21566 24019 21592
rect 24164 21566 24224 21592
rect 24282 21566 24342 21592
rect 24400 21306 24460 21592
rect 24324 21289 24460 21306
rect 24324 21234 24343 21289
rect 24401 21234 24460 21289
rect 24324 21219 24460 21234
rect 23374 21117 23901 21174
rect 23374 21018 23434 21117
rect 23364 21005 23445 21018
rect 23364 20950 23374 21005
rect 23432 20950 23445 21005
rect 23364 20939 23445 20950
rect 23374 20659 23434 20939
rect 24400 20907 24460 21219
rect 23566 20862 24460 20907
rect 25100 21443 25160 21592
rect 25218 21566 25278 21592
rect 25336 21566 25396 21592
rect 25573 21566 25633 21592
rect 25204 21443 25270 21446
rect 25100 21430 25270 21443
rect 25100 21396 25220 21430
rect 25254 21396 25270 21430
rect 25100 21383 25270 21396
rect 25100 20907 25160 21383
rect 25204 21380 25270 21383
rect 25691 21176 25751 21592
rect 25809 21566 25869 21592
rect 26046 21566 26106 21592
rect 26164 21267 26224 21592
rect 26282 21566 26342 21592
rect 26400 21566 26460 21592
rect 26518 21566 26578 21592
rect 26636 21566 26696 21592
rect 26867 21566 26927 21592
rect 26518 21406 26577 21566
rect 26514 21405 26577 21406
rect 26514 21389 26580 21405
rect 26514 21355 26530 21389
rect 26564 21355 26580 21389
rect 26514 21339 26580 21355
rect 26382 21290 26477 21305
rect 26382 21267 26400 21290
rect 26164 21235 26400 21267
rect 26458 21235 26477 21290
rect 26164 21218 26477 21235
rect 25691 21159 26229 21176
rect 25691 21125 26176 21159
rect 26210 21125 26229 21159
rect 25691 21119 26229 21125
rect 26160 21109 26229 21119
rect 26164 21107 26229 21109
rect 25100 20862 26028 20907
rect 23566 20659 23626 20862
rect 25968 20659 26028 20862
rect 26164 20659 26224 21107
rect 26279 20769 26345 20785
rect 26279 20735 26295 20769
rect 26329 20735 26345 20769
rect 26279 20719 26345 20735
rect 26282 20659 26342 20719
rect 26400 20659 26460 21218
rect 26985 21174 27045 21592
rect 27103 21566 27163 21592
rect 27308 21566 27368 21592
rect 27426 21566 27486 21592
rect 27544 21306 27604 21592
rect 27468 21289 27604 21306
rect 27468 21234 27487 21289
rect 27545 21234 27604 21289
rect 39655 21300 39951 21336
rect 39655 21279 39715 21300
rect 39773 21279 39833 21300
rect 39891 21279 39951 21300
rect 40009 21299 40305 21335
rect 40009 21279 40069 21299
rect 40127 21279 40187 21299
rect 40245 21279 40305 21299
rect 40363 21299 40659 21335
rect 40363 21279 40423 21299
rect 40481 21279 40541 21299
rect 40599 21279 40659 21299
rect 27468 21219 27604 21234
rect 26518 21117 27045 21174
rect 26518 21018 26578 21117
rect 26508 21005 26589 21018
rect 26508 20950 26518 21005
rect 26576 20950 26589 21005
rect 26508 20939 26589 20950
rect 26518 20659 26578 20939
rect 27544 20907 27604 21219
rect 41249 21146 41309 21844
rect 41551 21796 41847 21856
rect 41551 21773 41611 21796
rect 41669 21773 41729 21796
rect 41787 21773 41847 21796
rect 41905 21797 42201 21857
rect 42546 21856 42607 21876
rect 41905 21773 41965 21797
rect 42023 21773 42083 21797
rect 42141 21773 42201 21797
rect 42527 21840 42607 21856
rect 42527 21806 42542 21840
rect 42576 21806 42607 21840
rect 42527 21790 42607 21806
rect 42546 21767 42607 21790
rect 42547 21621 42607 21767
rect 42546 21448 42607 21621
rect 41551 21347 41611 21373
rect 41519 21206 41586 21213
rect 41669 21206 41729 21373
rect 41787 21347 41847 21373
rect 41905 21347 41965 21373
rect 41519 21197 41729 21206
rect 41519 21163 41535 21197
rect 41569 21163 41729 21197
rect 41519 21147 41729 21163
rect 41249 21130 41400 21146
rect 41249 21096 41350 21130
rect 41384 21096 41400 21130
rect 41249 21080 41400 21096
rect 39655 21053 39715 21079
rect 39773 21053 39833 21079
rect 39891 21053 39951 21079
rect 40009 21059 40069 21079
rect 40009 21053 40070 21059
rect 40127 21053 40187 21079
rect 40245 21053 40305 21079
rect 26710 20862 27604 20907
rect 39892 20868 39950 21053
rect 26710 20659 26770 20862
rect 39892 20842 39952 20868
rect 40010 20842 40070 21053
rect 40363 21047 40423 21079
rect 40481 21053 40541 21079
rect 40599 21053 40659 21079
rect 40360 21031 40426 21047
rect 41249 21041 41309 21080
rect 41669 21041 41729 21147
rect 42023 21206 42083 21373
rect 42141 21347 42201 21373
rect 42166 21206 42233 21213
rect 42023 21197 42233 21206
rect 42023 21163 42183 21197
rect 42217 21163 42233 21197
rect 42023 21147 42233 21163
rect 41785 21113 41851 21129
rect 41785 21079 41801 21113
rect 41835 21079 41851 21113
rect 41785 21063 41851 21079
rect 41903 21114 41969 21129
rect 41903 21080 41919 21114
rect 41953 21080 41969 21114
rect 41903 21064 41969 21080
rect 41787 21041 41847 21063
rect 41905 21041 41965 21064
rect 42023 21041 42083 21147
rect 42547 21145 42607 21448
rect 42457 21129 42607 21145
rect 42457 21095 42473 21129
rect 42507 21095 42607 21129
rect 42457 21079 42607 21095
rect 42547 21041 42607 21079
rect 43147 21340 43207 21998
rect 43860 21996 44403 22047
rect 44445 22040 44521 22047
rect 44579 22040 44639 22066
rect 47637 22263 47697 22289
rect 47755 22263 47815 22289
rect 47873 22263 47933 22289
rect 46763 22217 46823 22243
rect 44445 21996 44520 22040
rect 46410 22021 46470 22043
rect 46528 22027 46588 22043
rect 46407 22005 46473 22021
rect 43449 21796 43745 21856
rect 43449 21773 43509 21796
rect 43567 21773 43627 21796
rect 43685 21773 43745 21796
rect 43803 21797 44099 21857
rect 43803 21773 43863 21797
rect 43921 21773 43981 21797
rect 44039 21773 44099 21797
rect 44445 21843 44505 21996
rect 46407 21971 46423 22005
rect 46457 21971 46473 22005
rect 46407 21955 46473 21971
rect 46522 22005 46596 22027
rect 46522 21971 46541 22005
rect 46575 21971 46596 22005
rect 48958 22280 49254 22331
rect 48958 22263 49018 22280
rect 49076 22263 49136 22280
rect 49194 22263 49254 22280
rect 49535 22263 49595 22289
rect 49653 22263 49713 22289
rect 49771 22263 49831 22289
rect 52944 22438 53004 22464
rect 53062 22438 53122 22649
rect 53415 22643 53475 22675
rect 53533 22649 53593 22675
rect 53651 22649 53711 22675
rect 59265 22653 59325 22679
rect 59383 22653 59443 22679
rect 59501 22653 59561 22679
rect 59619 22659 59679 22679
rect 59619 22653 59680 22659
rect 59737 22653 59797 22679
rect 59855 22653 59915 22679
rect 53412 22627 53478 22643
rect 53412 22593 53428 22627
rect 53462 22593 53478 22627
rect 53412 22577 53478 22593
rect 53294 22510 53360 22526
rect 53294 22476 53310 22510
rect 53344 22476 53360 22510
rect 53294 22460 53360 22476
rect 54655 22473 54951 22524
rect 53297 22438 53357 22460
rect 54655 22458 54715 22473
rect 54773 22458 54833 22473
rect 54891 22458 54951 22473
rect 55009 22458 55069 22484
rect 55127 22458 55187 22484
rect 55245 22458 55305 22484
rect 56553 22473 56849 22524
rect 56553 22458 56613 22473
rect 56671 22458 56731 22473
rect 56789 22458 56849 22473
rect 56907 22458 56967 22484
rect 57025 22458 57085 22484
rect 57143 22458 57203 22484
rect 59502 22468 59560 22653
rect 50856 22280 51152 22331
rect 50856 22263 50916 22280
rect 50974 22263 51034 22280
rect 51092 22263 51152 22280
rect 47637 22046 47697 22063
rect 47755 22046 47815 22063
rect 47873 22046 47933 22063
rect 48121 22046 48181 22063
rect 47637 21995 48181 22046
rect 48239 22037 48299 22063
rect 48357 22037 48417 22063
rect 48475 22044 48535 22063
rect 48593 22044 48653 22063
rect 48711 22044 48771 22063
rect 48958 22044 49018 22063
rect 49076 22044 49136 22063
rect 46522 21914 46596 21971
rect 47762 21914 47822 21995
rect 48475 21993 49018 22044
rect 49060 22037 49136 22044
rect 49194 22037 49254 22063
rect 49535 22046 49595 22063
rect 49653 22046 49713 22063
rect 49771 22046 49831 22063
rect 50019 22046 50079 22063
rect 49060 21993 49135 22037
rect 49535 21995 50079 22046
rect 50137 22037 50197 22063
rect 50255 22037 50315 22063
rect 50373 22044 50433 22063
rect 50491 22044 50551 22063
rect 50609 22044 50669 22063
rect 50856 22044 50916 22063
rect 50974 22044 51034 22063
rect 46522 21889 47822 21914
rect 44445 21819 44699 21843
rect 46521 21841 47822 21889
rect 49060 21873 49120 21993
rect 44445 21785 44649 21819
rect 44683 21785 44699 21819
rect 44445 21769 44699 21785
rect 43449 21347 43509 21373
rect 43147 21324 43214 21340
rect 43147 21290 43163 21324
rect 43197 21290 43214 21324
rect 43147 21274 43214 21290
rect 43147 21146 43207 21274
rect 43417 21206 43484 21213
rect 43567 21206 43627 21373
rect 43685 21347 43745 21373
rect 43803 21347 43863 21373
rect 43417 21197 43627 21206
rect 43417 21163 43433 21197
rect 43467 21163 43627 21197
rect 43417 21147 43627 21163
rect 43147 21130 43298 21146
rect 43147 21096 43248 21130
rect 43282 21096 43298 21130
rect 43147 21080 43298 21096
rect 43147 21041 43207 21080
rect 43567 21041 43627 21147
rect 43921 21206 43981 21373
rect 44039 21347 44099 21373
rect 44062 21207 44129 21214
rect 44056 21206 44129 21207
rect 43921 21198 44129 21206
rect 43921 21164 44079 21198
rect 44113 21164 44129 21198
rect 43921 21148 44129 21164
rect 43921 21147 44118 21148
rect 43683 21113 43749 21129
rect 43683 21079 43699 21113
rect 43733 21079 43749 21113
rect 43683 21063 43749 21079
rect 43801 21114 43867 21129
rect 43801 21080 43817 21114
rect 43851 21080 43867 21114
rect 43801 21064 43867 21080
rect 43685 21041 43745 21063
rect 43803 21041 43863 21064
rect 43921 21041 43981 21147
rect 44445 21145 44505 21769
rect 46168 21297 46464 21333
rect 46168 21276 46228 21297
rect 46286 21276 46346 21297
rect 46404 21276 46464 21297
rect 46522 21296 46818 21332
rect 46522 21276 46582 21296
rect 46640 21276 46700 21296
rect 46758 21276 46818 21296
rect 46876 21296 47172 21332
rect 46876 21276 46936 21296
rect 46994 21276 47054 21296
rect 47112 21276 47172 21296
rect 44355 21129 44505 21145
rect 44355 21095 44371 21129
rect 44405 21095 44505 21129
rect 44355 21079 44505 21095
rect 44445 21041 44505 21079
rect 47762 21143 47822 21841
rect 48064 21793 48360 21853
rect 48064 21770 48124 21793
rect 48182 21770 48242 21793
rect 48300 21770 48360 21793
rect 48418 21794 48714 21854
rect 49059 21853 49120 21873
rect 48418 21770 48478 21794
rect 48536 21770 48596 21794
rect 48654 21770 48714 21794
rect 49040 21837 49120 21853
rect 49040 21803 49055 21837
rect 49089 21803 49120 21837
rect 49040 21787 49120 21803
rect 49059 21764 49120 21787
rect 49060 21618 49120 21764
rect 49059 21445 49120 21618
rect 48064 21344 48124 21370
rect 48032 21203 48099 21210
rect 48182 21203 48242 21370
rect 48300 21344 48360 21370
rect 48418 21344 48478 21370
rect 48032 21194 48242 21203
rect 48032 21160 48048 21194
rect 48082 21160 48242 21194
rect 48032 21144 48242 21160
rect 47762 21127 47913 21143
rect 47762 21093 47863 21127
rect 47897 21093 47913 21127
rect 47762 21077 47913 21093
rect 46168 21050 46228 21076
rect 46286 21050 46346 21076
rect 46404 21050 46464 21076
rect 46522 21056 46582 21076
rect 46522 21050 46583 21056
rect 46640 21050 46700 21076
rect 46758 21050 46818 21076
rect 40360 20997 40376 21031
rect 40410 20997 40426 21031
rect 40360 20981 40426 20997
rect 40242 20914 40308 20930
rect 40242 20880 40258 20914
rect 40292 20880 40308 20914
rect 40242 20864 40308 20880
rect 40245 20842 40305 20864
rect 20434 20437 20494 20463
rect 19888 20237 19948 20263
rect 20006 20237 20066 20263
rect 20124 20237 20184 20263
rect 20242 20237 20302 20263
rect 20061 20182 20127 20190
rect 19692 20174 20127 20182
rect 19692 20140 20077 20174
rect 20111 20140 20127 20174
rect 19692 20131 20127 20140
rect 10571 20120 10637 20127
rect 13715 20120 13781 20127
rect 16917 20124 16983 20131
rect 20061 20124 20127 20131
rect 22824 20178 22884 20459
rect 23566 20433 23626 20459
rect 23020 20233 23080 20259
rect 23138 20233 23198 20259
rect 23256 20233 23316 20259
rect 23374 20233 23434 20259
rect 23193 20178 23259 20186
rect 22824 20170 23259 20178
rect 22824 20136 23209 20170
rect 23243 20136 23259 20170
rect 22824 20127 23259 20136
rect 25968 20178 26028 20459
rect 26710 20433 26770 20459
rect 41249 20815 41309 20841
rect 40245 20616 40305 20642
rect 42547 20815 42607 20841
rect 43147 20815 43207 20841
rect 46405 20865 46463 21050
rect 44445 20815 44505 20841
rect 46405 20839 46465 20865
rect 46523 20839 46583 21050
rect 46876 21044 46936 21076
rect 46994 21050 47054 21076
rect 47112 21050 47172 21076
rect 46873 21028 46939 21044
rect 47762 21038 47822 21077
rect 48182 21038 48242 21144
rect 48536 21203 48596 21370
rect 48654 21344 48714 21370
rect 48679 21203 48746 21210
rect 48536 21194 48746 21203
rect 48536 21160 48696 21194
rect 48730 21160 48746 21194
rect 48536 21144 48746 21160
rect 48298 21110 48364 21126
rect 48298 21076 48314 21110
rect 48348 21076 48364 21110
rect 48298 21060 48364 21076
rect 48416 21111 48482 21126
rect 48416 21077 48432 21111
rect 48466 21077 48482 21111
rect 48416 21061 48482 21077
rect 48300 21038 48360 21060
rect 48418 21038 48478 21061
rect 48536 21038 48596 21144
rect 49060 21142 49120 21445
rect 48970 21126 49120 21142
rect 48970 21092 48986 21126
rect 49020 21092 49120 21126
rect 48970 21076 49120 21092
rect 49060 21038 49120 21076
rect 49660 21337 49720 21995
rect 50373 21993 50916 22044
rect 50958 22037 51034 22044
rect 51092 22037 51152 22063
rect 54171 22258 54231 22284
rect 54289 22258 54349 22284
rect 54407 22258 54467 22284
rect 53297 22212 53357 22238
rect 50958 21993 51033 22037
rect 52944 22016 53004 22038
rect 53062 22022 53122 22038
rect 52941 22000 53007 22016
rect 49962 21793 50258 21853
rect 49962 21770 50022 21793
rect 50080 21770 50140 21793
rect 50198 21770 50258 21793
rect 50316 21794 50612 21854
rect 50316 21770 50376 21794
rect 50434 21770 50494 21794
rect 50552 21770 50612 21794
rect 50958 21840 51018 21993
rect 52941 21966 52957 22000
rect 52991 21966 53007 22000
rect 52941 21950 53007 21966
rect 53056 22000 53130 22022
rect 53056 21966 53075 22000
rect 53109 21966 53130 22000
rect 55492 22275 55788 22326
rect 55492 22258 55552 22275
rect 55610 22258 55670 22275
rect 55728 22258 55788 22275
rect 56069 22258 56129 22284
rect 56187 22258 56247 22284
rect 56305 22258 56365 22284
rect 59502 22442 59562 22468
rect 59620 22442 59680 22653
rect 59973 22647 60033 22679
rect 60091 22653 60151 22679
rect 60209 22653 60269 22679
rect 59970 22631 60036 22647
rect 59970 22597 59986 22631
rect 60020 22597 60036 22631
rect 59970 22581 60036 22597
rect 59852 22514 59918 22530
rect 59852 22480 59868 22514
rect 59902 22480 59918 22514
rect 59852 22464 59918 22480
rect 61213 22477 61509 22528
rect 59855 22442 59915 22464
rect 61213 22462 61273 22477
rect 61331 22462 61391 22477
rect 61449 22462 61509 22477
rect 61567 22462 61627 22488
rect 61685 22462 61745 22488
rect 61803 22462 61863 22488
rect 63111 22477 63407 22528
rect 63111 22462 63171 22477
rect 63229 22462 63289 22477
rect 63347 22462 63407 22477
rect 63465 22462 63525 22488
rect 63583 22462 63643 22488
rect 63701 22462 63761 22488
rect 57390 22275 57686 22326
rect 57390 22258 57450 22275
rect 57508 22258 57568 22275
rect 57626 22258 57686 22275
rect 54171 22041 54231 22058
rect 54289 22041 54349 22058
rect 54407 22041 54467 22058
rect 54655 22041 54715 22058
rect 54171 21990 54715 22041
rect 54773 22032 54833 22058
rect 54891 22032 54951 22058
rect 55009 22039 55069 22058
rect 55127 22039 55187 22058
rect 55245 22039 55305 22058
rect 55492 22039 55552 22058
rect 55610 22039 55670 22058
rect 53056 21909 53130 21966
rect 54296 21909 54356 21990
rect 55009 21988 55552 22039
rect 55594 22032 55670 22039
rect 55728 22032 55788 22058
rect 56069 22041 56129 22058
rect 56187 22041 56247 22058
rect 56305 22041 56365 22058
rect 56553 22041 56613 22058
rect 55594 21988 55669 22032
rect 56069 21990 56613 22041
rect 56671 22032 56731 22058
rect 56789 22032 56849 22058
rect 56907 22039 56967 22058
rect 57025 22039 57085 22058
rect 57143 22039 57203 22058
rect 57390 22039 57450 22058
rect 57508 22039 57568 22058
rect 53056 21884 54356 21909
rect 50958 21816 51212 21840
rect 53055 21836 54356 21884
rect 55594 21868 55654 21988
rect 50958 21782 51162 21816
rect 51196 21782 51212 21816
rect 50958 21766 51212 21782
rect 49962 21344 50022 21370
rect 49660 21321 49727 21337
rect 49660 21287 49676 21321
rect 49710 21287 49727 21321
rect 49660 21271 49727 21287
rect 49660 21143 49720 21271
rect 49930 21203 49997 21210
rect 50080 21203 50140 21370
rect 50198 21344 50258 21370
rect 50316 21344 50376 21370
rect 49930 21194 50140 21203
rect 49930 21160 49946 21194
rect 49980 21160 50140 21194
rect 49930 21144 50140 21160
rect 49660 21127 49811 21143
rect 49660 21093 49761 21127
rect 49795 21093 49811 21127
rect 49660 21077 49811 21093
rect 49660 21038 49720 21077
rect 50080 21038 50140 21144
rect 50434 21203 50494 21370
rect 50552 21344 50612 21370
rect 50575 21204 50642 21211
rect 50569 21203 50642 21204
rect 50434 21195 50642 21203
rect 50434 21161 50592 21195
rect 50626 21161 50642 21195
rect 50434 21145 50642 21161
rect 50434 21144 50631 21145
rect 50196 21110 50262 21126
rect 50196 21076 50212 21110
rect 50246 21076 50262 21110
rect 50196 21060 50262 21076
rect 50314 21111 50380 21126
rect 50314 21077 50330 21111
rect 50364 21077 50380 21111
rect 50314 21061 50380 21077
rect 50198 21038 50258 21060
rect 50316 21038 50376 21061
rect 50434 21038 50494 21144
rect 50958 21142 51018 21766
rect 52702 21292 52998 21328
rect 52702 21271 52762 21292
rect 52820 21271 52880 21292
rect 52938 21271 52998 21292
rect 53056 21291 53352 21327
rect 53056 21271 53116 21291
rect 53174 21271 53234 21291
rect 53292 21271 53352 21291
rect 53410 21291 53706 21327
rect 53410 21271 53470 21291
rect 53528 21271 53588 21291
rect 53646 21271 53706 21291
rect 50868 21126 51018 21142
rect 50868 21092 50884 21126
rect 50918 21092 51018 21126
rect 50868 21076 51018 21092
rect 50958 21038 51018 21076
rect 54296 21138 54356 21836
rect 54598 21788 54894 21848
rect 54598 21765 54658 21788
rect 54716 21765 54776 21788
rect 54834 21765 54894 21788
rect 54952 21789 55248 21849
rect 55593 21848 55654 21868
rect 54952 21765 55012 21789
rect 55070 21765 55130 21789
rect 55188 21765 55248 21789
rect 55574 21832 55654 21848
rect 55574 21798 55589 21832
rect 55623 21798 55654 21832
rect 55574 21782 55654 21798
rect 55593 21759 55654 21782
rect 55594 21613 55654 21759
rect 55593 21440 55654 21613
rect 54598 21339 54658 21365
rect 54566 21198 54633 21205
rect 54716 21198 54776 21365
rect 54834 21339 54894 21365
rect 54952 21339 55012 21365
rect 54566 21189 54776 21198
rect 54566 21155 54582 21189
rect 54616 21155 54776 21189
rect 54566 21139 54776 21155
rect 54296 21122 54447 21138
rect 54296 21088 54397 21122
rect 54431 21088 54447 21122
rect 54296 21072 54447 21088
rect 52702 21045 52762 21071
rect 52820 21045 52880 21071
rect 52938 21045 52998 21071
rect 53056 21051 53116 21071
rect 53056 21045 53117 21051
rect 53174 21045 53234 21071
rect 53292 21045 53352 21071
rect 46873 20994 46889 21028
rect 46923 20994 46939 21028
rect 46873 20978 46939 20994
rect 46755 20911 46821 20927
rect 46755 20877 46771 20911
rect 46805 20877 46821 20911
rect 46755 20861 46821 20877
rect 46758 20839 46818 20861
rect 41669 20615 41729 20641
rect 41787 20615 41847 20641
rect 41905 20615 41965 20641
rect 42023 20615 42083 20641
rect 43567 20615 43627 20641
rect 43685 20615 43745 20641
rect 43803 20615 43863 20641
rect 43921 20615 43981 20641
rect 39892 20420 39952 20442
rect 40010 20420 40070 20442
rect 39889 20404 39955 20420
rect 39889 20370 39905 20404
rect 39939 20370 39955 20404
rect 39889 20354 39955 20370
rect 40007 20404 40073 20420
rect 40007 20370 40023 20404
rect 40057 20370 40073 20404
rect 47762 20812 47822 20838
rect 46758 20613 46818 20639
rect 49060 20812 49120 20838
rect 49660 20812 49720 20838
rect 52939 20860 52997 21045
rect 50958 20812 51018 20838
rect 52939 20834 52999 20860
rect 53057 20834 53117 21045
rect 53410 21039 53470 21071
rect 53528 21045 53588 21071
rect 53646 21045 53706 21071
rect 53407 21023 53473 21039
rect 54296 21033 54356 21072
rect 54716 21033 54776 21139
rect 55070 21198 55130 21365
rect 55188 21339 55248 21365
rect 55213 21198 55280 21205
rect 55070 21189 55280 21198
rect 55070 21155 55230 21189
rect 55264 21155 55280 21189
rect 55070 21139 55280 21155
rect 54832 21105 54898 21121
rect 54832 21071 54848 21105
rect 54882 21071 54898 21105
rect 54832 21055 54898 21071
rect 54950 21106 55016 21121
rect 54950 21072 54966 21106
rect 55000 21072 55016 21106
rect 54950 21056 55016 21072
rect 54834 21033 54894 21055
rect 54952 21033 55012 21056
rect 55070 21033 55130 21139
rect 55594 21137 55654 21440
rect 55504 21121 55654 21137
rect 55504 21087 55520 21121
rect 55554 21087 55654 21121
rect 55504 21071 55654 21087
rect 55594 21033 55654 21071
rect 56194 21332 56254 21990
rect 56907 21988 57450 22039
rect 57492 22032 57568 22039
rect 57626 22032 57686 22058
rect 60729 22262 60789 22288
rect 60847 22262 60907 22288
rect 60965 22262 61025 22288
rect 59855 22216 59915 22242
rect 57492 21988 57567 22032
rect 59502 22020 59562 22042
rect 59620 22026 59680 22042
rect 59499 22004 59565 22020
rect 56496 21788 56792 21848
rect 56496 21765 56556 21788
rect 56614 21765 56674 21788
rect 56732 21765 56792 21788
rect 56850 21789 57146 21849
rect 56850 21765 56910 21789
rect 56968 21765 57028 21789
rect 57086 21765 57146 21789
rect 57492 21835 57552 21988
rect 59499 21970 59515 22004
rect 59549 21970 59565 22004
rect 59499 21954 59565 21970
rect 59614 22004 59688 22026
rect 59614 21970 59633 22004
rect 59667 21970 59688 22004
rect 62050 22279 62346 22330
rect 62050 22262 62110 22279
rect 62168 22262 62228 22279
rect 62286 22262 62346 22279
rect 62627 22262 62687 22288
rect 62745 22262 62805 22288
rect 62863 22262 62923 22288
rect 63948 22279 64244 22330
rect 63948 22262 64008 22279
rect 64066 22262 64126 22279
rect 64184 22262 64244 22279
rect 60729 22045 60789 22062
rect 60847 22045 60907 22062
rect 60965 22045 61025 22062
rect 61213 22045 61273 22062
rect 60729 21994 61273 22045
rect 61331 22036 61391 22062
rect 61449 22036 61509 22062
rect 61567 22043 61627 22062
rect 61685 22043 61745 22062
rect 61803 22043 61863 22062
rect 62050 22043 62110 22062
rect 62168 22043 62228 22062
rect 59614 21913 59688 21970
rect 60854 21913 60914 21994
rect 61567 21992 62110 22043
rect 62152 22036 62228 22043
rect 62286 22036 62346 22062
rect 62627 22045 62687 22062
rect 62745 22045 62805 22062
rect 62863 22045 62923 22062
rect 63111 22045 63171 22062
rect 62152 21992 62227 22036
rect 62627 21994 63171 22045
rect 63229 22036 63289 22062
rect 63347 22036 63407 22062
rect 63465 22043 63525 22062
rect 63583 22043 63643 22062
rect 63701 22043 63761 22062
rect 63948 22043 64008 22062
rect 64066 22043 64126 22062
rect 59614 21888 60914 21913
rect 59613 21840 60914 21888
rect 62152 21872 62212 21992
rect 57492 21811 57746 21835
rect 57492 21777 57696 21811
rect 57730 21777 57746 21811
rect 57492 21761 57746 21777
rect 56496 21339 56556 21365
rect 56194 21316 56261 21332
rect 56194 21282 56210 21316
rect 56244 21282 56261 21316
rect 56194 21266 56261 21282
rect 56194 21138 56254 21266
rect 56464 21198 56531 21205
rect 56614 21198 56674 21365
rect 56732 21339 56792 21365
rect 56850 21339 56910 21365
rect 56464 21189 56674 21198
rect 56464 21155 56480 21189
rect 56514 21155 56674 21189
rect 56464 21139 56674 21155
rect 56194 21122 56345 21138
rect 56194 21088 56295 21122
rect 56329 21088 56345 21122
rect 56194 21072 56345 21088
rect 56194 21033 56254 21072
rect 56614 21033 56674 21139
rect 56968 21198 57028 21365
rect 57086 21339 57146 21365
rect 57109 21199 57176 21206
rect 57103 21198 57176 21199
rect 56968 21190 57176 21198
rect 56968 21156 57126 21190
rect 57160 21156 57176 21190
rect 56968 21140 57176 21156
rect 56968 21139 57165 21140
rect 56730 21105 56796 21121
rect 56730 21071 56746 21105
rect 56780 21071 56796 21105
rect 56730 21055 56796 21071
rect 56848 21106 56914 21121
rect 56848 21072 56864 21106
rect 56898 21072 56914 21106
rect 56848 21056 56914 21072
rect 56732 21033 56792 21055
rect 56850 21033 56910 21056
rect 56968 21033 57028 21139
rect 57492 21137 57552 21761
rect 59260 21296 59556 21332
rect 59260 21275 59320 21296
rect 59378 21275 59438 21296
rect 59496 21275 59556 21296
rect 59614 21295 59910 21331
rect 59614 21275 59674 21295
rect 59732 21275 59792 21295
rect 59850 21275 59910 21295
rect 59968 21295 60264 21331
rect 59968 21275 60028 21295
rect 60086 21275 60146 21295
rect 60204 21275 60264 21295
rect 57402 21121 57552 21137
rect 57402 21087 57418 21121
rect 57452 21087 57552 21121
rect 57402 21071 57552 21087
rect 60854 21142 60914 21840
rect 61156 21792 61452 21852
rect 61156 21769 61216 21792
rect 61274 21769 61334 21792
rect 61392 21769 61452 21792
rect 61510 21793 61806 21853
rect 62151 21852 62212 21872
rect 61510 21769 61570 21793
rect 61628 21769 61688 21793
rect 61746 21769 61806 21793
rect 62132 21836 62212 21852
rect 62132 21802 62147 21836
rect 62181 21802 62212 21836
rect 62132 21786 62212 21802
rect 62151 21763 62212 21786
rect 62152 21617 62212 21763
rect 62151 21444 62212 21617
rect 61156 21343 61216 21369
rect 61124 21202 61191 21209
rect 61274 21202 61334 21369
rect 61392 21343 61452 21369
rect 61510 21343 61570 21369
rect 61124 21193 61334 21202
rect 61124 21159 61140 21193
rect 61174 21159 61334 21193
rect 61124 21143 61334 21159
rect 60854 21126 61005 21142
rect 60854 21092 60955 21126
rect 60989 21092 61005 21126
rect 60854 21076 61005 21092
rect 57492 21033 57552 21071
rect 59260 21049 59320 21075
rect 59378 21049 59438 21075
rect 59496 21049 59556 21075
rect 59614 21055 59674 21075
rect 59614 21049 59675 21055
rect 59732 21049 59792 21075
rect 59850 21049 59910 21075
rect 53407 20989 53423 21023
rect 53457 20989 53473 21023
rect 53407 20973 53473 20989
rect 53289 20906 53355 20922
rect 53289 20872 53305 20906
rect 53339 20872 53355 20906
rect 53289 20856 53355 20872
rect 53292 20834 53352 20856
rect 48182 20612 48242 20638
rect 48300 20612 48360 20638
rect 48418 20612 48478 20638
rect 48536 20612 48596 20638
rect 50080 20612 50140 20638
rect 50198 20612 50258 20638
rect 50316 20612 50376 20638
rect 50434 20612 50494 20638
rect 46405 20417 46465 20439
rect 46523 20417 46583 20439
rect 46402 20401 46468 20417
rect 40007 20354 40073 20370
rect 46402 20367 46418 20401
rect 46452 20367 46468 20401
rect 46402 20351 46468 20367
rect 46520 20401 46586 20417
rect 46520 20367 46536 20401
rect 46570 20367 46586 20401
rect 54296 20807 54356 20833
rect 53292 20608 53352 20634
rect 55594 20807 55654 20833
rect 56194 20807 56254 20833
rect 59497 20864 59555 21049
rect 59497 20838 59557 20864
rect 59615 20838 59675 21049
rect 59968 21043 60028 21075
rect 60086 21049 60146 21075
rect 60204 21049 60264 21075
rect 59965 21027 60031 21043
rect 60854 21037 60914 21076
rect 61274 21037 61334 21143
rect 61628 21202 61688 21369
rect 61746 21343 61806 21369
rect 61771 21202 61838 21209
rect 61628 21193 61838 21202
rect 61628 21159 61788 21193
rect 61822 21159 61838 21193
rect 61628 21143 61838 21159
rect 61390 21109 61456 21125
rect 61390 21075 61406 21109
rect 61440 21075 61456 21109
rect 61390 21059 61456 21075
rect 61508 21110 61574 21125
rect 61508 21076 61524 21110
rect 61558 21076 61574 21110
rect 61508 21060 61574 21076
rect 61392 21037 61452 21059
rect 61510 21037 61570 21060
rect 61628 21037 61688 21143
rect 62152 21141 62212 21444
rect 62062 21125 62212 21141
rect 62062 21091 62078 21125
rect 62112 21091 62212 21125
rect 62062 21075 62212 21091
rect 62152 21037 62212 21075
rect 62752 21336 62812 21994
rect 63465 21992 64008 22043
rect 64050 22036 64126 22043
rect 64184 22036 64244 22062
rect 64050 21992 64125 22036
rect 63054 21792 63350 21852
rect 63054 21769 63114 21792
rect 63172 21769 63232 21792
rect 63290 21769 63350 21792
rect 63408 21793 63704 21853
rect 63408 21769 63468 21793
rect 63526 21769 63586 21793
rect 63644 21769 63704 21793
rect 64050 21839 64110 21992
rect 70658 21955 70713 22015
rect 70913 21956 71643 22015
rect 70913 21955 71216 21956
rect 70658 21897 70697 21955
rect 71199 21898 71216 21955
rect 71271 21955 71643 21956
rect 71271 21898 71286 21955
rect 64050 21815 64304 21839
rect 64050 21781 64254 21815
rect 64288 21781 64304 21815
rect 64050 21765 64304 21781
rect 70658 21837 70713 21897
rect 70913 21837 70939 21897
rect 71199 21879 71286 21898
rect 70658 21779 70697 21837
rect 63054 21343 63114 21369
rect 62752 21320 62819 21336
rect 62752 21286 62768 21320
rect 62802 21286 62819 21320
rect 62752 21270 62819 21286
rect 62752 21142 62812 21270
rect 63022 21202 63089 21209
rect 63172 21202 63232 21369
rect 63290 21343 63350 21369
rect 63408 21343 63468 21369
rect 63022 21193 63232 21202
rect 63022 21159 63038 21193
rect 63072 21159 63232 21193
rect 63022 21143 63232 21159
rect 62752 21126 62903 21142
rect 62752 21092 62853 21126
rect 62887 21092 62903 21126
rect 62752 21076 62903 21092
rect 62752 21037 62812 21076
rect 63172 21037 63232 21143
rect 63526 21202 63586 21369
rect 63644 21343 63704 21369
rect 63667 21203 63734 21210
rect 63661 21202 63734 21203
rect 63526 21194 63734 21202
rect 63526 21160 63684 21194
rect 63718 21160 63734 21194
rect 63526 21144 63734 21160
rect 63526 21143 63723 21144
rect 63288 21109 63354 21125
rect 63288 21075 63304 21109
rect 63338 21075 63354 21109
rect 63288 21059 63354 21075
rect 63406 21110 63472 21125
rect 63406 21076 63422 21110
rect 63456 21076 63472 21110
rect 63406 21060 63472 21076
rect 63290 21037 63350 21059
rect 63408 21037 63468 21060
rect 63526 21037 63586 21143
rect 64050 21141 64110 21765
rect 70658 21719 70713 21779
rect 70913 21719 70939 21779
rect 70459 21514 70513 21574
rect 70913 21514 70939 21574
rect 70459 21456 70498 21514
rect 70459 21396 70513 21456
rect 70913 21396 71388 21456
rect 70459 21338 70498 21396
rect 70459 21278 70513 21338
rect 70913 21278 70939 21338
rect 63960 21125 64110 21141
rect 63960 21091 63976 21125
rect 64010 21091 64110 21125
rect 63960 21075 64110 21091
rect 64050 21037 64110 21075
rect 70459 21047 70513 21107
rect 70913 21047 70939 21107
rect 59965 20993 59981 21027
rect 60015 20993 60031 21027
rect 59965 20977 60031 20993
rect 59847 20910 59913 20926
rect 59847 20876 59863 20910
rect 59897 20876 59913 20910
rect 59847 20860 59913 20876
rect 59850 20838 59910 20860
rect 57492 20807 57552 20833
rect 54716 20607 54776 20633
rect 54834 20607 54894 20633
rect 54952 20607 55012 20633
rect 55070 20607 55130 20633
rect 56614 20607 56674 20633
rect 56732 20607 56792 20633
rect 56850 20607 56910 20633
rect 56968 20607 57028 20633
rect 52939 20412 52999 20434
rect 53057 20412 53117 20434
rect 52936 20396 53002 20412
rect 46520 20351 46586 20367
rect 26164 20233 26224 20259
rect 26282 20233 26342 20259
rect 26400 20233 26460 20259
rect 26518 20233 26578 20259
rect 26337 20178 26403 20186
rect 25968 20170 26403 20178
rect 25968 20136 26353 20170
rect 26387 20136 26403 20170
rect 52936 20362 52952 20396
rect 52986 20362 53002 20396
rect 52936 20346 53002 20362
rect 53054 20396 53120 20412
rect 53054 20362 53070 20396
rect 53104 20362 53120 20396
rect 60854 20811 60914 20837
rect 59850 20612 59910 20638
rect 62152 20811 62212 20837
rect 62752 20811 62812 20837
rect 70459 20989 70498 21047
rect 70459 20929 70513 20989
rect 70913 20988 70939 20989
rect 71100 20988 71166 20991
rect 70913 20975 71166 20988
rect 70913 20941 71116 20975
rect 71150 20941 71166 20975
rect 70913 20929 71166 20941
rect 71331 20989 71388 21396
rect 71598 21181 71643 21955
rect 71598 21121 71846 21181
rect 72046 21121 72072 21181
rect 71487 20989 71566 21000
rect 71331 20987 71846 20989
rect 71331 20929 71500 20987
rect 71555 20929 71846 20987
rect 72246 20929 72272 20989
rect 64050 20811 64110 20837
rect 70459 20871 70498 20929
rect 71099 20925 71166 20929
rect 71487 20919 71566 20929
rect 71200 20871 71287 20888
rect 70459 20811 70513 20871
rect 70913 20811 70939 20871
rect 71200 20869 71846 20871
rect 71200 20811 71215 20869
rect 71270 20811 71846 20869
rect 72246 20811 72272 20871
rect 71200 20793 71287 20811
rect 61274 20611 61334 20637
rect 61392 20611 61452 20637
rect 61510 20611 61570 20637
rect 61628 20611 61688 20637
rect 63172 20611 63232 20637
rect 63290 20611 63350 20637
rect 63408 20611 63468 20637
rect 63526 20611 63586 20637
rect 70459 20693 70513 20753
rect 70913 20693 70939 20753
rect 70459 20635 70498 20693
rect 71238 20635 71287 20793
rect 71720 20753 71786 20756
rect 72319 20798 72385 20814
rect 72319 20764 72335 20798
rect 72369 20764 72385 20798
rect 71720 20740 71846 20753
rect 71720 20706 71736 20740
rect 71770 20706 71846 20740
rect 71720 20693 71846 20706
rect 72246 20693 72272 20753
rect 72319 20748 72385 20764
rect 71720 20690 71786 20693
rect 70459 20575 70513 20635
rect 70913 20575 71287 20635
rect 71329 20635 71398 20640
rect 71329 20621 71846 20635
rect 71329 20587 71346 20621
rect 71380 20587 71846 20621
rect 71329 20575 71846 20587
rect 72246 20575 72272 20635
rect 59497 20416 59557 20438
rect 59615 20416 59675 20438
rect 59494 20400 59560 20416
rect 53054 20346 53120 20362
rect 59494 20366 59510 20400
rect 59544 20366 59560 20400
rect 59494 20350 59560 20366
rect 59612 20400 59678 20416
rect 59612 20366 59628 20400
rect 59662 20366 59678 20400
rect 70459 20517 70498 20575
rect 71329 20571 71396 20575
rect 70459 20457 70513 20517
rect 70913 20457 70939 20517
rect 59612 20350 59678 20366
rect 70459 20220 70513 20280
rect 70913 20220 70939 20280
rect 70459 20162 70498 20220
rect 71329 20162 71386 20571
rect 72327 20439 72378 20748
rect 25968 20127 26403 20136
rect 23193 20120 23259 20127
rect 26337 20120 26403 20127
rect 70459 20102 70513 20162
rect 70913 20102 71386 20162
rect 71598 20379 71846 20439
rect 72046 20379 72378 20439
rect 70459 20044 70498 20102
rect 70459 19984 70513 20044
rect 70913 19984 70939 20044
rect 70658 19747 70713 19807
rect 70913 19747 70939 19807
rect 70658 19689 70697 19747
rect 70658 19629 70713 19689
rect 70913 19629 70939 19689
rect 71059 19665 71125 19681
rect 71059 19631 71075 19665
rect 71109 19631 71125 19665
rect 70658 19571 70697 19629
rect 71059 19615 71125 19631
rect 71062 19571 71122 19615
rect 71598 19571 71643 20379
rect 70658 19511 70713 19571
rect 70913 19511 71643 19571
rect 40430 19167 40496 19183
rect 40430 19158 40446 19167
rect 39909 19133 40446 19158
rect 40480 19133 40496 19167
rect 41560 19161 41626 19177
rect 41560 19154 41576 19161
rect 39909 19115 40496 19133
rect 41051 19127 41576 19154
rect 41610 19127 41626 19161
rect 39909 19063 39953 19115
rect 41051 19111 41626 19127
rect 39657 19022 39953 19063
rect 39657 19001 39717 19022
rect 39775 19001 39835 19022
rect 39893 19001 39953 19022
rect 40011 19047 40496 19063
rect 41051 19059 41095 19111
rect 46988 19163 47054 19179
rect 46988 19154 47004 19163
rect 46467 19129 47004 19154
rect 47038 19129 47054 19163
rect 48118 19157 48184 19173
rect 48118 19150 48134 19157
rect 46467 19111 47054 19129
rect 47609 19123 48134 19150
rect 48168 19123 48184 19157
rect 46467 19059 46511 19111
rect 47609 19107 48184 19123
rect 40011 19022 40446 19047
rect 40011 19001 40071 19022
rect 40129 19001 40189 19022
rect 40247 19021 40446 19022
rect 40247 19001 40307 19021
rect 40430 19013 40446 19021
rect 40480 19013 40496 19047
rect 40430 18997 40496 19013
rect 40799 19018 41095 19059
rect 40799 18997 40859 19018
rect 40917 18997 40977 19018
rect 41035 18997 41095 19018
rect 41153 19043 41626 19059
rect 41153 19018 41576 19043
rect 41153 18997 41213 19018
rect 41271 18997 41331 19018
rect 41389 19017 41576 19018
rect 41389 18997 41449 19017
rect 41560 19009 41576 19017
rect 41610 19009 41626 19043
rect 39657 18575 39717 18601
rect 39775 18575 39835 18601
rect 39893 18400 39953 18601
rect 40011 18575 40071 18601
rect 40129 18575 40189 18601
rect 40247 18584 40307 18601
rect 41560 18993 41626 19009
rect 46215 19018 46511 19059
rect 46215 18997 46275 19018
rect 46333 18997 46393 19018
rect 46451 18997 46511 19018
rect 46569 19043 47054 19059
rect 47609 19055 47653 19107
rect 53522 19168 53588 19184
rect 53522 19159 53538 19168
rect 53001 19134 53538 19159
rect 53572 19134 53588 19168
rect 54652 19162 54718 19178
rect 54652 19155 54668 19162
rect 53001 19116 53588 19134
rect 54143 19128 54668 19155
rect 54702 19128 54718 19162
rect 53001 19064 53045 19116
rect 54143 19112 54718 19128
rect 46569 19018 47004 19043
rect 46569 18997 46629 19018
rect 46687 18997 46747 19018
rect 46805 19017 47004 19018
rect 46805 18997 46865 19017
rect 46988 19009 47004 19017
rect 47038 19009 47054 19043
rect 42770 18945 43066 18981
rect 42770 18925 42830 18945
rect 42888 18925 42948 18945
rect 43006 18925 43066 18945
rect 43124 18945 43420 18981
rect 43124 18925 43184 18945
rect 43242 18925 43302 18945
rect 43360 18925 43420 18945
rect 43478 18946 43774 18982
rect 43478 18925 43538 18946
rect 43596 18925 43656 18946
rect 43714 18925 43774 18946
rect 42770 18699 42830 18725
rect 42888 18699 42948 18725
rect 43006 18693 43066 18725
rect 43124 18699 43184 18725
rect 43242 18699 43302 18725
rect 43360 18705 43420 18725
rect 43359 18699 43420 18705
rect 43478 18699 43538 18725
rect 43596 18699 43656 18725
rect 43714 18699 43774 18725
rect 43003 18677 43069 18693
rect 43003 18643 43019 18677
rect 43053 18643 43069 18677
rect 43003 18627 43069 18643
rect 40246 18495 40307 18584
rect 40799 18571 40859 18597
rect 40917 18571 40977 18597
rect 40246 18442 40397 18495
rect 39893 18349 40279 18400
rect 40098 18291 40164 18307
rect 40098 18257 40114 18291
rect 40148 18257 40164 18291
rect 39582 18218 39642 18244
rect 39700 18218 39760 18244
rect 39818 18218 39878 18244
rect 40098 18241 40164 18257
rect 40101 18218 40161 18241
rect 40219 18218 40279 18349
rect 40337 18218 40397 18442
rect 41035 18396 41095 18597
rect 41153 18571 41213 18597
rect 41271 18571 41331 18597
rect 41389 18580 41449 18597
rect 41388 18491 41449 18580
rect 43121 18560 43187 18576
rect 43121 18526 43137 18560
rect 43171 18526 43187 18560
rect 43121 18510 43187 18526
rect 41388 18438 41539 18491
rect 43124 18488 43184 18510
rect 43359 18488 43419 18699
rect 43479 18514 43537 18699
rect 46988 18993 47054 19009
rect 47357 19014 47653 19055
rect 47357 18993 47417 19014
rect 47475 18993 47535 19014
rect 47593 18993 47653 19014
rect 47711 19039 48184 19055
rect 47711 19014 48134 19039
rect 47711 18993 47771 19014
rect 47829 18993 47889 19014
rect 47947 19013 48134 19014
rect 47947 18993 48007 19013
rect 48118 19005 48134 19013
rect 48168 19005 48184 19039
rect 46215 18571 46275 18597
rect 46333 18571 46393 18597
rect 43477 18488 43537 18514
rect 41035 18345 41421 18396
rect 41240 18287 41306 18303
rect 41240 18253 41256 18287
rect 41290 18253 41306 18287
rect 40724 18214 40784 18240
rect 40842 18214 40902 18240
rect 40960 18214 41020 18240
rect 41240 18237 41306 18253
rect 41243 18214 41303 18237
rect 41361 18214 41421 18345
rect 41479 18214 41539 18438
rect 43124 18262 43184 18288
rect 39582 17986 39642 18018
rect 39700 17986 39760 18018
rect 39818 17986 39878 18018
rect 40101 17986 40161 18018
rect 40219 17992 40279 18018
rect 40337 17992 40397 18018
rect 46451 18396 46511 18597
rect 46569 18571 46629 18597
rect 46687 18571 46747 18597
rect 46805 18580 46865 18597
rect 48118 18989 48184 19005
rect 52749 19023 53045 19064
rect 52749 19002 52809 19023
rect 52867 19002 52927 19023
rect 52985 19002 53045 19023
rect 53103 19048 53588 19064
rect 54143 19060 54187 19112
rect 60035 19171 60101 19187
rect 60035 19162 60051 19171
rect 59514 19137 60051 19162
rect 60085 19137 60101 19171
rect 61165 19165 61231 19181
rect 61165 19158 61181 19165
rect 59514 19119 60101 19137
rect 60656 19131 61181 19158
rect 61215 19131 61231 19165
rect 59514 19067 59558 19119
rect 60656 19115 61231 19131
rect 53103 19023 53538 19048
rect 53103 19002 53163 19023
rect 53221 19002 53281 19023
rect 53339 19022 53538 19023
rect 53339 19002 53399 19022
rect 53522 19014 53538 19022
rect 53572 19014 53588 19048
rect 49328 18941 49624 18977
rect 49328 18921 49388 18941
rect 49446 18921 49506 18941
rect 49564 18921 49624 18941
rect 49682 18941 49978 18977
rect 49682 18921 49742 18941
rect 49800 18921 49860 18941
rect 49918 18921 49978 18941
rect 50036 18942 50332 18978
rect 50036 18921 50096 18942
rect 50154 18921 50214 18942
rect 50272 18921 50332 18942
rect 49328 18695 49388 18721
rect 49446 18695 49506 18721
rect 49564 18689 49624 18721
rect 49682 18695 49742 18721
rect 49800 18695 49860 18721
rect 49918 18701 49978 18721
rect 49917 18695 49978 18701
rect 50036 18695 50096 18721
rect 50154 18695 50214 18721
rect 50272 18695 50332 18721
rect 49561 18673 49627 18689
rect 49561 18639 49577 18673
rect 49611 18639 49627 18673
rect 49561 18623 49627 18639
rect 46804 18491 46865 18580
rect 47357 18567 47417 18593
rect 47475 18567 47535 18593
rect 46804 18438 46955 18491
rect 46451 18345 46837 18396
rect 46656 18287 46722 18303
rect 46656 18253 46672 18287
rect 46706 18253 46722 18287
rect 46140 18214 46200 18240
rect 46258 18214 46318 18240
rect 46376 18214 46436 18240
rect 46656 18237 46722 18253
rect 46659 18214 46719 18237
rect 46777 18214 46837 18345
rect 46895 18214 46955 18438
rect 47593 18392 47653 18593
rect 47711 18567 47771 18593
rect 47829 18567 47889 18593
rect 47947 18576 48007 18593
rect 47946 18487 48007 18576
rect 49679 18556 49745 18572
rect 49679 18522 49695 18556
rect 49729 18522 49745 18556
rect 49679 18506 49745 18522
rect 47946 18434 48097 18487
rect 49682 18484 49742 18506
rect 49917 18484 49977 18695
rect 50037 18510 50095 18695
rect 53522 18998 53588 19014
rect 53891 19019 54187 19060
rect 53891 18998 53951 19019
rect 54009 18998 54069 19019
rect 54127 18998 54187 19019
rect 54245 19044 54718 19060
rect 54245 19019 54668 19044
rect 54245 18998 54305 19019
rect 54363 18998 54423 19019
rect 54481 19018 54668 19019
rect 54481 18998 54541 19018
rect 54652 19010 54668 19018
rect 54702 19010 54718 19044
rect 52749 18576 52809 18602
rect 52867 18576 52927 18602
rect 50035 18484 50095 18510
rect 47593 18341 47979 18392
rect 47798 18283 47864 18299
rect 47798 18249 47814 18283
rect 47848 18249 47864 18283
rect 43359 18066 43419 18088
rect 43477 18066 43537 18088
rect 43356 18050 43422 18066
rect 43356 18016 43372 18050
rect 43406 18016 43422 18050
rect 39582 17945 40161 17986
rect 40724 17982 40784 18014
rect 40842 17982 40902 18014
rect 40960 17982 41020 18014
rect 41243 17982 41303 18014
rect 41361 17988 41421 18014
rect 41479 17988 41539 18014
rect 43356 18000 43422 18016
rect 43474 18050 43540 18066
rect 43474 18016 43490 18050
rect 43524 18016 43540 18050
rect 43474 18000 43540 18016
rect 47282 18210 47342 18236
rect 47400 18210 47460 18236
rect 47518 18210 47578 18236
rect 47798 18233 47864 18249
rect 47801 18210 47861 18233
rect 47919 18210 47979 18341
rect 48037 18210 48097 18434
rect 49682 18258 49742 18284
rect 40724 17941 41303 17982
rect 46140 17982 46200 18014
rect 46258 17982 46318 18014
rect 46376 17982 46436 18014
rect 46659 17982 46719 18014
rect 46777 17988 46837 18014
rect 46895 17988 46955 18014
rect 52985 18401 53045 18602
rect 53103 18576 53163 18602
rect 53221 18576 53281 18602
rect 53339 18585 53399 18602
rect 54652 18994 54718 19010
rect 59262 19026 59558 19067
rect 59262 19005 59322 19026
rect 59380 19005 59440 19026
rect 59498 19005 59558 19026
rect 59616 19051 60101 19067
rect 60656 19063 60700 19115
rect 59616 19026 60051 19051
rect 59616 19005 59676 19026
rect 59734 19005 59794 19026
rect 59852 19025 60051 19026
rect 59852 19005 59912 19025
rect 60035 19017 60051 19025
rect 60085 19017 60101 19051
rect 55862 18946 56158 18982
rect 55862 18926 55922 18946
rect 55980 18926 56040 18946
rect 56098 18926 56158 18946
rect 56216 18946 56512 18982
rect 56216 18926 56276 18946
rect 56334 18926 56394 18946
rect 56452 18926 56512 18946
rect 56570 18947 56866 18983
rect 56570 18926 56630 18947
rect 56688 18926 56748 18947
rect 56806 18926 56866 18947
rect 55862 18700 55922 18726
rect 55980 18700 56040 18726
rect 56098 18694 56158 18726
rect 56216 18700 56276 18726
rect 56334 18700 56394 18726
rect 56452 18706 56512 18726
rect 56451 18700 56512 18706
rect 56570 18700 56630 18726
rect 56688 18700 56748 18726
rect 56806 18700 56866 18726
rect 56095 18678 56161 18694
rect 56095 18644 56111 18678
rect 56145 18644 56161 18678
rect 56095 18628 56161 18644
rect 53338 18496 53399 18585
rect 53891 18572 53951 18598
rect 54009 18572 54069 18598
rect 53338 18443 53489 18496
rect 52985 18350 53371 18401
rect 53190 18292 53256 18308
rect 53190 18258 53206 18292
rect 53240 18258 53256 18292
rect 52674 18219 52734 18245
rect 52792 18219 52852 18245
rect 52910 18219 52970 18245
rect 53190 18242 53256 18258
rect 53193 18219 53253 18242
rect 53311 18219 53371 18350
rect 53429 18219 53489 18443
rect 54127 18397 54187 18598
rect 54245 18572 54305 18598
rect 54363 18572 54423 18598
rect 54481 18581 54541 18598
rect 54480 18492 54541 18581
rect 56213 18561 56279 18577
rect 56213 18527 56229 18561
rect 56263 18527 56279 18561
rect 56213 18511 56279 18527
rect 54480 18439 54631 18492
rect 56216 18489 56276 18511
rect 56451 18489 56511 18700
rect 56571 18515 56629 18700
rect 60035 19001 60101 19017
rect 60404 19022 60700 19063
rect 60404 19001 60464 19022
rect 60522 19001 60582 19022
rect 60640 19001 60700 19022
rect 60758 19047 61231 19063
rect 60758 19022 61181 19047
rect 60758 19001 60818 19022
rect 60876 19001 60936 19022
rect 60994 19021 61181 19022
rect 60994 19001 61054 19021
rect 61165 19013 61181 19021
rect 61215 19013 61231 19047
rect 59262 18579 59322 18605
rect 59380 18579 59440 18605
rect 56569 18489 56629 18515
rect 54127 18346 54513 18397
rect 54332 18288 54398 18304
rect 54332 18254 54348 18288
rect 54382 18254 54398 18288
rect 49917 18062 49977 18084
rect 50035 18062 50095 18084
rect 49914 18046 49980 18062
rect 49914 18012 49930 18046
rect 49964 18012 49980 18046
rect 46140 17941 46719 17982
rect 47282 17978 47342 18010
rect 47400 17978 47460 18010
rect 47518 17978 47578 18010
rect 47801 17978 47861 18010
rect 47919 17984 47979 18010
rect 48037 17984 48097 18010
rect 49914 17996 49980 18012
rect 50032 18046 50098 18062
rect 50032 18012 50048 18046
rect 50082 18012 50098 18046
rect 53816 18215 53876 18241
rect 53934 18215 53994 18241
rect 54052 18215 54112 18241
rect 54332 18238 54398 18254
rect 54335 18215 54395 18238
rect 54453 18215 54513 18346
rect 54571 18215 54631 18439
rect 56216 18263 56276 18289
rect 50032 17996 50098 18012
rect 52674 17987 52734 18019
rect 52792 17987 52852 18019
rect 52910 17987 52970 18019
rect 53193 17987 53253 18019
rect 53311 17993 53371 18019
rect 53429 17993 53489 18019
rect 59498 18404 59558 18605
rect 59616 18579 59676 18605
rect 59734 18579 59794 18605
rect 59852 18588 59912 18605
rect 61165 18997 61231 19013
rect 62375 18949 62671 18985
rect 62375 18929 62435 18949
rect 62493 18929 62553 18949
rect 62611 18929 62671 18949
rect 62729 18949 63025 18985
rect 62729 18929 62789 18949
rect 62847 18929 62907 18949
rect 62965 18929 63025 18949
rect 63083 18950 63379 18986
rect 63083 18929 63143 18950
rect 63201 18929 63261 18950
rect 63319 18929 63379 18950
rect 70658 18811 70713 18871
rect 70913 18812 71643 18871
rect 70913 18811 71216 18812
rect 70658 18753 70697 18811
rect 71199 18754 71216 18811
rect 71271 18811 71643 18812
rect 71271 18754 71286 18811
rect 62375 18703 62435 18729
rect 62493 18703 62553 18729
rect 62611 18697 62671 18729
rect 62729 18703 62789 18729
rect 62847 18703 62907 18729
rect 62965 18709 63025 18729
rect 62964 18703 63025 18709
rect 63083 18703 63143 18729
rect 63201 18703 63261 18729
rect 63319 18703 63379 18729
rect 62608 18681 62674 18697
rect 62608 18647 62624 18681
rect 62658 18647 62674 18681
rect 62608 18631 62674 18647
rect 59851 18499 59912 18588
rect 60404 18575 60464 18601
rect 60522 18575 60582 18601
rect 59851 18446 60002 18499
rect 59498 18353 59884 18404
rect 59703 18295 59769 18311
rect 59703 18261 59719 18295
rect 59753 18261 59769 18295
rect 59187 18222 59247 18248
rect 59305 18222 59365 18248
rect 59423 18222 59483 18248
rect 59703 18245 59769 18261
rect 59706 18222 59766 18245
rect 59824 18222 59884 18353
rect 59942 18222 60002 18446
rect 60640 18400 60700 18601
rect 60758 18575 60818 18601
rect 60876 18575 60936 18601
rect 60994 18584 61054 18601
rect 60993 18495 61054 18584
rect 62726 18564 62792 18580
rect 62726 18530 62742 18564
rect 62776 18530 62792 18564
rect 62726 18514 62792 18530
rect 60993 18442 61144 18495
rect 62729 18492 62789 18514
rect 62964 18492 63024 18703
rect 63084 18518 63142 18703
rect 70658 18693 70713 18753
rect 70913 18693 70939 18753
rect 71199 18735 71286 18754
rect 70658 18635 70697 18693
rect 70658 18575 70713 18635
rect 70913 18575 70939 18635
rect 63082 18492 63142 18518
rect 60640 18349 61026 18400
rect 60845 18291 60911 18307
rect 60845 18257 60861 18291
rect 60895 18257 60911 18291
rect 56451 18067 56511 18089
rect 56569 18067 56629 18089
rect 56448 18051 56514 18067
rect 56448 18017 56464 18051
rect 56498 18017 56514 18051
rect 47282 17937 47861 17978
rect 52674 17946 53253 17987
rect 53816 17983 53876 18015
rect 53934 17983 53994 18015
rect 54052 17983 54112 18015
rect 54335 17983 54395 18015
rect 54453 17989 54513 18015
rect 54571 17989 54631 18015
rect 56448 18001 56514 18017
rect 56566 18051 56632 18067
rect 56566 18017 56582 18051
rect 56616 18017 56632 18051
rect 60329 18218 60389 18244
rect 60447 18218 60507 18244
rect 60565 18218 60625 18244
rect 60845 18241 60911 18257
rect 60848 18218 60908 18241
rect 60966 18218 61026 18349
rect 61084 18218 61144 18442
rect 62729 18266 62789 18292
rect 56566 18001 56632 18017
rect 59187 17990 59247 18022
rect 59305 17990 59365 18022
rect 59423 17990 59483 18022
rect 59706 17990 59766 18022
rect 59824 17996 59884 18022
rect 59942 17996 60002 18022
rect 70459 18370 70513 18430
rect 70913 18370 70939 18430
rect 70459 18312 70498 18370
rect 70459 18252 70513 18312
rect 70913 18252 71388 18312
rect 70459 18194 70498 18252
rect 70459 18134 70513 18194
rect 70913 18134 70939 18194
rect 62964 18070 63024 18092
rect 63082 18070 63142 18092
rect 62961 18054 63027 18070
rect 62961 18020 62977 18054
rect 63011 18020 63027 18054
rect 53816 17942 54395 17983
rect 59187 17949 59766 17990
rect 60329 17986 60389 18018
rect 60447 17986 60507 18018
rect 60565 17986 60625 18018
rect 60848 17986 60908 18018
rect 60966 17992 61026 18018
rect 61084 17992 61144 18018
rect 62961 18004 63027 18020
rect 63079 18054 63145 18070
rect 63079 18020 63095 18054
rect 63129 18020 63145 18054
rect 63079 18004 63145 18020
rect 60329 17945 60908 17986
rect 70459 17903 70513 17963
rect 70913 17903 70939 17963
rect 70459 17845 70498 17903
rect 70459 17785 70513 17845
rect 70913 17844 70939 17845
rect 71100 17844 71166 17847
rect 70913 17831 71166 17844
rect 70913 17797 71116 17831
rect 71150 17797 71166 17831
rect 70913 17785 71166 17797
rect 71331 17845 71388 18252
rect 71598 18037 71643 18811
rect 71598 17977 71846 18037
rect 72046 17977 72072 18037
rect 71487 17845 71566 17856
rect 71331 17843 71846 17845
rect 71331 17785 71500 17843
rect 71555 17785 71846 17843
rect 72246 17785 72272 17845
rect 70459 17727 70498 17785
rect 71099 17781 71166 17785
rect 71487 17775 71566 17785
rect 71200 17727 71287 17744
rect 70459 17667 70513 17727
rect 70913 17667 70939 17727
rect 71200 17725 71846 17727
rect 71200 17667 71215 17725
rect 71270 17667 71846 17725
rect 72246 17667 72272 17727
rect 71200 17649 71287 17667
rect 70459 17549 70513 17609
rect 70913 17549 70939 17609
rect 70459 17491 70498 17549
rect 71238 17491 71287 17649
rect 71720 17609 71786 17612
rect 72319 17654 72385 17670
rect 72319 17620 72335 17654
rect 72369 17620 72385 17654
rect 71720 17596 71846 17609
rect 71720 17562 71736 17596
rect 71770 17562 71846 17596
rect 71720 17549 71846 17562
rect 72246 17549 72272 17609
rect 72319 17604 72385 17620
rect 71720 17546 71786 17549
rect 70459 17431 70513 17491
rect 70913 17431 71287 17491
rect 71329 17491 71398 17496
rect 71329 17477 71846 17491
rect 71329 17443 71346 17477
rect 71380 17443 71846 17477
rect 71329 17431 71846 17443
rect 72246 17431 72272 17491
rect 42756 17295 43052 17331
rect 42756 17275 42816 17295
rect 42874 17275 42934 17295
rect 42992 17275 43052 17295
rect 43110 17295 43406 17331
rect 43110 17275 43170 17295
rect 43228 17275 43288 17295
rect 43346 17275 43406 17295
rect 43464 17296 43760 17332
rect 43464 17275 43524 17296
rect 43582 17275 43642 17296
rect 43700 17275 43760 17296
rect 5302 16970 5368 16986
rect 5302 16966 5318 16970
rect 4818 16936 5318 16966
rect 5352 16936 5368 16970
rect 6470 16970 6536 16986
rect 6470 16966 6486 16970
rect 4818 16923 5368 16936
rect 4818 16871 4862 16923
rect 5302 16920 5368 16923
rect 5986 16936 6486 16966
rect 6520 16936 6536 16970
rect 7638 16970 7704 16986
rect 7638 16966 7654 16970
rect 5986 16923 6536 16936
rect 5302 16871 5368 16878
rect 5986 16871 6030 16923
rect 6470 16920 6536 16923
rect 7154 16936 7654 16966
rect 7688 16936 7704 16970
rect 8806 16970 8872 16986
rect 8806 16966 8822 16970
rect 7154 16923 7704 16936
rect 6470 16871 6536 16878
rect 7154 16871 7198 16923
rect 7638 16920 7704 16923
rect 8322 16936 8822 16966
rect 8856 16936 8872 16970
rect 9980 16968 10046 16984
rect 9980 16964 9996 16968
rect 8322 16923 8872 16936
rect 7638 16871 7704 16878
rect 8322 16871 8366 16923
rect 8806 16920 8872 16923
rect 9496 16934 9996 16964
rect 10030 16934 10046 16968
rect 11148 16968 11214 16984
rect 11148 16964 11164 16968
rect 9496 16921 10046 16934
rect 8806 16871 8872 16878
rect 4566 16830 4862 16871
rect 4566 16808 4626 16830
rect 4684 16808 4744 16830
rect 4802 16808 4862 16830
rect 4920 16862 5368 16871
rect 4920 16830 5318 16862
rect 4920 16808 4980 16830
rect 5038 16808 5098 16830
rect 5156 16829 5318 16830
rect 5156 16808 5216 16829
rect 5302 16828 5318 16829
rect 5352 16828 5368 16862
rect 5302 16812 5368 16828
rect 5734 16830 6030 16871
rect 5734 16810 5794 16830
rect 5852 16810 5912 16830
rect 5970 16810 6030 16830
rect 6088 16862 6536 16871
rect 6088 16830 6486 16862
rect 6088 16810 6148 16830
rect 6206 16810 6266 16830
rect 6324 16829 6486 16830
rect 6324 16810 6384 16829
rect 6470 16828 6486 16829
rect 6520 16828 6536 16862
rect 6470 16812 6536 16828
rect 6902 16830 7198 16871
rect 6902 16808 6962 16830
rect 7020 16808 7080 16830
rect 7138 16808 7198 16830
rect 7256 16862 7704 16871
rect 7256 16830 7654 16862
rect 7256 16808 7316 16830
rect 7374 16808 7434 16830
rect 7492 16829 7654 16830
rect 7492 16808 7552 16829
rect 7638 16828 7654 16829
rect 7688 16828 7704 16862
rect 7638 16812 7704 16828
rect 8070 16830 8366 16871
rect 8070 16810 8130 16830
rect 8188 16810 8248 16830
rect 8306 16810 8366 16830
rect 8424 16862 8872 16871
rect 9496 16869 9540 16921
rect 9980 16918 10046 16921
rect 10664 16934 11164 16964
rect 11198 16934 11214 16968
rect 49314 17291 49610 17327
rect 49314 17271 49374 17291
rect 49432 17271 49492 17291
rect 49550 17271 49610 17291
rect 49668 17291 49964 17327
rect 49668 17271 49728 17291
rect 49786 17271 49846 17291
rect 49904 17271 49964 17291
rect 50022 17292 50318 17328
rect 50022 17271 50082 17292
rect 50140 17271 50200 17292
rect 50258 17271 50318 17292
rect 42756 17049 42816 17075
rect 42874 17049 42934 17075
rect 12316 16968 12382 16984
rect 12316 16964 12332 16968
rect 10664 16921 11214 16934
rect 9980 16869 10046 16876
rect 10664 16869 10708 16921
rect 11148 16918 11214 16921
rect 11832 16934 12332 16964
rect 12366 16934 12382 16968
rect 42992 17043 43052 17075
rect 43110 17049 43170 17075
rect 43228 17049 43288 17075
rect 43346 17055 43406 17075
rect 43345 17049 43406 17055
rect 43464 17049 43524 17075
rect 43582 17049 43642 17075
rect 43700 17049 43760 17075
rect 55848 17296 56144 17332
rect 55848 17276 55908 17296
rect 55966 17276 56026 17296
rect 56084 17276 56144 17296
rect 56202 17296 56498 17332
rect 56202 17276 56262 17296
rect 56320 17276 56380 17296
rect 56438 17276 56498 17296
rect 56556 17297 56852 17333
rect 56556 17276 56616 17297
rect 56674 17276 56734 17297
rect 56792 17276 56852 17297
rect 70459 17373 70498 17431
rect 71329 17427 71396 17431
rect 62361 17299 62657 17335
rect 62361 17279 62421 17299
rect 62479 17279 62539 17299
rect 62597 17279 62657 17299
rect 62715 17299 63011 17335
rect 62715 17279 62775 17299
rect 62833 17279 62893 17299
rect 62951 17279 63011 17299
rect 63069 17300 63365 17336
rect 70459 17313 70513 17373
rect 70913 17313 70939 17373
rect 63069 17279 63129 17300
rect 63187 17279 63247 17300
rect 63305 17279 63365 17300
rect 42989 17027 43055 17043
rect 42989 16993 43005 17027
rect 43039 16993 43055 17027
rect 13484 16968 13550 16984
rect 42989 16977 43055 16993
rect 13484 16964 13500 16968
rect 11832 16921 12382 16934
rect 11148 16869 11214 16876
rect 11832 16869 11876 16921
rect 12316 16918 12382 16921
rect 13000 16934 13500 16964
rect 13534 16934 13550 16968
rect 13000 16921 13550 16934
rect 12316 16869 12382 16876
rect 13000 16869 13044 16921
rect 13484 16918 13550 16921
rect 13484 16869 13550 16876
rect 8424 16830 8822 16862
rect 8424 16810 8484 16830
rect 8542 16810 8602 16830
rect 8660 16829 8822 16830
rect 8660 16810 8720 16829
rect 8806 16828 8822 16829
rect 8856 16828 8872 16862
rect 8806 16812 8872 16828
rect 9244 16828 9540 16869
rect 4566 16382 4626 16408
rect 4684 16382 4744 16408
rect 4802 16208 4862 16408
rect 4920 16382 4980 16408
rect 5038 16382 5098 16408
rect 5156 16392 5216 16408
rect 5155 16303 5216 16392
rect 5734 16384 5794 16410
rect 5852 16384 5912 16410
rect 5155 16250 5306 16303
rect 4802 16157 5188 16208
rect 5007 16099 5073 16115
rect 5007 16065 5023 16099
rect 5057 16065 5073 16099
rect 5007 16049 5073 16065
rect 4491 16020 4551 16046
rect 4609 16020 4669 16046
rect 4727 16020 4787 16046
rect 5010 16026 5070 16049
rect 5128 16026 5188 16157
rect 5246 16026 5306 16250
rect 5970 16208 6030 16410
rect 6088 16384 6148 16410
rect 6206 16384 6266 16410
rect 6324 16392 6384 16410
rect 9244 16808 9304 16828
rect 9362 16808 9422 16828
rect 9480 16808 9540 16828
rect 9598 16860 10046 16869
rect 9598 16828 9996 16860
rect 9598 16808 9658 16828
rect 9716 16808 9776 16828
rect 9834 16827 9996 16828
rect 9834 16808 9894 16827
rect 9980 16826 9996 16827
rect 10030 16826 10046 16860
rect 9980 16810 10046 16826
rect 10412 16828 10708 16869
rect 6323 16303 6384 16392
rect 6902 16382 6962 16408
rect 7020 16382 7080 16408
rect 6323 16250 6474 16303
rect 5970 16157 6356 16208
rect 6175 16099 6241 16115
rect 6175 16065 6191 16099
rect 6225 16065 6241 16099
rect 6175 16049 6241 16065
rect 5659 16019 5719 16045
rect 5777 16019 5837 16045
rect 5895 16019 5955 16045
rect 6178 16026 6238 16049
rect 6296 16026 6356 16157
rect 6414 16026 6474 16250
rect 7138 16208 7198 16408
rect 7256 16382 7316 16408
rect 7374 16382 7434 16408
rect 7492 16392 7552 16408
rect 7491 16303 7552 16392
rect 8070 16384 8130 16410
rect 8188 16384 8248 16410
rect 7491 16250 7642 16303
rect 7138 16157 7524 16208
rect 7343 16099 7409 16115
rect 7343 16065 7359 16099
rect 7393 16065 7409 16099
rect 7343 16049 7409 16065
rect 4491 15794 4551 15820
rect 4609 15794 4669 15820
rect 4727 15794 4787 15820
rect 5010 15794 5070 15826
rect 5128 15800 5188 15826
rect 5246 15800 5306 15826
rect 6827 16019 6887 16045
rect 6945 16019 7005 16045
rect 7063 16019 7123 16045
rect 7346 16024 7406 16049
rect 7464 16024 7524 16157
rect 7582 16024 7642 16250
rect 8306 16208 8366 16410
rect 8424 16384 8484 16410
rect 8542 16384 8602 16410
rect 8660 16392 8720 16410
rect 10412 16806 10472 16828
rect 10530 16806 10590 16828
rect 10648 16806 10708 16828
rect 10766 16860 11214 16869
rect 10766 16828 11164 16860
rect 10766 16806 10826 16828
rect 10884 16806 10944 16828
rect 11002 16827 11164 16828
rect 11002 16806 11062 16827
rect 11148 16826 11164 16827
rect 11198 16826 11214 16860
rect 11148 16810 11214 16826
rect 11580 16828 11876 16869
rect 11580 16808 11640 16828
rect 11698 16808 11758 16828
rect 11816 16808 11876 16828
rect 11934 16860 12382 16869
rect 11934 16828 12332 16860
rect 11934 16808 11994 16828
rect 12052 16808 12112 16828
rect 12170 16827 12332 16828
rect 12170 16808 12230 16827
rect 12316 16826 12332 16827
rect 12366 16826 12382 16860
rect 12316 16810 12382 16826
rect 12748 16828 13044 16869
rect 12748 16808 12808 16828
rect 12866 16808 12926 16828
rect 12984 16808 13044 16828
rect 13102 16860 13550 16869
rect 13102 16828 13500 16860
rect 13102 16808 13162 16828
rect 13220 16808 13280 16828
rect 13338 16827 13500 16828
rect 13338 16808 13398 16827
rect 13484 16826 13500 16827
rect 13534 16826 13550 16860
rect 13484 16810 13550 16826
rect 8659 16303 8720 16392
rect 9244 16382 9304 16408
rect 9362 16382 9422 16408
rect 8659 16250 8810 16303
rect 8306 16157 8692 16208
rect 8511 16099 8577 16115
rect 8511 16065 8527 16099
rect 8561 16065 8577 16099
rect 8511 16049 8577 16065
rect 4491 15753 5070 15794
rect 5659 15794 5719 15819
rect 5777 15794 5837 15819
rect 5895 15794 5955 15819
rect 6178 15794 6238 15826
rect 6296 15800 6356 15826
rect 6414 15800 6474 15826
rect 7996 16020 8056 16046
rect 8114 16020 8174 16046
rect 8232 16020 8292 16046
rect 8514 16024 8574 16049
rect 8632 16024 8692 16157
rect 8750 16024 8810 16250
rect 9480 16206 9540 16408
rect 9598 16382 9658 16408
rect 9716 16382 9776 16408
rect 9834 16390 9894 16408
rect 39264 16858 39324 16884
rect 39382 16858 39442 16884
rect 39500 16858 39560 16884
rect 39618 16873 39914 16924
rect 39618 16858 39678 16873
rect 39736 16858 39796 16873
rect 39854 16858 39914 16873
rect 41162 16858 41222 16884
rect 41280 16858 41340 16884
rect 41398 16858 41458 16884
rect 41516 16873 41812 16924
rect 41516 16858 41576 16873
rect 41634 16858 41694 16873
rect 41752 16858 41812 16873
rect 43107 16910 43173 16926
rect 43107 16876 43123 16910
rect 43157 16876 43173 16910
rect 43107 16860 43173 16876
rect 38781 16675 39077 16726
rect 13849 16633 14145 16669
rect 13849 16613 13909 16633
rect 13967 16613 14027 16633
rect 14085 16613 14145 16633
rect 14203 16633 14499 16669
rect 14203 16613 14263 16633
rect 14321 16613 14381 16633
rect 14439 16613 14499 16633
rect 14557 16634 14853 16670
rect 14557 16613 14617 16634
rect 14675 16613 14735 16634
rect 14793 16613 14853 16634
rect 15297 16633 15593 16669
rect 15297 16613 15357 16633
rect 15415 16613 15475 16633
rect 15533 16613 15593 16633
rect 15651 16633 15947 16669
rect 15651 16613 15711 16633
rect 15769 16613 15829 16633
rect 15887 16613 15947 16633
rect 16005 16634 16301 16670
rect 16005 16613 16065 16634
rect 16123 16613 16183 16634
rect 16241 16613 16301 16634
rect 16795 16631 17091 16667
rect 16795 16611 16855 16631
rect 16913 16611 16973 16631
rect 17031 16611 17091 16631
rect 17149 16631 17445 16667
rect 17149 16611 17209 16631
rect 17267 16611 17327 16631
rect 17385 16611 17445 16631
rect 17503 16632 17799 16668
rect 17503 16611 17563 16632
rect 17621 16611 17681 16632
rect 17739 16611 17799 16632
rect 18243 16631 18539 16667
rect 18243 16611 18303 16631
rect 18361 16611 18421 16631
rect 18479 16611 18539 16631
rect 18597 16631 18893 16667
rect 18597 16611 18657 16631
rect 18715 16611 18775 16631
rect 18833 16611 18893 16631
rect 18951 16632 19247 16668
rect 18951 16611 19011 16632
rect 19069 16611 19129 16632
rect 19187 16611 19247 16632
rect 19763 16633 20059 16669
rect 19763 16613 19823 16633
rect 19881 16613 19941 16633
rect 19999 16613 20059 16633
rect 20117 16633 20413 16669
rect 20117 16613 20177 16633
rect 20235 16613 20295 16633
rect 20353 16613 20413 16633
rect 20471 16634 20767 16670
rect 20471 16613 20531 16634
rect 20589 16613 20649 16634
rect 20707 16613 20767 16634
rect 21211 16633 21507 16669
rect 21211 16613 21271 16633
rect 21329 16613 21389 16633
rect 21447 16613 21507 16633
rect 21565 16633 21861 16669
rect 21565 16613 21625 16633
rect 21683 16613 21743 16633
rect 21801 16613 21861 16633
rect 21919 16634 22215 16670
rect 21919 16613 21979 16634
rect 22037 16613 22097 16634
rect 22155 16613 22215 16634
rect 22709 16631 23005 16667
rect 9833 16301 9894 16390
rect 10412 16380 10472 16406
rect 10530 16380 10590 16406
rect 9833 16248 9984 16301
rect 9480 16155 9866 16206
rect 9685 16097 9751 16113
rect 9685 16063 9701 16097
rect 9735 16063 9751 16097
rect 9168 16024 9228 16050
rect 9286 16024 9346 16050
rect 9404 16024 9464 16050
rect 9685 16047 9751 16063
rect 9688 16024 9748 16047
rect 9806 16024 9866 16155
rect 9924 16024 9984 16248
rect 10648 16206 10708 16406
rect 10766 16380 10826 16406
rect 10884 16380 10944 16406
rect 11002 16390 11062 16406
rect 11001 16301 11062 16390
rect 11580 16382 11640 16408
rect 11698 16382 11758 16408
rect 11001 16248 11152 16301
rect 10648 16155 11034 16206
rect 10853 16097 10919 16113
rect 10853 16063 10869 16097
rect 10903 16063 10919 16097
rect 10337 16024 10397 16050
rect 10455 16024 10515 16050
rect 10573 16024 10633 16050
rect 10853 16047 10919 16063
rect 10856 16024 10916 16047
rect 10974 16024 11034 16155
rect 11092 16024 11152 16248
rect 11816 16206 11876 16408
rect 11934 16382 11994 16408
rect 12052 16382 12112 16408
rect 12170 16390 12230 16408
rect 12169 16301 12230 16390
rect 12748 16382 12808 16408
rect 12866 16382 12926 16408
rect 12169 16248 12320 16301
rect 11816 16155 12202 16206
rect 12021 16097 12087 16113
rect 12021 16063 12037 16097
rect 12071 16063 12087 16097
rect 11505 16024 11565 16050
rect 11623 16024 11683 16050
rect 11741 16024 11801 16050
rect 12021 16047 12087 16063
rect 12024 16024 12084 16047
rect 12142 16024 12202 16155
rect 12260 16024 12320 16248
rect 12984 16206 13044 16408
rect 13102 16382 13162 16408
rect 13220 16382 13280 16408
rect 13338 16390 13398 16408
rect 13337 16301 13398 16390
rect 13849 16387 13909 16413
rect 13967 16387 14027 16413
rect 14085 16381 14145 16413
rect 14203 16387 14263 16413
rect 14321 16387 14381 16413
rect 14439 16393 14499 16413
rect 14438 16387 14499 16393
rect 14557 16387 14617 16413
rect 14675 16387 14735 16413
rect 14793 16387 14853 16413
rect 15297 16387 15357 16413
rect 15415 16387 15475 16413
rect 14082 16365 14148 16381
rect 14082 16331 14098 16365
rect 14132 16331 14148 16365
rect 14082 16315 14148 16331
rect 13337 16248 13488 16301
rect 12984 16155 13370 16206
rect 13189 16097 13255 16113
rect 13189 16063 13205 16097
rect 13239 16063 13255 16097
rect 13189 16047 13255 16063
rect 5659 15753 6238 15794
rect 6827 15794 6887 15819
rect 6945 15794 7005 15819
rect 7063 15794 7123 15819
rect 7346 15794 7406 15824
rect 7464 15798 7524 15824
rect 7582 15798 7642 15824
rect 12672 16018 12732 16044
rect 12790 16018 12850 16044
rect 12908 16018 12968 16044
rect 13192 16022 13252 16047
rect 13310 16022 13370 16155
rect 13428 16022 13488 16248
rect 14200 16248 14266 16264
rect 14200 16214 14216 16248
rect 14250 16214 14266 16248
rect 14200 16198 14266 16214
rect 14203 16176 14263 16198
rect 14438 16176 14498 16387
rect 14558 16202 14616 16387
rect 15533 16381 15593 16413
rect 15651 16387 15711 16413
rect 15769 16387 15829 16413
rect 15887 16393 15947 16413
rect 15886 16387 15947 16393
rect 16005 16387 16065 16413
rect 16123 16387 16183 16413
rect 16241 16387 16301 16413
rect 22709 16611 22769 16631
rect 22827 16611 22887 16631
rect 22945 16611 23005 16631
rect 23063 16631 23359 16667
rect 23063 16611 23123 16631
rect 23181 16611 23241 16631
rect 23299 16611 23359 16631
rect 23417 16632 23713 16668
rect 23417 16611 23477 16632
rect 23535 16611 23595 16632
rect 23653 16611 23713 16632
rect 24157 16631 24453 16667
rect 24157 16611 24217 16631
rect 24275 16611 24335 16631
rect 24393 16611 24453 16631
rect 24511 16631 24807 16667
rect 24511 16611 24571 16631
rect 24629 16611 24689 16631
rect 24747 16611 24807 16631
rect 24865 16632 25161 16668
rect 38781 16658 38841 16675
rect 38899 16658 38959 16675
rect 39017 16658 39077 16675
rect 24865 16611 24925 16632
rect 24983 16611 25043 16632
rect 25101 16611 25161 16632
rect 15530 16365 15596 16381
rect 15530 16331 15546 16365
rect 15580 16331 15596 16365
rect 15530 16315 15596 16331
rect 14556 16176 14616 16202
rect 15648 16248 15714 16264
rect 15648 16214 15664 16248
rect 15698 16214 15714 16248
rect 15648 16198 15714 16214
rect 15651 16176 15711 16198
rect 15886 16176 15946 16387
rect 16006 16202 16064 16387
rect 16795 16385 16855 16411
rect 16913 16385 16973 16411
rect 17031 16379 17091 16411
rect 17149 16385 17209 16411
rect 17267 16385 17327 16411
rect 17385 16391 17445 16411
rect 17384 16385 17445 16391
rect 17503 16385 17563 16411
rect 17621 16385 17681 16411
rect 17739 16385 17799 16411
rect 18243 16385 18303 16411
rect 18361 16385 18421 16411
rect 17028 16363 17094 16379
rect 17028 16329 17044 16363
rect 17078 16329 17094 16363
rect 17028 16313 17094 16329
rect 16004 16176 16064 16202
rect 17146 16246 17212 16262
rect 17146 16212 17162 16246
rect 17196 16212 17212 16246
rect 17146 16196 17212 16212
rect 6827 15753 7406 15794
rect 7996 15794 8056 15820
rect 8114 15794 8174 15820
rect 8232 15794 8292 15820
rect 8514 15794 8574 15824
rect 8632 15798 8692 15824
rect 8750 15798 8810 15824
rect 9168 15798 9228 15824
rect 7996 15788 8574 15794
rect 7995 15753 8574 15788
rect 9169 15792 9228 15798
rect 9286 15792 9346 15824
rect 9404 15792 9464 15824
rect 9688 15792 9748 15824
rect 9806 15798 9866 15824
rect 9924 15798 9984 15824
rect 9169 15751 9748 15792
rect 10337 15792 10397 15824
rect 10455 15792 10515 15824
rect 10573 15792 10633 15824
rect 10856 15792 10916 15824
rect 10974 15798 11034 15824
rect 11092 15798 11152 15824
rect 10337 15751 10916 15792
rect 11505 15792 11565 15824
rect 11623 15792 11683 15824
rect 11741 15792 11801 15824
rect 12024 15792 12084 15824
rect 12142 15798 12202 15824
rect 12260 15798 12320 15824
rect 14203 15950 14263 15976
rect 12672 15792 12732 15818
rect 12790 15792 12850 15818
rect 12908 15792 12968 15818
rect 13192 15792 13252 15822
rect 13310 15796 13370 15822
rect 13428 15796 13488 15822
rect 11505 15751 12084 15792
rect 12673 15751 13252 15792
rect 15651 15950 15711 15976
rect 17149 16174 17209 16196
rect 17384 16174 17444 16385
rect 17504 16200 17562 16385
rect 18479 16379 18539 16411
rect 18597 16385 18657 16411
rect 18715 16385 18775 16411
rect 18833 16391 18893 16411
rect 18832 16385 18893 16391
rect 18951 16385 19011 16411
rect 19069 16385 19129 16411
rect 19187 16385 19247 16411
rect 19763 16387 19823 16413
rect 19881 16387 19941 16413
rect 18476 16363 18542 16379
rect 18476 16329 18492 16363
rect 18526 16329 18542 16363
rect 18476 16313 18542 16329
rect 17502 16174 17562 16200
rect 18594 16246 18660 16262
rect 18594 16212 18610 16246
rect 18644 16212 18660 16246
rect 18594 16196 18660 16212
rect 18597 16174 18657 16196
rect 18832 16174 18892 16385
rect 18952 16200 19010 16385
rect 19999 16381 20059 16413
rect 20117 16387 20177 16413
rect 20235 16387 20295 16413
rect 20353 16393 20413 16413
rect 20352 16387 20413 16393
rect 20471 16387 20531 16413
rect 20589 16387 20649 16413
rect 20707 16387 20767 16413
rect 21211 16387 21271 16413
rect 21329 16387 21389 16413
rect 19996 16365 20062 16381
rect 19996 16331 20012 16365
rect 20046 16331 20062 16365
rect 19996 16315 20062 16331
rect 18950 16174 19010 16200
rect 20114 16248 20180 16264
rect 20114 16214 20130 16248
rect 20164 16214 20180 16248
rect 20114 16198 20180 16214
rect 20117 16176 20177 16198
rect 20352 16176 20412 16387
rect 20472 16202 20530 16387
rect 21447 16381 21507 16413
rect 21565 16387 21625 16413
rect 21683 16387 21743 16413
rect 21801 16393 21861 16413
rect 21800 16387 21861 16393
rect 21919 16387 21979 16413
rect 22037 16387 22097 16413
rect 22155 16387 22215 16413
rect 40102 16658 40162 16684
rect 40220 16658 40280 16684
rect 40338 16658 40398 16684
rect 40679 16675 40975 16726
rect 40679 16658 40739 16675
rect 40797 16658 40857 16675
rect 40915 16658 40975 16675
rect 43110 16838 43170 16860
rect 43345 16838 43405 17049
rect 43465 16864 43523 17049
rect 49314 17045 49374 17071
rect 49432 17045 49492 17071
rect 49550 17039 49610 17071
rect 49668 17045 49728 17071
rect 49786 17045 49846 17071
rect 49904 17051 49964 17071
rect 49903 17045 49964 17051
rect 50022 17045 50082 17071
rect 50140 17045 50200 17071
rect 50258 17045 50318 17071
rect 55848 17050 55908 17076
rect 55966 17050 56026 17076
rect 49547 17023 49613 17039
rect 49547 16989 49563 17023
rect 49597 16989 49613 17023
rect 49547 16973 49613 16989
rect 43463 16838 43523 16864
rect 45822 16854 45882 16880
rect 45940 16854 46000 16880
rect 46058 16854 46118 16880
rect 46176 16869 46472 16920
rect 46176 16854 46236 16869
rect 46294 16854 46354 16869
rect 46412 16854 46472 16869
rect 47720 16854 47780 16880
rect 47838 16854 47898 16880
rect 47956 16854 48016 16880
rect 48074 16869 48370 16920
rect 48074 16854 48134 16869
rect 48192 16854 48252 16869
rect 48310 16854 48370 16869
rect 49665 16906 49731 16922
rect 49665 16872 49681 16906
rect 49715 16872 49731 16906
rect 49665 16856 49731 16872
rect 42000 16658 42060 16684
rect 42118 16658 42178 16684
rect 42236 16658 42296 16684
rect 43110 16612 43170 16638
rect 38781 16432 38841 16458
rect 38899 16439 38959 16458
rect 39017 16439 39077 16458
rect 39264 16439 39324 16458
rect 39382 16439 39442 16458
rect 39500 16439 39560 16458
rect 38899 16432 38975 16439
rect 21444 16365 21510 16381
rect 21444 16331 21460 16365
rect 21494 16331 21510 16365
rect 21444 16315 21510 16331
rect 20470 16176 20530 16202
rect 21562 16248 21628 16264
rect 21562 16214 21578 16248
rect 21612 16214 21628 16248
rect 21562 16198 21628 16214
rect 21565 16176 21625 16198
rect 21800 16176 21860 16387
rect 21920 16202 21978 16387
rect 22709 16385 22769 16411
rect 22827 16385 22887 16411
rect 22945 16379 23005 16411
rect 23063 16385 23123 16411
rect 23181 16385 23241 16411
rect 23299 16391 23359 16411
rect 23298 16385 23359 16391
rect 23417 16385 23477 16411
rect 23535 16385 23595 16411
rect 23653 16385 23713 16411
rect 24157 16385 24217 16411
rect 24275 16385 24335 16411
rect 22942 16363 23008 16379
rect 22942 16329 22958 16363
rect 22992 16329 23008 16363
rect 22942 16313 23008 16329
rect 21918 16176 21978 16202
rect 23060 16246 23126 16262
rect 23060 16212 23076 16246
rect 23110 16212 23126 16246
rect 23060 16196 23126 16212
rect 17149 15948 17209 15974
rect 14438 15754 14498 15776
rect 14556 15754 14616 15776
rect 15886 15754 15946 15776
rect 16004 15754 16064 15776
rect 18597 15948 18657 15974
rect 20117 15950 20177 15976
rect 21565 15950 21625 15976
rect 23063 16174 23123 16196
rect 23298 16174 23358 16385
rect 23418 16200 23476 16385
rect 24393 16379 24453 16411
rect 24511 16385 24571 16411
rect 24629 16385 24689 16411
rect 24747 16391 24807 16411
rect 24746 16385 24807 16391
rect 24865 16385 24925 16411
rect 24983 16385 25043 16411
rect 25101 16385 25161 16411
rect 38900 16388 38975 16432
rect 39017 16388 39560 16439
rect 39618 16432 39678 16458
rect 39736 16432 39796 16458
rect 39854 16441 39914 16458
rect 40102 16441 40162 16458
rect 40220 16441 40280 16458
rect 40338 16441 40398 16458
rect 39854 16390 40398 16441
rect 40679 16432 40739 16458
rect 40797 16439 40857 16458
rect 40915 16439 40975 16458
rect 41162 16439 41222 16458
rect 41280 16439 41340 16458
rect 41398 16439 41458 16458
rect 40797 16432 40873 16439
rect 24390 16363 24456 16379
rect 24390 16329 24406 16363
rect 24440 16329 24456 16363
rect 24390 16313 24456 16329
rect 23416 16174 23476 16200
rect 24508 16246 24574 16262
rect 24508 16212 24524 16246
rect 24558 16212 24574 16246
rect 24508 16196 24574 16212
rect 24511 16174 24571 16196
rect 24746 16174 24806 16385
rect 24866 16200 24924 16385
rect 38915 16235 38975 16388
rect 24864 16174 24924 16200
rect 38721 16211 38975 16235
rect 38721 16177 38737 16211
rect 38771 16177 38975 16211
rect 23063 15948 23123 15974
rect 14435 15738 14501 15754
rect 14435 15704 14451 15738
rect 14485 15704 14501 15738
rect 14435 15688 14501 15704
rect 14553 15738 14619 15754
rect 14553 15704 14569 15738
rect 14603 15704 14619 15738
rect 14553 15688 14619 15704
rect 15883 15738 15949 15754
rect 15883 15704 15899 15738
rect 15933 15704 15949 15738
rect 15883 15688 15949 15704
rect 16001 15738 16067 15754
rect 17384 15752 17444 15774
rect 17502 15752 17562 15774
rect 18832 15752 18892 15774
rect 18950 15752 19010 15774
rect 20352 15754 20412 15776
rect 20470 15754 20530 15776
rect 21800 15754 21860 15776
rect 21918 15754 21978 15776
rect 24511 15948 24571 15974
rect 38721 16161 38975 16177
rect 39321 16189 39617 16249
rect 39321 16165 39381 16189
rect 39439 16165 39499 16189
rect 39557 16165 39617 16189
rect 39675 16188 39971 16248
rect 39675 16165 39735 16188
rect 39793 16165 39853 16188
rect 39911 16165 39971 16188
rect 16001 15704 16017 15738
rect 16051 15704 16067 15738
rect 16001 15688 16067 15704
rect 17381 15736 17447 15752
rect 17381 15702 17397 15736
rect 17431 15702 17447 15736
rect 17381 15686 17447 15702
rect 17499 15736 17565 15752
rect 17499 15702 17515 15736
rect 17549 15702 17565 15736
rect 17499 15686 17565 15702
rect 18829 15736 18895 15752
rect 18829 15702 18845 15736
rect 18879 15702 18895 15736
rect 18829 15686 18895 15702
rect 18947 15736 19013 15752
rect 18947 15702 18963 15736
rect 18997 15702 19013 15736
rect 18947 15686 19013 15702
rect 20349 15738 20415 15754
rect 20349 15704 20365 15738
rect 20399 15704 20415 15738
rect 20349 15688 20415 15704
rect 20467 15738 20533 15754
rect 20467 15704 20483 15738
rect 20517 15704 20533 15738
rect 20467 15688 20533 15704
rect 21797 15738 21863 15754
rect 21797 15704 21813 15738
rect 21847 15704 21863 15738
rect 21797 15688 21863 15704
rect 21915 15738 21981 15754
rect 23298 15752 23358 15774
rect 23416 15752 23476 15774
rect 24746 15752 24806 15774
rect 24864 15752 24924 15774
rect 21915 15704 21931 15738
rect 21965 15704 21981 15738
rect 21915 15688 21981 15704
rect 23295 15736 23361 15752
rect 23295 15702 23311 15736
rect 23345 15702 23361 15736
rect 23295 15686 23361 15702
rect 23413 15736 23479 15752
rect 23413 15702 23429 15736
rect 23463 15702 23479 15736
rect 23413 15686 23479 15702
rect 24743 15736 24809 15752
rect 24743 15702 24759 15736
rect 24793 15702 24809 15736
rect 24743 15686 24809 15702
rect 24861 15736 24927 15752
rect 24861 15702 24877 15736
rect 24911 15702 24927 15736
rect 24861 15686 24927 15702
rect 38915 15537 38975 16161
rect 39321 15739 39381 15765
rect 39291 15599 39358 15606
rect 39291 15598 39364 15599
rect 39439 15598 39499 15765
rect 39557 15739 39617 15765
rect 39675 15739 39735 15765
rect 39291 15590 39499 15598
rect 39291 15556 39307 15590
rect 39341 15556 39499 15590
rect 39291 15540 39499 15556
rect 39302 15539 39499 15540
rect 38915 15521 39065 15537
rect 38915 15487 39015 15521
rect 39049 15487 39065 15521
rect 38915 15471 39065 15487
rect 38915 15433 38975 15471
rect 39439 15433 39499 15539
rect 39793 15598 39853 15765
rect 39911 15739 39971 15765
rect 40213 15732 40273 16390
rect 40798 16388 40873 16432
rect 40915 16388 41458 16439
rect 41516 16432 41576 16458
rect 41634 16432 41694 16458
rect 41752 16441 41812 16458
rect 42000 16441 42060 16458
rect 42118 16441 42178 16458
rect 42236 16441 42296 16458
rect 41752 16390 42296 16441
rect 45339 16671 45635 16722
rect 45339 16654 45399 16671
rect 45457 16654 45517 16671
rect 45575 16654 45635 16671
rect 46660 16654 46720 16680
rect 46778 16654 46838 16680
rect 46896 16654 46956 16680
rect 47237 16671 47533 16722
rect 47237 16654 47297 16671
rect 47355 16654 47415 16671
rect 47473 16654 47533 16671
rect 49668 16834 49728 16856
rect 49903 16834 49963 17045
rect 50023 16860 50081 17045
rect 56084 17044 56144 17076
rect 56202 17050 56262 17076
rect 56320 17050 56380 17076
rect 56438 17056 56498 17076
rect 56437 17050 56498 17056
rect 56556 17050 56616 17076
rect 56674 17050 56734 17076
rect 56792 17050 56852 17076
rect 62361 17053 62421 17079
rect 62479 17053 62539 17079
rect 56081 17028 56147 17044
rect 56081 16994 56097 17028
rect 56131 16994 56147 17028
rect 56081 16978 56147 16994
rect 50021 16834 50081 16860
rect 52356 16859 52416 16885
rect 52474 16859 52534 16885
rect 52592 16859 52652 16885
rect 52710 16874 53006 16925
rect 52710 16859 52770 16874
rect 52828 16859 52888 16874
rect 52946 16859 53006 16874
rect 54254 16859 54314 16885
rect 54372 16859 54432 16885
rect 54490 16859 54550 16885
rect 54608 16874 54904 16925
rect 54608 16859 54668 16874
rect 54726 16859 54786 16874
rect 54844 16859 54904 16874
rect 56199 16911 56265 16927
rect 56199 16877 56215 16911
rect 56249 16877 56265 16911
rect 56199 16861 56265 16877
rect 48558 16654 48618 16680
rect 48676 16654 48736 16680
rect 48794 16654 48854 16680
rect 49668 16608 49728 16634
rect 43345 16422 43405 16438
rect 40206 15716 40273 15732
rect 40206 15682 40223 15716
rect 40257 15682 40273 15716
rect 40206 15666 40273 15682
rect 39936 15598 40003 15605
rect 39793 15589 40003 15598
rect 39793 15555 39953 15589
rect 39987 15555 40003 15589
rect 39793 15539 40003 15555
rect 39553 15506 39619 15521
rect 39553 15472 39569 15506
rect 39603 15472 39619 15506
rect 39553 15456 39619 15472
rect 39671 15505 39737 15521
rect 39671 15471 39687 15505
rect 39721 15471 39737 15505
rect 39557 15433 39617 15456
rect 39671 15455 39737 15471
rect 39675 15433 39735 15455
rect 39793 15433 39853 15539
rect 40213 15538 40273 15666
rect 40122 15522 40273 15538
rect 40122 15488 40138 15522
rect 40172 15488 40273 15522
rect 40122 15472 40273 15488
rect 40213 15433 40273 15472
rect 40813 16268 40873 16388
rect 42111 16309 42171 16390
rect 43337 16400 43411 16422
rect 43463 16416 43523 16438
rect 45339 16428 45399 16454
rect 45457 16435 45517 16454
rect 45575 16435 45635 16454
rect 45822 16435 45882 16454
rect 45940 16435 46000 16454
rect 46058 16435 46118 16454
rect 45457 16428 45533 16435
rect 43337 16366 43358 16400
rect 43392 16366 43411 16400
rect 43337 16309 43411 16366
rect 43460 16400 43526 16416
rect 43460 16366 43476 16400
rect 43510 16366 43526 16400
rect 45458 16384 45533 16428
rect 45575 16384 46118 16435
rect 46176 16428 46236 16454
rect 46294 16428 46354 16454
rect 46412 16437 46472 16454
rect 46660 16437 46720 16454
rect 46778 16437 46838 16454
rect 46896 16437 46956 16454
rect 46412 16386 46956 16437
rect 47237 16428 47297 16454
rect 47355 16435 47415 16454
rect 47473 16435 47533 16454
rect 47720 16435 47780 16454
rect 47838 16435 47898 16454
rect 47956 16435 48016 16454
rect 47355 16428 47431 16435
rect 43460 16350 43526 16366
rect 42111 16284 43411 16309
rect 40813 16248 40874 16268
rect 40813 16232 40893 16248
rect 40813 16198 40844 16232
rect 40878 16198 40893 16232
rect 40813 16182 40893 16198
rect 41219 16189 41515 16249
rect 40813 16159 40874 16182
rect 41219 16165 41279 16189
rect 41337 16165 41397 16189
rect 41455 16165 41515 16189
rect 41573 16188 41869 16248
rect 41573 16165 41633 16188
rect 41691 16165 41751 16188
rect 41809 16165 41869 16188
rect 42111 16236 43412 16284
rect 40813 16013 40873 16159
rect 40813 15840 40874 16013
rect 40813 15537 40873 15840
rect 41219 15739 41279 15765
rect 41187 15598 41254 15605
rect 41337 15598 41397 15765
rect 41455 15739 41515 15765
rect 41573 15739 41633 15765
rect 41187 15589 41397 15598
rect 41187 15555 41203 15589
rect 41237 15555 41397 15589
rect 41187 15539 41397 15555
rect 40813 15521 40963 15537
rect 40813 15487 40913 15521
rect 40947 15487 40963 15521
rect 40813 15471 40963 15487
rect 40813 15433 40873 15471
rect 41337 15433 41397 15539
rect 41691 15598 41751 15765
rect 41809 15739 41869 15765
rect 41834 15598 41901 15605
rect 41691 15589 41901 15598
rect 41691 15555 41851 15589
rect 41885 15555 41901 15589
rect 41691 15539 41901 15555
rect 41451 15506 41517 15521
rect 41451 15472 41467 15506
rect 41501 15472 41517 15506
rect 41451 15456 41517 15472
rect 41569 15505 41635 15521
rect 41569 15471 41585 15505
rect 41619 15471 41635 15505
rect 41455 15433 41515 15456
rect 41569 15455 41635 15471
rect 41573 15433 41633 15455
rect 41691 15433 41751 15539
rect 42111 15538 42171 16236
rect 45473 16231 45533 16384
rect 45279 16207 45533 16231
rect 45279 16173 45295 16207
rect 45329 16173 45533 16207
rect 45279 16157 45533 16173
rect 45879 16185 46175 16245
rect 45879 16161 45939 16185
rect 45997 16161 46057 16185
rect 46115 16161 46175 16185
rect 46233 16184 46529 16244
rect 46233 16161 46293 16184
rect 46351 16161 46411 16184
rect 46469 16161 46529 16184
rect 42761 15691 43057 15727
rect 42761 15671 42821 15691
rect 42879 15671 42939 15691
rect 42997 15671 43057 15691
rect 43115 15691 43411 15727
rect 43115 15671 43175 15691
rect 43233 15671 43293 15691
rect 43351 15671 43411 15691
rect 43469 15692 43765 15728
rect 43469 15671 43529 15692
rect 43587 15671 43647 15692
rect 43705 15671 43765 15692
rect 42020 15522 42171 15538
rect 42020 15488 42036 15522
rect 42070 15488 42171 15522
rect 42020 15472 42171 15488
rect 42111 15433 42171 15472
rect 45473 15533 45533 16157
rect 45879 15735 45939 15761
rect 45849 15595 45916 15602
rect 45849 15594 45922 15595
rect 45997 15594 46057 15761
rect 46115 15735 46175 15761
rect 46233 15735 46293 15761
rect 45849 15586 46057 15594
rect 45849 15552 45865 15586
rect 45899 15552 46057 15586
rect 45849 15536 46057 15552
rect 45860 15535 46057 15536
rect 45473 15517 45623 15533
rect 45473 15483 45573 15517
rect 45607 15483 45623 15517
rect 42761 15445 42821 15471
rect 42879 15445 42939 15471
rect 42997 15439 43057 15471
rect 43115 15445 43175 15471
rect 43233 15445 43293 15471
rect 43351 15451 43411 15471
rect 43350 15445 43411 15451
rect 43469 15445 43529 15471
rect 43587 15445 43647 15471
rect 43705 15445 43765 15471
rect 45473 15467 45623 15483
rect 38915 15207 38975 15233
rect 40213 15207 40273 15233
rect 40813 15207 40873 15233
rect 42994 15423 43060 15439
rect 42994 15389 43010 15423
rect 43044 15389 43060 15423
rect 42994 15373 43060 15389
rect 43112 15306 43178 15322
rect 43112 15272 43128 15306
rect 43162 15272 43178 15306
rect 43112 15256 43178 15272
rect 43115 15234 43175 15256
rect 43350 15234 43410 15445
rect 43470 15260 43528 15445
rect 45473 15429 45533 15467
rect 45997 15429 46057 15535
rect 46351 15594 46411 15761
rect 46469 15735 46529 15761
rect 46771 15728 46831 16386
rect 47356 16384 47431 16428
rect 47473 16384 48016 16435
rect 48074 16428 48134 16454
rect 48192 16428 48252 16454
rect 48310 16437 48370 16454
rect 48558 16437 48618 16454
rect 48676 16437 48736 16454
rect 48794 16437 48854 16454
rect 48310 16386 48854 16437
rect 51873 16676 52169 16727
rect 51873 16659 51933 16676
rect 51991 16659 52051 16676
rect 52109 16659 52169 16676
rect 53194 16659 53254 16685
rect 53312 16659 53372 16685
rect 53430 16659 53490 16685
rect 53771 16676 54067 16727
rect 53771 16659 53831 16676
rect 53889 16659 53949 16676
rect 54007 16659 54067 16676
rect 56202 16839 56262 16861
rect 56437 16839 56497 17050
rect 56557 16865 56615 17050
rect 62597 17047 62657 17079
rect 62715 17053 62775 17079
rect 62833 17053 62893 17079
rect 62951 17059 63011 17079
rect 62950 17053 63011 17059
rect 63069 17053 63129 17079
rect 63187 17053 63247 17079
rect 63305 17053 63365 17079
rect 70459 17076 70513 17136
rect 70913 17076 70939 17136
rect 62594 17031 62660 17047
rect 62594 16997 62610 17031
rect 62644 16997 62660 17031
rect 62594 16981 62660 16997
rect 56555 16839 56615 16865
rect 58869 16862 58929 16888
rect 58987 16862 59047 16888
rect 59105 16862 59165 16888
rect 59223 16877 59519 16928
rect 59223 16862 59283 16877
rect 59341 16862 59401 16877
rect 59459 16862 59519 16877
rect 60767 16862 60827 16888
rect 60885 16862 60945 16888
rect 61003 16862 61063 16888
rect 61121 16877 61417 16928
rect 61121 16862 61181 16877
rect 61239 16862 61299 16877
rect 61357 16862 61417 16877
rect 62712 16914 62778 16930
rect 62712 16880 62728 16914
rect 62762 16880 62778 16914
rect 62712 16864 62778 16880
rect 55092 16659 55152 16685
rect 55210 16659 55270 16685
rect 55328 16659 55388 16685
rect 56202 16613 56262 16639
rect 49903 16418 49963 16434
rect 46764 15712 46831 15728
rect 46764 15678 46781 15712
rect 46815 15678 46831 15712
rect 46764 15662 46831 15678
rect 46494 15594 46561 15601
rect 46351 15585 46561 15594
rect 46351 15551 46511 15585
rect 46545 15551 46561 15585
rect 46351 15535 46561 15551
rect 46111 15502 46177 15517
rect 46111 15468 46127 15502
rect 46161 15468 46177 15502
rect 46111 15452 46177 15468
rect 46229 15501 46295 15517
rect 46229 15467 46245 15501
rect 46279 15467 46295 15501
rect 46115 15429 46175 15452
rect 46229 15451 46295 15467
rect 46233 15429 46293 15451
rect 46351 15429 46411 15535
rect 46771 15534 46831 15662
rect 46680 15518 46831 15534
rect 46680 15484 46696 15518
rect 46730 15484 46831 15518
rect 46680 15468 46831 15484
rect 46771 15429 46831 15468
rect 47371 16264 47431 16384
rect 48669 16305 48729 16386
rect 49895 16396 49969 16418
rect 50021 16412 50081 16434
rect 51873 16433 51933 16459
rect 51991 16440 52051 16459
rect 52109 16440 52169 16459
rect 52356 16440 52416 16459
rect 52474 16440 52534 16459
rect 52592 16440 52652 16459
rect 51991 16433 52067 16440
rect 49895 16362 49916 16396
rect 49950 16362 49969 16396
rect 49895 16305 49969 16362
rect 50018 16396 50084 16412
rect 50018 16362 50034 16396
rect 50068 16362 50084 16396
rect 51992 16389 52067 16433
rect 52109 16389 52652 16440
rect 52710 16433 52770 16459
rect 52828 16433 52888 16459
rect 52946 16442 53006 16459
rect 53194 16442 53254 16459
rect 53312 16442 53372 16459
rect 53430 16442 53490 16459
rect 52946 16391 53490 16442
rect 53771 16433 53831 16459
rect 53889 16440 53949 16459
rect 54007 16440 54067 16459
rect 54254 16440 54314 16459
rect 54372 16440 54432 16459
rect 54490 16440 54550 16459
rect 53889 16433 53965 16440
rect 50018 16346 50084 16362
rect 48669 16280 49969 16305
rect 47371 16244 47432 16264
rect 47371 16228 47451 16244
rect 47371 16194 47402 16228
rect 47436 16194 47451 16228
rect 47371 16178 47451 16194
rect 47777 16185 48073 16245
rect 47371 16155 47432 16178
rect 47777 16161 47837 16185
rect 47895 16161 47955 16185
rect 48013 16161 48073 16185
rect 48131 16184 48427 16244
rect 48131 16161 48191 16184
rect 48249 16161 48309 16184
rect 48367 16161 48427 16184
rect 48669 16232 49970 16280
rect 52007 16236 52067 16389
rect 47371 16009 47431 16155
rect 47371 15836 47432 16009
rect 47371 15533 47431 15836
rect 47777 15735 47837 15761
rect 47745 15594 47812 15601
rect 47895 15594 47955 15761
rect 48013 15735 48073 15761
rect 48131 15735 48191 15761
rect 47745 15585 47955 15594
rect 47745 15551 47761 15585
rect 47795 15551 47955 15585
rect 47745 15535 47955 15551
rect 47371 15517 47521 15533
rect 47371 15483 47471 15517
rect 47505 15483 47521 15517
rect 47371 15467 47521 15483
rect 47371 15429 47431 15467
rect 47895 15429 47955 15535
rect 48249 15594 48309 15761
rect 48367 15735 48427 15761
rect 48392 15594 48459 15601
rect 48249 15585 48459 15594
rect 48249 15551 48409 15585
rect 48443 15551 48459 15585
rect 48249 15535 48459 15551
rect 48009 15502 48075 15517
rect 48009 15468 48025 15502
rect 48059 15468 48075 15502
rect 48009 15452 48075 15468
rect 48127 15501 48193 15517
rect 48127 15467 48143 15501
rect 48177 15467 48193 15501
rect 48013 15429 48073 15452
rect 48127 15451 48193 15467
rect 48131 15429 48191 15451
rect 48249 15429 48309 15535
rect 48669 15534 48729 16232
rect 51813 16212 52067 16236
rect 51813 16178 51829 16212
rect 51863 16178 52067 16212
rect 51813 16162 52067 16178
rect 52413 16190 52709 16250
rect 52413 16166 52473 16190
rect 52531 16166 52591 16190
rect 52649 16166 52709 16190
rect 52767 16189 53063 16249
rect 52767 16166 52827 16189
rect 52885 16166 52945 16189
rect 53003 16166 53063 16189
rect 49319 15687 49615 15723
rect 49319 15667 49379 15687
rect 49437 15667 49497 15687
rect 49555 15667 49615 15687
rect 49673 15687 49969 15723
rect 49673 15667 49733 15687
rect 49791 15667 49851 15687
rect 49909 15667 49969 15687
rect 50027 15688 50323 15724
rect 50027 15667 50087 15688
rect 50145 15667 50205 15688
rect 50263 15667 50323 15688
rect 48578 15518 48729 15534
rect 48578 15484 48594 15518
rect 48628 15484 48729 15518
rect 48578 15468 48729 15484
rect 48669 15429 48729 15468
rect 52007 15538 52067 16162
rect 52413 15740 52473 15766
rect 52383 15600 52450 15607
rect 52383 15599 52456 15600
rect 52531 15599 52591 15766
rect 52649 15740 52709 15766
rect 52767 15740 52827 15766
rect 52383 15591 52591 15599
rect 52383 15557 52399 15591
rect 52433 15557 52591 15591
rect 52383 15541 52591 15557
rect 52394 15540 52591 15541
rect 52007 15522 52157 15538
rect 52007 15488 52107 15522
rect 52141 15488 52157 15522
rect 52007 15472 52157 15488
rect 49319 15441 49379 15467
rect 49437 15441 49497 15467
rect 49555 15435 49615 15467
rect 49673 15441 49733 15467
rect 49791 15441 49851 15467
rect 49909 15447 49969 15467
rect 49908 15441 49969 15447
rect 50027 15441 50087 15467
rect 50145 15441 50205 15467
rect 50263 15441 50323 15467
rect 43468 15234 43528 15260
rect 42111 15207 42171 15233
rect 39439 15007 39499 15033
rect 39557 15007 39617 15033
rect 39675 15007 39735 15033
rect 39793 15007 39853 15033
rect 41337 15007 41397 15033
rect 41455 15007 41515 15033
rect 41573 15007 41633 15033
rect 41691 15007 41751 15033
rect 43115 15008 43175 15034
rect 1029 14873 1325 14912
rect 1029 14858 1089 14873
rect 1147 14858 1207 14873
rect 1265 14858 1325 14873
rect 1502 14873 1798 14912
rect 1502 14858 1562 14873
rect 1620 14858 1680 14873
rect 1738 14858 1798 14873
rect 1856 14873 2152 14912
rect 1856 14858 1916 14873
rect 1974 14858 2034 14873
rect 2092 14858 2152 14873
rect 2323 14873 2619 14912
rect 2323 14858 2383 14873
rect 2441 14858 2501 14873
rect 2559 14858 2619 14873
rect 4173 14873 4469 14912
rect 4173 14858 4233 14873
rect 4291 14858 4351 14873
rect 4409 14858 4469 14873
rect 4646 14873 4942 14912
rect 4646 14858 4706 14873
rect 4764 14858 4824 14873
rect 4882 14858 4942 14873
rect 5000 14873 5296 14912
rect 5000 14858 5060 14873
rect 5118 14858 5178 14873
rect 5236 14858 5296 14873
rect 5467 14873 5763 14912
rect 5467 14858 5527 14873
rect 5585 14858 5645 14873
rect 5703 14858 5763 14873
rect 7305 14869 7601 14908
rect 556 14674 852 14713
rect 556 14658 616 14674
rect 674 14658 734 14674
rect 792 14658 852 14674
rect 2764 14674 3060 14713
rect 2764 14658 2824 14674
rect 2882 14658 2942 14674
rect 3000 14658 3060 14674
rect 3700 14674 3996 14713
rect 3700 14658 3760 14674
rect 3818 14658 3878 14674
rect 3936 14658 3996 14674
rect 7305 14854 7365 14869
rect 7423 14854 7483 14869
rect 7541 14854 7601 14869
rect 7778 14869 8074 14908
rect 7778 14854 7838 14869
rect 7896 14854 7956 14869
rect 8014 14854 8074 14869
rect 8132 14869 8428 14908
rect 8132 14854 8192 14869
rect 8250 14854 8310 14869
rect 8368 14854 8428 14869
rect 8599 14869 8895 14908
rect 8599 14854 8659 14869
rect 8717 14854 8777 14869
rect 8835 14854 8895 14869
rect 10449 14869 10745 14908
rect 10449 14854 10509 14869
rect 10567 14854 10627 14869
rect 10685 14854 10745 14869
rect 10922 14869 11218 14908
rect 10922 14854 10982 14869
rect 11040 14854 11100 14869
rect 11158 14854 11218 14869
rect 11276 14869 11572 14908
rect 11276 14854 11336 14869
rect 11394 14854 11454 14869
rect 11512 14854 11572 14869
rect 11743 14869 12039 14908
rect 11743 14854 11803 14869
rect 11861 14854 11921 14869
rect 11979 14854 12039 14869
rect 13651 14873 13947 14912
rect 13651 14858 13711 14873
rect 13769 14858 13829 14873
rect 13887 14858 13947 14873
rect 14124 14873 14420 14912
rect 14124 14858 14184 14873
rect 14242 14858 14302 14873
rect 14360 14858 14420 14873
rect 14478 14873 14774 14912
rect 14478 14858 14538 14873
rect 14596 14858 14656 14873
rect 14714 14858 14774 14873
rect 14945 14873 15241 14912
rect 14945 14858 15005 14873
rect 15063 14858 15123 14873
rect 15181 14858 15241 14873
rect 16795 14873 17091 14912
rect 16795 14858 16855 14873
rect 16913 14858 16973 14873
rect 17031 14858 17091 14873
rect 17268 14873 17564 14912
rect 17268 14858 17328 14873
rect 17386 14858 17446 14873
rect 17504 14858 17564 14873
rect 17622 14873 17918 14912
rect 17622 14858 17682 14873
rect 17740 14858 17800 14873
rect 17858 14858 17918 14873
rect 18089 14873 18385 14912
rect 18089 14858 18149 14873
rect 18207 14858 18267 14873
rect 18325 14858 18385 14873
rect 19927 14869 20223 14908
rect 5908 14674 6204 14713
rect 5908 14658 5968 14674
rect 6026 14658 6086 14674
rect 6144 14658 6204 14674
rect 6832 14670 7128 14709
rect 6832 14654 6892 14670
rect 6950 14654 7010 14670
rect 7068 14654 7128 14670
rect 556 14309 616 14458
rect 674 14432 734 14458
rect 792 14432 852 14458
rect 1029 14432 1089 14458
rect 660 14309 726 14312
rect 556 14296 726 14309
rect 556 14262 676 14296
rect 710 14262 726 14296
rect 556 14249 726 14262
rect 556 13773 616 14249
rect 660 14246 726 14249
rect 1147 14042 1207 14458
rect 1265 14432 1325 14458
rect 1502 14432 1562 14458
rect 1620 14133 1680 14458
rect 1738 14432 1798 14458
rect 1856 14432 1916 14458
rect 1974 14432 2034 14458
rect 2092 14432 2152 14458
rect 2323 14432 2383 14458
rect 1974 14272 2033 14432
rect 1970 14271 2033 14272
rect 1970 14255 2036 14271
rect 1970 14221 1986 14255
rect 2020 14221 2036 14255
rect 1970 14205 2036 14221
rect 1838 14156 1933 14171
rect 1838 14133 1856 14156
rect 1620 14101 1856 14133
rect 1914 14101 1933 14156
rect 1620 14084 1933 14101
rect 1147 14025 1685 14042
rect 1147 13991 1632 14025
rect 1666 13991 1685 14025
rect 1147 13985 1685 13991
rect 1616 13975 1685 13985
rect 1620 13973 1685 13975
rect 556 13728 1484 13773
rect 1424 13525 1484 13728
rect 1620 13525 1680 13973
rect 1735 13635 1801 13651
rect 1735 13601 1751 13635
rect 1785 13601 1801 13635
rect 1735 13585 1801 13601
rect 1738 13525 1798 13585
rect 1856 13525 1916 14084
rect 2441 14040 2501 14458
rect 2559 14432 2619 14458
rect 2764 14432 2824 14458
rect 2882 14432 2942 14458
rect 3000 14172 3060 14458
rect 2924 14155 3060 14172
rect 2924 14100 2943 14155
rect 3001 14100 3060 14155
rect 2924 14085 3060 14100
rect 1974 13983 2501 14040
rect 1974 13884 2034 13983
rect 1964 13871 2045 13884
rect 1964 13816 1974 13871
rect 2032 13816 2045 13871
rect 1964 13805 2045 13816
rect 1974 13525 2034 13805
rect 3000 13773 3060 14085
rect 2166 13728 3060 13773
rect 3700 14309 3760 14458
rect 3818 14432 3878 14458
rect 3936 14432 3996 14458
rect 4173 14432 4233 14458
rect 3804 14309 3870 14312
rect 3700 14296 3870 14309
rect 3700 14262 3820 14296
rect 3854 14262 3870 14296
rect 3700 14249 3870 14262
rect 3700 13773 3760 14249
rect 3804 14246 3870 14249
rect 4291 14042 4351 14458
rect 4409 14432 4469 14458
rect 4646 14432 4706 14458
rect 4764 14133 4824 14458
rect 4882 14432 4942 14458
rect 5000 14432 5060 14458
rect 5118 14432 5178 14458
rect 5236 14432 5296 14458
rect 5467 14432 5527 14458
rect 5118 14272 5177 14432
rect 5114 14271 5177 14272
rect 5114 14255 5180 14271
rect 5114 14221 5130 14255
rect 5164 14221 5180 14255
rect 5114 14205 5180 14221
rect 4982 14156 5077 14171
rect 4982 14133 5000 14156
rect 4764 14101 5000 14133
rect 5058 14101 5077 14156
rect 4764 14084 5077 14101
rect 4291 14025 4829 14042
rect 4291 13991 4776 14025
rect 4810 13991 4829 14025
rect 4291 13985 4829 13991
rect 4760 13975 4829 13985
rect 4764 13973 4829 13975
rect 3700 13728 4628 13773
rect 2166 13525 2226 13728
rect 4568 13525 4628 13728
rect 4764 13525 4824 13973
rect 4879 13635 4945 13651
rect 4879 13601 4895 13635
rect 4929 13601 4945 13635
rect 4879 13585 4945 13601
rect 4882 13525 4942 13585
rect 5000 13525 5060 14084
rect 5585 14040 5645 14458
rect 5703 14432 5763 14458
rect 5908 14432 5968 14458
rect 6026 14432 6086 14458
rect 6144 14172 6204 14458
rect 9040 14670 9336 14709
rect 9040 14654 9100 14670
rect 9158 14654 9218 14670
rect 9276 14654 9336 14670
rect 9976 14670 10272 14709
rect 9976 14654 10036 14670
rect 10094 14654 10154 14670
rect 10212 14654 10272 14670
rect 12184 14670 12480 14709
rect 12184 14654 12244 14670
rect 12302 14654 12362 14670
rect 12420 14654 12480 14670
rect 13178 14674 13474 14713
rect 13178 14658 13238 14674
rect 13296 14658 13356 14674
rect 13414 14658 13474 14674
rect 15386 14674 15682 14713
rect 15386 14658 15446 14674
rect 15504 14658 15564 14674
rect 15622 14658 15682 14674
rect 16322 14674 16618 14713
rect 16322 14658 16382 14674
rect 16440 14658 16500 14674
rect 16558 14658 16618 14674
rect 19927 14854 19987 14869
rect 20045 14854 20105 14869
rect 20163 14854 20223 14869
rect 20400 14869 20696 14908
rect 20400 14854 20460 14869
rect 20518 14854 20578 14869
rect 20636 14854 20696 14869
rect 20754 14869 21050 14908
rect 20754 14854 20814 14869
rect 20872 14854 20932 14869
rect 20990 14854 21050 14869
rect 21221 14869 21517 14908
rect 21221 14854 21281 14869
rect 21339 14854 21399 14869
rect 21457 14854 21517 14869
rect 23071 14869 23367 14908
rect 23071 14854 23131 14869
rect 23189 14854 23249 14869
rect 23307 14854 23367 14869
rect 23544 14869 23840 14908
rect 23544 14854 23604 14869
rect 23662 14854 23722 14869
rect 23780 14854 23840 14869
rect 23898 14869 24194 14908
rect 23898 14854 23958 14869
rect 24016 14854 24076 14869
rect 24134 14854 24194 14869
rect 24365 14869 24661 14908
rect 24365 14854 24425 14869
rect 24483 14854 24543 14869
rect 24601 14854 24661 14869
rect 18530 14674 18826 14713
rect 18530 14658 18590 14674
rect 18648 14658 18708 14674
rect 18766 14658 18826 14674
rect 19454 14670 19750 14709
rect 19454 14654 19514 14670
rect 19572 14654 19632 14670
rect 19690 14654 19750 14670
rect 6068 14155 6204 14172
rect 6068 14100 6087 14155
rect 6145 14100 6204 14155
rect 6068 14085 6204 14100
rect 5118 13983 5645 14040
rect 5118 13884 5178 13983
rect 5108 13871 5189 13884
rect 5108 13816 5118 13871
rect 5176 13816 5189 13871
rect 5108 13805 5189 13816
rect 5118 13525 5178 13805
rect 6144 13773 6204 14085
rect 5310 13728 6204 13773
rect 6832 14305 6892 14454
rect 6950 14428 7010 14454
rect 7068 14428 7128 14454
rect 7305 14428 7365 14454
rect 6936 14305 7002 14308
rect 6832 14292 7002 14305
rect 6832 14258 6952 14292
rect 6986 14258 7002 14292
rect 6832 14245 7002 14258
rect 6832 13769 6892 14245
rect 6936 14242 7002 14245
rect 7423 14038 7483 14454
rect 7541 14428 7601 14454
rect 7778 14428 7838 14454
rect 7896 14129 7956 14454
rect 8014 14428 8074 14454
rect 8132 14428 8192 14454
rect 8250 14428 8310 14454
rect 8368 14428 8428 14454
rect 8599 14428 8659 14454
rect 8250 14268 8309 14428
rect 8246 14267 8309 14268
rect 8246 14251 8312 14267
rect 8246 14217 8262 14251
rect 8296 14217 8312 14251
rect 8246 14201 8312 14217
rect 8114 14152 8209 14167
rect 8114 14129 8132 14152
rect 7896 14097 8132 14129
rect 8190 14097 8209 14152
rect 7896 14080 8209 14097
rect 7423 14021 7961 14038
rect 7423 13987 7908 14021
rect 7942 13987 7961 14021
rect 7423 13981 7961 13987
rect 7892 13971 7961 13981
rect 7896 13969 7961 13971
rect 5310 13525 5370 13728
rect 6832 13724 7760 13769
rect 1424 13044 1484 13325
rect 2166 13299 2226 13325
rect 1620 13099 1680 13125
rect 1738 13099 1798 13125
rect 1856 13099 1916 13125
rect 1974 13099 2034 13125
rect 1793 13044 1859 13052
rect 1424 13036 1859 13044
rect 1424 13002 1809 13036
rect 1843 13002 1859 13036
rect 1424 12993 1859 13002
rect 4568 13044 4628 13325
rect 7700 13521 7760 13724
rect 7896 13521 7956 13969
rect 8011 13631 8077 13647
rect 8011 13597 8027 13631
rect 8061 13597 8077 13631
rect 8011 13581 8077 13597
rect 8014 13521 8074 13581
rect 8132 13521 8192 14080
rect 8717 14036 8777 14454
rect 8835 14428 8895 14454
rect 9040 14428 9100 14454
rect 9158 14428 9218 14454
rect 9276 14168 9336 14454
rect 9200 14151 9336 14168
rect 9200 14096 9219 14151
rect 9277 14096 9336 14151
rect 9200 14081 9336 14096
rect 8250 13979 8777 14036
rect 8250 13880 8310 13979
rect 8240 13867 8321 13880
rect 8240 13812 8250 13867
rect 8308 13812 8321 13867
rect 8240 13801 8321 13812
rect 8250 13521 8310 13801
rect 9276 13769 9336 14081
rect 8442 13724 9336 13769
rect 9976 14305 10036 14454
rect 10094 14428 10154 14454
rect 10212 14428 10272 14454
rect 10449 14428 10509 14454
rect 10080 14305 10146 14308
rect 9976 14292 10146 14305
rect 9976 14258 10096 14292
rect 10130 14258 10146 14292
rect 9976 14245 10146 14258
rect 9976 13769 10036 14245
rect 10080 14242 10146 14245
rect 10567 14038 10627 14454
rect 10685 14428 10745 14454
rect 10922 14428 10982 14454
rect 11040 14129 11100 14454
rect 11158 14428 11218 14454
rect 11276 14428 11336 14454
rect 11394 14428 11454 14454
rect 11512 14428 11572 14454
rect 11743 14428 11803 14454
rect 11394 14268 11453 14428
rect 11390 14267 11453 14268
rect 11390 14251 11456 14267
rect 11390 14217 11406 14251
rect 11440 14217 11456 14251
rect 11390 14201 11456 14217
rect 11258 14152 11353 14167
rect 11258 14129 11276 14152
rect 11040 14097 11276 14129
rect 11334 14097 11353 14152
rect 11040 14080 11353 14097
rect 10567 14021 11105 14038
rect 10567 13987 11052 14021
rect 11086 13987 11105 14021
rect 10567 13981 11105 13987
rect 11036 13971 11105 13981
rect 11040 13969 11105 13971
rect 9976 13724 10904 13769
rect 8442 13521 8502 13724
rect 10844 13521 10904 13724
rect 11040 13521 11100 13969
rect 11155 13631 11221 13647
rect 11155 13597 11171 13631
rect 11205 13597 11221 13631
rect 11155 13581 11221 13597
rect 11158 13521 11218 13581
rect 11276 13521 11336 14080
rect 11861 14036 11921 14454
rect 11979 14428 12039 14454
rect 12184 14428 12244 14454
rect 12302 14428 12362 14454
rect 12420 14168 12480 14454
rect 12344 14151 12480 14168
rect 12344 14096 12363 14151
rect 12421 14096 12480 14151
rect 12344 14081 12480 14096
rect 11394 13979 11921 14036
rect 11394 13880 11454 13979
rect 11384 13867 11465 13880
rect 11384 13812 11394 13867
rect 11452 13812 11465 13867
rect 11384 13801 11465 13812
rect 11394 13521 11454 13801
rect 12420 13769 12480 14081
rect 11586 13724 12480 13769
rect 13178 14309 13238 14458
rect 13296 14432 13356 14458
rect 13414 14432 13474 14458
rect 13651 14432 13711 14458
rect 13282 14309 13348 14312
rect 13178 14296 13348 14309
rect 13178 14262 13298 14296
rect 13332 14262 13348 14296
rect 13178 14249 13348 14262
rect 13178 13773 13238 14249
rect 13282 14246 13348 14249
rect 13769 14042 13829 14458
rect 13887 14432 13947 14458
rect 14124 14432 14184 14458
rect 14242 14133 14302 14458
rect 14360 14432 14420 14458
rect 14478 14432 14538 14458
rect 14596 14432 14656 14458
rect 14714 14432 14774 14458
rect 14945 14432 15005 14458
rect 14596 14272 14655 14432
rect 14592 14271 14655 14272
rect 14592 14255 14658 14271
rect 14592 14221 14608 14255
rect 14642 14221 14658 14255
rect 14592 14205 14658 14221
rect 14460 14156 14555 14171
rect 14460 14133 14478 14156
rect 14242 14101 14478 14133
rect 14536 14101 14555 14156
rect 14242 14084 14555 14101
rect 13769 14025 14307 14042
rect 13769 13991 14254 14025
rect 14288 13991 14307 14025
rect 13769 13985 14307 13991
rect 14238 13975 14307 13985
rect 14242 13973 14307 13975
rect 13178 13728 14106 13773
rect 11586 13521 11646 13724
rect 14046 13525 14106 13728
rect 14242 13525 14302 13973
rect 14357 13635 14423 13651
rect 14357 13601 14373 13635
rect 14407 13601 14423 13635
rect 14357 13585 14423 13601
rect 14360 13525 14420 13585
rect 14478 13525 14538 14084
rect 15063 14040 15123 14458
rect 15181 14432 15241 14458
rect 15386 14432 15446 14458
rect 15504 14432 15564 14458
rect 15622 14172 15682 14458
rect 15546 14155 15682 14172
rect 15546 14100 15565 14155
rect 15623 14100 15682 14155
rect 15546 14085 15682 14100
rect 14596 13983 15123 14040
rect 14596 13884 14656 13983
rect 14586 13871 14667 13884
rect 14586 13816 14596 13871
rect 14654 13816 14667 13871
rect 14586 13805 14667 13816
rect 14596 13525 14656 13805
rect 15622 13773 15682 14085
rect 14788 13728 15682 13773
rect 16322 14309 16382 14458
rect 16440 14432 16500 14458
rect 16558 14432 16618 14458
rect 16795 14432 16855 14458
rect 16426 14309 16492 14312
rect 16322 14296 16492 14309
rect 16322 14262 16442 14296
rect 16476 14262 16492 14296
rect 16322 14249 16492 14262
rect 16322 13773 16382 14249
rect 16426 14246 16492 14249
rect 16913 14042 16973 14458
rect 17031 14432 17091 14458
rect 17268 14432 17328 14458
rect 17386 14133 17446 14458
rect 17504 14432 17564 14458
rect 17622 14432 17682 14458
rect 17740 14432 17800 14458
rect 17858 14432 17918 14458
rect 18089 14432 18149 14458
rect 17740 14272 17799 14432
rect 17736 14271 17799 14272
rect 17736 14255 17802 14271
rect 17736 14221 17752 14255
rect 17786 14221 17802 14255
rect 17736 14205 17802 14221
rect 17604 14156 17699 14171
rect 17604 14133 17622 14156
rect 17386 14101 17622 14133
rect 17680 14101 17699 14156
rect 17386 14084 17699 14101
rect 16913 14025 17451 14042
rect 16913 13991 17398 14025
rect 17432 13991 17451 14025
rect 16913 13985 17451 13991
rect 17382 13975 17451 13985
rect 17386 13973 17451 13975
rect 16322 13728 17250 13773
rect 14788 13525 14848 13728
rect 17190 13525 17250 13728
rect 17386 13525 17446 13973
rect 17501 13635 17567 13651
rect 17501 13601 17517 13635
rect 17551 13601 17567 13635
rect 17501 13585 17567 13601
rect 17504 13525 17564 13585
rect 17622 13525 17682 14084
rect 18207 14040 18267 14458
rect 18325 14432 18385 14458
rect 18530 14432 18590 14458
rect 18648 14432 18708 14458
rect 18766 14172 18826 14458
rect 21662 14670 21958 14709
rect 21662 14654 21722 14670
rect 21780 14654 21840 14670
rect 21898 14654 21958 14670
rect 22598 14670 22894 14709
rect 22598 14654 22658 14670
rect 22716 14654 22776 14670
rect 22834 14654 22894 14670
rect 45473 15203 45533 15229
rect 46771 15203 46831 15229
rect 47371 15203 47431 15229
rect 49552 15419 49618 15435
rect 49552 15385 49568 15419
rect 49602 15385 49618 15419
rect 49552 15369 49618 15385
rect 49670 15302 49736 15318
rect 49670 15268 49686 15302
rect 49720 15268 49736 15302
rect 49670 15252 49736 15268
rect 49673 15230 49733 15252
rect 49908 15230 49968 15441
rect 50028 15256 50086 15441
rect 52007 15434 52067 15472
rect 52531 15434 52591 15540
rect 52885 15599 52945 15766
rect 53003 15740 53063 15766
rect 53305 15733 53365 16391
rect 53890 16389 53965 16433
rect 54007 16389 54550 16440
rect 54608 16433 54668 16459
rect 54726 16433 54786 16459
rect 54844 16442 54904 16459
rect 55092 16442 55152 16459
rect 55210 16442 55270 16459
rect 55328 16442 55388 16459
rect 54844 16391 55388 16442
rect 58386 16679 58682 16730
rect 58386 16662 58446 16679
rect 58504 16662 58564 16679
rect 58622 16662 58682 16679
rect 59707 16662 59767 16688
rect 59825 16662 59885 16688
rect 59943 16662 60003 16688
rect 60284 16679 60580 16730
rect 60284 16662 60344 16679
rect 60402 16662 60462 16679
rect 60520 16662 60580 16679
rect 62715 16842 62775 16864
rect 62950 16842 63010 17053
rect 63070 16868 63128 17053
rect 63068 16842 63128 16868
rect 70459 17018 70498 17076
rect 71329 17018 71386 17427
rect 72327 17295 72378 17604
rect 70459 16958 70513 17018
rect 70913 16958 71386 17018
rect 71598 17235 71846 17295
rect 72046 17235 72378 17295
rect 70459 16900 70498 16958
rect 61605 16662 61665 16688
rect 61723 16662 61783 16688
rect 61841 16662 61901 16688
rect 62715 16616 62775 16642
rect 56437 16423 56497 16439
rect 53298 15717 53365 15733
rect 53298 15683 53315 15717
rect 53349 15683 53365 15717
rect 53298 15667 53365 15683
rect 53028 15599 53095 15606
rect 52885 15590 53095 15599
rect 52885 15556 53045 15590
rect 53079 15556 53095 15590
rect 52885 15540 53095 15556
rect 52645 15507 52711 15522
rect 52645 15473 52661 15507
rect 52695 15473 52711 15507
rect 52645 15457 52711 15473
rect 52763 15506 52829 15522
rect 52763 15472 52779 15506
rect 52813 15472 52829 15506
rect 52649 15434 52709 15457
rect 52763 15456 52829 15472
rect 52767 15434 52827 15456
rect 52885 15434 52945 15540
rect 53305 15539 53365 15667
rect 53214 15523 53365 15539
rect 53214 15489 53230 15523
rect 53264 15489 53365 15523
rect 53214 15473 53365 15489
rect 53305 15434 53365 15473
rect 53905 16269 53965 16389
rect 55203 16310 55263 16391
rect 56429 16401 56503 16423
rect 56555 16417 56615 16439
rect 58386 16436 58446 16462
rect 58504 16443 58564 16462
rect 58622 16443 58682 16462
rect 58869 16443 58929 16462
rect 58987 16443 59047 16462
rect 59105 16443 59165 16462
rect 58504 16436 58580 16443
rect 56429 16367 56450 16401
rect 56484 16367 56503 16401
rect 56429 16310 56503 16367
rect 56552 16401 56618 16417
rect 56552 16367 56568 16401
rect 56602 16367 56618 16401
rect 58505 16392 58580 16436
rect 58622 16392 59165 16443
rect 59223 16436 59283 16462
rect 59341 16436 59401 16462
rect 59459 16445 59519 16462
rect 59707 16445 59767 16462
rect 59825 16445 59885 16462
rect 59943 16445 60003 16462
rect 59459 16394 60003 16445
rect 60284 16436 60344 16462
rect 60402 16443 60462 16462
rect 60520 16443 60580 16462
rect 60767 16443 60827 16462
rect 60885 16443 60945 16462
rect 61003 16443 61063 16462
rect 60402 16436 60478 16443
rect 56552 16351 56618 16367
rect 55203 16285 56503 16310
rect 53905 16249 53966 16269
rect 53905 16233 53985 16249
rect 53905 16199 53936 16233
rect 53970 16199 53985 16233
rect 53905 16183 53985 16199
rect 54311 16190 54607 16250
rect 53905 16160 53966 16183
rect 54311 16166 54371 16190
rect 54429 16166 54489 16190
rect 54547 16166 54607 16190
rect 54665 16189 54961 16249
rect 54665 16166 54725 16189
rect 54783 16166 54843 16189
rect 54901 16166 54961 16189
rect 55203 16237 56504 16285
rect 58520 16239 58580 16392
rect 53905 16014 53965 16160
rect 53905 15841 53966 16014
rect 53905 15538 53965 15841
rect 54311 15740 54371 15766
rect 54279 15599 54346 15606
rect 54429 15599 54489 15766
rect 54547 15740 54607 15766
rect 54665 15740 54725 15766
rect 54279 15590 54489 15599
rect 54279 15556 54295 15590
rect 54329 15556 54489 15590
rect 54279 15540 54489 15556
rect 53905 15522 54055 15538
rect 53905 15488 54005 15522
rect 54039 15488 54055 15522
rect 53905 15472 54055 15488
rect 53905 15434 53965 15472
rect 54429 15434 54489 15540
rect 54783 15599 54843 15766
rect 54901 15740 54961 15766
rect 54926 15599 54993 15606
rect 54783 15590 54993 15599
rect 54783 15556 54943 15590
rect 54977 15556 54993 15590
rect 54783 15540 54993 15556
rect 54543 15507 54609 15522
rect 54543 15473 54559 15507
rect 54593 15473 54609 15507
rect 54543 15457 54609 15473
rect 54661 15506 54727 15522
rect 54661 15472 54677 15506
rect 54711 15472 54727 15506
rect 54547 15434 54607 15457
rect 54661 15456 54727 15472
rect 54665 15434 54725 15456
rect 54783 15434 54843 15540
rect 55203 15539 55263 16237
rect 58326 16215 58580 16239
rect 58326 16181 58342 16215
rect 58376 16181 58580 16215
rect 58326 16165 58580 16181
rect 58926 16193 59222 16253
rect 58926 16169 58986 16193
rect 59044 16169 59104 16193
rect 59162 16169 59222 16193
rect 59280 16192 59576 16252
rect 59280 16169 59340 16192
rect 59398 16169 59458 16192
rect 59516 16169 59576 16192
rect 55853 15692 56149 15728
rect 55853 15672 55913 15692
rect 55971 15672 56031 15692
rect 56089 15672 56149 15692
rect 56207 15692 56503 15728
rect 56207 15672 56267 15692
rect 56325 15672 56385 15692
rect 56443 15672 56503 15692
rect 56561 15693 56857 15729
rect 56561 15672 56621 15693
rect 56679 15672 56739 15693
rect 56797 15672 56857 15693
rect 55112 15523 55263 15539
rect 55112 15489 55128 15523
rect 55162 15489 55263 15523
rect 55112 15473 55263 15489
rect 55203 15434 55263 15473
rect 58520 15541 58580 16165
rect 58926 15743 58986 15769
rect 58896 15603 58963 15610
rect 58896 15602 58969 15603
rect 59044 15602 59104 15769
rect 59162 15743 59222 15769
rect 59280 15743 59340 15769
rect 58896 15594 59104 15602
rect 58896 15560 58912 15594
rect 58946 15560 59104 15594
rect 58896 15544 59104 15560
rect 58907 15543 59104 15544
rect 58520 15525 58670 15541
rect 58520 15491 58620 15525
rect 58654 15491 58670 15525
rect 58520 15475 58670 15491
rect 55853 15446 55913 15472
rect 55971 15446 56031 15472
rect 56089 15440 56149 15472
rect 56207 15446 56267 15472
rect 56325 15446 56385 15472
rect 56443 15452 56503 15472
rect 56442 15446 56503 15452
rect 56561 15446 56621 15472
rect 56679 15446 56739 15472
rect 56797 15446 56857 15472
rect 50026 15230 50086 15256
rect 48669 15203 48729 15229
rect 45997 15003 46057 15029
rect 46115 15003 46175 15029
rect 46233 15003 46293 15029
rect 46351 15003 46411 15029
rect 47895 15003 47955 15029
rect 48013 15003 48073 15029
rect 48131 15003 48191 15029
rect 48249 15003 48309 15029
rect 49673 15004 49733 15030
rect 43350 14812 43410 14834
rect 43468 14812 43528 14834
rect 43347 14796 43413 14812
rect 43347 14762 43363 14796
rect 43397 14762 43413 14796
rect 43347 14746 43413 14762
rect 43465 14796 43531 14812
rect 43465 14762 43481 14796
rect 43515 14762 43531 14796
rect 52007 15208 52067 15234
rect 53305 15208 53365 15234
rect 53905 15208 53965 15234
rect 56086 15424 56152 15440
rect 56086 15390 56102 15424
rect 56136 15390 56152 15424
rect 56086 15374 56152 15390
rect 56204 15307 56270 15323
rect 56204 15273 56220 15307
rect 56254 15273 56270 15307
rect 56204 15257 56270 15273
rect 56207 15235 56267 15257
rect 56442 15235 56502 15446
rect 56562 15261 56620 15446
rect 58520 15437 58580 15475
rect 59044 15437 59104 15543
rect 59398 15602 59458 15769
rect 59516 15743 59576 15769
rect 59818 15736 59878 16394
rect 60403 16392 60478 16436
rect 60520 16392 61063 16443
rect 61121 16436 61181 16462
rect 61239 16436 61299 16462
rect 61357 16445 61417 16462
rect 61605 16445 61665 16462
rect 61723 16445 61783 16462
rect 61841 16445 61901 16462
rect 61357 16394 61901 16445
rect 70459 16840 70513 16900
rect 70913 16840 70939 16900
rect 70658 16603 70713 16663
rect 70913 16603 70939 16663
rect 70658 16545 70697 16603
rect 70658 16485 70713 16545
rect 70913 16485 70939 16545
rect 71059 16521 71125 16537
rect 71059 16487 71075 16521
rect 71109 16487 71125 16521
rect 62950 16426 63010 16442
rect 59811 15720 59878 15736
rect 59811 15686 59828 15720
rect 59862 15686 59878 15720
rect 59811 15670 59878 15686
rect 59541 15602 59608 15609
rect 59398 15593 59608 15602
rect 59398 15559 59558 15593
rect 59592 15559 59608 15593
rect 59398 15543 59608 15559
rect 59158 15510 59224 15525
rect 59158 15476 59174 15510
rect 59208 15476 59224 15510
rect 59158 15460 59224 15476
rect 59276 15509 59342 15525
rect 59276 15475 59292 15509
rect 59326 15475 59342 15509
rect 59162 15437 59222 15460
rect 59276 15459 59342 15475
rect 59280 15437 59340 15459
rect 59398 15437 59458 15543
rect 59818 15542 59878 15670
rect 59727 15526 59878 15542
rect 59727 15492 59743 15526
rect 59777 15492 59878 15526
rect 59727 15476 59878 15492
rect 59818 15437 59878 15476
rect 60418 16272 60478 16392
rect 61716 16313 61776 16394
rect 62942 16404 63016 16426
rect 63068 16420 63128 16442
rect 70658 16427 70697 16485
rect 71059 16471 71125 16487
rect 71062 16427 71122 16471
rect 71598 16427 71643 17235
rect 62942 16370 62963 16404
rect 62997 16370 63016 16404
rect 62942 16313 63016 16370
rect 63065 16404 63131 16420
rect 63065 16370 63081 16404
rect 63115 16370 63131 16404
rect 63065 16354 63131 16370
rect 70658 16367 70713 16427
rect 70913 16367 71643 16427
rect 61716 16288 63016 16313
rect 60418 16252 60479 16272
rect 60418 16236 60498 16252
rect 60418 16202 60449 16236
rect 60483 16202 60498 16236
rect 60418 16186 60498 16202
rect 60824 16193 61120 16253
rect 60418 16163 60479 16186
rect 60824 16169 60884 16193
rect 60942 16169 61002 16193
rect 61060 16169 61120 16193
rect 61178 16192 61474 16252
rect 61178 16169 61238 16192
rect 61296 16169 61356 16192
rect 61414 16169 61474 16192
rect 61716 16240 63017 16288
rect 60418 16017 60478 16163
rect 60418 15844 60479 16017
rect 60418 15541 60478 15844
rect 60824 15743 60884 15769
rect 60792 15602 60859 15609
rect 60942 15602 61002 15769
rect 61060 15743 61120 15769
rect 61178 15743 61238 15769
rect 60792 15593 61002 15602
rect 60792 15559 60808 15593
rect 60842 15559 61002 15593
rect 60792 15543 61002 15559
rect 60418 15525 60568 15541
rect 60418 15491 60518 15525
rect 60552 15491 60568 15525
rect 60418 15475 60568 15491
rect 60418 15437 60478 15475
rect 60942 15437 61002 15543
rect 61296 15602 61356 15769
rect 61414 15743 61474 15769
rect 61439 15602 61506 15609
rect 61296 15593 61506 15602
rect 61296 15559 61456 15593
rect 61490 15559 61506 15593
rect 61296 15543 61506 15559
rect 61056 15510 61122 15525
rect 61056 15476 61072 15510
rect 61106 15476 61122 15510
rect 61056 15460 61122 15476
rect 61174 15509 61240 15525
rect 61174 15475 61190 15509
rect 61224 15475 61240 15509
rect 61060 15437 61120 15460
rect 61174 15459 61240 15475
rect 61178 15437 61238 15459
rect 61296 15437 61356 15543
rect 61716 15542 61776 16240
rect 62366 15695 62662 15731
rect 62366 15675 62426 15695
rect 62484 15675 62544 15695
rect 62602 15675 62662 15695
rect 62720 15695 63016 15731
rect 62720 15675 62780 15695
rect 62838 15675 62898 15695
rect 62956 15675 63016 15695
rect 63074 15696 63370 15732
rect 63074 15675 63134 15696
rect 63192 15675 63252 15696
rect 63310 15675 63370 15696
rect 70654 15679 70709 15739
rect 70909 15680 71639 15739
rect 70909 15679 71212 15680
rect 61625 15526 61776 15542
rect 61625 15492 61641 15526
rect 61675 15492 61776 15526
rect 61625 15476 61776 15492
rect 61716 15437 61776 15476
rect 70654 15621 70693 15679
rect 71195 15622 71212 15679
rect 71267 15679 71639 15680
rect 71267 15622 71282 15679
rect 70654 15561 70709 15621
rect 70909 15561 70935 15621
rect 71195 15603 71282 15622
rect 70654 15503 70693 15561
rect 62366 15449 62426 15475
rect 62484 15449 62544 15475
rect 62602 15443 62662 15475
rect 62720 15449 62780 15475
rect 62838 15449 62898 15475
rect 62956 15455 63016 15475
rect 62955 15449 63016 15455
rect 63074 15449 63134 15475
rect 63192 15449 63252 15475
rect 63310 15449 63370 15475
rect 56560 15235 56620 15261
rect 55203 15208 55263 15234
rect 52531 15008 52591 15034
rect 52649 15008 52709 15034
rect 52767 15008 52827 15034
rect 52885 15008 52945 15034
rect 54429 15008 54489 15034
rect 54547 15008 54607 15034
rect 54665 15008 54725 15034
rect 54783 15008 54843 15034
rect 56207 15009 56267 15035
rect 49908 14808 49968 14830
rect 50026 14808 50086 14830
rect 43465 14746 43531 14762
rect 24806 14670 25102 14709
rect 24806 14654 24866 14670
rect 24924 14654 24984 14670
rect 25042 14654 25102 14670
rect 49905 14792 49971 14808
rect 49905 14758 49921 14792
rect 49955 14758 49971 14792
rect 49905 14742 49971 14758
rect 50023 14792 50089 14808
rect 50023 14758 50039 14792
rect 50073 14758 50089 14792
rect 58520 15211 58580 15237
rect 59818 15211 59878 15237
rect 60418 15211 60478 15237
rect 62599 15427 62665 15443
rect 62599 15393 62615 15427
rect 62649 15393 62665 15427
rect 62599 15377 62665 15393
rect 62717 15310 62783 15326
rect 62717 15276 62733 15310
rect 62767 15276 62783 15310
rect 62717 15260 62783 15276
rect 62720 15238 62780 15260
rect 62955 15238 63015 15449
rect 63075 15264 63133 15449
rect 70654 15443 70709 15503
rect 70909 15443 70935 15503
rect 63073 15238 63133 15264
rect 70455 15238 70509 15298
rect 70909 15238 70935 15298
rect 61716 15211 61776 15237
rect 59044 15011 59104 15037
rect 59162 15011 59222 15037
rect 59280 15011 59340 15037
rect 59398 15011 59458 15037
rect 60942 15011 61002 15037
rect 61060 15011 61120 15037
rect 61178 15011 61238 15037
rect 61296 15011 61356 15037
rect 62720 15012 62780 15038
rect 56442 14813 56502 14835
rect 56560 14813 56620 14835
rect 50023 14742 50089 14758
rect 56439 14797 56505 14813
rect 56439 14763 56455 14797
rect 56489 14763 56505 14797
rect 56439 14747 56505 14763
rect 56557 14797 56623 14813
rect 56557 14763 56573 14797
rect 56607 14763 56623 14797
rect 70455 15180 70494 15238
rect 70455 15120 70509 15180
rect 70909 15120 71384 15180
rect 70455 15062 70494 15120
rect 70455 15002 70509 15062
rect 70909 15002 70935 15062
rect 62955 14816 63015 14838
rect 63073 14816 63133 14838
rect 56557 14747 56623 14763
rect 62952 14800 63018 14816
rect 62952 14766 62968 14800
rect 63002 14766 63018 14800
rect 62952 14750 63018 14766
rect 63070 14800 63136 14816
rect 63070 14766 63086 14800
rect 63120 14766 63136 14800
rect 63070 14750 63136 14766
rect 70455 14771 70509 14831
rect 70909 14771 70935 14831
rect 70455 14713 70494 14771
rect 70455 14653 70509 14713
rect 70909 14712 70935 14713
rect 71096 14712 71162 14715
rect 70909 14699 71162 14712
rect 70909 14665 71112 14699
rect 71146 14665 71162 14699
rect 70909 14653 71162 14665
rect 71327 14713 71384 15120
rect 71594 14905 71639 15679
rect 71594 14845 71842 14905
rect 72042 14845 72068 14905
rect 71483 14713 71562 14724
rect 71327 14711 71842 14713
rect 71327 14653 71496 14711
rect 71551 14653 71842 14711
rect 72242 14653 72268 14713
rect 18690 14155 18826 14172
rect 18690 14100 18709 14155
rect 18767 14100 18826 14155
rect 18690 14085 18826 14100
rect 17740 13983 18267 14040
rect 17740 13884 17800 13983
rect 17730 13871 17811 13884
rect 17730 13816 17740 13871
rect 17798 13816 17811 13871
rect 17730 13805 17811 13816
rect 17740 13525 17800 13805
rect 18766 13773 18826 14085
rect 17932 13728 18826 13773
rect 19454 14305 19514 14454
rect 19572 14428 19632 14454
rect 19690 14428 19750 14454
rect 19927 14428 19987 14454
rect 19558 14305 19624 14308
rect 19454 14292 19624 14305
rect 19454 14258 19574 14292
rect 19608 14258 19624 14292
rect 19454 14245 19624 14258
rect 19454 13769 19514 14245
rect 19558 14242 19624 14245
rect 20045 14038 20105 14454
rect 20163 14428 20223 14454
rect 20400 14428 20460 14454
rect 20518 14129 20578 14454
rect 20636 14428 20696 14454
rect 20754 14428 20814 14454
rect 20872 14428 20932 14454
rect 20990 14428 21050 14454
rect 21221 14428 21281 14454
rect 20872 14268 20931 14428
rect 20868 14267 20931 14268
rect 20868 14251 20934 14267
rect 20868 14217 20884 14251
rect 20918 14217 20934 14251
rect 20868 14201 20934 14217
rect 20736 14152 20831 14167
rect 20736 14129 20754 14152
rect 20518 14097 20754 14129
rect 20812 14097 20831 14152
rect 20518 14080 20831 14097
rect 20045 14021 20583 14038
rect 20045 13987 20530 14021
rect 20564 13987 20583 14021
rect 20045 13981 20583 13987
rect 20514 13971 20583 13981
rect 20518 13969 20583 13971
rect 17932 13525 17992 13728
rect 19454 13724 20382 13769
rect 5310 13299 5370 13325
rect 4764 13099 4824 13125
rect 4882 13099 4942 13125
rect 5000 13099 5060 13125
rect 5118 13099 5178 13125
rect 4937 13044 5003 13052
rect 4568 13036 5003 13044
rect 4568 13002 4953 13036
rect 4987 13002 5003 13036
rect 4568 12993 5003 13002
rect 1793 12986 1859 12993
rect 4937 12986 5003 12993
rect 7700 13040 7760 13321
rect 8442 13295 8502 13321
rect 7896 13095 7956 13121
rect 8014 13095 8074 13121
rect 8132 13095 8192 13121
rect 8250 13095 8310 13121
rect 8069 13040 8135 13048
rect 7700 13032 8135 13040
rect 7700 12998 8085 13032
rect 8119 12998 8135 13032
rect 7700 12989 8135 12998
rect 10844 13040 10904 13321
rect 11586 13295 11646 13321
rect 11040 13095 11100 13121
rect 11158 13095 11218 13121
rect 11276 13095 11336 13121
rect 11394 13095 11454 13121
rect 11213 13040 11279 13048
rect 10844 13032 11279 13040
rect 10844 12998 11229 13032
rect 11263 12998 11279 13032
rect 10844 12989 11279 12998
rect 14046 13044 14106 13325
rect 14788 13299 14848 13325
rect 14242 13099 14302 13125
rect 14360 13099 14420 13125
rect 14478 13099 14538 13125
rect 14596 13099 14656 13125
rect 14415 13044 14481 13052
rect 14046 13036 14481 13044
rect 14046 13002 14431 13036
rect 14465 13002 14481 13036
rect 14046 12993 14481 13002
rect 17190 13044 17250 13325
rect 20322 13521 20382 13724
rect 20518 13521 20578 13969
rect 20633 13631 20699 13647
rect 20633 13597 20649 13631
rect 20683 13597 20699 13631
rect 20633 13581 20699 13597
rect 20636 13521 20696 13581
rect 20754 13521 20814 14080
rect 21339 14036 21399 14454
rect 21457 14428 21517 14454
rect 21662 14428 21722 14454
rect 21780 14428 21840 14454
rect 21898 14168 21958 14454
rect 21822 14151 21958 14168
rect 21822 14096 21841 14151
rect 21899 14096 21958 14151
rect 21822 14081 21958 14096
rect 20872 13979 21399 14036
rect 20872 13880 20932 13979
rect 20862 13867 20943 13880
rect 20862 13812 20872 13867
rect 20930 13812 20943 13867
rect 20862 13801 20943 13812
rect 20872 13521 20932 13801
rect 21898 13769 21958 14081
rect 21064 13724 21958 13769
rect 22598 14305 22658 14454
rect 22716 14428 22776 14454
rect 22834 14428 22894 14454
rect 23071 14428 23131 14454
rect 22702 14305 22768 14308
rect 22598 14292 22768 14305
rect 22598 14258 22718 14292
rect 22752 14258 22768 14292
rect 22598 14245 22768 14258
rect 22598 13769 22658 14245
rect 22702 14242 22768 14245
rect 23189 14038 23249 14454
rect 23307 14428 23367 14454
rect 23544 14428 23604 14454
rect 23662 14129 23722 14454
rect 23780 14428 23840 14454
rect 23898 14428 23958 14454
rect 24016 14428 24076 14454
rect 24134 14428 24194 14454
rect 24365 14428 24425 14454
rect 24016 14268 24075 14428
rect 24012 14267 24075 14268
rect 24012 14251 24078 14267
rect 24012 14217 24028 14251
rect 24062 14217 24078 14251
rect 24012 14201 24078 14217
rect 23880 14152 23975 14167
rect 23880 14129 23898 14152
rect 23662 14097 23898 14129
rect 23956 14097 23975 14152
rect 23662 14080 23975 14097
rect 23189 14021 23727 14038
rect 23189 13987 23674 14021
rect 23708 13987 23727 14021
rect 23189 13981 23727 13987
rect 23658 13971 23727 13981
rect 23662 13969 23727 13971
rect 22598 13724 23526 13769
rect 21064 13521 21124 13724
rect 23466 13521 23526 13724
rect 23662 13521 23722 13969
rect 23777 13631 23843 13647
rect 23777 13597 23793 13631
rect 23827 13597 23843 13631
rect 23777 13581 23843 13597
rect 23780 13521 23840 13581
rect 23898 13521 23958 14080
rect 24483 14036 24543 14454
rect 24601 14428 24661 14454
rect 24806 14428 24866 14454
rect 24924 14428 24984 14454
rect 25042 14168 25102 14454
rect 70455 14595 70494 14653
rect 71095 14649 71162 14653
rect 71483 14643 71562 14653
rect 71196 14595 71283 14612
rect 70455 14535 70509 14595
rect 70909 14535 70935 14595
rect 71196 14593 71842 14595
rect 71196 14535 71211 14593
rect 71266 14535 71842 14593
rect 72242 14535 72268 14595
rect 71196 14517 71283 14535
rect 70455 14417 70509 14477
rect 70909 14417 70935 14477
rect 70455 14359 70494 14417
rect 71234 14359 71283 14517
rect 71716 14477 71782 14480
rect 72315 14522 72381 14538
rect 72315 14488 72331 14522
rect 72365 14488 72381 14522
rect 71716 14464 71842 14477
rect 71716 14430 71732 14464
rect 71766 14430 71842 14464
rect 71716 14417 71842 14430
rect 72242 14417 72268 14477
rect 72315 14472 72381 14488
rect 71716 14414 71782 14417
rect 70455 14299 70509 14359
rect 70909 14299 71283 14359
rect 71325 14359 71394 14364
rect 71325 14345 71842 14359
rect 71325 14311 71342 14345
rect 71376 14311 71842 14345
rect 71325 14299 71842 14311
rect 72242 14299 72268 14359
rect 70455 14241 70494 14299
rect 71325 14295 71392 14299
rect 70455 14181 70509 14241
rect 70909 14181 70935 14241
rect 24966 14151 25102 14168
rect 24966 14096 24985 14151
rect 25043 14096 25102 14151
rect 24966 14081 25102 14096
rect 24016 13979 24543 14036
rect 24016 13880 24076 13979
rect 24006 13867 24087 13880
rect 24006 13812 24016 13867
rect 24074 13812 24087 13867
rect 24006 13801 24087 13812
rect 24016 13521 24076 13801
rect 25042 13769 25102 14081
rect 24208 13724 25102 13769
rect 70455 13944 70509 14004
rect 70909 13944 70935 14004
rect 70455 13886 70494 13944
rect 71325 13886 71382 14295
rect 72323 14163 72374 14472
rect 70455 13826 70509 13886
rect 70909 13826 71382 13886
rect 71594 14103 71842 14163
rect 72042 14103 72374 14163
rect 70455 13768 70494 13826
rect 24208 13521 24268 13724
rect 70455 13708 70509 13768
rect 70909 13708 70935 13768
rect 17932 13299 17992 13325
rect 17386 13099 17446 13125
rect 17504 13099 17564 13125
rect 17622 13099 17682 13125
rect 17740 13099 17800 13125
rect 17559 13044 17625 13052
rect 17190 13036 17625 13044
rect 17190 13002 17575 13036
rect 17609 13002 17625 13036
rect 17190 12993 17625 13002
rect 8069 12982 8135 12989
rect 11213 12982 11279 12989
rect 14415 12986 14481 12993
rect 17559 12986 17625 12993
rect 20322 13040 20382 13321
rect 21064 13295 21124 13321
rect 20518 13095 20578 13121
rect 20636 13095 20696 13121
rect 20754 13095 20814 13121
rect 20872 13095 20932 13121
rect 20691 13040 20757 13048
rect 20322 13032 20757 13040
rect 20322 12998 20707 13032
rect 20741 12998 20757 13032
rect 20322 12989 20757 12998
rect 23466 13040 23526 13321
rect 70654 13471 70709 13531
rect 70909 13471 70935 13531
rect 70654 13413 70693 13471
rect 70654 13353 70709 13413
rect 70909 13353 70935 13413
rect 71055 13389 71121 13405
rect 71055 13355 71071 13389
rect 71105 13355 71121 13389
rect 24208 13295 24268 13321
rect 70654 13295 70693 13353
rect 71055 13339 71121 13355
rect 71058 13295 71118 13339
rect 71594 13295 71639 14103
rect 70654 13235 70709 13295
rect 70909 13235 71639 13295
rect 30701 13145 30761 13161
rect 23662 13095 23722 13121
rect 23780 13095 23840 13121
rect 23898 13095 23958 13121
rect 24016 13095 24076 13121
rect 30128 13062 30154 13122
rect 30354 13062 30422 13122
rect 23835 13040 23901 13048
rect 23466 13032 23901 13040
rect 23466 12998 23851 13032
rect 23885 12998 23901 13032
rect 30371 13004 30422 13062
rect 23466 12989 23901 12998
rect 20691 12982 20757 12989
rect 23835 12982 23901 12989
rect 30128 12944 30154 13004
rect 30354 12997 30422 13004
rect 30701 13111 30715 13145
rect 30749 13111 30761 13145
rect 30701 12997 30761 13111
rect 30354 12944 31379 12997
rect 30371 12937 31379 12944
rect 31579 12937 31605 12997
rect 30371 12886 30422 12937
rect 30128 12826 30154 12886
rect 30354 12826 30422 12886
rect 31274 12896 31340 12937
rect 31274 12862 31290 12896
rect 31324 12862 31340 12896
rect 31274 12846 31340 12862
rect 30371 12638 30422 12826
rect 31207 12711 31273 12727
rect 29888 12578 29954 12638
rect 30354 12578 30422 12638
rect 30564 12635 30647 12695
rect 31047 12635 31073 12695
rect 31207 12677 31223 12711
rect 31257 12677 31273 12711
rect 31207 12660 31273 12677
rect 29888 12520 29939 12578
rect 30564 12577 30624 12635
rect 31214 12577 31273 12660
rect 29888 12460 29954 12520
rect 30354 12460 30380 12520
rect 30564 12517 30647 12577
rect 31047 12517 31379 12577
rect 31779 12517 31805 12577
rect 70654 12535 70709 12595
rect 70909 12536 71639 12595
rect 70909 12535 71212 12536
rect 29888 12402 29939 12460
rect 30564 12459 30624 12517
rect 31291 12459 31357 12461
rect 29888 12342 29954 12402
rect 30354 12342 30380 12402
rect 30564 12399 30647 12459
rect 31047 12399 31073 12459
rect 31291 12445 31379 12459
rect 31291 12411 31307 12445
rect 31341 12411 31379 12445
rect 31291 12399 31379 12411
rect 31779 12399 31805 12459
rect 70654 12477 70693 12535
rect 71195 12478 71212 12535
rect 71267 12535 71639 12536
rect 71267 12478 71282 12535
rect 31291 12395 31357 12399
rect 31291 12341 31356 12343
rect 1029 12139 1325 12178
rect 1029 12124 1089 12139
rect 1147 12124 1207 12139
rect 1265 12124 1325 12139
rect 1502 12139 1798 12178
rect 1502 12124 1562 12139
rect 1620 12124 1680 12139
rect 1738 12124 1798 12139
rect 1856 12139 2152 12178
rect 1856 12124 1916 12139
rect 1974 12124 2034 12139
rect 2092 12124 2152 12139
rect 2323 12139 2619 12178
rect 2323 12124 2383 12139
rect 2441 12124 2501 12139
rect 2559 12124 2619 12139
rect 4173 12139 4469 12178
rect 4173 12124 4233 12139
rect 4291 12124 4351 12139
rect 4409 12124 4469 12139
rect 4646 12139 4942 12178
rect 4646 12124 4706 12139
rect 4764 12124 4824 12139
rect 4882 12124 4942 12139
rect 5000 12139 5296 12178
rect 5000 12124 5060 12139
rect 5118 12124 5178 12139
rect 5236 12124 5296 12139
rect 5467 12139 5763 12178
rect 5467 12124 5527 12139
rect 5585 12124 5645 12139
rect 5703 12124 5763 12139
rect 7305 12135 7601 12174
rect 556 11940 852 11979
rect 556 11924 616 11940
rect 674 11924 734 11940
rect 792 11924 852 11940
rect 2764 11940 3060 11979
rect 2764 11924 2824 11940
rect 2882 11924 2942 11940
rect 3000 11924 3060 11940
rect 3700 11940 3996 11979
rect 3700 11924 3760 11940
rect 3818 11924 3878 11940
rect 3936 11924 3996 11940
rect 7305 12120 7365 12135
rect 7423 12120 7483 12135
rect 7541 12120 7601 12135
rect 7778 12135 8074 12174
rect 7778 12120 7838 12135
rect 7896 12120 7956 12135
rect 8014 12120 8074 12135
rect 8132 12135 8428 12174
rect 8132 12120 8192 12135
rect 8250 12120 8310 12135
rect 8368 12120 8428 12135
rect 8599 12135 8895 12174
rect 8599 12120 8659 12135
rect 8717 12120 8777 12135
rect 8835 12120 8895 12135
rect 10449 12135 10745 12174
rect 10449 12120 10509 12135
rect 10567 12120 10627 12135
rect 10685 12120 10745 12135
rect 10922 12135 11218 12174
rect 10922 12120 10982 12135
rect 11040 12120 11100 12135
rect 11158 12120 11218 12135
rect 11276 12135 11572 12174
rect 11276 12120 11336 12135
rect 11394 12120 11454 12135
rect 11512 12120 11572 12135
rect 11743 12135 12039 12174
rect 11743 12120 11803 12135
rect 11861 12120 11921 12135
rect 11979 12120 12039 12135
rect 13651 12139 13947 12178
rect 13651 12124 13711 12139
rect 13769 12124 13829 12139
rect 13887 12124 13947 12139
rect 14124 12139 14420 12178
rect 14124 12124 14184 12139
rect 14242 12124 14302 12139
rect 14360 12124 14420 12139
rect 14478 12139 14774 12178
rect 14478 12124 14538 12139
rect 14596 12124 14656 12139
rect 14714 12124 14774 12139
rect 14945 12139 15241 12178
rect 14945 12124 15005 12139
rect 15063 12124 15123 12139
rect 15181 12124 15241 12139
rect 16795 12139 17091 12178
rect 16795 12124 16855 12139
rect 16913 12124 16973 12139
rect 17031 12124 17091 12139
rect 17268 12139 17564 12178
rect 17268 12124 17328 12139
rect 17386 12124 17446 12139
rect 17504 12124 17564 12139
rect 17622 12139 17918 12178
rect 17622 12124 17682 12139
rect 17740 12124 17800 12139
rect 17858 12124 17918 12139
rect 18089 12139 18385 12178
rect 18089 12124 18149 12139
rect 18207 12124 18267 12139
rect 18325 12124 18385 12139
rect 19927 12135 20223 12174
rect 5908 11940 6204 11979
rect 5908 11924 5968 11940
rect 6026 11924 6086 11940
rect 6144 11924 6204 11940
rect 6832 11936 7128 11975
rect 6832 11920 6892 11936
rect 6950 11920 7010 11936
rect 7068 11920 7128 11936
rect 556 11575 616 11724
rect 674 11698 734 11724
rect 792 11698 852 11724
rect 1029 11698 1089 11724
rect 660 11575 726 11578
rect 556 11562 726 11575
rect 556 11528 676 11562
rect 710 11528 726 11562
rect 556 11515 726 11528
rect 556 11039 616 11515
rect 660 11512 726 11515
rect 1147 11308 1207 11724
rect 1265 11698 1325 11724
rect 1502 11698 1562 11724
rect 1620 11399 1680 11724
rect 1738 11698 1798 11724
rect 1856 11698 1916 11724
rect 1974 11698 2034 11724
rect 2092 11698 2152 11724
rect 2323 11698 2383 11724
rect 1974 11538 2033 11698
rect 1970 11537 2033 11538
rect 1970 11521 2036 11537
rect 1970 11487 1986 11521
rect 2020 11487 2036 11521
rect 1970 11471 2036 11487
rect 1838 11422 1933 11437
rect 1838 11399 1856 11422
rect 1620 11367 1856 11399
rect 1914 11367 1933 11422
rect 1620 11350 1933 11367
rect 1147 11291 1685 11308
rect 1147 11257 1632 11291
rect 1666 11257 1685 11291
rect 1147 11251 1685 11257
rect 1616 11241 1685 11251
rect 1620 11239 1685 11241
rect 556 10994 1484 11039
rect 1424 10791 1484 10994
rect 1620 10791 1680 11239
rect 1735 10901 1801 10917
rect 1735 10867 1751 10901
rect 1785 10867 1801 10901
rect 1735 10851 1801 10867
rect 1738 10791 1798 10851
rect 1856 10791 1916 11350
rect 2441 11306 2501 11724
rect 2559 11698 2619 11724
rect 2764 11698 2824 11724
rect 2882 11698 2942 11724
rect 3000 11438 3060 11724
rect 2924 11421 3060 11438
rect 2924 11366 2943 11421
rect 3001 11366 3060 11421
rect 2924 11351 3060 11366
rect 1974 11249 2501 11306
rect 1974 11150 2034 11249
rect 1964 11137 2045 11150
rect 1964 11082 1974 11137
rect 2032 11082 2045 11137
rect 1964 11071 2045 11082
rect 1974 10791 2034 11071
rect 3000 11039 3060 11351
rect 2166 10994 3060 11039
rect 3700 11575 3760 11724
rect 3818 11698 3878 11724
rect 3936 11698 3996 11724
rect 4173 11698 4233 11724
rect 3804 11575 3870 11578
rect 3700 11562 3870 11575
rect 3700 11528 3820 11562
rect 3854 11528 3870 11562
rect 3700 11515 3870 11528
rect 3700 11039 3760 11515
rect 3804 11512 3870 11515
rect 4291 11308 4351 11724
rect 4409 11698 4469 11724
rect 4646 11698 4706 11724
rect 4764 11399 4824 11724
rect 4882 11698 4942 11724
rect 5000 11698 5060 11724
rect 5118 11698 5178 11724
rect 5236 11698 5296 11724
rect 5467 11698 5527 11724
rect 5118 11538 5177 11698
rect 5114 11537 5177 11538
rect 5114 11521 5180 11537
rect 5114 11487 5130 11521
rect 5164 11487 5180 11521
rect 5114 11471 5180 11487
rect 4982 11422 5077 11437
rect 4982 11399 5000 11422
rect 4764 11367 5000 11399
rect 5058 11367 5077 11422
rect 4764 11350 5077 11367
rect 4291 11291 4829 11308
rect 4291 11257 4776 11291
rect 4810 11257 4829 11291
rect 4291 11251 4829 11257
rect 4760 11241 4829 11251
rect 4764 11239 4829 11241
rect 3700 10994 4628 11039
rect 2166 10791 2226 10994
rect 4568 10791 4628 10994
rect 4764 10791 4824 11239
rect 4879 10901 4945 10917
rect 4879 10867 4895 10901
rect 4929 10867 4945 10901
rect 4879 10851 4945 10867
rect 4882 10791 4942 10851
rect 5000 10791 5060 11350
rect 5585 11306 5645 11724
rect 5703 11698 5763 11724
rect 5908 11698 5968 11724
rect 6026 11698 6086 11724
rect 6144 11438 6204 11724
rect 9040 11936 9336 11975
rect 9040 11920 9100 11936
rect 9158 11920 9218 11936
rect 9276 11920 9336 11936
rect 9976 11936 10272 11975
rect 9976 11920 10036 11936
rect 10094 11920 10154 11936
rect 10212 11920 10272 11936
rect 12184 11936 12480 11975
rect 12184 11920 12244 11936
rect 12302 11920 12362 11936
rect 12420 11920 12480 11936
rect 13178 11940 13474 11979
rect 13178 11924 13238 11940
rect 13296 11924 13356 11940
rect 13414 11924 13474 11940
rect 15386 11940 15682 11979
rect 15386 11924 15446 11940
rect 15504 11924 15564 11940
rect 15622 11924 15682 11940
rect 16322 11940 16618 11979
rect 16322 11924 16382 11940
rect 16440 11924 16500 11940
rect 16558 11924 16618 11940
rect 19927 12120 19987 12135
rect 20045 12120 20105 12135
rect 20163 12120 20223 12135
rect 20400 12135 20696 12174
rect 20400 12120 20460 12135
rect 20518 12120 20578 12135
rect 20636 12120 20696 12135
rect 20754 12135 21050 12174
rect 20754 12120 20814 12135
rect 20872 12120 20932 12135
rect 20990 12120 21050 12135
rect 21221 12135 21517 12174
rect 21221 12120 21281 12135
rect 21339 12120 21399 12135
rect 21457 12120 21517 12135
rect 23071 12135 23367 12174
rect 23071 12120 23131 12135
rect 23189 12120 23249 12135
rect 23307 12120 23367 12135
rect 23544 12135 23840 12174
rect 23544 12120 23604 12135
rect 23662 12120 23722 12135
rect 23780 12120 23840 12135
rect 23898 12135 24194 12174
rect 23898 12120 23958 12135
rect 24016 12120 24076 12135
rect 24134 12120 24194 12135
rect 24365 12135 24661 12174
rect 24365 12120 24425 12135
rect 24483 12120 24543 12135
rect 24601 12120 24661 12135
rect 18530 11940 18826 11979
rect 18530 11924 18590 11940
rect 18648 11924 18708 11940
rect 18766 11924 18826 11940
rect 19454 11936 19750 11975
rect 19454 11920 19514 11936
rect 19572 11920 19632 11936
rect 19690 11920 19750 11936
rect 6068 11421 6204 11438
rect 6068 11366 6087 11421
rect 6145 11366 6204 11421
rect 6068 11351 6204 11366
rect 5118 11249 5645 11306
rect 5118 11150 5178 11249
rect 5108 11137 5189 11150
rect 5108 11082 5118 11137
rect 5176 11082 5189 11137
rect 5108 11071 5189 11082
rect 5118 10791 5178 11071
rect 6144 11039 6204 11351
rect 5310 10994 6204 11039
rect 6832 11571 6892 11720
rect 6950 11694 7010 11720
rect 7068 11694 7128 11720
rect 7305 11694 7365 11720
rect 6936 11571 7002 11574
rect 6832 11558 7002 11571
rect 6832 11524 6952 11558
rect 6986 11524 7002 11558
rect 6832 11511 7002 11524
rect 6832 11035 6892 11511
rect 6936 11508 7002 11511
rect 7423 11304 7483 11720
rect 7541 11694 7601 11720
rect 7778 11694 7838 11720
rect 7896 11395 7956 11720
rect 8014 11694 8074 11720
rect 8132 11694 8192 11720
rect 8250 11694 8310 11720
rect 8368 11694 8428 11720
rect 8599 11694 8659 11720
rect 8250 11534 8309 11694
rect 8246 11533 8309 11534
rect 8246 11517 8312 11533
rect 8246 11483 8262 11517
rect 8296 11483 8312 11517
rect 8246 11467 8312 11483
rect 8114 11418 8209 11433
rect 8114 11395 8132 11418
rect 7896 11363 8132 11395
rect 8190 11363 8209 11418
rect 7896 11346 8209 11363
rect 7423 11287 7961 11304
rect 7423 11253 7908 11287
rect 7942 11253 7961 11287
rect 7423 11247 7961 11253
rect 7892 11237 7961 11247
rect 7896 11235 7961 11237
rect 5310 10791 5370 10994
rect 6832 10990 7760 11035
rect 1424 10310 1484 10591
rect 2166 10565 2226 10591
rect 1620 10365 1680 10391
rect 1738 10365 1798 10391
rect 1856 10365 1916 10391
rect 1974 10365 2034 10391
rect 1793 10310 1859 10318
rect 1424 10302 1859 10310
rect 1424 10268 1809 10302
rect 1843 10268 1859 10302
rect 1424 10259 1859 10268
rect 4568 10310 4628 10591
rect 7700 10787 7760 10990
rect 7896 10787 7956 11235
rect 8011 10897 8077 10913
rect 8011 10863 8027 10897
rect 8061 10863 8077 10897
rect 8011 10847 8077 10863
rect 8014 10787 8074 10847
rect 8132 10787 8192 11346
rect 8717 11302 8777 11720
rect 8835 11694 8895 11720
rect 9040 11694 9100 11720
rect 9158 11694 9218 11720
rect 9276 11434 9336 11720
rect 9200 11417 9336 11434
rect 9200 11362 9219 11417
rect 9277 11362 9336 11417
rect 9200 11347 9336 11362
rect 8250 11245 8777 11302
rect 8250 11146 8310 11245
rect 8240 11133 8321 11146
rect 8240 11078 8250 11133
rect 8308 11078 8321 11133
rect 8240 11067 8321 11078
rect 8250 10787 8310 11067
rect 9276 11035 9336 11347
rect 8442 10990 9336 11035
rect 9976 11571 10036 11720
rect 10094 11694 10154 11720
rect 10212 11694 10272 11720
rect 10449 11694 10509 11720
rect 10080 11571 10146 11574
rect 9976 11558 10146 11571
rect 9976 11524 10096 11558
rect 10130 11524 10146 11558
rect 9976 11511 10146 11524
rect 9976 11035 10036 11511
rect 10080 11508 10146 11511
rect 10567 11304 10627 11720
rect 10685 11694 10745 11720
rect 10922 11694 10982 11720
rect 11040 11395 11100 11720
rect 11158 11694 11218 11720
rect 11276 11694 11336 11720
rect 11394 11694 11454 11720
rect 11512 11694 11572 11720
rect 11743 11694 11803 11720
rect 11394 11534 11453 11694
rect 11390 11533 11453 11534
rect 11390 11517 11456 11533
rect 11390 11483 11406 11517
rect 11440 11483 11456 11517
rect 11390 11467 11456 11483
rect 11258 11418 11353 11433
rect 11258 11395 11276 11418
rect 11040 11363 11276 11395
rect 11334 11363 11353 11418
rect 11040 11346 11353 11363
rect 10567 11287 11105 11304
rect 10567 11253 11052 11287
rect 11086 11253 11105 11287
rect 10567 11247 11105 11253
rect 11036 11237 11105 11247
rect 11040 11235 11105 11237
rect 9976 10990 10904 11035
rect 8442 10787 8502 10990
rect 10844 10787 10904 10990
rect 11040 10787 11100 11235
rect 11155 10897 11221 10913
rect 11155 10863 11171 10897
rect 11205 10863 11221 10897
rect 11155 10847 11221 10863
rect 11158 10787 11218 10847
rect 11276 10787 11336 11346
rect 11861 11302 11921 11720
rect 11979 11694 12039 11720
rect 12184 11694 12244 11720
rect 12302 11694 12362 11720
rect 12420 11434 12480 11720
rect 12344 11417 12480 11434
rect 12344 11362 12363 11417
rect 12421 11362 12480 11417
rect 12344 11347 12480 11362
rect 11394 11245 11921 11302
rect 11394 11146 11454 11245
rect 11384 11133 11465 11146
rect 11384 11078 11394 11133
rect 11452 11078 11465 11133
rect 11384 11067 11465 11078
rect 11394 10787 11454 11067
rect 12420 11035 12480 11347
rect 11586 10990 12480 11035
rect 13178 11575 13238 11724
rect 13296 11698 13356 11724
rect 13414 11698 13474 11724
rect 13651 11698 13711 11724
rect 13282 11575 13348 11578
rect 13178 11562 13348 11575
rect 13178 11528 13298 11562
rect 13332 11528 13348 11562
rect 13178 11515 13348 11528
rect 13178 11039 13238 11515
rect 13282 11512 13348 11515
rect 13769 11308 13829 11724
rect 13887 11698 13947 11724
rect 14124 11698 14184 11724
rect 14242 11399 14302 11724
rect 14360 11698 14420 11724
rect 14478 11698 14538 11724
rect 14596 11698 14656 11724
rect 14714 11698 14774 11724
rect 14945 11698 15005 11724
rect 14596 11538 14655 11698
rect 14592 11537 14655 11538
rect 14592 11521 14658 11537
rect 14592 11487 14608 11521
rect 14642 11487 14658 11521
rect 14592 11471 14658 11487
rect 14460 11422 14555 11437
rect 14460 11399 14478 11422
rect 14242 11367 14478 11399
rect 14536 11367 14555 11422
rect 14242 11350 14555 11367
rect 13769 11291 14307 11308
rect 13769 11257 14254 11291
rect 14288 11257 14307 11291
rect 13769 11251 14307 11257
rect 14238 11241 14307 11251
rect 14242 11239 14307 11241
rect 13178 10994 14106 11039
rect 11586 10787 11646 10990
rect 14046 10791 14106 10994
rect 14242 10791 14302 11239
rect 14357 10901 14423 10917
rect 14357 10867 14373 10901
rect 14407 10867 14423 10901
rect 14357 10851 14423 10867
rect 14360 10791 14420 10851
rect 14478 10791 14538 11350
rect 15063 11306 15123 11724
rect 15181 11698 15241 11724
rect 15386 11698 15446 11724
rect 15504 11698 15564 11724
rect 15622 11438 15682 11724
rect 15546 11421 15682 11438
rect 15546 11366 15565 11421
rect 15623 11366 15682 11421
rect 15546 11351 15682 11366
rect 14596 11249 15123 11306
rect 14596 11150 14656 11249
rect 14586 11137 14667 11150
rect 14586 11082 14596 11137
rect 14654 11082 14667 11137
rect 14586 11071 14667 11082
rect 14596 10791 14656 11071
rect 15622 11039 15682 11351
rect 14788 10994 15682 11039
rect 16322 11575 16382 11724
rect 16440 11698 16500 11724
rect 16558 11698 16618 11724
rect 16795 11698 16855 11724
rect 16426 11575 16492 11578
rect 16322 11562 16492 11575
rect 16322 11528 16442 11562
rect 16476 11528 16492 11562
rect 16322 11515 16492 11528
rect 16322 11039 16382 11515
rect 16426 11512 16492 11515
rect 16913 11308 16973 11724
rect 17031 11698 17091 11724
rect 17268 11698 17328 11724
rect 17386 11399 17446 11724
rect 17504 11698 17564 11724
rect 17622 11698 17682 11724
rect 17740 11698 17800 11724
rect 17858 11698 17918 11724
rect 18089 11698 18149 11724
rect 17740 11538 17799 11698
rect 17736 11537 17799 11538
rect 17736 11521 17802 11537
rect 17736 11487 17752 11521
rect 17786 11487 17802 11521
rect 17736 11471 17802 11487
rect 17604 11422 17699 11437
rect 17604 11399 17622 11422
rect 17386 11367 17622 11399
rect 17680 11367 17699 11422
rect 17386 11350 17699 11367
rect 16913 11291 17451 11308
rect 16913 11257 17398 11291
rect 17432 11257 17451 11291
rect 16913 11251 17451 11257
rect 17382 11241 17451 11251
rect 17386 11239 17451 11241
rect 16322 10994 17250 11039
rect 14788 10791 14848 10994
rect 17190 10791 17250 10994
rect 17386 10791 17446 11239
rect 17501 10901 17567 10917
rect 17501 10867 17517 10901
rect 17551 10867 17567 10901
rect 17501 10851 17567 10867
rect 17504 10791 17564 10851
rect 17622 10791 17682 11350
rect 18207 11306 18267 11724
rect 18325 11698 18385 11724
rect 18530 11698 18590 11724
rect 18648 11698 18708 11724
rect 18766 11438 18826 11724
rect 21662 11936 21958 11975
rect 21662 11920 21722 11936
rect 21780 11920 21840 11936
rect 21898 11920 21958 11936
rect 22598 11936 22894 11975
rect 22598 11920 22658 11936
rect 22716 11920 22776 11936
rect 22834 11920 22894 11936
rect 29928 12224 29954 12284
rect 30354 12224 30424 12284
rect 30373 12166 30424 12224
rect 29928 12106 29954 12166
rect 30354 12106 30424 12166
rect 30373 12048 30424 12106
rect 29928 11988 29954 12048
rect 30354 11988 30424 12048
rect 30563 12281 30647 12341
rect 31047 12281 31073 12341
rect 31291 12327 31379 12341
rect 31291 12293 31306 12327
rect 31340 12293 31379 12327
rect 31291 12281 31379 12293
rect 31779 12281 31805 12341
rect 30563 12223 30623 12281
rect 31291 12277 31356 12281
rect 70654 12417 70709 12477
rect 70909 12417 70935 12477
rect 71195 12459 71282 12478
rect 70654 12359 70693 12417
rect 70654 12299 70709 12359
rect 70909 12299 70935 12359
rect 30563 12163 30647 12223
rect 31047 12163 31379 12223
rect 31779 12163 31805 12223
rect 41616 12170 41912 12206
rect 30563 12105 30623 12163
rect 30563 12045 30647 12105
rect 31047 12045 31073 12105
rect 31214 12080 31273 12163
rect 41616 12149 41676 12170
rect 41734 12149 41794 12170
rect 41852 12149 41912 12170
rect 41970 12169 42266 12205
rect 41970 12149 42030 12169
rect 42088 12149 42148 12169
rect 42206 12149 42266 12169
rect 42324 12169 42620 12205
rect 42324 12149 42384 12169
rect 42442 12149 42502 12169
rect 42560 12149 42620 12169
rect 48165 12169 48461 12205
rect 31207 12063 31273 12080
rect 24806 11936 25102 11975
rect 24806 11920 24866 11936
rect 24924 11920 24984 11936
rect 25042 11920 25102 11936
rect 30373 11801 30424 11988
rect 31207 12029 31223 12063
rect 31257 12029 31273 12063
rect 31207 12013 31273 12029
rect 48165 12148 48225 12169
rect 48283 12148 48343 12169
rect 48401 12148 48461 12169
rect 48519 12168 48815 12204
rect 48519 12148 48579 12168
rect 48637 12148 48697 12168
rect 48755 12148 48815 12168
rect 48873 12168 49169 12204
rect 54819 12190 55115 12226
rect 54819 12169 54879 12190
rect 54937 12169 54997 12190
rect 55055 12169 55115 12190
rect 55173 12189 55469 12225
rect 55173 12169 55233 12189
rect 55291 12169 55351 12189
rect 55409 12169 55469 12189
rect 55527 12189 55823 12225
rect 55527 12169 55587 12189
rect 55645 12169 55705 12189
rect 55763 12169 55823 12189
rect 48873 12148 48933 12168
rect 48991 12148 49051 12168
rect 49109 12148 49169 12168
rect 41616 11923 41676 11949
rect 41734 11923 41794 11949
rect 41852 11923 41912 11949
rect 41970 11929 42030 11949
rect 41970 11923 42031 11929
rect 42088 11923 42148 11949
rect 42206 11923 42266 11949
rect 30086 11741 30154 11801
rect 30354 11741 30424 11801
rect 31275 11773 31341 11789
rect 30511 11751 30565 11767
rect 18690 11421 18826 11438
rect 18690 11366 18709 11421
rect 18767 11366 18826 11421
rect 18690 11351 18826 11366
rect 17740 11249 18267 11306
rect 17740 11150 17800 11249
rect 17730 11137 17811 11150
rect 17730 11082 17740 11137
rect 17798 11082 17811 11137
rect 17730 11071 17811 11082
rect 17740 10791 17800 11071
rect 18766 11039 18826 11351
rect 17932 10994 18826 11039
rect 19454 11571 19514 11720
rect 19572 11694 19632 11720
rect 19690 11694 19750 11720
rect 19927 11694 19987 11720
rect 19558 11571 19624 11574
rect 19454 11558 19624 11571
rect 19454 11524 19574 11558
rect 19608 11524 19624 11558
rect 19454 11511 19624 11524
rect 19454 11035 19514 11511
rect 19558 11508 19624 11511
rect 20045 11304 20105 11720
rect 20163 11694 20223 11720
rect 20400 11694 20460 11720
rect 20518 11395 20578 11720
rect 20636 11694 20696 11720
rect 20754 11694 20814 11720
rect 20872 11694 20932 11720
rect 20990 11694 21050 11720
rect 21221 11694 21281 11720
rect 20872 11534 20931 11694
rect 20868 11533 20931 11534
rect 20868 11517 20934 11533
rect 20868 11483 20884 11517
rect 20918 11483 20934 11517
rect 20868 11467 20934 11483
rect 20736 11418 20831 11433
rect 20736 11395 20754 11418
rect 20518 11363 20754 11395
rect 20812 11363 20831 11418
rect 20518 11346 20831 11363
rect 20045 11287 20583 11304
rect 20045 11253 20530 11287
rect 20564 11253 20583 11287
rect 20045 11247 20583 11253
rect 20514 11237 20583 11247
rect 20518 11235 20583 11237
rect 17932 10791 17992 10994
rect 19454 10990 20382 11035
rect 5310 10565 5370 10591
rect 4764 10365 4824 10391
rect 4882 10365 4942 10391
rect 5000 10365 5060 10391
rect 5118 10365 5178 10391
rect 4937 10310 5003 10318
rect 4568 10302 5003 10310
rect 4568 10268 4953 10302
rect 4987 10268 5003 10302
rect 4568 10259 5003 10268
rect 1793 10252 1859 10259
rect 4937 10252 5003 10259
rect 7700 10306 7760 10587
rect 8442 10561 8502 10587
rect 7896 10361 7956 10387
rect 8014 10361 8074 10387
rect 8132 10361 8192 10387
rect 8250 10361 8310 10387
rect 8069 10306 8135 10314
rect 7700 10298 8135 10306
rect 7700 10264 8085 10298
rect 8119 10264 8135 10298
rect 7700 10255 8135 10264
rect 10844 10306 10904 10587
rect 11586 10561 11646 10587
rect 11040 10361 11100 10387
rect 11158 10361 11218 10387
rect 11276 10361 11336 10387
rect 11394 10361 11454 10387
rect 11213 10306 11279 10314
rect 10844 10298 11279 10306
rect 10844 10264 11229 10298
rect 11263 10264 11279 10298
rect 10844 10255 11279 10264
rect 14046 10310 14106 10591
rect 14788 10565 14848 10591
rect 14242 10365 14302 10391
rect 14360 10365 14420 10391
rect 14478 10365 14538 10391
rect 14596 10365 14656 10391
rect 14415 10310 14481 10318
rect 14046 10302 14481 10310
rect 14046 10268 14431 10302
rect 14465 10268 14481 10302
rect 14046 10259 14481 10268
rect 17190 10310 17250 10591
rect 20322 10787 20382 10990
rect 20518 10787 20578 11235
rect 20633 10897 20699 10913
rect 20633 10863 20649 10897
rect 20683 10863 20699 10897
rect 20633 10847 20699 10863
rect 20636 10787 20696 10847
rect 20754 10787 20814 11346
rect 21339 11302 21399 11720
rect 21457 11694 21517 11720
rect 21662 11694 21722 11720
rect 21780 11694 21840 11720
rect 21898 11434 21958 11720
rect 21822 11417 21958 11434
rect 21822 11362 21841 11417
rect 21899 11362 21958 11417
rect 21822 11347 21958 11362
rect 20872 11245 21399 11302
rect 20872 11146 20932 11245
rect 20862 11133 20943 11146
rect 20862 11078 20872 11133
rect 20930 11078 20943 11133
rect 20862 11067 20943 11078
rect 20872 10787 20932 11067
rect 21898 11035 21958 11347
rect 21064 10990 21958 11035
rect 22598 11571 22658 11720
rect 22716 11694 22776 11720
rect 22834 11694 22894 11720
rect 23071 11694 23131 11720
rect 22702 11571 22768 11574
rect 22598 11558 22768 11571
rect 22598 11524 22718 11558
rect 22752 11524 22768 11558
rect 22598 11511 22768 11524
rect 22598 11035 22658 11511
rect 22702 11508 22768 11511
rect 23189 11304 23249 11720
rect 23307 11694 23367 11720
rect 23544 11694 23604 11720
rect 23662 11395 23722 11720
rect 23780 11694 23840 11720
rect 23898 11694 23958 11720
rect 24016 11694 24076 11720
rect 24134 11694 24194 11720
rect 24365 11694 24425 11720
rect 24016 11534 24075 11694
rect 24012 11533 24075 11534
rect 24012 11517 24078 11533
rect 24012 11483 24028 11517
rect 24062 11483 24078 11517
rect 24012 11467 24078 11483
rect 23880 11418 23975 11433
rect 23880 11395 23898 11418
rect 23662 11363 23898 11395
rect 23956 11363 23975 11418
rect 23662 11346 23975 11363
rect 23189 11287 23727 11304
rect 23189 11253 23674 11287
rect 23708 11253 23727 11287
rect 23189 11247 23727 11253
rect 23658 11237 23727 11247
rect 23662 11235 23727 11237
rect 22598 10990 23526 11035
rect 21064 10787 21124 10990
rect 23466 10787 23526 10990
rect 23662 10787 23722 11235
rect 23777 10897 23843 10913
rect 23777 10863 23793 10897
rect 23827 10863 23843 10897
rect 23777 10847 23843 10863
rect 23780 10787 23840 10847
rect 23898 10787 23958 11346
rect 24483 11302 24543 11720
rect 24601 11694 24661 11720
rect 24806 11694 24866 11720
rect 24924 11694 24984 11720
rect 25042 11434 25102 11720
rect 30086 11683 30137 11741
rect 30511 11717 30521 11751
rect 30555 11717 30565 11751
rect 30511 11699 30565 11717
rect 31275 11739 31291 11773
rect 31325 11739 31341 11773
rect 31275 11699 31341 11739
rect 41853 11738 41911 11923
rect 41853 11712 41913 11738
rect 41971 11712 42031 11923
rect 42324 11917 42384 11949
rect 42442 11923 42502 11949
rect 42560 11923 42620 11949
rect 70455 12094 70509 12154
rect 70909 12094 70935 12154
rect 63472 12023 63768 12059
rect 63472 12002 63532 12023
rect 63590 12002 63650 12023
rect 63708 12002 63768 12023
rect 63826 12022 64122 12058
rect 63826 12002 63886 12022
rect 63944 12002 64004 12022
rect 64062 12002 64122 12022
rect 64180 12022 64476 12058
rect 64180 12002 64240 12022
rect 64298 12002 64358 12022
rect 64416 12002 64476 12022
rect 70455 12036 70494 12094
rect 48165 11922 48225 11948
rect 48283 11922 48343 11948
rect 48401 11922 48461 11948
rect 48519 11928 48579 11948
rect 48519 11922 48580 11928
rect 48637 11922 48697 11948
rect 48755 11922 48815 11948
rect 42321 11901 42387 11917
rect 42321 11867 42337 11901
rect 42371 11867 42387 11901
rect 42321 11851 42387 11867
rect 42203 11784 42269 11800
rect 42203 11750 42219 11784
rect 42253 11750 42269 11784
rect 42203 11734 42269 11750
rect 48402 11737 48460 11922
rect 42206 11712 42266 11734
rect 30373 11683 31379 11699
rect 30086 11623 30154 11683
rect 30354 11639 31379 11683
rect 31579 11639 31605 11699
rect 30354 11624 30424 11639
rect 30354 11623 30380 11624
rect 30086 11565 30137 11623
rect 30086 11505 30154 11565
rect 30354 11505 30380 11565
rect 24966 11417 25102 11434
rect 24966 11362 24985 11417
rect 25043 11362 25102 11417
rect 24966 11347 25102 11362
rect 24016 11245 24543 11302
rect 24016 11146 24076 11245
rect 24006 11133 24087 11146
rect 24006 11078 24016 11133
rect 24074 11078 24087 11133
rect 24006 11067 24087 11078
rect 24016 10787 24076 11067
rect 25042 11035 25102 11347
rect 48402 11711 48462 11737
rect 48520 11711 48580 11922
rect 48873 11916 48933 11948
rect 48991 11922 49051 11948
rect 49109 11922 49169 11948
rect 54819 11943 54879 11969
rect 54937 11943 54997 11969
rect 55055 11943 55115 11969
rect 55173 11949 55233 11969
rect 55173 11943 55234 11949
rect 55291 11943 55351 11969
rect 55409 11943 55469 11969
rect 48870 11900 48936 11916
rect 48870 11866 48886 11900
rect 48920 11866 48936 11900
rect 48870 11850 48936 11866
rect 48752 11783 48818 11799
rect 48752 11749 48768 11783
rect 48802 11749 48818 11783
rect 48752 11733 48818 11749
rect 55056 11758 55114 11943
rect 48755 11711 48815 11733
rect 55056 11732 55116 11758
rect 55174 11732 55234 11943
rect 55527 11937 55587 11969
rect 55645 11943 55705 11969
rect 55763 11943 55823 11969
rect 55524 11921 55590 11937
rect 55524 11887 55540 11921
rect 55574 11887 55590 11921
rect 55524 11871 55590 11887
rect 55406 11804 55472 11820
rect 55406 11770 55422 11804
rect 55456 11770 55472 11804
rect 70455 11976 70509 12036
rect 70909 11976 71384 12036
rect 70455 11918 70494 11976
rect 65764 11812 66060 11863
rect 63472 11776 63532 11802
rect 63590 11776 63650 11802
rect 63708 11776 63768 11802
rect 63826 11782 63886 11802
rect 63826 11776 63887 11782
rect 63944 11776 64004 11802
rect 64062 11776 64122 11802
rect 55406 11754 55472 11770
rect 55409 11732 55469 11754
rect 42206 11486 42266 11512
rect 41853 11290 41913 11312
rect 41971 11290 42031 11312
rect 48755 11485 48815 11511
rect 63709 11591 63767 11776
rect 63709 11565 63769 11591
rect 63827 11565 63887 11776
rect 64180 11770 64240 11802
rect 64298 11776 64358 11802
rect 64416 11776 64476 11802
rect 65764 11797 65824 11812
rect 65882 11797 65942 11812
rect 66000 11797 66060 11812
rect 66118 11797 66178 11823
rect 66236 11797 66296 11823
rect 66354 11797 66414 11823
rect 70455 11858 70509 11918
rect 70909 11858 70935 11918
rect 64177 11754 64243 11770
rect 64177 11720 64193 11754
rect 64227 11720 64243 11754
rect 64177 11704 64243 11720
rect 64059 11637 64125 11653
rect 64059 11603 64075 11637
rect 64109 11603 64125 11637
rect 64059 11587 64125 11603
rect 65280 11597 65340 11623
rect 65398 11597 65458 11623
rect 65516 11597 65576 11623
rect 64062 11565 64122 11587
rect 55409 11506 55469 11532
rect 41850 11274 41916 11290
rect 41850 11240 41866 11274
rect 41900 11240 41916 11274
rect 41850 11224 41916 11240
rect 41968 11274 42034 11290
rect 48402 11289 48462 11311
rect 48520 11289 48580 11311
rect 55056 11310 55116 11332
rect 55174 11310 55234 11332
rect 55053 11294 55119 11310
rect 41968 11240 41984 11274
rect 42018 11240 42034 11274
rect 41968 11224 42034 11240
rect 48399 11273 48465 11289
rect 48399 11239 48415 11273
rect 48449 11239 48465 11273
rect 48399 11223 48465 11239
rect 48517 11273 48583 11289
rect 48517 11239 48533 11273
rect 48567 11239 48583 11273
rect 55053 11260 55069 11294
rect 55103 11260 55119 11294
rect 55053 11244 55119 11260
rect 55171 11294 55237 11310
rect 55171 11260 55187 11294
rect 55221 11260 55237 11294
rect 55171 11244 55237 11260
rect 48517 11223 48583 11239
rect 30699 11077 30759 11093
rect 66601 11614 66897 11665
rect 66601 11597 66661 11614
rect 66719 11597 66779 11614
rect 66837 11597 66897 11614
rect 67073 11615 67369 11651
rect 67073 11594 67133 11615
rect 67191 11594 67251 11615
rect 67309 11594 67369 11615
rect 67427 11614 67723 11650
rect 67427 11594 67487 11614
rect 67545 11594 67605 11614
rect 67663 11594 67723 11614
rect 67781 11614 68077 11650
rect 67781 11594 67841 11614
rect 67899 11594 67959 11614
rect 68017 11594 68077 11614
rect 70455 11627 70509 11687
rect 70909 11627 70935 11687
rect 65280 11380 65340 11397
rect 65398 11380 65458 11397
rect 65516 11380 65576 11397
rect 65764 11380 65824 11397
rect 64062 11339 64122 11365
rect 65280 11329 65824 11380
rect 65882 11371 65942 11397
rect 66000 11371 66060 11397
rect 66118 11378 66178 11397
rect 66236 11378 66296 11397
rect 66354 11378 66414 11397
rect 66601 11378 66661 11397
rect 66719 11378 66779 11397
rect 63709 11143 63769 11165
rect 63827 11143 63887 11165
rect 63706 11127 63772 11143
rect 63706 11093 63722 11127
rect 63756 11093 63772 11127
rect 63706 11077 63772 11093
rect 63824 11127 63890 11143
rect 63824 11093 63840 11127
rect 63874 11093 63890 11127
rect 63824 11077 63890 11093
rect 65405 11125 65465 11329
rect 66118 11327 66661 11378
rect 66703 11371 66779 11378
rect 66837 11371 66897 11397
rect 70455 11569 70494 11627
rect 70455 11509 70509 11569
rect 70909 11568 70935 11569
rect 71096 11568 71162 11571
rect 70909 11555 71162 11568
rect 70909 11521 71112 11555
rect 71146 11521 71162 11555
rect 70909 11509 71162 11521
rect 71327 11569 71384 11976
rect 71594 11761 71639 12535
rect 71594 11701 71842 11761
rect 72042 11701 72068 11761
rect 71483 11569 71562 11580
rect 71327 11567 71842 11569
rect 71327 11509 71496 11567
rect 71551 11509 71842 11567
rect 72242 11509 72268 11569
rect 66703 11327 66778 11371
rect 67073 11368 67133 11394
rect 67191 11368 67251 11394
rect 67309 11368 67369 11394
rect 67427 11374 67487 11394
rect 67427 11368 67488 11374
rect 67545 11368 67605 11394
rect 67663 11368 67723 11394
rect 66703 11245 66763 11327
rect 66703 11227 66937 11245
rect 66703 11193 66886 11227
rect 66920 11193 66937 11227
rect 65707 11127 66003 11187
rect 65405 11108 65536 11125
rect 24208 10990 25102 11035
rect 30126 10994 30152 11054
rect 30352 10994 30420 11054
rect 24208 10787 24268 10990
rect 30369 10936 30420 10994
rect 30126 10876 30152 10936
rect 30352 10929 30420 10936
rect 30699 11043 30713 11077
rect 30747 11043 30759 11077
rect 65405 11074 65486 11108
rect 65520 11074 65536 11108
rect 65707 11104 65767 11127
rect 65825 11104 65885 11127
rect 65943 11104 66003 11127
rect 66061 11128 66357 11188
rect 66061 11104 66121 11128
rect 66179 11104 66239 11128
rect 66297 11104 66357 11128
rect 66703 11177 66937 11193
rect 67310 11183 67368 11368
rect 65405 11057 65536 11074
rect 30699 10929 30759 11043
rect 30352 10876 31377 10929
rect 30369 10869 31377 10876
rect 31577 10869 31603 10929
rect 30369 10818 30420 10869
rect 17932 10565 17992 10591
rect 17386 10365 17446 10391
rect 17504 10365 17564 10391
rect 17622 10365 17682 10391
rect 17740 10365 17800 10391
rect 17559 10310 17625 10318
rect 17190 10302 17625 10310
rect 17190 10268 17575 10302
rect 17609 10268 17625 10302
rect 17190 10259 17625 10268
rect 8069 10248 8135 10255
rect 11213 10248 11279 10255
rect 14415 10252 14481 10259
rect 17559 10252 17625 10259
rect 20322 10306 20382 10587
rect 21064 10561 21124 10587
rect 20518 10361 20578 10387
rect 20636 10361 20696 10387
rect 20754 10361 20814 10387
rect 20872 10361 20932 10387
rect 20691 10306 20757 10314
rect 20322 10298 20757 10306
rect 20322 10264 20707 10298
rect 20741 10264 20757 10298
rect 20322 10255 20757 10264
rect 23466 10306 23526 10587
rect 30126 10758 30152 10818
rect 30352 10758 30420 10818
rect 31272 10828 31338 10869
rect 31272 10794 31288 10828
rect 31322 10794 31338 10828
rect 31272 10778 31338 10794
rect 24208 10561 24268 10587
rect 30369 10570 30420 10758
rect 31205 10643 31271 10659
rect 29886 10510 29952 10570
rect 30352 10510 30420 10570
rect 30562 10567 30645 10627
rect 31045 10567 31071 10627
rect 31205 10609 31221 10643
rect 31255 10609 31271 10643
rect 31205 10592 31271 10609
rect 29886 10452 29937 10510
rect 30562 10509 30622 10567
rect 31212 10509 31271 10592
rect 23662 10361 23722 10387
rect 23780 10361 23840 10387
rect 23898 10361 23958 10387
rect 24016 10361 24076 10387
rect 23835 10306 23901 10314
rect 23466 10298 23901 10306
rect 23466 10264 23851 10298
rect 23885 10264 23901 10298
rect 23466 10255 23901 10264
rect 20691 10248 20757 10255
rect 23835 10248 23901 10255
rect 29886 10392 29952 10452
rect 30352 10392 30378 10452
rect 30562 10449 30645 10509
rect 31045 10449 31377 10509
rect 31777 10449 31803 10509
rect 29886 10334 29937 10392
rect 30562 10391 30622 10449
rect 31289 10391 31355 10393
rect 29886 10274 29952 10334
rect 30352 10274 30378 10334
rect 30562 10331 30645 10391
rect 31045 10331 31071 10391
rect 31289 10377 31377 10391
rect 31289 10343 31305 10377
rect 31339 10343 31377 10377
rect 31289 10331 31377 10343
rect 31777 10331 31803 10391
rect 31289 10327 31355 10331
rect 31289 10273 31354 10275
rect 29926 10156 29952 10216
rect 30352 10156 30422 10216
rect 30371 10098 30422 10156
rect 29926 10038 29952 10098
rect 30352 10038 30422 10098
rect 30371 9980 30422 10038
rect 29926 9920 29952 9980
rect 30352 9920 30422 9980
rect 30561 10213 30645 10273
rect 31045 10213 31071 10273
rect 31289 10259 31377 10273
rect 31289 10225 31304 10259
rect 31338 10225 31377 10259
rect 31289 10213 31377 10225
rect 31777 10213 31803 10273
rect 34952 10270 35248 10306
rect 34952 10249 35012 10270
rect 35070 10249 35130 10270
rect 35188 10249 35248 10270
rect 35306 10269 35602 10305
rect 35306 10249 35366 10269
rect 35424 10249 35484 10269
rect 35542 10249 35602 10269
rect 35660 10269 35956 10305
rect 35660 10249 35720 10269
rect 35778 10249 35838 10269
rect 35896 10249 35956 10269
rect 30561 10155 30621 10213
rect 31289 10209 31354 10213
rect 30561 10095 30645 10155
rect 31045 10095 31377 10155
rect 31777 10095 31803 10155
rect 30561 10037 30621 10095
rect 30561 9977 30645 10037
rect 31045 9977 31071 10037
rect 31212 10012 31271 10095
rect 39990 10218 40056 10234
rect 41120 10224 41186 10240
rect 39990 10184 40006 10218
rect 40040 10211 40056 10218
rect 40040 10184 40565 10211
rect 39990 10168 40565 10184
rect 41120 10190 41136 10224
rect 41170 10215 41186 10224
rect 46539 10306 46605 10322
rect 47669 10312 47735 10328
rect 46539 10272 46555 10306
rect 46589 10299 46605 10306
rect 46589 10272 47114 10299
rect 46539 10256 47114 10272
rect 47669 10278 47685 10312
rect 47719 10303 47735 10312
rect 47719 10278 48256 10303
rect 47669 10260 48256 10278
rect 41170 10190 41707 10215
rect 47070 10204 47114 10256
rect 48212 10208 48256 10260
rect 41120 10172 41707 10190
rect 40521 10116 40565 10168
rect 41663 10120 41707 10172
rect 46539 10188 47012 10204
rect 46539 10154 46555 10188
rect 46589 10163 47012 10188
rect 46589 10162 46776 10163
rect 46589 10154 46605 10162
rect 46539 10138 46605 10154
rect 46716 10142 46776 10162
rect 46834 10142 46894 10163
rect 46952 10142 47012 10163
rect 47070 10163 47366 10204
rect 47070 10142 47130 10163
rect 47188 10142 47248 10163
rect 47306 10142 47366 10163
rect 47669 10192 48154 10208
rect 47669 10158 47685 10192
rect 47719 10167 48154 10192
rect 47719 10166 47918 10167
rect 47719 10158 47735 10166
rect 47669 10142 47735 10158
rect 47858 10146 47918 10166
rect 47976 10146 48036 10167
rect 48094 10146 48154 10167
rect 48212 10167 48508 10208
rect 53193 10238 53259 10254
rect 54323 10244 54389 10260
rect 53193 10204 53209 10238
rect 53243 10231 53259 10238
rect 53243 10204 53768 10231
rect 53193 10188 53768 10204
rect 54323 10210 54339 10244
rect 54373 10235 54389 10244
rect 59818 10306 59884 10322
rect 60948 10312 61014 10328
rect 59818 10272 59834 10306
rect 59868 10299 59884 10306
rect 59868 10272 60393 10299
rect 59818 10256 60393 10272
rect 60948 10278 60964 10312
rect 60998 10303 61014 10312
rect 65405 10477 65465 11057
rect 65707 10678 65767 10704
rect 65675 10537 65742 10544
rect 65825 10537 65885 10704
rect 65943 10678 66003 10704
rect 66061 10678 66121 10704
rect 65675 10528 65885 10537
rect 65675 10494 65691 10528
rect 65725 10494 65885 10528
rect 65675 10478 65885 10494
rect 65405 10461 65556 10477
rect 65405 10427 65506 10461
rect 65540 10427 65556 10461
rect 65405 10411 65556 10427
rect 65405 10372 65465 10411
rect 65825 10372 65885 10478
rect 66179 10537 66239 10704
rect 66297 10678 66357 10704
rect 66322 10537 66389 10544
rect 66179 10528 66389 10537
rect 66179 10494 66339 10528
rect 66373 10494 66389 10528
rect 66179 10478 66389 10494
rect 65941 10444 66007 10460
rect 65941 10410 65957 10444
rect 65991 10410 66007 10444
rect 65941 10394 66007 10410
rect 66059 10445 66125 10460
rect 66059 10411 66075 10445
rect 66109 10411 66125 10445
rect 66059 10395 66125 10411
rect 65943 10372 66003 10394
rect 66061 10372 66121 10395
rect 66179 10372 66239 10478
rect 66703 10476 66763 11177
rect 67310 11157 67370 11183
rect 67428 11157 67488 11368
rect 67781 11362 67841 11394
rect 67899 11368 67959 11394
rect 68017 11368 68077 11394
rect 67778 11346 67844 11362
rect 67778 11312 67794 11346
rect 67828 11312 67844 11346
rect 67778 11296 67844 11312
rect 70455 11451 70494 11509
rect 71095 11505 71162 11509
rect 71483 11499 71562 11509
rect 71196 11451 71283 11468
rect 70455 11391 70509 11451
rect 70909 11391 70935 11451
rect 71196 11449 71842 11451
rect 71196 11391 71211 11449
rect 71266 11391 71842 11449
rect 72242 11391 72268 11451
rect 71196 11373 71283 11391
rect 67660 11229 67726 11245
rect 67660 11195 67676 11229
rect 67710 11195 67726 11229
rect 70455 11273 70509 11333
rect 70909 11273 70935 11333
rect 70455 11215 70494 11273
rect 71234 11215 71283 11373
rect 71716 11333 71782 11336
rect 72315 11378 72381 11394
rect 72315 11344 72331 11378
rect 72365 11344 72381 11378
rect 71716 11320 71842 11333
rect 71716 11286 71732 11320
rect 71766 11286 71842 11320
rect 71716 11273 71842 11286
rect 72242 11273 72268 11333
rect 72315 11328 72381 11344
rect 71716 11270 71782 11273
rect 67660 11179 67726 11195
rect 67663 11157 67723 11179
rect 70455 11155 70509 11215
rect 70909 11155 71283 11215
rect 71325 11215 71394 11220
rect 71325 11201 71842 11215
rect 71325 11167 71342 11201
rect 71376 11167 71842 11201
rect 71325 11155 71842 11167
rect 72242 11155 72268 11215
rect 70455 11097 70494 11155
rect 71325 11151 71392 11155
rect 70455 11037 70509 11097
rect 70909 11037 70935 11097
rect 67663 10931 67723 10957
rect 70455 10800 70509 10860
rect 70909 10800 70935 10860
rect 67310 10735 67370 10757
rect 67428 10735 67488 10757
rect 70455 10742 70494 10800
rect 71325 10742 71382 11151
rect 72323 11019 72374 11328
rect 67307 10719 67373 10735
rect 67307 10685 67323 10719
rect 67357 10685 67373 10719
rect 67307 10669 67373 10685
rect 67425 10719 67491 10735
rect 67425 10685 67441 10719
rect 67475 10685 67491 10719
rect 67425 10669 67491 10685
rect 70455 10682 70509 10742
rect 70909 10682 71382 10742
rect 71594 10959 71842 11019
rect 72042 10959 72374 11019
rect 70455 10624 70494 10682
rect 70455 10564 70509 10624
rect 70909 10564 70935 10624
rect 66613 10460 66763 10476
rect 66613 10426 66629 10460
rect 66663 10426 66763 10460
rect 66613 10410 66763 10426
rect 66703 10372 66763 10410
rect 60998 10278 61535 10303
rect 60948 10260 61535 10278
rect 54373 10210 54910 10235
rect 54323 10192 54910 10210
rect 60349 10204 60393 10256
rect 61491 10208 61535 10260
rect 48212 10146 48272 10167
rect 48330 10146 48390 10167
rect 48448 10146 48508 10167
rect 39990 10100 40463 10116
rect 39990 10066 40006 10100
rect 40040 10075 40463 10100
rect 40040 10074 40227 10075
rect 40040 10066 40056 10074
rect 39990 10050 40056 10066
rect 40167 10054 40227 10074
rect 40285 10054 40345 10075
rect 40403 10054 40463 10075
rect 40521 10075 40817 10116
rect 40521 10054 40581 10075
rect 40639 10054 40699 10075
rect 40757 10054 40817 10075
rect 41120 10104 41605 10120
rect 41120 10070 41136 10104
rect 41170 10079 41605 10104
rect 41170 10078 41369 10079
rect 41170 10070 41186 10078
rect 41120 10054 41186 10070
rect 41309 10058 41369 10078
rect 41427 10058 41487 10079
rect 41545 10058 41605 10079
rect 41663 10079 41959 10120
rect 41663 10058 41723 10079
rect 41781 10058 41841 10079
rect 41899 10058 41959 10079
rect 44391 10091 44687 10127
rect 44391 10070 44451 10091
rect 44509 10070 44569 10091
rect 44627 10070 44687 10091
rect 44745 10090 45041 10126
rect 44745 10070 44805 10090
rect 44863 10070 44923 10090
rect 44981 10070 45041 10090
rect 45099 10090 45395 10126
rect 45099 10070 45159 10090
rect 45217 10070 45277 10090
rect 45335 10070 45395 10090
rect 34952 10023 35012 10049
rect 35070 10023 35130 10049
rect 35188 10023 35248 10049
rect 35306 10029 35366 10049
rect 35306 10023 35367 10029
rect 35424 10023 35484 10049
rect 35542 10023 35602 10049
rect 31205 9995 31271 10012
rect 30371 9733 30422 9920
rect 31205 9961 31221 9995
rect 31255 9961 31271 9995
rect 31205 9945 31271 9961
rect 35189 9838 35247 10023
rect 35189 9812 35249 9838
rect 35307 9812 35367 10023
rect 35660 10017 35720 10049
rect 35778 10023 35838 10049
rect 35896 10023 35956 10049
rect 35657 10001 35723 10017
rect 35657 9967 35673 10001
rect 35707 9967 35723 10001
rect 37842 10003 38138 10039
rect 37842 9982 37902 10003
rect 37960 9982 38020 10003
rect 38078 9982 38138 10003
rect 38196 10002 38492 10038
rect 38196 9982 38256 10002
rect 38314 9982 38374 10002
rect 38432 9982 38492 10002
rect 38550 10002 38846 10038
rect 38550 9982 38610 10002
rect 38668 9982 38728 10002
rect 38786 9982 38846 10002
rect 35657 9951 35723 9967
rect 35539 9884 35605 9900
rect 35539 9850 35555 9884
rect 35589 9850 35605 9884
rect 35539 9834 35605 9850
rect 35542 9812 35602 9834
rect 30084 9673 30152 9733
rect 30352 9673 30422 9733
rect 31273 9705 31339 9721
rect 30509 9683 30563 9699
rect 30084 9615 30135 9673
rect 30509 9649 30519 9683
rect 30553 9649 30563 9683
rect 30509 9631 30563 9649
rect 31273 9671 31289 9705
rect 31323 9671 31339 9705
rect 31273 9631 31339 9671
rect 30371 9615 31377 9631
rect 30084 9555 30152 9615
rect 30352 9571 31377 9615
rect 31577 9571 31603 9631
rect 30352 9556 30422 9571
rect 30352 9555 30378 9556
rect 30084 9497 30135 9555
rect 1039 9407 1335 9446
rect 1039 9392 1099 9407
rect 1157 9392 1217 9407
rect 1275 9392 1335 9407
rect 1512 9407 1808 9446
rect 1512 9392 1572 9407
rect 1630 9392 1690 9407
rect 1748 9392 1808 9407
rect 1866 9407 2162 9446
rect 1866 9392 1926 9407
rect 1984 9392 2044 9407
rect 2102 9392 2162 9407
rect 2333 9407 2629 9446
rect 2333 9392 2393 9407
rect 2451 9392 2511 9407
rect 2569 9392 2629 9407
rect 4183 9407 4479 9446
rect 4183 9392 4243 9407
rect 4301 9392 4361 9407
rect 4419 9392 4479 9407
rect 4656 9407 4952 9446
rect 4656 9392 4716 9407
rect 4774 9392 4834 9407
rect 4892 9392 4952 9407
rect 5010 9407 5306 9446
rect 5010 9392 5070 9407
rect 5128 9392 5188 9407
rect 5246 9392 5306 9407
rect 5477 9407 5773 9446
rect 5477 9392 5537 9407
rect 5595 9392 5655 9407
rect 5713 9392 5773 9407
rect 7315 9403 7611 9442
rect 566 9208 862 9247
rect 566 9192 626 9208
rect 684 9192 744 9208
rect 802 9192 862 9208
rect 2774 9208 3070 9247
rect 2774 9192 2834 9208
rect 2892 9192 2952 9208
rect 3010 9192 3070 9208
rect 3710 9208 4006 9247
rect 3710 9192 3770 9208
rect 3828 9192 3888 9208
rect 3946 9192 4006 9208
rect 7315 9388 7375 9403
rect 7433 9388 7493 9403
rect 7551 9388 7611 9403
rect 7788 9403 8084 9442
rect 7788 9388 7848 9403
rect 7906 9388 7966 9403
rect 8024 9388 8084 9403
rect 8142 9403 8438 9442
rect 8142 9388 8202 9403
rect 8260 9388 8320 9403
rect 8378 9388 8438 9403
rect 8609 9403 8905 9442
rect 8609 9388 8669 9403
rect 8727 9388 8787 9403
rect 8845 9388 8905 9403
rect 10459 9403 10755 9442
rect 10459 9388 10519 9403
rect 10577 9388 10637 9403
rect 10695 9388 10755 9403
rect 10932 9403 11228 9442
rect 10932 9388 10992 9403
rect 11050 9388 11110 9403
rect 11168 9388 11228 9403
rect 11286 9403 11582 9442
rect 11286 9388 11346 9403
rect 11404 9388 11464 9403
rect 11522 9388 11582 9403
rect 11753 9403 12049 9442
rect 11753 9388 11813 9403
rect 11871 9388 11931 9403
rect 11989 9388 12049 9403
rect 13661 9407 13957 9446
rect 13661 9392 13721 9407
rect 13779 9392 13839 9407
rect 13897 9392 13957 9407
rect 14134 9407 14430 9446
rect 14134 9392 14194 9407
rect 14252 9392 14312 9407
rect 14370 9392 14430 9407
rect 14488 9407 14784 9446
rect 14488 9392 14548 9407
rect 14606 9392 14666 9407
rect 14724 9392 14784 9407
rect 14955 9407 15251 9446
rect 14955 9392 15015 9407
rect 15073 9392 15133 9407
rect 15191 9392 15251 9407
rect 16805 9407 17101 9446
rect 16805 9392 16865 9407
rect 16923 9392 16983 9407
rect 17041 9392 17101 9407
rect 17278 9407 17574 9446
rect 17278 9392 17338 9407
rect 17396 9392 17456 9407
rect 17514 9392 17574 9407
rect 17632 9407 17928 9446
rect 17632 9392 17692 9407
rect 17750 9392 17810 9407
rect 17868 9392 17928 9407
rect 18099 9407 18395 9446
rect 18099 9392 18159 9407
rect 18217 9392 18277 9407
rect 18335 9392 18395 9407
rect 19937 9403 20233 9442
rect 5918 9208 6214 9247
rect 5918 9192 5978 9208
rect 6036 9192 6096 9208
rect 6154 9192 6214 9208
rect 6842 9204 7138 9243
rect 6842 9188 6902 9204
rect 6960 9188 7020 9204
rect 7078 9188 7138 9204
rect 566 8843 626 8992
rect 684 8966 744 8992
rect 802 8966 862 8992
rect 1039 8966 1099 8992
rect 670 8843 736 8846
rect 566 8830 736 8843
rect 566 8796 686 8830
rect 720 8796 736 8830
rect 566 8783 736 8796
rect 566 8307 626 8783
rect 670 8780 736 8783
rect 1157 8576 1217 8992
rect 1275 8966 1335 8992
rect 1512 8966 1572 8992
rect 1630 8667 1690 8992
rect 1748 8966 1808 8992
rect 1866 8966 1926 8992
rect 1984 8966 2044 8992
rect 2102 8966 2162 8992
rect 2333 8966 2393 8992
rect 1984 8806 2043 8966
rect 1980 8805 2043 8806
rect 1980 8789 2046 8805
rect 1980 8755 1996 8789
rect 2030 8755 2046 8789
rect 1980 8739 2046 8755
rect 1848 8690 1943 8705
rect 1848 8667 1866 8690
rect 1630 8635 1866 8667
rect 1924 8635 1943 8690
rect 1630 8618 1943 8635
rect 1157 8559 1695 8576
rect 1157 8525 1642 8559
rect 1676 8525 1695 8559
rect 1157 8519 1695 8525
rect 1626 8509 1695 8519
rect 1630 8507 1695 8509
rect 566 8262 1494 8307
rect 1434 8059 1494 8262
rect 1630 8059 1690 8507
rect 1745 8169 1811 8185
rect 1745 8135 1761 8169
rect 1795 8135 1811 8169
rect 1745 8119 1811 8135
rect 1748 8059 1808 8119
rect 1866 8059 1926 8618
rect 2451 8574 2511 8992
rect 2569 8966 2629 8992
rect 2774 8966 2834 8992
rect 2892 8966 2952 8992
rect 3010 8706 3070 8992
rect 2934 8689 3070 8706
rect 2934 8634 2953 8689
rect 3011 8634 3070 8689
rect 2934 8619 3070 8634
rect 1984 8517 2511 8574
rect 1984 8418 2044 8517
rect 1974 8405 2055 8418
rect 1974 8350 1984 8405
rect 2042 8350 2055 8405
rect 1974 8339 2055 8350
rect 1984 8059 2044 8339
rect 3010 8307 3070 8619
rect 2176 8262 3070 8307
rect 3710 8843 3770 8992
rect 3828 8966 3888 8992
rect 3946 8966 4006 8992
rect 4183 8966 4243 8992
rect 3814 8843 3880 8846
rect 3710 8830 3880 8843
rect 3710 8796 3830 8830
rect 3864 8796 3880 8830
rect 3710 8783 3880 8796
rect 3710 8307 3770 8783
rect 3814 8780 3880 8783
rect 4301 8576 4361 8992
rect 4419 8966 4479 8992
rect 4656 8966 4716 8992
rect 4774 8667 4834 8992
rect 4892 8966 4952 8992
rect 5010 8966 5070 8992
rect 5128 8966 5188 8992
rect 5246 8966 5306 8992
rect 5477 8966 5537 8992
rect 5128 8806 5187 8966
rect 5124 8805 5187 8806
rect 5124 8789 5190 8805
rect 5124 8755 5140 8789
rect 5174 8755 5190 8789
rect 5124 8739 5190 8755
rect 4992 8690 5087 8705
rect 4992 8667 5010 8690
rect 4774 8635 5010 8667
rect 5068 8635 5087 8690
rect 4774 8618 5087 8635
rect 4301 8559 4839 8576
rect 4301 8525 4786 8559
rect 4820 8525 4839 8559
rect 4301 8519 4839 8525
rect 4770 8509 4839 8519
rect 4774 8507 4839 8509
rect 3710 8262 4638 8307
rect 2176 8059 2236 8262
rect 4578 8059 4638 8262
rect 4774 8059 4834 8507
rect 4889 8169 4955 8185
rect 4889 8135 4905 8169
rect 4939 8135 4955 8169
rect 4889 8119 4955 8135
rect 4892 8059 4952 8119
rect 5010 8059 5070 8618
rect 5595 8574 5655 8992
rect 5713 8966 5773 8992
rect 5918 8966 5978 8992
rect 6036 8966 6096 8992
rect 6154 8706 6214 8992
rect 9050 9204 9346 9243
rect 9050 9188 9110 9204
rect 9168 9188 9228 9204
rect 9286 9188 9346 9204
rect 9986 9204 10282 9243
rect 9986 9188 10046 9204
rect 10104 9188 10164 9204
rect 10222 9188 10282 9204
rect 12194 9204 12490 9243
rect 12194 9188 12254 9204
rect 12312 9188 12372 9204
rect 12430 9188 12490 9204
rect 13188 9208 13484 9247
rect 13188 9192 13248 9208
rect 13306 9192 13366 9208
rect 13424 9192 13484 9208
rect 15396 9208 15692 9247
rect 15396 9192 15456 9208
rect 15514 9192 15574 9208
rect 15632 9192 15692 9208
rect 16332 9208 16628 9247
rect 16332 9192 16392 9208
rect 16450 9192 16510 9208
rect 16568 9192 16628 9208
rect 19937 9388 19997 9403
rect 20055 9388 20115 9403
rect 20173 9388 20233 9403
rect 20410 9403 20706 9442
rect 20410 9388 20470 9403
rect 20528 9388 20588 9403
rect 20646 9388 20706 9403
rect 20764 9403 21060 9442
rect 20764 9388 20824 9403
rect 20882 9388 20942 9403
rect 21000 9388 21060 9403
rect 21231 9403 21527 9442
rect 21231 9388 21291 9403
rect 21349 9388 21409 9403
rect 21467 9388 21527 9403
rect 23081 9403 23377 9442
rect 23081 9388 23141 9403
rect 23199 9388 23259 9403
rect 23317 9388 23377 9403
rect 23554 9403 23850 9442
rect 23554 9388 23614 9403
rect 23672 9388 23732 9403
rect 23790 9388 23850 9403
rect 23908 9403 24204 9442
rect 23908 9388 23968 9403
rect 24026 9388 24086 9403
rect 24144 9388 24204 9403
rect 24375 9403 24671 9442
rect 30084 9437 30152 9497
rect 30352 9437 30378 9497
rect 24375 9388 24435 9403
rect 24493 9388 24553 9403
rect 24611 9388 24671 9403
rect 37842 9756 37902 9782
rect 37960 9756 38020 9782
rect 38078 9756 38138 9782
rect 38196 9762 38256 9782
rect 38196 9756 38257 9762
rect 38314 9756 38374 9782
rect 38432 9756 38492 9782
rect 35542 9586 35602 9612
rect 38079 9571 38137 9756
rect 38079 9545 38139 9571
rect 38197 9545 38257 9756
rect 38550 9750 38610 9782
rect 38668 9756 38728 9782
rect 38786 9756 38846 9782
rect 38547 9734 38613 9750
rect 38547 9700 38563 9734
rect 38597 9700 38613 9734
rect 38547 9684 38613 9700
rect 44391 9844 44451 9870
rect 44509 9844 44569 9870
rect 44627 9844 44687 9870
rect 44745 9850 44805 9870
rect 44745 9844 44806 9850
rect 44863 9844 44923 9870
rect 44981 9844 45041 9870
rect 44628 9659 44686 9844
rect 40167 9637 40227 9654
rect 38429 9617 38495 9633
rect 38429 9583 38445 9617
rect 38479 9583 38495 9617
rect 38429 9567 38495 9583
rect 38432 9545 38492 9567
rect 40167 9548 40228 9637
rect 40285 9628 40345 9654
rect 40403 9628 40463 9654
rect 18540 9208 18836 9247
rect 18540 9192 18600 9208
rect 18658 9192 18718 9208
rect 18776 9192 18836 9208
rect 19464 9204 19760 9243
rect 19464 9188 19524 9204
rect 19582 9188 19642 9204
rect 19700 9188 19760 9204
rect 6078 8689 6214 8706
rect 6078 8634 6097 8689
rect 6155 8634 6214 8689
rect 6078 8619 6214 8634
rect 5128 8517 5655 8574
rect 5128 8418 5188 8517
rect 5118 8405 5199 8418
rect 5118 8350 5128 8405
rect 5186 8350 5199 8405
rect 5118 8339 5199 8350
rect 5128 8059 5188 8339
rect 6154 8307 6214 8619
rect 5320 8262 6214 8307
rect 6842 8839 6902 8988
rect 6960 8962 7020 8988
rect 7078 8962 7138 8988
rect 7315 8962 7375 8988
rect 6946 8839 7012 8842
rect 6842 8826 7012 8839
rect 6842 8792 6962 8826
rect 6996 8792 7012 8826
rect 6842 8779 7012 8792
rect 6842 8303 6902 8779
rect 6946 8776 7012 8779
rect 7433 8572 7493 8988
rect 7551 8962 7611 8988
rect 7788 8962 7848 8988
rect 7906 8663 7966 8988
rect 8024 8962 8084 8988
rect 8142 8962 8202 8988
rect 8260 8962 8320 8988
rect 8378 8962 8438 8988
rect 8609 8962 8669 8988
rect 8260 8802 8319 8962
rect 8256 8801 8319 8802
rect 8256 8785 8322 8801
rect 8256 8751 8272 8785
rect 8306 8751 8322 8785
rect 8256 8735 8322 8751
rect 8124 8686 8219 8701
rect 8124 8663 8142 8686
rect 7906 8631 8142 8663
rect 8200 8631 8219 8686
rect 7906 8614 8219 8631
rect 7433 8555 7971 8572
rect 7433 8521 7918 8555
rect 7952 8521 7971 8555
rect 7433 8515 7971 8521
rect 7902 8505 7971 8515
rect 7906 8503 7971 8505
rect 5320 8059 5380 8262
rect 6842 8258 7770 8303
rect 1434 7578 1494 7859
rect 2176 7833 2236 7859
rect 1630 7633 1690 7659
rect 1748 7633 1808 7659
rect 1866 7633 1926 7659
rect 1984 7633 2044 7659
rect 1803 7578 1869 7586
rect 1434 7570 1869 7578
rect 1434 7536 1819 7570
rect 1853 7536 1869 7570
rect 1434 7527 1869 7536
rect 4578 7578 4638 7859
rect 7710 8055 7770 8258
rect 7906 8055 7966 8503
rect 8021 8165 8087 8181
rect 8021 8131 8037 8165
rect 8071 8131 8087 8165
rect 8021 8115 8087 8131
rect 8024 8055 8084 8115
rect 8142 8055 8202 8614
rect 8727 8570 8787 8988
rect 8845 8962 8905 8988
rect 9050 8962 9110 8988
rect 9168 8962 9228 8988
rect 9286 8702 9346 8988
rect 9210 8685 9346 8702
rect 9210 8630 9229 8685
rect 9287 8630 9346 8685
rect 9210 8615 9346 8630
rect 8260 8513 8787 8570
rect 8260 8414 8320 8513
rect 8250 8401 8331 8414
rect 8250 8346 8260 8401
rect 8318 8346 8331 8401
rect 8250 8335 8331 8346
rect 8260 8055 8320 8335
rect 9286 8303 9346 8615
rect 8452 8258 9346 8303
rect 9986 8839 10046 8988
rect 10104 8962 10164 8988
rect 10222 8962 10282 8988
rect 10459 8962 10519 8988
rect 10090 8839 10156 8842
rect 9986 8826 10156 8839
rect 9986 8792 10106 8826
rect 10140 8792 10156 8826
rect 9986 8779 10156 8792
rect 9986 8303 10046 8779
rect 10090 8776 10156 8779
rect 10577 8572 10637 8988
rect 10695 8962 10755 8988
rect 10932 8962 10992 8988
rect 11050 8663 11110 8988
rect 11168 8962 11228 8988
rect 11286 8962 11346 8988
rect 11404 8962 11464 8988
rect 11522 8962 11582 8988
rect 11753 8962 11813 8988
rect 11404 8802 11463 8962
rect 11400 8801 11463 8802
rect 11400 8785 11466 8801
rect 11400 8751 11416 8785
rect 11450 8751 11466 8785
rect 11400 8735 11466 8751
rect 11268 8686 11363 8701
rect 11268 8663 11286 8686
rect 11050 8631 11286 8663
rect 11344 8631 11363 8686
rect 11050 8614 11363 8631
rect 10577 8555 11115 8572
rect 10577 8521 11062 8555
rect 11096 8521 11115 8555
rect 10577 8515 11115 8521
rect 11046 8505 11115 8515
rect 11050 8503 11115 8505
rect 9986 8258 10914 8303
rect 8452 8055 8512 8258
rect 10854 8055 10914 8258
rect 11050 8055 11110 8503
rect 11165 8165 11231 8181
rect 11165 8131 11181 8165
rect 11215 8131 11231 8165
rect 11165 8115 11231 8131
rect 11168 8055 11228 8115
rect 11286 8055 11346 8614
rect 11871 8570 11931 8988
rect 11989 8962 12049 8988
rect 12194 8962 12254 8988
rect 12312 8962 12372 8988
rect 12430 8702 12490 8988
rect 12354 8685 12490 8702
rect 12354 8630 12373 8685
rect 12431 8630 12490 8685
rect 12354 8615 12490 8630
rect 11404 8513 11931 8570
rect 11404 8414 11464 8513
rect 11394 8401 11475 8414
rect 11394 8346 11404 8401
rect 11462 8346 11475 8401
rect 11394 8335 11475 8346
rect 11404 8055 11464 8335
rect 12430 8303 12490 8615
rect 11596 8258 12490 8303
rect 13188 8843 13248 8992
rect 13306 8966 13366 8992
rect 13424 8966 13484 8992
rect 13661 8966 13721 8992
rect 13292 8843 13358 8846
rect 13188 8830 13358 8843
rect 13188 8796 13308 8830
rect 13342 8796 13358 8830
rect 13188 8783 13358 8796
rect 13188 8307 13248 8783
rect 13292 8780 13358 8783
rect 13779 8576 13839 8992
rect 13897 8966 13957 8992
rect 14134 8966 14194 8992
rect 14252 8667 14312 8992
rect 14370 8966 14430 8992
rect 14488 8966 14548 8992
rect 14606 8966 14666 8992
rect 14724 8966 14784 8992
rect 14955 8966 15015 8992
rect 14606 8806 14665 8966
rect 14602 8805 14665 8806
rect 14602 8789 14668 8805
rect 14602 8755 14618 8789
rect 14652 8755 14668 8789
rect 14602 8739 14668 8755
rect 14470 8690 14565 8705
rect 14470 8667 14488 8690
rect 14252 8635 14488 8667
rect 14546 8635 14565 8690
rect 14252 8618 14565 8635
rect 13779 8559 14317 8576
rect 13779 8525 14264 8559
rect 14298 8525 14317 8559
rect 13779 8519 14317 8525
rect 14248 8509 14317 8519
rect 14252 8507 14317 8509
rect 13188 8262 14116 8307
rect 11596 8055 11656 8258
rect 14056 8059 14116 8262
rect 14252 8059 14312 8507
rect 14367 8169 14433 8185
rect 14367 8135 14383 8169
rect 14417 8135 14433 8169
rect 14367 8119 14433 8135
rect 14370 8059 14430 8119
rect 14488 8059 14548 8618
rect 15073 8574 15133 8992
rect 15191 8966 15251 8992
rect 15396 8966 15456 8992
rect 15514 8966 15574 8992
rect 15632 8706 15692 8992
rect 15556 8689 15692 8706
rect 15556 8634 15575 8689
rect 15633 8634 15692 8689
rect 15556 8619 15692 8634
rect 14606 8517 15133 8574
rect 14606 8418 14666 8517
rect 14596 8405 14677 8418
rect 14596 8350 14606 8405
rect 14664 8350 14677 8405
rect 14596 8339 14677 8350
rect 14606 8059 14666 8339
rect 15632 8307 15692 8619
rect 14798 8262 15692 8307
rect 16332 8843 16392 8992
rect 16450 8966 16510 8992
rect 16568 8966 16628 8992
rect 16805 8966 16865 8992
rect 16436 8843 16502 8846
rect 16332 8830 16502 8843
rect 16332 8796 16452 8830
rect 16486 8796 16502 8830
rect 16332 8783 16502 8796
rect 16332 8307 16392 8783
rect 16436 8780 16502 8783
rect 16923 8576 16983 8992
rect 17041 8966 17101 8992
rect 17278 8966 17338 8992
rect 17396 8667 17456 8992
rect 17514 8966 17574 8992
rect 17632 8966 17692 8992
rect 17750 8966 17810 8992
rect 17868 8966 17928 8992
rect 18099 8966 18159 8992
rect 17750 8806 17809 8966
rect 17746 8805 17809 8806
rect 17746 8789 17812 8805
rect 17746 8755 17762 8789
rect 17796 8755 17812 8789
rect 17746 8739 17812 8755
rect 17614 8690 17709 8705
rect 17614 8667 17632 8690
rect 17396 8635 17632 8667
rect 17690 8635 17709 8690
rect 17396 8618 17709 8635
rect 16923 8559 17461 8576
rect 16923 8525 17408 8559
rect 17442 8525 17461 8559
rect 16923 8519 17461 8525
rect 17392 8509 17461 8519
rect 17396 8507 17461 8509
rect 16332 8262 17260 8307
rect 14798 8059 14858 8262
rect 17200 8059 17260 8262
rect 17396 8059 17456 8507
rect 17511 8169 17577 8185
rect 17511 8135 17527 8169
rect 17561 8135 17577 8169
rect 17511 8119 17577 8135
rect 17514 8059 17574 8119
rect 17632 8059 17692 8618
rect 18217 8574 18277 8992
rect 18335 8966 18395 8992
rect 18540 8966 18600 8992
rect 18658 8966 18718 8992
rect 18776 8706 18836 8992
rect 21672 9204 21968 9243
rect 21672 9188 21732 9204
rect 21790 9188 21850 9204
rect 21908 9188 21968 9204
rect 22608 9204 22904 9243
rect 22608 9188 22668 9204
rect 22726 9188 22786 9204
rect 22844 9188 22904 9204
rect 35189 9390 35249 9412
rect 35307 9390 35367 9412
rect 35186 9374 35252 9390
rect 35186 9340 35202 9374
rect 35236 9340 35252 9374
rect 35186 9324 35252 9340
rect 35304 9374 35370 9390
rect 35304 9340 35320 9374
rect 35354 9340 35370 9374
rect 35304 9324 35370 9340
rect 24816 9204 25112 9243
rect 24816 9188 24876 9204
rect 24934 9188 24994 9204
rect 25052 9188 25112 9204
rect 40077 9495 40228 9548
rect 38432 9319 38492 9345
rect 40077 9271 40137 9495
rect 40521 9453 40581 9654
rect 40639 9628 40699 9654
rect 40757 9628 40817 9654
rect 41309 9641 41369 9658
rect 41309 9552 41370 9641
rect 41427 9632 41487 9658
rect 41545 9632 41605 9658
rect 40195 9402 40581 9453
rect 41219 9499 41370 9552
rect 40195 9271 40255 9402
rect 40310 9344 40376 9360
rect 40310 9310 40326 9344
rect 40360 9310 40376 9344
rect 40310 9294 40376 9310
rect 40313 9271 40373 9294
rect 40596 9271 40656 9297
rect 40714 9271 40774 9297
rect 40832 9271 40892 9297
rect 41219 9275 41279 9499
rect 41663 9457 41723 9658
rect 41781 9632 41841 9658
rect 41899 9632 41959 9658
rect 44628 9633 44688 9659
rect 44746 9633 44806 9844
rect 45099 9838 45159 9870
rect 45217 9844 45277 9870
rect 45335 9844 45395 9870
rect 45096 9822 45162 9838
rect 45096 9788 45112 9822
rect 45146 9788 45162 9822
rect 45096 9772 45162 9788
rect 53724 10136 53768 10188
rect 54866 10140 54910 10192
rect 59818 10188 60291 10204
rect 59818 10154 59834 10188
rect 59868 10163 60291 10188
rect 59868 10162 60055 10163
rect 59868 10154 59884 10162
rect 53193 10120 53666 10136
rect 53193 10086 53209 10120
rect 53243 10095 53666 10120
rect 53243 10094 53430 10095
rect 53243 10086 53259 10094
rect 53193 10070 53259 10086
rect 53370 10074 53430 10094
rect 53488 10074 53548 10095
rect 53606 10074 53666 10095
rect 53724 10095 54020 10136
rect 53724 10074 53784 10095
rect 53842 10074 53902 10095
rect 53960 10074 54020 10095
rect 54323 10124 54808 10140
rect 54323 10090 54339 10124
rect 54373 10099 54808 10124
rect 54373 10098 54572 10099
rect 54373 10090 54389 10098
rect 54323 10074 54389 10090
rect 54512 10078 54572 10098
rect 54630 10078 54690 10099
rect 54748 10078 54808 10099
rect 54866 10099 55162 10140
rect 59818 10138 59884 10154
rect 59995 10142 60055 10162
rect 60113 10142 60173 10163
rect 60231 10142 60291 10163
rect 60349 10163 60645 10204
rect 60349 10142 60409 10163
rect 60467 10142 60527 10163
rect 60585 10142 60645 10163
rect 60948 10192 61433 10208
rect 60948 10158 60964 10192
rect 60998 10167 61433 10192
rect 60998 10166 61197 10167
rect 60998 10158 61014 10166
rect 60948 10142 61014 10158
rect 61137 10146 61197 10166
rect 61255 10146 61315 10167
rect 61373 10146 61433 10167
rect 61491 10167 61787 10208
rect 61491 10146 61551 10167
rect 61609 10146 61669 10167
rect 61727 10146 61787 10167
rect 65405 10146 65465 10172
rect 54866 10078 54926 10099
rect 54984 10078 55044 10099
rect 55102 10078 55162 10099
rect 57670 10091 57966 10127
rect 51045 10023 51341 10059
rect 51045 10002 51105 10023
rect 51163 10002 51223 10023
rect 51281 10002 51341 10023
rect 51399 10022 51695 10058
rect 51399 10002 51459 10022
rect 51517 10002 51577 10022
rect 51635 10002 51695 10022
rect 51753 10022 52049 10058
rect 51753 10002 51813 10022
rect 51871 10002 51931 10022
rect 51989 10002 52049 10022
rect 51045 9776 51105 9802
rect 51163 9776 51223 9802
rect 51281 9776 51341 9802
rect 51399 9782 51459 9802
rect 51399 9776 51460 9782
rect 51517 9776 51577 9802
rect 51635 9776 51695 9802
rect 46716 9725 46776 9742
rect 44978 9705 45044 9721
rect 44978 9671 44994 9705
rect 45028 9671 45044 9705
rect 44978 9655 45044 9671
rect 44981 9633 45041 9655
rect 46716 9636 46777 9725
rect 46834 9716 46894 9742
rect 46952 9716 47012 9742
rect 41337 9406 41723 9457
rect 41337 9275 41397 9406
rect 41452 9348 41518 9364
rect 41452 9314 41468 9348
rect 41502 9314 41518 9348
rect 41452 9298 41518 9314
rect 41455 9275 41515 9298
rect 41738 9275 41798 9301
rect 41856 9275 41916 9301
rect 41974 9275 42034 9301
rect 38079 9123 38139 9145
rect 38197 9123 38257 9145
rect 38076 9107 38142 9123
rect 38076 9073 38092 9107
rect 38126 9073 38142 9107
rect 38076 9057 38142 9073
rect 38194 9107 38260 9123
rect 38194 9073 38210 9107
rect 38244 9073 38260 9107
rect 38194 9057 38260 9073
rect 46626 9583 46777 9636
rect 44981 9407 45041 9433
rect 46626 9359 46686 9583
rect 47070 9541 47130 9742
rect 47188 9716 47248 9742
rect 47306 9716 47366 9742
rect 47858 9729 47918 9746
rect 47858 9640 47919 9729
rect 47976 9720 48036 9746
rect 48094 9720 48154 9746
rect 46744 9490 47130 9541
rect 47768 9587 47919 9640
rect 46744 9359 46804 9490
rect 46859 9432 46925 9448
rect 46859 9398 46875 9432
rect 46909 9398 46925 9432
rect 46859 9382 46925 9398
rect 46862 9359 46922 9382
rect 47145 9359 47205 9385
rect 47263 9359 47323 9385
rect 47381 9359 47441 9385
rect 47768 9363 47828 9587
rect 48212 9545 48272 9746
rect 48330 9720 48390 9746
rect 48448 9720 48508 9746
rect 51282 9591 51340 9776
rect 51282 9565 51342 9591
rect 51400 9565 51460 9776
rect 51753 9770 51813 9802
rect 51871 9776 51931 9802
rect 51989 9776 52049 9802
rect 51750 9754 51816 9770
rect 51750 9720 51766 9754
rect 51800 9720 51816 9754
rect 51750 9704 51816 9720
rect 57670 10070 57730 10091
rect 57788 10070 57848 10091
rect 57906 10070 57966 10091
rect 58024 10090 58320 10126
rect 58024 10070 58084 10090
rect 58142 10070 58202 10090
rect 58260 10070 58320 10090
rect 58378 10090 58674 10126
rect 58378 10070 58438 10090
rect 58496 10070 58556 10090
rect 58614 10070 58674 10090
rect 57670 9844 57730 9870
rect 57788 9844 57848 9870
rect 57906 9844 57966 9870
rect 58024 9850 58084 9870
rect 58024 9844 58085 9850
rect 58142 9844 58202 9870
rect 58260 9844 58320 9870
rect 53370 9657 53430 9674
rect 51632 9637 51698 9653
rect 51632 9603 51648 9637
rect 51682 9603 51698 9637
rect 51632 9587 51698 9603
rect 51635 9565 51695 9587
rect 53370 9568 53431 9657
rect 53488 9648 53548 9674
rect 53606 9648 53666 9674
rect 47886 9494 48272 9545
rect 47886 9363 47946 9494
rect 48001 9436 48067 9452
rect 48001 9402 48017 9436
rect 48051 9402 48067 9436
rect 48001 9386 48067 9402
rect 48004 9363 48064 9386
rect 48287 9363 48347 9389
rect 48405 9363 48465 9389
rect 48523 9363 48583 9389
rect 44628 9211 44688 9233
rect 44746 9211 44806 9233
rect 44625 9195 44691 9211
rect 44625 9161 44641 9195
rect 44675 9161 44691 9195
rect 44625 9145 44691 9161
rect 44743 9195 44809 9211
rect 44743 9161 44759 9195
rect 44793 9161 44809 9195
rect 44743 9145 44809 9161
rect 53280 9515 53431 9568
rect 51635 9339 51695 9365
rect 53280 9291 53340 9515
rect 53724 9473 53784 9674
rect 53842 9648 53902 9674
rect 53960 9648 54020 9674
rect 54512 9661 54572 9678
rect 54512 9572 54573 9661
rect 54630 9652 54690 9678
rect 54748 9652 54808 9678
rect 53398 9422 53784 9473
rect 54422 9519 54573 9572
rect 53398 9291 53458 9422
rect 53513 9364 53579 9380
rect 53513 9330 53529 9364
rect 53563 9330 53579 9364
rect 53513 9314 53579 9330
rect 53516 9291 53576 9314
rect 53799 9291 53859 9317
rect 53917 9291 53977 9317
rect 54035 9291 54095 9317
rect 54422 9295 54482 9519
rect 54866 9477 54926 9678
rect 54984 9652 55044 9678
rect 55102 9652 55162 9678
rect 57907 9659 57965 9844
rect 57907 9633 57967 9659
rect 58025 9633 58085 9844
rect 58378 9838 58438 9870
rect 58496 9844 58556 9870
rect 58614 9844 58674 9870
rect 58375 9822 58441 9838
rect 58375 9788 58391 9822
rect 58425 9788 58441 9822
rect 58375 9772 58441 9788
rect 70654 10327 70709 10387
rect 70909 10327 70935 10387
rect 70654 10269 70693 10327
rect 70654 10209 70709 10269
rect 70909 10209 70935 10269
rect 71055 10245 71121 10261
rect 71055 10211 71071 10245
rect 71105 10211 71121 10245
rect 66703 10146 66763 10172
rect 70654 10151 70693 10209
rect 71055 10195 71121 10211
rect 71058 10151 71118 10195
rect 71594 10151 71639 10959
rect 70654 10091 70709 10151
rect 70909 10091 71639 10151
rect 65825 9946 65885 9972
rect 65943 9946 66003 9972
rect 66061 9946 66121 9972
rect 66179 9946 66239 9972
rect 59995 9725 60055 9742
rect 58257 9705 58323 9721
rect 58257 9671 58273 9705
rect 58307 9671 58323 9705
rect 58257 9655 58323 9671
rect 58260 9633 58320 9655
rect 59995 9636 60056 9725
rect 60113 9716 60173 9742
rect 60231 9716 60291 9742
rect 54540 9426 54926 9477
rect 54540 9295 54600 9426
rect 54655 9368 54721 9384
rect 54655 9334 54671 9368
rect 54705 9334 54721 9368
rect 54655 9318 54721 9334
rect 54658 9295 54718 9318
rect 54941 9295 55001 9321
rect 55059 9295 55119 9321
rect 55177 9295 55237 9321
rect 46626 9133 46686 9159
rect 46744 9133 46804 9159
rect 46862 9127 46922 9159
rect 47145 9127 47205 9159
rect 47263 9127 47323 9159
rect 47381 9127 47441 9159
rect 47768 9137 47828 9163
rect 47886 9137 47946 9163
rect 46862 9086 47441 9127
rect 48004 9131 48064 9163
rect 48287 9131 48347 9163
rect 48405 9131 48465 9163
rect 48523 9131 48583 9163
rect 51282 9143 51342 9165
rect 51400 9143 51460 9165
rect 48004 9090 48583 9131
rect 51279 9127 51345 9143
rect 51279 9093 51295 9127
rect 51329 9093 51345 9127
rect 51279 9077 51345 9093
rect 51397 9127 51463 9143
rect 51397 9093 51413 9127
rect 51447 9093 51463 9127
rect 51397 9077 51463 9093
rect 59905 9583 60056 9636
rect 58260 9407 58320 9433
rect 59905 9359 59965 9583
rect 60349 9541 60409 9742
rect 60467 9716 60527 9742
rect 60585 9716 60645 9742
rect 61137 9729 61197 9746
rect 61137 9640 61198 9729
rect 61255 9720 61315 9746
rect 61373 9720 61433 9746
rect 60023 9490 60409 9541
rect 61047 9587 61198 9640
rect 60023 9359 60083 9490
rect 60138 9432 60204 9448
rect 60138 9398 60154 9432
rect 60188 9398 60204 9432
rect 60138 9382 60204 9398
rect 60141 9359 60201 9382
rect 60424 9359 60484 9385
rect 60542 9359 60602 9385
rect 60660 9359 60720 9385
rect 61047 9363 61107 9587
rect 61491 9545 61551 9746
rect 61609 9720 61669 9746
rect 61727 9720 61787 9746
rect 61165 9494 61551 9545
rect 61165 9363 61225 9494
rect 63467 9452 63763 9488
rect 61280 9436 61346 9452
rect 61280 9402 61296 9436
rect 61330 9402 61346 9436
rect 63467 9431 63527 9452
rect 63585 9431 63645 9452
rect 63703 9431 63763 9452
rect 63821 9451 64117 9487
rect 63821 9431 63881 9451
rect 63939 9431 63999 9451
rect 64057 9431 64117 9451
rect 64175 9451 64471 9487
rect 64175 9431 64235 9451
rect 64293 9431 64353 9451
rect 64411 9431 64471 9451
rect 61280 9386 61346 9402
rect 61283 9363 61343 9386
rect 61566 9363 61626 9389
rect 61684 9363 61744 9389
rect 61802 9363 61862 9389
rect 57907 9211 57967 9233
rect 58025 9211 58085 9233
rect 57904 9195 57970 9211
rect 57904 9161 57920 9195
rect 57954 9161 57970 9195
rect 57904 9145 57970 9161
rect 58022 9195 58088 9211
rect 58022 9161 58038 9195
rect 58072 9161 58088 9195
rect 58022 9145 58088 9161
rect 70658 9333 70713 9393
rect 70913 9334 71643 9393
rect 70913 9333 71216 9334
rect 70658 9275 70697 9333
rect 71199 9276 71216 9333
rect 71271 9333 71643 9334
rect 71271 9276 71286 9333
rect 63467 9205 63527 9231
rect 63585 9205 63645 9231
rect 63703 9205 63763 9231
rect 63821 9211 63881 9231
rect 63821 9205 63882 9211
rect 63939 9205 63999 9231
rect 64057 9205 64117 9231
rect 59905 9133 59965 9159
rect 60023 9133 60083 9159
rect 60141 9127 60201 9159
rect 60424 9127 60484 9159
rect 60542 9127 60602 9159
rect 60660 9127 60720 9159
rect 61047 9137 61107 9163
rect 61165 9137 61225 9163
rect 40077 9045 40137 9071
rect 40195 9045 40255 9071
rect 40313 9039 40373 9071
rect 40596 9039 40656 9071
rect 40714 9039 40774 9071
rect 40832 9039 40892 9071
rect 41219 9049 41279 9075
rect 41337 9049 41397 9075
rect 18700 8689 18836 8706
rect 18700 8634 18719 8689
rect 18777 8634 18836 8689
rect 18700 8619 18836 8634
rect 17750 8517 18277 8574
rect 17750 8418 17810 8517
rect 17740 8405 17821 8418
rect 17740 8350 17750 8405
rect 17808 8350 17821 8405
rect 17740 8339 17821 8350
rect 17750 8059 17810 8339
rect 18776 8307 18836 8619
rect 17942 8262 18836 8307
rect 19464 8839 19524 8988
rect 19582 8962 19642 8988
rect 19700 8962 19760 8988
rect 19937 8962 19997 8988
rect 19568 8839 19634 8842
rect 19464 8826 19634 8839
rect 19464 8792 19584 8826
rect 19618 8792 19634 8826
rect 19464 8779 19634 8792
rect 19464 8303 19524 8779
rect 19568 8776 19634 8779
rect 20055 8572 20115 8988
rect 20173 8962 20233 8988
rect 20410 8962 20470 8988
rect 20528 8663 20588 8988
rect 20646 8962 20706 8988
rect 20764 8962 20824 8988
rect 20882 8962 20942 8988
rect 21000 8962 21060 8988
rect 21231 8962 21291 8988
rect 20882 8802 20941 8962
rect 20878 8801 20941 8802
rect 20878 8785 20944 8801
rect 20878 8751 20894 8785
rect 20928 8751 20944 8785
rect 20878 8735 20944 8751
rect 20746 8686 20841 8701
rect 20746 8663 20764 8686
rect 20528 8631 20764 8663
rect 20822 8631 20841 8686
rect 20528 8614 20841 8631
rect 20055 8555 20593 8572
rect 20055 8521 20540 8555
rect 20574 8521 20593 8555
rect 20055 8515 20593 8521
rect 20524 8505 20593 8515
rect 20528 8503 20593 8505
rect 17942 8059 18002 8262
rect 19464 8258 20392 8303
rect 5320 7833 5380 7859
rect 4774 7633 4834 7659
rect 4892 7633 4952 7659
rect 5010 7633 5070 7659
rect 5128 7633 5188 7659
rect 4947 7578 5013 7586
rect 4578 7570 5013 7578
rect 4578 7536 4963 7570
rect 4997 7536 5013 7570
rect 4578 7527 5013 7536
rect 1803 7520 1869 7527
rect 4947 7520 5013 7527
rect 7710 7574 7770 7855
rect 8452 7829 8512 7855
rect 7906 7629 7966 7655
rect 8024 7629 8084 7655
rect 8142 7629 8202 7655
rect 8260 7629 8320 7655
rect 8079 7574 8145 7582
rect 7710 7566 8145 7574
rect 7710 7532 8095 7566
rect 8129 7532 8145 7566
rect 7710 7523 8145 7532
rect 10854 7574 10914 7855
rect 11596 7829 11656 7855
rect 11050 7629 11110 7655
rect 11168 7629 11228 7655
rect 11286 7629 11346 7655
rect 11404 7629 11464 7655
rect 11223 7574 11289 7582
rect 10854 7566 11289 7574
rect 10854 7532 11239 7566
rect 11273 7532 11289 7566
rect 10854 7523 11289 7532
rect 14056 7578 14116 7859
rect 14798 7833 14858 7859
rect 14252 7633 14312 7659
rect 14370 7633 14430 7659
rect 14488 7633 14548 7659
rect 14606 7633 14666 7659
rect 14425 7578 14491 7586
rect 14056 7570 14491 7578
rect 14056 7536 14441 7570
rect 14475 7536 14491 7570
rect 14056 7527 14491 7536
rect 17200 7578 17260 7859
rect 20332 8055 20392 8258
rect 20528 8055 20588 8503
rect 20643 8165 20709 8181
rect 20643 8131 20659 8165
rect 20693 8131 20709 8165
rect 20643 8115 20709 8131
rect 20646 8055 20706 8115
rect 20764 8055 20824 8614
rect 21349 8570 21409 8988
rect 21467 8962 21527 8988
rect 21672 8962 21732 8988
rect 21790 8962 21850 8988
rect 21908 8702 21968 8988
rect 21832 8685 21968 8702
rect 21832 8630 21851 8685
rect 21909 8630 21968 8685
rect 21832 8615 21968 8630
rect 20882 8513 21409 8570
rect 20882 8414 20942 8513
rect 20872 8401 20953 8414
rect 20872 8346 20882 8401
rect 20940 8346 20953 8401
rect 20872 8335 20953 8346
rect 20882 8055 20942 8335
rect 21908 8303 21968 8615
rect 21074 8258 21968 8303
rect 22608 8839 22668 8988
rect 22726 8962 22786 8988
rect 22844 8962 22904 8988
rect 23081 8962 23141 8988
rect 22712 8839 22778 8842
rect 22608 8826 22778 8839
rect 22608 8792 22728 8826
rect 22762 8792 22778 8826
rect 22608 8779 22778 8792
rect 22608 8303 22668 8779
rect 22712 8776 22778 8779
rect 23199 8572 23259 8988
rect 23317 8962 23377 8988
rect 23554 8962 23614 8988
rect 23672 8663 23732 8988
rect 23790 8962 23850 8988
rect 23908 8962 23968 8988
rect 24026 8962 24086 8988
rect 24144 8962 24204 8988
rect 24375 8962 24435 8988
rect 24026 8802 24085 8962
rect 24022 8801 24085 8802
rect 24022 8785 24088 8801
rect 24022 8751 24038 8785
rect 24072 8751 24088 8785
rect 24022 8735 24088 8751
rect 23890 8686 23985 8701
rect 23890 8663 23908 8686
rect 23672 8631 23908 8663
rect 23966 8631 23985 8686
rect 23672 8614 23985 8631
rect 23199 8555 23737 8572
rect 23199 8521 23684 8555
rect 23718 8521 23737 8555
rect 23199 8515 23737 8521
rect 23668 8505 23737 8515
rect 23672 8503 23737 8505
rect 22608 8258 23536 8303
rect 21074 8055 21134 8258
rect 23476 8055 23536 8258
rect 23672 8055 23732 8503
rect 23787 8165 23853 8181
rect 23787 8131 23803 8165
rect 23837 8131 23853 8165
rect 23787 8115 23853 8131
rect 23790 8055 23850 8115
rect 23908 8055 23968 8614
rect 24493 8570 24553 8988
rect 24611 8962 24671 8988
rect 24816 8962 24876 8988
rect 24934 8962 24994 8988
rect 25052 8702 25112 8988
rect 30701 9008 30761 9024
rect 30128 8925 30154 8985
rect 30354 8925 30422 8985
rect 30371 8867 30422 8925
rect 30128 8807 30154 8867
rect 30354 8860 30422 8867
rect 30701 8974 30715 9008
rect 30749 8974 30761 9008
rect 40313 8998 40892 9039
rect 41455 9043 41515 9075
rect 41738 9043 41798 9075
rect 41856 9043 41916 9075
rect 41974 9043 42034 9075
rect 53280 9065 53340 9091
rect 53398 9065 53458 9091
rect 41455 9002 42034 9043
rect 53516 9059 53576 9091
rect 53799 9059 53859 9091
rect 53917 9059 53977 9091
rect 54035 9059 54095 9091
rect 54422 9069 54482 9095
rect 54540 9069 54600 9095
rect 53516 9018 54095 9059
rect 54658 9063 54718 9095
rect 54941 9063 55001 9095
rect 55059 9063 55119 9095
rect 55177 9063 55237 9095
rect 60141 9086 60720 9127
rect 61283 9131 61343 9163
rect 61566 9131 61626 9163
rect 61684 9131 61744 9163
rect 61802 9131 61862 9163
rect 61283 9090 61862 9131
rect 54658 9022 55237 9063
rect 63704 9020 63762 9205
rect 63704 8994 63764 9020
rect 63822 8994 63882 9205
rect 64175 9199 64235 9231
rect 64293 9205 64353 9231
rect 64411 9205 64471 9231
rect 70658 9215 70713 9275
rect 70913 9215 70939 9275
rect 71199 9257 71286 9276
rect 64172 9183 64238 9199
rect 64172 9149 64188 9183
rect 64222 9149 64238 9183
rect 64172 9133 64238 9149
rect 70658 9157 70697 9215
rect 70658 9097 70713 9157
rect 70913 9097 70939 9157
rect 64054 9066 64120 9082
rect 64054 9032 64070 9066
rect 64104 9032 64120 9066
rect 64054 9016 64120 9032
rect 64057 8994 64117 9016
rect 30701 8860 30761 8974
rect 30354 8807 31379 8860
rect 30371 8800 31379 8807
rect 31579 8800 31605 8860
rect 30371 8749 30422 8800
rect 24976 8685 25112 8702
rect 30128 8689 30154 8749
rect 30354 8689 30422 8749
rect 31274 8759 31340 8800
rect 31274 8725 31290 8759
rect 31324 8725 31340 8759
rect 31274 8709 31340 8725
rect 24976 8630 24995 8685
rect 25053 8630 25112 8685
rect 24976 8615 25112 8630
rect 24026 8513 24553 8570
rect 24026 8414 24086 8513
rect 24016 8401 24097 8414
rect 24016 8346 24026 8401
rect 24084 8346 24097 8401
rect 24016 8335 24097 8346
rect 24026 8055 24086 8335
rect 25052 8303 25112 8615
rect 30371 8501 30422 8689
rect 31207 8574 31273 8590
rect 29888 8441 29954 8501
rect 30354 8441 30422 8501
rect 30564 8498 30647 8558
rect 31047 8498 31073 8558
rect 31207 8540 31223 8574
rect 31257 8540 31273 8574
rect 31207 8523 31273 8540
rect 29888 8383 29939 8441
rect 30564 8440 30624 8498
rect 31214 8440 31273 8523
rect 70459 8892 70513 8952
rect 70913 8892 70939 8952
rect 70459 8834 70498 8892
rect 64057 8768 64117 8794
rect 70459 8774 70513 8834
rect 70913 8774 71388 8834
rect 70459 8716 70498 8774
rect 70459 8656 70513 8716
rect 70913 8656 70939 8716
rect 63704 8572 63764 8594
rect 63822 8572 63882 8594
rect 63701 8556 63767 8572
rect 63701 8522 63717 8556
rect 63751 8522 63767 8556
rect 44405 8441 44701 8477
rect 24218 8258 25112 8303
rect 24218 8055 24278 8258
rect 29888 8323 29954 8383
rect 30354 8323 30380 8383
rect 30564 8380 30647 8440
rect 31047 8380 31379 8440
rect 31779 8380 31805 8440
rect 44405 8420 44465 8441
rect 44523 8420 44583 8441
rect 44641 8420 44701 8441
rect 44759 8440 45055 8476
rect 44759 8420 44819 8440
rect 44877 8420 44937 8440
rect 44995 8420 45055 8440
rect 45113 8440 45409 8476
rect 45113 8420 45173 8440
rect 45231 8420 45291 8440
rect 45349 8420 45409 8440
rect 29888 8265 29939 8323
rect 30564 8322 30624 8380
rect 31291 8322 31357 8324
rect 29888 8205 29954 8265
rect 30354 8205 30380 8265
rect 30564 8262 30647 8322
rect 31047 8262 31073 8322
rect 31291 8308 31379 8322
rect 31291 8274 31307 8308
rect 31341 8274 31379 8308
rect 31291 8262 31379 8274
rect 31779 8262 31805 8322
rect 37856 8353 38152 8389
rect 37856 8332 37916 8353
rect 37974 8332 38034 8353
rect 38092 8332 38152 8353
rect 38210 8352 38506 8388
rect 38210 8332 38270 8352
rect 38328 8332 38388 8352
rect 38446 8332 38506 8352
rect 38564 8352 38860 8388
rect 38564 8332 38624 8352
rect 38682 8332 38742 8352
rect 38800 8332 38860 8352
rect 31291 8258 31357 8262
rect 31291 8204 31356 8206
rect 17942 7833 18002 7859
rect 17396 7633 17456 7659
rect 17514 7633 17574 7659
rect 17632 7633 17692 7659
rect 17750 7633 17810 7659
rect 17569 7578 17635 7586
rect 17200 7570 17635 7578
rect 17200 7536 17585 7570
rect 17619 7536 17635 7570
rect 17200 7527 17635 7536
rect 8079 7516 8145 7523
rect 11223 7516 11289 7523
rect 14425 7520 14491 7527
rect 17569 7520 17635 7527
rect 20332 7574 20392 7855
rect 21074 7829 21134 7855
rect 20528 7629 20588 7655
rect 20646 7629 20706 7655
rect 20764 7629 20824 7655
rect 20882 7629 20942 7655
rect 20701 7574 20767 7582
rect 20332 7566 20767 7574
rect 20332 7532 20717 7566
rect 20751 7532 20767 7566
rect 20332 7523 20767 7532
rect 23476 7574 23536 7855
rect 29928 8087 29954 8147
rect 30354 8087 30424 8147
rect 30373 8029 30424 8087
rect 29928 7969 29954 8029
rect 30354 7969 30424 8029
rect 30373 7911 30424 7969
rect 24218 7829 24278 7855
rect 29928 7851 29954 7911
rect 30354 7851 30424 7911
rect 30563 8144 30647 8204
rect 31047 8144 31073 8204
rect 31291 8190 31379 8204
rect 31291 8156 31306 8190
rect 31340 8156 31379 8190
rect 31291 8144 31379 8156
rect 31779 8144 31805 8204
rect 30563 8086 30623 8144
rect 31291 8140 31356 8144
rect 63701 8506 63767 8522
rect 63819 8556 63885 8572
rect 63819 8522 63835 8556
rect 63869 8522 63885 8556
rect 63819 8506 63885 8522
rect 57684 8441 57980 8477
rect 57684 8420 57744 8441
rect 57802 8420 57862 8441
rect 57920 8420 57980 8441
rect 58038 8440 58334 8476
rect 58038 8420 58098 8440
rect 58156 8420 58216 8440
rect 58274 8420 58334 8440
rect 58392 8440 58688 8476
rect 58392 8420 58452 8440
rect 58510 8420 58570 8440
rect 58628 8420 58688 8440
rect 51059 8373 51355 8409
rect 51059 8352 51119 8373
rect 51177 8352 51237 8373
rect 51295 8352 51355 8373
rect 51413 8372 51709 8408
rect 51413 8352 51473 8372
rect 51531 8352 51591 8372
rect 51649 8352 51709 8372
rect 51767 8372 52063 8408
rect 51767 8352 51827 8372
rect 51885 8352 51945 8372
rect 52003 8352 52063 8372
rect 44405 8194 44465 8220
rect 44523 8194 44583 8220
rect 44641 8194 44701 8220
rect 44759 8200 44819 8220
rect 44759 8194 44820 8200
rect 44877 8194 44937 8220
rect 44995 8194 45055 8220
rect 37856 8106 37916 8132
rect 37974 8106 38034 8132
rect 38092 8106 38152 8132
rect 38210 8112 38270 8132
rect 38210 8106 38271 8112
rect 38328 8106 38388 8132
rect 38446 8106 38506 8132
rect 30563 8026 30647 8086
rect 31047 8026 31379 8086
rect 31779 8026 31805 8086
rect 30563 7968 30623 8026
rect 30563 7908 30647 7968
rect 31047 7908 31073 7968
rect 31214 7943 31273 8026
rect 31207 7926 31273 7943
rect 30373 7664 30424 7851
rect 31207 7892 31223 7926
rect 31257 7892 31273 7926
rect 31207 7876 31273 7892
rect 38093 7921 38151 8106
rect 38093 7895 38153 7921
rect 38211 7895 38271 8106
rect 38564 8100 38624 8132
rect 38682 8106 38742 8132
rect 38800 8106 38860 8132
rect 38561 8084 38627 8100
rect 38561 8050 38577 8084
rect 38611 8050 38627 8084
rect 38561 8034 38627 8050
rect 44642 8009 44700 8194
rect 44642 7983 44702 8009
rect 44760 7983 44820 8194
rect 45113 8188 45173 8220
rect 45231 8194 45291 8220
rect 45349 8194 45409 8220
rect 45110 8172 45176 8188
rect 45110 8138 45126 8172
rect 45160 8138 45176 8172
rect 70459 8425 70513 8485
rect 70913 8425 70939 8485
rect 70459 8367 70498 8425
rect 70459 8307 70513 8367
rect 70913 8366 70939 8367
rect 71100 8366 71166 8369
rect 70913 8353 71166 8366
rect 70913 8319 71116 8353
rect 71150 8319 71166 8353
rect 70913 8307 71166 8319
rect 71331 8367 71388 8774
rect 71598 8559 71643 9333
rect 71598 8499 71846 8559
rect 72046 8499 72072 8559
rect 71487 8367 71566 8378
rect 71331 8365 71846 8367
rect 71331 8307 71500 8365
rect 71555 8307 71846 8365
rect 72246 8307 72272 8367
rect 57684 8194 57744 8220
rect 57802 8194 57862 8220
rect 57920 8194 57980 8220
rect 58038 8200 58098 8220
rect 58038 8194 58099 8200
rect 58156 8194 58216 8220
rect 58274 8194 58334 8220
rect 45110 8122 45176 8138
rect 51059 8126 51119 8152
rect 51177 8126 51237 8152
rect 51295 8126 51355 8152
rect 51413 8132 51473 8152
rect 51413 8126 51474 8132
rect 51531 8126 51591 8152
rect 51649 8126 51709 8152
rect 44992 8055 45058 8071
rect 44992 8021 45008 8055
rect 45042 8021 45058 8055
rect 44992 8005 45058 8021
rect 46353 8018 46649 8069
rect 44995 7983 45055 8005
rect 46353 8003 46413 8018
rect 46471 8003 46531 8018
rect 46589 8003 46649 8018
rect 46707 8003 46767 8029
rect 46825 8003 46885 8029
rect 46943 8003 47003 8029
rect 48251 8018 48547 8069
rect 48251 8003 48311 8018
rect 48369 8003 48429 8018
rect 48487 8003 48547 8018
rect 48605 8003 48665 8029
rect 48723 8003 48783 8029
rect 48841 8003 48901 8029
rect 38443 7967 38509 7983
rect 38443 7933 38459 7967
rect 38493 7933 38509 7967
rect 38443 7917 38509 7933
rect 39804 7930 40100 7981
rect 38446 7895 38506 7917
rect 39804 7915 39864 7930
rect 39922 7915 39982 7930
rect 40040 7915 40100 7930
rect 40158 7915 40218 7941
rect 40276 7915 40336 7941
rect 40394 7915 40454 7941
rect 41702 7930 41998 7981
rect 41702 7915 41762 7930
rect 41820 7915 41880 7930
rect 41938 7915 41998 7930
rect 42056 7915 42116 7941
rect 42174 7915 42234 7941
rect 42292 7915 42352 7941
rect 34944 7685 35240 7721
rect 34944 7664 35004 7685
rect 35062 7664 35122 7685
rect 35180 7664 35240 7685
rect 35298 7684 35594 7720
rect 35298 7664 35358 7684
rect 35416 7664 35476 7684
rect 35534 7664 35594 7684
rect 35652 7684 35948 7720
rect 35652 7664 35712 7684
rect 35770 7664 35830 7684
rect 35888 7664 35948 7684
rect 23672 7629 23732 7655
rect 23790 7629 23850 7655
rect 23908 7629 23968 7655
rect 24026 7629 24086 7655
rect 30086 7604 30154 7664
rect 30354 7604 30424 7664
rect 31275 7636 31341 7652
rect 30511 7614 30565 7630
rect 23845 7574 23911 7582
rect 23476 7566 23911 7574
rect 23476 7532 23861 7566
rect 23895 7532 23911 7566
rect 23476 7523 23911 7532
rect 20701 7516 20767 7523
rect 23845 7516 23911 7523
rect 30086 7546 30137 7604
rect 30511 7580 30521 7614
rect 30555 7580 30565 7614
rect 30511 7562 30565 7580
rect 31275 7602 31291 7636
rect 31325 7602 31341 7636
rect 31275 7562 31341 7602
rect 30373 7546 31379 7562
rect 30086 7486 30154 7546
rect 30354 7502 31379 7546
rect 31579 7502 31605 7562
rect 30354 7487 30424 7502
rect 30354 7486 30380 7487
rect 30086 7428 30137 7486
rect 39320 7715 39380 7741
rect 39438 7715 39498 7741
rect 39556 7715 39616 7741
rect 38446 7669 38506 7695
rect 38093 7473 38153 7495
rect 38211 7479 38271 7495
rect 34944 7438 35004 7464
rect 35062 7438 35122 7464
rect 35180 7438 35240 7464
rect 35298 7444 35358 7464
rect 35298 7438 35359 7444
rect 35416 7438 35476 7464
rect 35534 7438 35594 7464
rect 30086 7368 30154 7428
rect 30354 7368 30380 7428
rect 35181 7253 35239 7438
rect 35181 7227 35241 7253
rect 35299 7227 35359 7438
rect 35652 7432 35712 7464
rect 35770 7438 35830 7464
rect 35888 7438 35948 7464
rect 38090 7457 38156 7473
rect 35649 7416 35715 7432
rect 35649 7382 35665 7416
rect 35699 7382 35715 7416
rect 38090 7423 38106 7457
rect 38140 7423 38156 7457
rect 38090 7407 38156 7423
rect 38205 7457 38279 7479
rect 38205 7423 38224 7457
rect 38258 7423 38279 7457
rect 40641 7732 40937 7783
rect 40641 7715 40701 7732
rect 40759 7715 40819 7732
rect 40877 7715 40937 7732
rect 41218 7715 41278 7741
rect 41336 7715 41396 7741
rect 41454 7715 41514 7741
rect 42539 7732 42835 7783
rect 42539 7715 42599 7732
rect 42657 7715 42717 7732
rect 42775 7715 42835 7732
rect 45869 7803 45929 7829
rect 45987 7803 46047 7829
rect 46105 7803 46165 7829
rect 44995 7757 45055 7783
rect 44642 7561 44702 7583
rect 44760 7567 44820 7583
rect 44639 7545 44705 7561
rect 39320 7498 39380 7515
rect 39438 7498 39498 7515
rect 39556 7498 39616 7515
rect 39804 7498 39864 7515
rect 39320 7447 39864 7498
rect 39922 7489 39982 7515
rect 40040 7489 40100 7515
rect 40158 7496 40218 7515
rect 40276 7496 40336 7515
rect 40394 7496 40454 7515
rect 40641 7496 40701 7515
rect 40759 7496 40819 7515
rect 35649 7366 35715 7382
rect 38205 7366 38279 7423
rect 39445 7366 39505 7447
rect 40158 7445 40701 7496
rect 40743 7489 40819 7496
rect 40877 7489 40937 7515
rect 41218 7498 41278 7515
rect 41336 7498 41396 7515
rect 41454 7498 41514 7515
rect 41702 7498 41762 7515
rect 40743 7445 40818 7489
rect 41218 7447 41762 7498
rect 41820 7489 41880 7515
rect 41938 7489 41998 7515
rect 42056 7496 42116 7515
rect 42174 7496 42234 7515
rect 42292 7496 42352 7515
rect 42539 7496 42599 7515
rect 42657 7496 42717 7515
rect 38205 7341 39505 7366
rect 35531 7299 35597 7315
rect 35531 7265 35547 7299
rect 35581 7265 35597 7299
rect 38204 7293 39505 7341
rect 40743 7325 40803 7445
rect 35531 7249 35597 7265
rect 35534 7227 35594 7249
rect 30699 6940 30759 6956
rect 30126 6857 30152 6917
rect 30352 6857 30420 6917
rect 30369 6799 30420 6857
rect 30126 6739 30152 6799
rect 30352 6792 30420 6799
rect 30699 6906 30713 6940
rect 30747 6906 30759 6940
rect 30699 6792 30759 6906
rect 35534 7001 35594 7027
rect 35181 6805 35241 6827
rect 35299 6805 35359 6827
rect 30352 6739 31377 6792
rect 30369 6732 31377 6739
rect 31577 6732 31603 6792
rect 35178 6789 35244 6805
rect 35178 6755 35194 6789
rect 35228 6755 35244 6789
rect 35178 6739 35244 6755
rect 35296 6789 35362 6805
rect 35296 6755 35312 6789
rect 35346 6755 35362 6789
rect 35296 6739 35362 6755
rect 37851 6749 38147 6785
rect 30369 6681 30420 6732
rect 30126 6621 30152 6681
rect 30352 6621 30420 6681
rect 31272 6691 31338 6732
rect 31272 6657 31288 6691
rect 31322 6657 31338 6691
rect 37851 6728 37911 6749
rect 37969 6728 38029 6749
rect 38087 6728 38147 6749
rect 38205 6748 38501 6784
rect 38205 6728 38265 6748
rect 38323 6728 38383 6748
rect 38441 6728 38501 6748
rect 38559 6748 38855 6784
rect 38559 6728 38619 6748
rect 38677 6728 38737 6748
rect 38795 6728 38855 6748
rect 31272 6641 31338 6657
rect 3175 6557 3235 6583
rect 3293 6557 3353 6583
rect 3411 6557 3471 6583
rect 3913 6557 3973 6583
rect 4031 6557 4091 6583
rect 4149 6557 4209 6583
rect 4651 6557 4711 6583
rect 4769 6557 4829 6583
rect 4887 6557 4947 6583
rect 5389 6557 5449 6583
rect 5507 6557 5567 6583
rect 5625 6557 5685 6583
rect 6129 6557 6189 6583
rect 6247 6557 6307 6583
rect 6365 6557 6425 6583
rect 6871 6559 6931 6585
rect 6989 6559 7049 6585
rect 7107 6559 7167 6585
rect 7609 6563 7669 6589
rect 7727 6563 7787 6589
rect 7845 6563 7905 6589
rect 8347 6559 8407 6585
rect 8465 6559 8525 6585
rect 8583 6559 8643 6585
rect 3175 6341 3235 6357
rect 3293 6341 3353 6357
rect 3411 6341 3471 6357
rect 3175 6305 3471 6341
rect 3913 6341 3973 6357
rect 4031 6341 4091 6357
rect 4149 6341 4209 6357
rect 3913 6305 4209 6341
rect 4651 6341 4711 6357
rect 4769 6341 4829 6357
rect 4887 6341 4947 6357
rect 4651 6305 4947 6341
rect 5389 6341 5449 6357
rect 5507 6341 5567 6357
rect 5625 6341 5685 6357
rect 5389 6305 5685 6341
rect 6129 6341 6189 6357
rect 6247 6341 6307 6357
rect 6365 6341 6425 6357
rect 6129 6305 6425 6341
rect 6871 6341 6931 6359
rect 6989 6341 7049 6359
rect 7107 6341 7167 6359
rect 6871 6305 7167 6341
rect 7609 6341 7669 6363
rect 7727 6341 7787 6363
rect 7845 6341 7905 6363
rect 9762 6447 9822 6473
rect 9880 6447 9940 6473
rect 9998 6447 10058 6473
rect 10116 6462 10412 6513
rect 10116 6447 10176 6462
rect 10234 6447 10294 6462
rect 10352 6447 10412 6462
rect 7609 6305 7905 6341
rect 8347 6343 8407 6359
rect 8465 6343 8525 6359
rect 8583 6343 8643 6359
rect 8347 6307 8643 6343
rect 3293 6263 3353 6305
rect 3293 6229 3307 6263
rect 3341 6229 3353 6263
rect 3293 6175 3353 6229
rect 4031 6263 4091 6305
rect 4031 6229 4045 6263
rect 4079 6229 4091 6263
rect 4031 6175 4091 6229
rect 4769 6263 4829 6305
rect 4769 6229 4783 6263
rect 4817 6229 4829 6263
rect 4769 6171 4829 6229
rect 5507 6263 5567 6305
rect 5507 6229 5521 6263
rect 5555 6229 5567 6263
rect 5507 6171 5567 6229
rect 6247 6263 6307 6305
rect 6247 6229 6261 6263
rect 6295 6229 6307 6263
rect 6247 6171 6307 6229
rect 6989 6263 7049 6305
rect 6989 6229 7003 6263
rect 7037 6229 7049 6263
rect 6989 6171 7049 6229
rect 7727 6263 7787 6305
rect 7727 6229 7741 6263
rect 7775 6229 7787 6263
rect 7727 6175 7787 6229
rect 8465 6265 8525 6307
rect 8465 6231 8479 6265
rect 8513 6231 8525 6265
rect 9279 6264 9575 6315
rect 9279 6247 9339 6264
rect 9397 6247 9457 6264
rect 9515 6247 9575 6264
rect 3293 5949 3353 5975
rect 4031 5949 4091 5975
rect 8465 6173 8525 6231
rect 4769 5945 4829 5971
rect 5507 5945 5567 5971
rect 6247 5945 6307 5971
rect 6989 5945 7049 5971
rect 7727 5949 7787 5975
rect 11830 6445 11890 6471
rect 11948 6445 12008 6471
rect 12066 6445 12126 6471
rect 12184 6460 12480 6511
rect 12184 6445 12244 6460
rect 12302 6445 12362 6460
rect 12420 6445 12480 6460
rect 13899 6447 13959 6473
rect 14017 6447 14077 6473
rect 14135 6447 14195 6473
rect 14253 6462 14549 6513
rect 14253 6447 14313 6462
rect 14371 6447 14431 6462
rect 14489 6447 14549 6462
rect 10600 6247 10660 6273
rect 10718 6247 10778 6273
rect 10836 6247 10896 6273
rect 11347 6262 11643 6313
rect 11347 6245 11407 6262
rect 11465 6245 11525 6262
rect 11583 6245 11643 6262
rect 9279 6021 9339 6047
rect 9397 6028 9457 6047
rect 9515 6028 9575 6047
rect 9762 6028 9822 6047
rect 9880 6028 9940 6047
rect 9998 6028 10058 6047
rect 9397 6021 9473 6028
rect 9398 5977 9473 6021
rect 9515 5977 10058 6028
rect 10116 6021 10176 6047
rect 10234 6021 10294 6047
rect 10352 6030 10412 6047
rect 10600 6030 10660 6047
rect 10718 6030 10778 6047
rect 10836 6030 10896 6047
rect 12668 6245 12728 6271
rect 12786 6245 12846 6271
rect 12904 6245 12964 6271
rect 13416 6264 13712 6315
rect 13416 6247 13476 6264
rect 13534 6247 13594 6264
rect 13652 6247 13712 6264
rect 15967 6445 16027 6471
rect 16085 6445 16145 6471
rect 16203 6445 16263 6471
rect 16321 6460 16617 6511
rect 16321 6445 16381 6460
rect 16439 6445 16499 6460
rect 16557 6445 16617 6460
rect 18036 6445 18096 6471
rect 18154 6445 18214 6471
rect 18272 6445 18332 6471
rect 18390 6460 18686 6511
rect 18390 6445 18450 6460
rect 18508 6445 18568 6460
rect 18626 6445 18686 6460
rect 14737 6247 14797 6273
rect 14855 6247 14915 6273
rect 14973 6247 15033 6273
rect 15484 6262 15780 6313
rect 15484 6245 15544 6262
rect 15602 6245 15662 6262
rect 15720 6245 15780 6262
rect 10352 5979 10896 6030
rect 11347 6019 11407 6045
rect 11465 6026 11525 6045
rect 11583 6026 11643 6045
rect 11830 6026 11890 6045
rect 11948 6026 12008 6045
rect 12066 6026 12126 6045
rect 11465 6019 11541 6026
rect 8465 5947 8525 5973
rect 9413 5890 9473 5977
rect 9413 5880 9541 5890
rect 9413 5846 9491 5880
rect 9525 5846 9541 5880
rect 9413 5836 9541 5846
rect 9413 5126 9473 5836
rect 9819 5778 10115 5838
rect 9819 5754 9879 5778
rect 9937 5754 9997 5778
rect 10055 5754 10115 5778
rect 10173 5777 10469 5837
rect 10173 5754 10233 5777
rect 10291 5754 10351 5777
rect 10409 5754 10469 5777
rect 10711 5700 10771 5979
rect 11466 5975 11541 6019
rect 11583 5975 12126 6026
rect 12184 6019 12244 6045
rect 12302 6019 12362 6045
rect 12420 6028 12480 6045
rect 12668 6028 12728 6045
rect 12786 6028 12846 6045
rect 12904 6028 12964 6045
rect 12420 5977 12964 6028
rect 13416 6021 13476 6047
rect 13534 6028 13594 6047
rect 13652 6028 13712 6047
rect 13899 6028 13959 6047
rect 14017 6028 14077 6047
rect 14135 6028 14195 6047
rect 13534 6021 13610 6028
rect 13535 5977 13610 6021
rect 13652 5977 14195 6028
rect 14253 6021 14313 6047
rect 14371 6021 14431 6047
rect 14489 6030 14549 6047
rect 14737 6030 14797 6047
rect 14855 6030 14915 6047
rect 14973 6030 15033 6047
rect 16805 6245 16865 6271
rect 16923 6245 16983 6271
rect 17041 6245 17101 6271
rect 17553 6262 17849 6313
rect 17553 6245 17613 6262
rect 17671 6245 17731 6262
rect 17789 6245 17849 6262
rect 20104 6443 20164 6469
rect 20222 6443 20282 6469
rect 20340 6443 20400 6469
rect 20458 6458 20754 6509
rect 20458 6443 20518 6458
rect 20576 6443 20636 6458
rect 20694 6443 20754 6458
rect 22173 6445 22233 6471
rect 22291 6445 22351 6471
rect 22409 6445 22469 6471
rect 22527 6460 22823 6511
rect 22527 6445 22587 6460
rect 22645 6445 22705 6460
rect 22763 6445 22823 6460
rect 18874 6245 18934 6271
rect 18992 6245 19052 6271
rect 19110 6245 19170 6271
rect 19621 6260 19917 6311
rect 19621 6243 19681 6260
rect 19739 6243 19799 6260
rect 19857 6243 19917 6260
rect 14489 5979 15033 6030
rect 15484 6019 15544 6045
rect 15602 6026 15662 6045
rect 15720 6026 15780 6045
rect 15967 6026 16027 6045
rect 16085 6026 16145 6045
rect 16203 6026 16263 6045
rect 15602 6019 15678 6026
rect 11481 5888 11541 5975
rect 11481 5878 11609 5888
rect 11481 5844 11559 5878
rect 11593 5844 11609 5878
rect 11481 5834 11609 5844
rect 10711 5686 10935 5700
rect 10711 5652 10885 5686
rect 10919 5652 10935 5686
rect 10711 5640 10935 5652
rect 9819 5328 9879 5354
rect 9787 5187 9854 5194
rect 9937 5187 9997 5354
rect 10055 5328 10115 5354
rect 10173 5328 10233 5354
rect 9787 5178 9997 5187
rect 9787 5144 9803 5178
rect 9837 5144 9997 5178
rect 9787 5128 9997 5144
rect 9413 5110 9563 5126
rect 9413 5076 9513 5110
rect 9547 5076 9563 5110
rect 9413 5060 9563 5076
rect 9413 5022 9473 5060
rect 9937 5022 9997 5128
rect 10291 5187 10351 5354
rect 10409 5328 10469 5354
rect 10434 5187 10501 5194
rect 10291 5178 10501 5187
rect 10291 5144 10451 5178
rect 10485 5144 10501 5178
rect 10291 5128 10501 5144
rect 10051 5095 10117 5110
rect 10051 5061 10067 5095
rect 10101 5061 10117 5095
rect 10051 5045 10117 5061
rect 10169 5094 10235 5110
rect 10169 5060 10185 5094
rect 10219 5060 10235 5094
rect 10055 5022 10115 5045
rect 10169 5044 10235 5060
rect 10173 5022 10233 5044
rect 10291 5022 10351 5128
rect 10711 5127 10771 5640
rect 10620 5111 10771 5127
rect 10620 5077 10636 5111
rect 10670 5077 10771 5111
rect 10620 5061 10771 5077
rect 10711 5022 10771 5061
rect 11481 5124 11541 5834
rect 11887 5776 12183 5836
rect 11887 5752 11947 5776
rect 12005 5752 12065 5776
rect 12123 5752 12183 5776
rect 12241 5775 12537 5835
rect 12241 5752 12301 5775
rect 12359 5752 12419 5775
rect 12477 5752 12537 5775
rect 12779 5698 12839 5977
rect 13550 5890 13610 5977
rect 13550 5880 13678 5890
rect 13550 5846 13628 5880
rect 13662 5846 13678 5880
rect 13550 5836 13678 5846
rect 12779 5684 13003 5698
rect 12779 5650 12953 5684
rect 12987 5650 13003 5684
rect 12779 5638 13003 5650
rect 11887 5326 11947 5352
rect 11855 5185 11922 5192
rect 12005 5185 12065 5352
rect 12123 5326 12183 5352
rect 12241 5326 12301 5352
rect 11855 5176 12065 5185
rect 11855 5142 11871 5176
rect 11905 5142 12065 5176
rect 11855 5126 12065 5142
rect 11481 5108 11631 5124
rect 11481 5074 11581 5108
rect 11615 5074 11631 5108
rect 11481 5058 11631 5074
rect 9413 4796 9473 4822
rect 11481 5020 11541 5058
rect 12005 5020 12065 5126
rect 12359 5185 12419 5352
rect 12477 5326 12537 5352
rect 12502 5185 12569 5192
rect 12359 5176 12569 5185
rect 12359 5142 12519 5176
rect 12553 5142 12569 5176
rect 12359 5126 12569 5142
rect 12119 5093 12185 5108
rect 12119 5059 12135 5093
rect 12169 5059 12185 5093
rect 12119 5043 12185 5059
rect 12237 5092 12303 5108
rect 12237 5058 12253 5092
rect 12287 5058 12303 5092
rect 12123 5020 12183 5043
rect 12237 5042 12303 5058
rect 12241 5020 12301 5042
rect 12359 5020 12419 5126
rect 12779 5125 12839 5638
rect 12688 5109 12839 5125
rect 12688 5075 12704 5109
rect 12738 5075 12839 5109
rect 12688 5059 12839 5075
rect 12779 5020 12839 5059
rect 13550 5126 13610 5836
rect 13956 5778 14252 5838
rect 13956 5754 14016 5778
rect 14074 5754 14134 5778
rect 14192 5754 14252 5778
rect 14310 5777 14606 5837
rect 14310 5754 14370 5777
rect 14428 5754 14488 5777
rect 14546 5754 14606 5777
rect 14848 5700 14908 5979
rect 15603 5975 15678 6019
rect 15720 5975 16263 6026
rect 16321 6019 16381 6045
rect 16439 6019 16499 6045
rect 16557 6028 16617 6045
rect 16805 6028 16865 6045
rect 16923 6028 16983 6045
rect 17041 6028 17101 6045
rect 16557 5977 17101 6028
rect 17553 6019 17613 6045
rect 17671 6026 17731 6045
rect 17789 6026 17849 6045
rect 18036 6026 18096 6045
rect 18154 6026 18214 6045
rect 18272 6026 18332 6045
rect 17671 6019 17747 6026
rect 15618 5888 15678 5975
rect 15618 5878 15746 5888
rect 15618 5844 15696 5878
rect 15730 5844 15746 5878
rect 15618 5834 15746 5844
rect 14848 5686 15072 5700
rect 14848 5652 15022 5686
rect 15056 5652 15072 5686
rect 14848 5640 15072 5652
rect 13956 5328 14016 5354
rect 13924 5187 13991 5194
rect 14074 5187 14134 5354
rect 14192 5328 14252 5354
rect 14310 5328 14370 5354
rect 13924 5178 14134 5187
rect 13924 5144 13940 5178
rect 13974 5144 14134 5178
rect 13924 5128 14134 5144
rect 13550 5110 13700 5126
rect 13550 5076 13650 5110
rect 13684 5076 13700 5110
rect 13550 5060 13700 5076
rect 13550 5022 13610 5060
rect 14074 5022 14134 5128
rect 14428 5187 14488 5354
rect 14546 5328 14606 5354
rect 14571 5187 14638 5194
rect 14428 5178 14638 5187
rect 14428 5144 14588 5178
rect 14622 5144 14638 5178
rect 14428 5128 14638 5144
rect 14188 5095 14254 5110
rect 14188 5061 14204 5095
rect 14238 5061 14254 5095
rect 14188 5045 14254 5061
rect 14306 5094 14372 5110
rect 14306 5060 14322 5094
rect 14356 5060 14372 5094
rect 14192 5022 14252 5045
rect 14306 5044 14372 5060
rect 14310 5022 14370 5044
rect 14428 5022 14488 5128
rect 14848 5127 14908 5640
rect 14757 5111 14908 5127
rect 14757 5077 14773 5111
rect 14807 5077 14908 5111
rect 14757 5061 14908 5077
rect 14848 5022 14908 5061
rect 15618 5124 15678 5834
rect 16024 5776 16320 5836
rect 16024 5752 16084 5776
rect 16142 5752 16202 5776
rect 16260 5752 16320 5776
rect 16378 5775 16674 5835
rect 16378 5752 16438 5775
rect 16496 5752 16556 5775
rect 16614 5752 16674 5775
rect 16916 5698 16976 5977
rect 17672 5975 17747 6019
rect 17789 5975 18332 6026
rect 18390 6019 18450 6045
rect 18508 6019 18568 6045
rect 18626 6028 18686 6045
rect 18874 6028 18934 6045
rect 18992 6028 19052 6045
rect 19110 6028 19170 6045
rect 20942 6243 21002 6269
rect 21060 6243 21120 6269
rect 21178 6243 21238 6269
rect 21690 6262 21986 6313
rect 21690 6245 21750 6262
rect 21808 6245 21868 6262
rect 21926 6245 21986 6262
rect 24241 6443 24301 6469
rect 24359 6443 24419 6469
rect 24477 6443 24537 6469
rect 24595 6458 24891 6509
rect 24595 6443 24655 6458
rect 24713 6443 24773 6458
rect 24831 6443 24891 6458
rect 23011 6245 23071 6271
rect 23129 6245 23189 6271
rect 23247 6245 23307 6271
rect 23758 6260 24054 6311
rect 23758 6243 23818 6260
rect 23876 6243 23936 6260
rect 23994 6243 24054 6260
rect 18626 5977 19170 6028
rect 19621 6017 19681 6043
rect 19739 6024 19799 6043
rect 19857 6024 19917 6043
rect 20104 6024 20164 6043
rect 20222 6024 20282 6043
rect 20340 6024 20400 6043
rect 19739 6017 19815 6024
rect 17687 5888 17747 5975
rect 17687 5878 17815 5888
rect 17687 5844 17765 5878
rect 17799 5844 17815 5878
rect 17687 5834 17815 5844
rect 16916 5684 17140 5698
rect 16916 5650 17090 5684
rect 17124 5650 17140 5684
rect 16916 5638 17140 5650
rect 16024 5326 16084 5352
rect 15992 5185 16059 5192
rect 16142 5185 16202 5352
rect 16260 5326 16320 5352
rect 16378 5326 16438 5352
rect 15992 5176 16202 5185
rect 15992 5142 16008 5176
rect 16042 5142 16202 5176
rect 15992 5126 16202 5142
rect 15618 5108 15768 5124
rect 15618 5074 15718 5108
rect 15752 5074 15768 5108
rect 15618 5058 15768 5074
rect 10711 4796 10771 4822
rect 11481 4794 11541 4820
rect 9937 4596 9997 4622
rect 10055 4596 10115 4622
rect 10173 4596 10233 4622
rect 10291 4596 10351 4622
rect 12779 4794 12839 4820
rect 13550 4796 13610 4822
rect 15618 5020 15678 5058
rect 16142 5020 16202 5126
rect 16496 5185 16556 5352
rect 16614 5326 16674 5352
rect 16639 5185 16706 5192
rect 16496 5176 16706 5185
rect 16496 5142 16656 5176
rect 16690 5142 16706 5176
rect 16496 5126 16706 5142
rect 16256 5093 16322 5108
rect 16256 5059 16272 5093
rect 16306 5059 16322 5093
rect 16256 5043 16322 5059
rect 16374 5092 16440 5108
rect 16374 5058 16390 5092
rect 16424 5058 16440 5092
rect 16260 5020 16320 5043
rect 16374 5042 16440 5058
rect 16378 5020 16438 5042
rect 16496 5020 16556 5126
rect 16916 5125 16976 5638
rect 16825 5109 16976 5125
rect 16825 5075 16841 5109
rect 16875 5075 16976 5109
rect 16825 5059 16976 5075
rect 16916 5020 16976 5059
rect 17687 5124 17747 5834
rect 18093 5776 18389 5836
rect 18093 5752 18153 5776
rect 18211 5752 18271 5776
rect 18329 5752 18389 5776
rect 18447 5775 18743 5835
rect 18447 5752 18507 5775
rect 18565 5752 18625 5775
rect 18683 5752 18743 5775
rect 18985 5698 19045 5977
rect 19740 5973 19815 6017
rect 19857 5973 20400 6024
rect 20458 6017 20518 6043
rect 20576 6017 20636 6043
rect 20694 6026 20754 6043
rect 20942 6026 21002 6043
rect 21060 6026 21120 6043
rect 21178 6026 21238 6043
rect 20694 5975 21238 6026
rect 21690 6019 21750 6045
rect 21808 6026 21868 6045
rect 21926 6026 21986 6045
rect 22173 6026 22233 6045
rect 22291 6026 22351 6045
rect 22409 6026 22469 6045
rect 21808 6019 21884 6026
rect 21809 5975 21884 6019
rect 21926 5975 22469 6026
rect 22527 6019 22587 6045
rect 22645 6019 22705 6045
rect 22763 6028 22823 6045
rect 23011 6028 23071 6045
rect 23129 6028 23189 6045
rect 23247 6028 23307 6045
rect 30369 6433 30420 6621
rect 39445 6595 39505 7293
rect 39747 7245 40043 7305
rect 39747 7222 39807 7245
rect 39865 7222 39925 7245
rect 39983 7222 40043 7245
rect 40101 7246 40397 7306
rect 40742 7305 40803 7325
rect 40101 7222 40161 7246
rect 40219 7222 40279 7246
rect 40337 7222 40397 7246
rect 40723 7289 40803 7305
rect 40723 7255 40738 7289
rect 40772 7255 40803 7289
rect 40723 7239 40803 7255
rect 40742 7216 40803 7239
rect 40743 7070 40803 7216
rect 40742 6897 40803 7070
rect 39747 6796 39807 6822
rect 39715 6655 39782 6662
rect 39865 6655 39925 6822
rect 39983 6796 40043 6822
rect 40101 6796 40161 6822
rect 39715 6646 39925 6655
rect 39715 6612 39731 6646
rect 39765 6612 39925 6646
rect 39715 6596 39925 6612
rect 39445 6579 39596 6595
rect 39445 6545 39546 6579
rect 39580 6545 39596 6579
rect 39445 6529 39596 6545
rect 31205 6506 31271 6522
rect 29886 6373 29952 6433
rect 30352 6373 30420 6433
rect 30562 6430 30645 6490
rect 31045 6430 31071 6490
rect 31205 6472 31221 6506
rect 31255 6472 31271 6506
rect 37851 6502 37911 6528
rect 37969 6502 38029 6528
rect 38087 6502 38147 6528
rect 38205 6508 38265 6528
rect 38205 6502 38266 6508
rect 38323 6502 38383 6528
rect 38441 6502 38501 6528
rect 31205 6455 31271 6472
rect 29886 6315 29937 6373
rect 30562 6372 30622 6430
rect 31212 6372 31271 6455
rect 25079 6243 25139 6269
rect 25197 6243 25257 6269
rect 25315 6243 25375 6269
rect 29886 6255 29952 6315
rect 30352 6255 30378 6315
rect 30562 6312 30645 6372
rect 31045 6312 31377 6372
rect 31777 6312 31803 6372
rect 38088 6317 38146 6502
rect 29886 6197 29937 6255
rect 30562 6254 30622 6312
rect 38088 6291 38148 6317
rect 38206 6291 38266 6502
rect 38559 6496 38619 6528
rect 38677 6502 38737 6528
rect 38795 6502 38855 6528
rect 38556 6480 38622 6496
rect 39445 6490 39505 6529
rect 39865 6490 39925 6596
rect 40219 6655 40279 6822
rect 40337 6796 40397 6822
rect 40362 6655 40429 6662
rect 40219 6646 40429 6655
rect 40219 6612 40379 6646
rect 40413 6612 40429 6646
rect 40219 6596 40429 6612
rect 39981 6562 40047 6578
rect 39981 6528 39997 6562
rect 40031 6528 40047 6562
rect 39981 6512 40047 6528
rect 40099 6563 40165 6578
rect 40099 6529 40115 6563
rect 40149 6529 40165 6563
rect 40099 6513 40165 6529
rect 39983 6490 40043 6512
rect 40101 6490 40161 6513
rect 40219 6490 40279 6596
rect 40743 6594 40803 6897
rect 40653 6578 40803 6594
rect 40653 6544 40669 6578
rect 40703 6544 40803 6578
rect 40653 6528 40803 6544
rect 40743 6490 40803 6528
rect 41343 6789 41403 7447
rect 42056 7445 42599 7496
rect 42641 7489 42717 7496
rect 42775 7489 42835 7515
rect 44639 7511 44655 7545
rect 44689 7511 44705 7545
rect 44639 7495 44705 7511
rect 44754 7545 44828 7567
rect 44754 7511 44773 7545
rect 44807 7511 44828 7545
rect 47190 7820 47486 7871
rect 47190 7803 47250 7820
rect 47308 7803 47368 7820
rect 47426 7803 47486 7820
rect 47767 7803 47827 7829
rect 47885 7803 47945 7829
rect 48003 7803 48063 7829
rect 51296 7941 51354 8126
rect 51296 7915 51356 7941
rect 51414 7915 51474 8126
rect 51767 8120 51827 8152
rect 51885 8126 51945 8152
rect 52003 8126 52063 8152
rect 51764 8104 51830 8120
rect 51764 8070 51780 8104
rect 51814 8070 51830 8104
rect 51764 8054 51830 8070
rect 57921 8009 57979 8194
rect 51646 7987 51712 8003
rect 51646 7953 51662 7987
rect 51696 7953 51712 7987
rect 51646 7937 51712 7953
rect 53007 7950 53303 8001
rect 51649 7915 51709 7937
rect 53007 7935 53067 7950
rect 53125 7935 53185 7950
rect 53243 7935 53303 7950
rect 53361 7935 53421 7961
rect 53479 7935 53539 7961
rect 53597 7935 53657 7961
rect 54905 7950 55201 8001
rect 57921 7983 57981 8009
rect 58039 7983 58099 8194
rect 58392 8188 58452 8220
rect 58510 8194 58570 8220
rect 58628 8194 58688 8220
rect 58389 8172 58455 8188
rect 58389 8138 58405 8172
rect 58439 8138 58455 8172
rect 58389 8122 58455 8138
rect 58271 8055 58337 8071
rect 58271 8021 58287 8055
rect 58321 8021 58337 8055
rect 58271 8005 58337 8021
rect 59632 8018 59928 8069
rect 58274 7983 58334 8005
rect 59632 8003 59692 8018
rect 59750 8003 59810 8018
rect 59868 8003 59928 8018
rect 59986 8003 60046 8029
rect 60104 8003 60164 8029
rect 60222 8003 60282 8029
rect 61530 8018 61826 8069
rect 70459 8249 70498 8307
rect 71099 8303 71166 8307
rect 71487 8297 71566 8307
rect 71200 8249 71287 8266
rect 70459 8189 70513 8249
rect 70913 8189 70939 8249
rect 71200 8247 71846 8249
rect 71200 8189 71215 8247
rect 71270 8189 71846 8247
rect 72246 8189 72272 8249
rect 71200 8171 71287 8189
rect 61530 8003 61590 8018
rect 61648 8003 61708 8018
rect 61766 8003 61826 8018
rect 61884 8003 61944 8029
rect 62002 8003 62062 8029
rect 62120 8003 62180 8029
rect 70459 8071 70513 8131
rect 70913 8071 70939 8131
rect 70459 8013 70498 8071
rect 71238 8013 71287 8171
rect 71720 8131 71786 8134
rect 72319 8176 72385 8192
rect 72319 8142 72335 8176
rect 72369 8142 72385 8176
rect 71720 8118 71846 8131
rect 71720 8084 71736 8118
rect 71770 8084 71846 8118
rect 71720 8071 71846 8084
rect 72246 8071 72272 8131
rect 72319 8126 72385 8142
rect 71720 8068 71786 8071
rect 54905 7935 54965 7950
rect 55023 7935 55083 7950
rect 55141 7935 55201 7950
rect 55259 7935 55319 7961
rect 55377 7935 55437 7961
rect 55495 7935 55555 7961
rect 49088 7820 49384 7871
rect 49088 7803 49148 7820
rect 49206 7803 49266 7820
rect 49324 7803 49384 7820
rect 45869 7586 45929 7603
rect 45987 7586 46047 7603
rect 46105 7586 46165 7603
rect 46353 7586 46413 7603
rect 45869 7535 46413 7586
rect 46471 7577 46531 7603
rect 46589 7577 46649 7603
rect 46707 7584 46767 7603
rect 46825 7584 46885 7603
rect 46943 7584 47003 7603
rect 47190 7584 47250 7603
rect 47308 7584 47368 7603
rect 42641 7445 42716 7489
rect 44754 7454 44828 7511
rect 45994 7454 46054 7535
rect 46707 7533 47250 7584
rect 47292 7577 47368 7584
rect 47426 7577 47486 7603
rect 47767 7586 47827 7603
rect 47885 7586 47945 7603
rect 48003 7586 48063 7603
rect 48251 7586 48311 7603
rect 47292 7533 47367 7577
rect 47767 7535 48311 7586
rect 48369 7577 48429 7603
rect 48487 7577 48547 7603
rect 48605 7584 48665 7603
rect 48723 7584 48783 7603
rect 48841 7584 48901 7603
rect 49088 7584 49148 7603
rect 49206 7584 49266 7603
rect 41645 7245 41941 7305
rect 41645 7222 41705 7245
rect 41763 7222 41823 7245
rect 41881 7222 41941 7245
rect 41999 7246 42295 7306
rect 41999 7222 42059 7246
rect 42117 7222 42177 7246
rect 42235 7222 42295 7246
rect 42641 7292 42701 7445
rect 44754 7429 46054 7454
rect 44753 7381 46054 7429
rect 47292 7413 47352 7533
rect 42641 7268 42895 7292
rect 42641 7234 42845 7268
rect 42879 7234 42895 7268
rect 42641 7218 42895 7234
rect 41645 6796 41705 6822
rect 41343 6773 41410 6789
rect 41343 6739 41359 6773
rect 41393 6739 41410 6773
rect 41343 6723 41410 6739
rect 41343 6595 41403 6723
rect 41613 6655 41680 6662
rect 41763 6655 41823 6822
rect 41881 6796 41941 6822
rect 41999 6796 42059 6822
rect 41613 6646 41823 6655
rect 41613 6612 41629 6646
rect 41663 6612 41823 6646
rect 41613 6596 41823 6612
rect 41343 6579 41494 6595
rect 41343 6545 41444 6579
rect 41478 6545 41494 6579
rect 41343 6529 41494 6545
rect 41343 6490 41403 6529
rect 41763 6490 41823 6596
rect 42117 6655 42177 6822
rect 42235 6796 42295 6822
rect 42258 6656 42325 6663
rect 42252 6655 42325 6656
rect 42117 6647 42325 6655
rect 42117 6613 42275 6647
rect 42309 6613 42325 6647
rect 42117 6597 42325 6613
rect 42117 6596 42314 6597
rect 41879 6562 41945 6578
rect 41879 6528 41895 6562
rect 41929 6528 41945 6562
rect 41879 6512 41945 6528
rect 41997 6563 42063 6578
rect 41997 6529 42013 6563
rect 42047 6529 42063 6563
rect 41997 6513 42063 6529
rect 41881 6490 41941 6512
rect 41999 6490 42059 6513
rect 42117 6490 42177 6596
rect 42641 6594 42701 7218
rect 44400 6837 44696 6873
rect 44400 6816 44460 6837
rect 44518 6816 44578 6837
rect 44636 6816 44696 6837
rect 44754 6836 45050 6872
rect 44754 6816 44814 6836
rect 44872 6816 44932 6836
rect 44990 6816 45050 6836
rect 45108 6836 45404 6872
rect 45108 6816 45168 6836
rect 45226 6816 45286 6836
rect 45344 6816 45404 6836
rect 45994 6683 46054 7381
rect 46296 7333 46592 7393
rect 46296 7310 46356 7333
rect 46414 7310 46474 7333
rect 46532 7310 46592 7333
rect 46650 7334 46946 7394
rect 47291 7393 47352 7413
rect 46650 7310 46710 7334
rect 46768 7310 46828 7334
rect 46886 7310 46946 7334
rect 47272 7377 47352 7393
rect 47272 7343 47287 7377
rect 47321 7343 47352 7377
rect 47272 7327 47352 7343
rect 47291 7304 47352 7327
rect 47292 7158 47352 7304
rect 47291 6985 47352 7158
rect 46296 6884 46356 6910
rect 46264 6743 46331 6750
rect 46414 6743 46474 6910
rect 46532 6884 46592 6910
rect 46650 6884 46710 6910
rect 46264 6734 46474 6743
rect 46264 6700 46280 6734
rect 46314 6700 46474 6734
rect 46264 6684 46474 6700
rect 45994 6667 46145 6683
rect 45994 6633 46095 6667
rect 46129 6633 46145 6667
rect 45994 6617 46145 6633
rect 42551 6578 42701 6594
rect 44400 6590 44460 6616
rect 44518 6590 44578 6616
rect 44636 6590 44696 6616
rect 44754 6596 44814 6616
rect 44754 6590 44815 6596
rect 44872 6590 44932 6616
rect 44990 6590 45050 6616
rect 42551 6544 42567 6578
rect 42601 6544 42701 6578
rect 42551 6528 42701 6544
rect 42641 6490 42701 6528
rect 38556 6446 38572 6480
rect 38606 6446 38622 6480
rect 38556 6430 38622 6446
rect 38438 6363 38504 6379
rect 38438 6329 38454 6363
rect 38488 6329 38504 6363
rect 38438 6313 38504 6329
rect 38441 6291 38501 6313
rect 31289 6254 31355 6256
rect 29886 6137 29952 6197
rect 30352 6137 30378 6197
rect 30562 6194 30645 6254
rect 31045 6194 31071 6254
rect 31289 6240 31377 6254
rect 31289 6206 31305 6240
rect 31339 6206 31377 6240
rect 31289 6194 31377 6206
rect 31777 6194 31803 6254
rect 31289 6190 31355 6194
rect 31289 6136 31354 6138
rect 22763 5977 23307 6028
rect 23758 6017 23818 6043
rect 23876 6024 23936 6043
rect 23994 6024 24054 6043
rect 24241 6024 24301 6043
rect 24359 6024 24419 6043
rect 24477 6024 24537 6043
rect 23876 6017 23952 6024
rect 19755 5886 19815 5973
rect 19755 5876 19883 5886
rect 19755 5842 19833 5876
rect 19867 5842 19883 5876
rect 19755 5832 19883 5842
rect 18985 5684 19209 5698
rect 18985 5650 19159 5684
rect 19193 5650 19209 5684
rect 18985 5638 19209 5650
rect 18093 5326 18153 5352
rect 18061 5185 18128 5192
rect 18211 5185 18271 5352
rect 18329 5326 18389 5352
rect 18447 5326 18507 5352
rect 18061 5176 18271 5185
rect 18061 5142 18077 5176
rect 18111 5142 18271 5176
rect 18061 5126 18271 5142
rect 17687 5108 17837 5124
rect 17687 5074 17787 5108
rect 17821 5074 17837 5108
rect 17687 5058 17837 5074
rect 17687 5020 17747 5058
rect 18211 5020 18271 5126
rect 18565 5185 18625 5352
rect 18683 5326 18743 5352
rect 18708 5185 18775 5192
rect 18565 5176 18775 5185
rect 18565 5142 18725 5176
rect 18759 5142 18775 5176
rect 18565 5126 18775 5142
rect 18325 5093 18391 5108
rect 18325 5059 18341 5093
rect 18375 5059 18391 5093
rect 18325 5043 18391 5059
rect 18443 5092 18509 5108
rect 18443 5058 18459 5092
rect 18493 5058 18509 5092
rect 18329 5020 18389 5043
rect 18443 5042 18509 5058
rect 18447 5020 18507 5042
rect 18565 5020 18625 5126
rect 18985 5125 19045 5638
rect 18894 5109 19045 5125
rect 18894 5075 18910 5109
rect 18944 5075 19045 5109
rect 18894 5059 19045 5075
rect 18985 5020 19045 5059
rect 19755 5122 19815 5832
rect 20161 5774 20457 5834
rect 20161 5750 20221 5774
rect 20279 5750 20339 5774
rect 20397 5750 20457 5774
rect 20515 5773 20811 5833
rect 20515 5750 20575 5773
rect 20633 5750 20693 5773
rect 20751 5750 20811 5773
rect 21053 5696 21113 5975
rect 21824 5888 21884 5975
rect 21824 5878 21952 5888
rect 21824 5844 21902 5878
rect 21936 5844 21952 5878
rect 21824 5834 21952 5844
rect 21053 5682 21277 5696
rect 21053 5648 21227 5682
rect 21261 5648 21277 5682
rect 21053 5636 21277 5648
rect 20161 5324 20221 5350
rect 20129 5183 20196 5190
rect 20279 5183 20339 5350
rect 20397 5324 20457 5350
rect 20515 5324 20575 5350
rect 20129 5174 20339 5183
rect 20129 5140 20145 5174
rect 20179 5140 20339 5174
rect 20129 5124 20339 5140
rect 19755 5106 19905 5122
rect 19755 5072 19855 5106
rect 19889 5072 19905 5106
rect 19755 5056 19905 5072
rect 14848 4796 14908 4822
rect 15618 4794 15678 4820
rect 12005 4594 12065 4620
rect 12123 4594 12183 4620
rect 12241 4594 12301 4620
rect 12359 4594 12419 4620
rect 14074 4596 14134 4622
rect 14192 4596 14252 4622
rect 14310 4596 14370 4622
rect 14428 4596 14488 4622
rect 16916 4794 16976 4820
rect 17687 4794 17747 4820
rect 19755 5018 19815 5056
rect 20279 5018 20339 5124
rect 20633 5183 20693 5350
rect 20751 5324 20811 5350
rect 20776 5183 20843 5190
rect 20633 5174 20843 5183
rect 20633 5140 20793 5174
rect 20827 5140 20843 5174
rect 20633 5124 20843 5140
rect 20393 5091 20459 5106
rect 20393 5057 20409 5091
rect 20443 5057 20459 5091
rect 20393 5041 20459 5057
rect 20511 5090 20577 5106
rect 20511 5056 20527 5090
rect 20561 5056 20577 5090
rect 20397 5018 20457 5041
rect 20511 5040 20577 5056
rect 20515 5018 20575 5040
rect 20633 5018 20693 5124
rect 21053 5123 21113 5636
rect 20962 5107 21113 5123
rect 20962 5073 20978 5107
rect 21012 5073 21113 5107
rect 20962 5057 21113 5073
rect 21053 5018 21113 5057
rect 21824 5124 21884 5834
rect 22230 5776 22526 5836
rect 22230 5752 22290 5776
rect 22348 5752 22408 5776
rect 22466 5752 22526 5776
rect 22584 5775 22880 5835
rect 22584 5752 22644 5775
rect 22702 5752 22762 5775
rect 22820 5752 22880 5775
rect 23122 5698 23182 5977
rect 23877 5973 23952 6017
rect 23994 5973 24537 6024
rect 24595 6017 24655 6043
rect 24713 6017 24773 6043
rect 24831 6026 24891 6043
rect 25079 6026 25139 6043
rect 25197 6026 25257 6043
rect 25315 6026 25375 6043
rect 24831 5975 25375 6026
rect 23892 5886 23952 5973
rect 23892 5876 24020 5886
rect 23892 5842 23970 5876
rect 24004 5842 24020 5876
rect 23892 5832 24020 5842
rect 23122 5684 23346 5698
rect 23122 5650 23296 5684
rect 23330 5650 23346 5684
rect 23122 5638 23346 5650
rect 22230 5326 22290 5352
rect 22198 5185 22265 5192
rect 22348 5185 22408 5352
rect 22466 5326 22526 5352
rect 22584 5326 22644 5352
rect 22198 5176 22408 5185
rect 22198 5142 22214 5176
rect 22248 5142 22408 5176
rect 22198 5126 22408 5142
rect 21824 5108 21974 5124
rect 21824 5074 21924 5108
rect 21958 5074 21974 5108
rect 21824 5058 21974 5074
rect 21824 5020 21884 5058
rect 22348 5020 22408 5126
rect 22702 5185 22762 5352
rect 22820 5326 22880 5352
rect 22845 5185 22912 5192
rect 22702 5176 22912 5185
rect 22702 5142 22862 5176
rect 22896 5142 22912 5176
rect 22702 5126 22912 5142
rect 22462 5093 22528 5108
rect 22462 5059 22478 5093
rect 22512 5059 22528 5093
rect 22462 5043 22528 5059
rect 22580 5092 22646 5108
rect 22580 5058 22596 5092
rect 22630 5058 22646 5092
rect 22466 5020 22526 5043
rect 22580 5042 22646 5058
rect 22584 5020 22644 5042
rect 22702 5020 22762 5126
rect 23122 5125 23182 5638
rect 23031 5109 23182 5125
rect 23031 5075 23047 5109
rect 23081 5075 23182 5109
rect 23031 5059 23182 5075
rect 23122 5020 23182 5059
rect 23892 5122 23952 5832
rect 24298 5774 24594 5834
rect 24298 5750 24358 5774
rect 24416 5750 24476 5774
rect 24534 5750 24594 5774
rect 24652 5773 24948 5833
rect 24652 5750 24712 5773
rect 24770 5750 24830 5773
rect 24888 5750 24948 5773
rect 25190 5696 25250 5975
rect 29926 6019 29952 6079
rect 30352 6019 30422 6079
rect 30371 5961 30422 6019
rect 29926 5901 29952 5961
rect 30352 5901 30422 5961
rect 30371 5843 30422 5901
rect 29926 5783 29952 5843
rect 30352 5783 30422 5843
rect 30561 6076 30645 6136
rect 31045 6076 31071 6136
rect 31289 6122 31377 6136
rect 31289 6088 31304 6122
rect 31338 6088 31377 6122
rect 31289 6076 31377 6088
rect 31777 6076 31803 6136
rect 30561 6018 30621 6076
rect 31289 6072 31354 6076
rect 30561 5958 30645 6018
rect 31045 5958 31377 6018
rect 31777 5958 31803 6018
rect 30561 5900 30621 5958
rect 30561 5840 30645 5900
rect 31045 5840 31071 5900
rect 31212 5875 31271 5958
rect 39445 6264 39505 6290
rect 38441 6065 38501 6091
rect 40743 6264 40803 6290
rect 41343 6264 41403 6290
rect 44637 6405 44695 6590
rect 44637 6379 44697 6405
rect 44755 6379 44815 6590
rect 45108 6584 45168 6616
rect 45226 6590 45286 6616
rect 45344 6590 45404 6616
rect 45105 6568 45171 6584
rect 45994 6578 46054 6617
rect 46414 6578 46474 6684
rect 46768 6743 46828 6910
rect 46886 6884 46946 6910
rect 46911 6743 46978 6750
rect 46768 6734 46978 6743
rect 46768 6700 46928 6734
rect 46962 6700 46978 6734
rect 46768 6684 46978 6700
rect 46530 6650 46596 6666
rect 46530 6616 46546 6650
rect 46580 6616 46596 6650
rect 46530 6600 46596 6616
rect 46648 6651 46714 6666
rect 46648 6617 46664 6651
rect 46698 6617 46714 6651
rect 46648 6601 46714 6617
rect 46532 6578 46592 6600
rect 46650 6578 46710 6601
rect 46768 6578 46828 6684
rect 47292 6682 47352 6985
rect 47202 6666 47352 6682
rect 47202 6632 47218 6666
rect 47252 6632 47352 6666
rect 47202 6616 47352 6632
rect 47292 6578 47352 6616
rect 47892 6877 47952 7535
rect 48605 7533 49148 7584
rect 49190 7577 49266 7584
rect 49324 7577 49384 7603
rect 49190 7533 49265 7577
rect 48194 7333 48490 7393
rect 48194 7310 48254 7333
rect 48312 7310 48372 7333
rect 48430 7310 48490 7333
rect 48548 7334 48844 7394
rect 48548 7310 48608 7334
rect 48666 7310 48726 7334
rect 48784 7310 48844 7334
rect 49190 7380 49250 7533
rect 52523 7735 52583 7761
rect 52641 7735 52701 7761
rect 52759 7735 52819 7761
rect 51649 7689 51709 7715
rect 51296 7493 51356 7515
rect 51414 7499 51474 7515
rect 51293 7477 51359 7493
rect 51293 7443 51309 7477
rect 51343 7443 51359 7477
rect 51293 7427 51359 7443
rect 51408 7477 51482 7499
rect 51408 7443 51427 7477
rect 51461 7443 51482 7477
rect 53844 7752 54140 7803
rect 53844 7735 53904 7752
rect 53962 7735 54022 7752
rect 54080 7735 54140 7752
rect 54421 7735 54481 7761
rect 54539 7735 54599 7761
rect 54657 7735 54717 7761
rect 55742 7752 56038 7803
rect 55742 7735 55802 7752
rect 55860 7735 55920 7752
rect 55978 7735 56038 7752
rect 59148 7803 59208 7829
rect 59266 7803 59326 7829
rect 59384 7803 59444 7829
rect 58274 7757 58334 7783
rect 57921 7561 57981 7583
rect 58039 7567 58099 7583
rect 57918 7545 57984 7561
rect 52523 7518 52583 7535
rect 52641 7518 52701 7535
rect 52759 7518 52819 7535
rect 53007 7518 53067 7535
rect 52523 7467 53067 7518
rect 53125 7509 53185 7535
rect 53243 7509 53303 7535
rect 53361 7516 53421 7535
rect 53479 7516 53539 7535
rect 53597 7516 53657 7535
rect 53844 7516 53904 7535
rect 53962 7516 54022 7535
rect 51408 7386 51482 7443
rect 52648 7386 52708 7467
rect 53361 7465 53904 7516
rect 53946 7509 54022 7516
rect 54080 7509 54140 7535
rect 54421 7518 54481 7535
rect 54539 7518 54599 7535
rect 54657 7518 54717 7535
rect 54905 7518 54965 7535
rect 53946 7465 54021 7509
rect 54421 7467 54965 7518
rect 55023 7509 55083 7535
rect 55141 7509 55201 7535
rect 55259 7516 55319 7535
rect 55377 7516 55437 7535
rect 55495 7516 55555 7535
rect 55742 7516 55802 7535
rect 55860 7516 55920 7535
rect 49190 7356 49444 7380
rect 51408 7361 52708 7386
rect 49190 7322 49394 7356
rect 49428 7322 49444 7356
rect 49190 7306 49444 7322
rect 51407 7313 52708 7361
rect 53946 7345 54006 7465
rect 48194 6884 48254 6910
rect 47892 6861 47959 6877
rect 47892 6827 47908 6861
rect 47942 6827 47959 6861
rect 47892 6811 47959 6827
rect 47892 6683 47952 6811
rect 48162 6743 48229 6750
rect 48312 6743 48372 6910
rect 48430 6884 48490 6910
rect 48548 6884 48608 6910
rect 48162 6734 48372 6743
rect 48162 6700 48178 6734
rect 48212 6700 48372 6734
rect 48162 6684 48372 6700
rect 47892 6667 48043 6683
rect 47892 6633 47993 6667
rect 48027 6633 48043 6667
rect 47892 6617 48043 6633
rect 47892 6578 47952 6617
rect 48312 6578 48372 6684
rect 48666 6743 48726 6910
rect 48784 6884 48844 6910
rect 48807 6744 48874 6751
rect 48801 6743 48874 6744
rect 48666 6735 48874 6743
rect 48666 6701 48824 6735
rect 48858 6701 48874 6735
rect 48666 6685 48874 6701
rect 48666 6684 48863 6685
rect 48428 6650 48494 6666
rect 48428 6616 48444 6650
rect 48478 6616 48494 6650
rect 48428 6600 48494 6616
rect 48546 6651 48612 6666
rect 48546 6617 48562 6651
rect 48596 6617 48612 6651
rect 48546 6601 48612 6617
rect 48430 6578 48490 6600
rect 48548 6578 48608 6601
rect 48666 6578 48726 6684
rect 49190 6682 49250 7306
rect 51054 6769 51350 6805
rect 51054 6748 51114 6769
rect 51172 6748 51232 6769
rect 51290 6748 51350 6769
rect 51408 6768 51704 6804
rect 51408 6748 51468 6768
rect 51526 6748 51586 6768
rect 51644 6748 51704 6768
rect 51762 6768 52058 6804
rect 51762 6748 51822 6768
rect 51880 6748 51940 6768
rect 51998 6748 52058 6768
rect 49100 6666 49250 6682
rect 49100 6632 49116 6666
rect 49150 6632 49250 6666
rect 49100 6616 49250 6632
rect 49190 6578 49250 6616
rect 45105 6534 45121 6568
rect 45155 6534 45171 6568
rect 45105 6518 45171 6534
rect 44987 6451 45053 6467
rect 44987 6417 45003 6451
rect 45037 6417 45053 6451
rect 44987 6401 45053 6417
rect 44990 6379 45050 6401
rect 42641 6264 42701 6290
rect 39865 6064 39925 6090
rect 39983 6064 40043 6090
rect 40101 6064 40161 6090
rect 40219 6064 40279 6090
rect 41763 6064 41823 6090
rect 41881 6064 41941 6090
rect 41999 6064 42059 6090
rect 42117 6064 42177 6090
rect 45994 6352 46054 6378
rect 44990 6153 45050 6179
rect 47292 6352 47352 6378
rect 47892 6352 47952 6378
rect 52648 6615 52708 7313
rect 52950 7265 53246 7325
rect 52950 7242 53010 7265
rect 53068 7242 53128 7265
rect 53186 7242 53246 7265
rect 53304 7266 53600 7326
rect 53945 7325 54006 7345
rect 53304 7242 53364 7266
rect 53422 7242 53482 7266
rect 53540 7242 53600 7266
rect 53926 7309 54006 7325
rect 53926 7275 53941 7309
rect 53975 7275 54006 7309
rect 53926 7259 54006 7275
rect 53945 7236 54006 7259
rect 53946 7090 54006 7236
rect 53945 6917 54006 7090
rect 52950 6816 53010 6842
rect 52918 6675 52985 6682
rect 53068 6675 53128 6842
rect 53186 6816 53246 6842
rect 53304 6816 53364 6842
rect 52918 6666 53128 6675
rect 52918 6632 52934 6666
rect 52968 6632 53128 6666
rect 52918 6616 53128 6632
rect 52648 6599 52799 6615
rect 52648 6565 52749 6599
rect 52783 6565 52799 6599
rect 52648 6549 52799 6565
rect 51054 6522 51114 6548
rect 51172 6522 51232 6548
rect 51290 6522 51350 6548
rect 51408 6528 51468 6548
rect 51408 6522 51469 6528
rect 51526 6522 51586 6548
rect 51644 6522 51704 6548
rect 49190 6352 49250 6378
rect 51291 6337 51349 6522
rect 51291 6311 51351 6337
rect 51409 6311 51469 6522
rect 51762 6516 51822 6548
rect 51880 6522 51940 6548
rect 51998 6522 52058 6548
rect 51759 6500 51825 6516
rect 52648 6510 52708 6549
rect 53068 6510 53128 6616
rect 53422 6675 53482 6842
rect 53540 6816 53600 6842
rect 53565 6675 53632 6682
rect 53422 6666 53632 6675
rect 53422 6632 53582 6666
rect 53616 6632 53632 6666
rect 53422 6616 53632 6632
rect 53184 6582 53250 6598
rect 53184 6548 53200 6582
rect 53234 6548 53250 6582
rect 53184 6532 53250 6548
rect 53302 6583 53368 6598
rect 53302 6549 53318 6583
rect 53352 6549 53368 6583
rect 53302 6533 53368 6549
rect 53186 6510 53246 6532
rect 53304 6510 53364 6533
rect 53422 6510 53482 6616
rect 53946 6614 54006 6917
rect 53856 6598 54006 6614
rect 53856 6564 53872 6598
rect 53906 6564 54006 6598
rect 53856 6548 54006 6564
rect 53946 6510 54006 6548
rect 54546 6809 54606 7467
rect 55259 7465 55802 7516
rect 55844 7509 55920 7516
rect 55978 7509 56038 7535
rect 57918 7511 57934 7545
rect 57968 7511 57984 7545
rect 55844 7465 55919 7509
rect 57918 7495 57984 7511
rect 58033 7545 58107 7567
rect 58033 7511 58052 7545
rect 58086 7511 58107 7545
rect 60469 7820 60765 7871
rect 60469 7803 60529 7820
rect 60587 7803 60647 7820
rect 60705 7803 60765 7820
rect 61046 7803 61106 7829
rect 61164 7803 61224 7829
rect 61282 7803 61342 7829
rect 70459 7953 70513 8013
rect 70913 7953 71287 8013
rect 71329 8013 71398 8018
rect 71329 7999 71846 8013
rect 71329 7965 71346 7999
rect 71380 7965 71846 7999
rect 71329 7953 71846 7965
rect 72246 7953 72272 8013
rect 70459 7895 70498 7953
rect 71329 7949 71396 7953
rect 62367 7820 62663 7871
rect 70459 7835 70513 7895
rect 70913 7835 70939 7895
rect 62367 7803 62427 7820
rect 62485 7803 62545 7820
rect 62603 7803 62663 7820
rect 65766 7721 66062 7772
rect 65766 7706 65826 7721
rect 65884 7706 65944 7721
rect 66002 7706 66062 7721
rect 66120 7706 66180 7732
rect 66238 7706 66298 7732
rect 66356 7706 66416 7732
rect 59148 7586 59208 7603
rect 59266 7586 59326 7603
rect 59384 7586 59444 7603
rect 59632 7586 59692 7603
rect 59148 7535 59692 7586
rect 59750 7577 59810 7603
rect 59868 7577 59928 7603
rect 59986 7584 60046 7603
rect 60104 7584 60164 7603
rect 60222 7584 60282 7603
rect 60469 7584 60529 7603
rect 60587 7584 60647 7603
rect 54848 7265 55144 7325
rect 54848 7242 54908 7265
rect 54966 7242 55026 7265
rect 55084 7242 55144 7265
rect 55202 7266 55498 7326
rect 55202 7242 55262 7266
rect 55320 7242 55380 7266
rect 55438 7242 55498 7266
rect 55844 7312 55904 7465
rect 58033 7454 58107 7511
rect 59273 7454 59333 7535
rect 59986 7533 60529 7584
rect 60571 7577 60647 7584
rect 60705 7577 60765 7603
rect 61046 7586 61106 7603
rect 61164 7586 61224 7603
rect 61282 7586 61342 7603
rect 61530 7586 61590 7603
rect 60571 7533 60646 7577
rect 61046 7535 61590 7586
rect 61648 7577 61708 7603
rect 61766 7577 61826 7603
rect 61884 7584 61944 7603
rect 62002 7584 62062 7603
rect 62120 7584 62180 7603
rect 62367 7584 62427 7603
rect 62485 7584 62545 7603
rect 58033 7429 59333 7454
rect 58032 7381 59333 7429
rect 60571 7413 60631 7533
rect 55844 7288 56098 7312
rect 55844 7254 56048 7288
rect 56082 7254 56098 7288
rect 55844 7238 56098 7254
rect 54848 6816 54908 6842
rect 54546 6793 54613 6809
rect 54546 6759 54562 6793
rect 54596 6759 54613 6793
rect 54546 6743 54613 6759
rect 54546 6615 54606 6743
rect 54816 6675 54883 6682
rect 54966 6675 55026 6842
rect 55084 6816 55144 6842
rect 55202 6816 55262 6842
rect 54816 6666 55026 6675
rect 54816 6632 54832 6666
rect 54866 6632 55026 6666
rect 54816 6616 55026 6632
rect 54546 6599 54697 6615
rect 54546 6565 54647 6599
rect 54681 6565 54697 6599
rect 54546 6549 54697 6565
rect 54546 6510 54606 6549
rect 54966 6510 55026 6616
rect 55320 6675 55380 6842
rect 55438 6816 55498 6842
rect 55461 6676 55528 6683
rect 55455 6675 55528 6676
rect 55320 6667 55528 6675
rect 55320 6633 55478 6667
rect 55512 6633 55528 6667
rect 55320 6617 55528 6633
rect 55320 6616 55517 6617
rect 55082 6582 55148 6598
rect 55082 6548 55098 6582
rect 55132 6548 55148 6582
rect 55082 6532 55148 6548
rect 55200 6583 55266 6598
rect 55200 6549 55216 6583
rect 55250 6549 55266 6583
rect 55200 6533 55266 6549
rect 55084 6510 55144 6532
rect 55202 6510 55262 6533
rect 55320 6510 55380 6616
rect 55844 6614 55904 7238
rect 57679 6837 57975 6873
rect 57679 6816 57739 6837
rect 57797 6816 57857 6837
rect 57915 6816 57975 6837
rect 58033 6836 58329 6872
rect 58033 6816 58093 6836
rect 58151 6816 58211 6836
rect 58269 6816 58329 6836
rect 58387 6836 58683 6872
rect 58387 6816 58447 6836
rect 58505 6816 58565 6836
rect 58623 6816 58683 6836
rect 59273 6683 59333 7381
rect 59575 7333 59871 7393
rect 59575 7310 59635 7333
rect 59693 7310 59753 7333
rect 59811 7310 59871 7333
rect 59929 7334 60225 7394
rect 60570 7393 60631 7413
rect 59929 7310 59989 7334
rect 60047 7310 60107 7334
rect 60165 7310 60225 7334
rect 60551 7377 60631 7393
rect 60551 7343 60566 7377
rect 60600 7343 60631 7377
rect 60551 7327 60631 7343
rect 60570 7304 60631 7327
rect 60571 7158 60631 7304
rect 60570 6985 60631 7158
rect 59575 6884 59635 6910
rect 59543 6743 59610 6750
rect 59693 6743 59753 6910
rect 59811 6884 59871 6910
rect 59929 6884 59989 6910
rect 59543 6734 59753 6743
rect 59543 6700 59559 6734
rect 59593 6700 59753 6734
rect 59543 6684 59753 6700
rect 59273 6667 59424 6683
rect 59273 6633 59374 6667
rect 59408 6633 59424 6667
rect 59273 6617 59424 6633
rect 55754 6598 55904 6614
rect 55754 6564 55770 6598
rect 55804 6564 55904 6598
rect 57679 6590 57739 6616
rect 57797 6590 57857 6616
rect 57915 6590 57975 6616
rect 58033 6596 58093 6616
rect 58033 6590 58094 6596
rect 58151 6590 58211 6616
rect 58269 6590 58329 6616
rect 55754 6548 55904 6564
rect 55844 6510 55904 6548
rect 51759 6466 51775 6500
rect 51809 6466 51825 6500
rect 51759 6450 51825 6466
rect 51641 6383 51707 6399
rect 51641 6349 51657 6383
rect 51691 6349 51707 6383
rect 51641 6333 51707 6349
rect 51644 6311 51704 6333
rect 46414 6152 46474 6178
rect 46532 6152 46592 6178
rect 46650 6152 46710 6178
rect 46768 6152 46828 6178
rect 48312 6152 48372 6178
rect 48430 6152 48490 6178
rect 48548 6152 48608 6178
rect 48666 6152 48726 6178
rect 44637 5957 44697 5979
rect 44755 5957 44815 5979
rect 31205 5858 31271 5875
rect 38088 5869 38148 5891
rect 38206 5869 38266 5891
rect 25190 5682 25414 5696
rect 25190 5648 25364 5682
rect 25398 5648 25414 5682
rect 25190 5636 25414 5648
rect 24298 5324 24358 5350
rect 24266 5183 24333 5190
rect 24416 5183 24476 5350
rect 24534 5324 24594 5350
rect 24652 5324 24712 5350
rect 24266 5174 24476 5183
rect 24266 5140 24282 5174
rect 24316 5140 24476 5174
rect 24266 5124 24476 5140
rect 23892 5106 24042 5122
rect 23892 5072 23992 5106
rect 24026 5072 24042 5106
rect 23892 5056 24042 5072
rect 18985 4794 19045 4820
rect 19755 4792 19815 4818
rect 16142 4594 16202 4620
rect 16260 4594 16320 4620
rect 16378 4594 16438 4620
rect 16496 4594 16556 4620
rect 18211 4594 18271 4620
rect 18329 4594 18389 4620
rect 18447 4594 18507 4620
rect 18565 4594 18625 4620
rect 21053 4792 21113 4818
rect 21824 4794 21884 4820
rect 23892 5018 23952 5056
rect 24416 5018 24476 5124
rect 24770 5183 24830 5350
rect 24888 5324 24948 5350
rect 24913 5183 24980 5190
rect 24770 5174 24980 5183
rect 24770 5140 24930 5174
rect 24964 5140 24980 5174
rect 24770 5124 24980 5140
rect 24530 5091 24596 5106
rect 24530 5057 24546 5091
rect 24580 5057 24596 5091
rect 24530 5041 24596 5057
rect 24648 5090 24714 5106
rect 24648 5056 24664 5090
rect 24698 5056 24714 5090
rect 24534 5018 24594 5041
rect 24648 5040 24714 5056
rect 24652 5018 24712 5040
rect 24770 5018 24830 5124
rect 25190 5123 25250 5636
rect 30371 5596 30422 5783
rect 31205 5824 31221 5858
rect 31255 5824 31271 5858
rect 31205 5808 31271 5824
rect 38085 5853 38151 5869
rect 38085 5819 38101 5853
rect 38135 5819 38151 5853
rect 38085 5803 38151 5819
rect 38203 5853 38269 5869
rect 38203 5819 38219 5853
rect 38253 5819 38269 5853
rect 44634 5941 44700 5957
rect 44634 5907 44650 5941
rect 44684 5907 44700 5941
rect 44634 5891 44700 5907
rect 44752 5941 44818 5957
rect 44752 5907 44768 5941
rect 44802 5907 44818 5941
rect 44752 5891 44818 5907
rect 52648 6284 52708 6310
rect 51644 6085 51704 6111
rect 53946 6284 54006 6310
rect 54546 6284 54606 6310
rect 57916 6405 57974 6590
rect 57916 6379 57976 6405
rect 58034 6379 58094 6590
rect 58387 6584 58447 6616
rect 58505 6590 58565 6616
rect 58623 6590 58683 6616
rect 58384 6568 58450 6584
rect 59273 6578 59333 6617
rect 59693 6578 59753 6684
rect 60047 6743 60107 6910
rect 60165 6884 60225 6910
rect 60190 6743 60257 6750
rect 60047 6734 60257 6743
rect 60047 6700 60207 6734
rect 60241 6700 60257 6734
rect 60047 6684 60257 6700
rect 59809 6650 59875 6666
rect 59809 6616 59825 6650
rect 59859 6616 59875 6650
rect 59809 6600 59875 6616
rect 59927 6651 59993 6666
rect 59927 6617 59943 6651
rect 59977 6617 59993 6651
rect 59927 6601 59993 6617
rect 59811 6578 59871 6600
rect 59929 6578 59989 6601
rect 60047 6578 60107 6684
rect 60571 6682 60631 6985
rect 60481 6666 60631 6682
rect 60481 6632 60497 6666
rect 60531 6632 60631 6666
rect 60481 6616 60631 6632
rect 60571 6578 60631 6616
rect 61171 6877 61231 7535
rect 61884 7533 62427 7584
rect 62469 7577 62545 7584
rect 62603 7577 62663 7603
rect 62469 7533 62544 7577
rect 61473 7333 61769 7393
rect 61473 7310 61533 7333
rect 61591 7310 61651 7333
rect 61709 7310 61769 7333
rect 61827 7334 62123 7394
rect 61827 7310 61887 7334
rect 61945 7310 62005 7334
rect 62063 7310 62123 7334
rect 62469 7380 62529 7533
rect 65282 7506 65342 7532
rect 65400 7506 65460 7532
rect 65518 7506 65578 7532
rect 62469 7356 62723 7380
rect 62469 7322 62673 7356
rect 62707 7322 62723 7356
rect 62469 7306 62723 7322
rect 70459 7598 70513 7658
rect 70913 7598 70939 7658
rect 66603 7523 66899 7574
rect 66603 7506 66663 7523
rect 66721 7506 66781 7523
rect 66839 7506 66899 7523
rect 67075 7524 67371 7560
rect 67075 7503 67135 7524
rect 67193 7503 67253 7524
rect 67311 7503 67371 7524
rect 67429 7523 67725 7559
rect 67429 7503 67489 7523
rect 67547 7503 67607 7523
rect 67665 7503 67725 7523
rect 67783 7523 68079 7559
rect 67783 7503 67843 7523
rect 67901 7503 67961 7523
rect 68019 7503 68079 7523
rect 70459 7540 70498 7598
rect 71329 7540 71386 7949
rect 72327 7817 72378 8126
rect 61473 6884 61533 6910
rect 61171 6861 61238 6877
rect 61171 6827 61187 6861
rect 61221 6827 61238 6861
rect 61171 6811 61238 6827
rect 61171 6683 61231 6811
rect 61441 6743 61508 6750
rect 61591 6743 61651 6910
rect 61709 6884 61769 6910
rect 61827 6884 61887 6910
rect 61441 6734 61651 6743
rect 61441 6700 61457 6734
rect 61491 6700 61651 6734
rect 61441 6684 61651 6700
rect 61171 6667 61322 6683
rect 61171 6633 61272 6667
rect 61306 6633 61322 6667
rect 61171 6617 61322 6633
rect 61171 6578 61231 6617
rect 61591 6578 61651 6684
rect 61945 6743 62005 6910
rect 62063 6884 62123 6910
rect 62086 6744 62153 6751
rect 62080 6743 62153 6744
rect 61945 6735 62153 6743
rect 61945 6701 62103 6735
rect 62137 6701 62153 6735
rect 61945 6685 62153 6701
rect 61945 6684 62142 6685
rect 61707 6650 61773 6666
rect 61707 6616 61723 6650
rect 61757 6616 61773 6650
rect 61707 6600 61773 6616
rect 61825 6651 61891 6666
rect 61825 6617 61841 6651
rect 61875 6617 61891 6651
rect 61825 6601 61891 6617
rect 61709 6578 61769 6600
rect 61827 6578 61887 6601
rect 61945 6578 62005 6684
rect 62469 6682 62529 7306
rect 65282 7289 65342 7306
rect 65400 7289 65460 7306
rect 65518 7289 65578 7306
rect 65766 7289 65826 7306
rect 65282 7238 65826 7289
rect 65884 7280 65944 7306
rect 66002 7280 66062 7306
rect 66120 7287 66180 7306
rect 66238 7287 66298 7306
rect 66356 7287 66416 7306
rect 66603 7287 66663 7306
rect 66721 7287 66781 7306
rect 62379 6666 62529 6682
rect 62379 6632 62395 6666
rect 62429 6632 62529 6666
rect 65407 7034 65467 7238
rect 66120 7236 66663 7287
rect 66705 7280 66781 7287
rect 66839 7280 66899 7306
rect 70459 7480 70513 7540
rect 70913 7480 71386 7540
rect 71598 7757 71846 7817
rect 72046 7757 72378 7817
rect 70459 7422 70498 7480
rect 70459 7362 70513 7422
rect 70913 7362 70939 7422
rect 66705 7236 66780 7280
rect 67075 7277 67135 7303
rect 67193 7277 67253 7303
rect 67311 7277 67371 7303
rect 67429 7283 67489 7303
rect 67429 7277 67490 7283
rect 67547 7277 67607 7303
rect 67665 7277 67725 7303
rect 66705 7154 66765 7236
rect 66705 7136 66939 7154
rect 66705 7102 66888 7136
rect 66922 7102 66939 7136
rect 65709 7036 66005 7096
rect 65407 7017 65538 7034
rect 65407 6983 65488 7017
rect 65522 6983 65538 7017
rect 65709 7013 65769 7036
rect 65827 7013 65887 7036
rect 65945 7013 66005 7036
rect 66063 7037 66359 7097
rect 66063 7013 66123 7037
rect 66181 7013 66241 7037
rect 66299 7013 66359 7037
rect 66705 7086 66939 7102
rect 67312 7092 67370 7277
rect 65407 6966 65538 6983
rect 62379 6616 62529 6632
rect 62469 6578 62529 6616
rect 58384 6534 58400 6568
rect 58434 6534 58450 6568
rect 58384 6518 58450 6534
rect 58266 6451 58332 6467
rect 58266 6417 58282 6451
rect 58316 6417 58332 6451
rect 58266 6401 58332 6417
rect 58269 6379 58329 6401
rect 55844 6284 55904 6310
rect 53068 6084 53128 6110
rect 53186 6084 53246 6110
rect 53304 6084 53364 6110
rect 53422 6084 53482 6110
rect 54966 6084 55026 6110
rect 55084 6084 55144 6110
rect 55202 6084 55262 6110
rect 55320 6084 55380 6110
rect 59273 6352 59333 6378
rect 58269 6153 58329 6179
rect 60571 6352 60631 6378
rect 61171 6352 61231 6378
rect 63467 6419 63763 6455
rect 63467 6398 63527 6419
rect 63585 6398 63645 6419
rect 63703 6398 63763 6419
rect 63821 6418 64117 6454
rect 63821 6398 63881 6418
rect 63939 6398 63999 6418
rect 64057 6398 64117 6418
rect 64175 6418 64471 6454
rect 64175 6398 64235 6418
rect 64293 6398 64353 6418
rect 64411 6398 64471 6418
rect 62469 6352 62529 6378
rect 65407 6386 65467 6966
rect 65709 6587 65769 6613
rect 65677 6446 65744 6453
rect 65827 6446 65887 6613
rect 65945 6587 66005 6613
rect 66063 6587 66123 6613
rect 65677 6437 65887 6446
rect 65677 6403 65693 6437
rect 65727 6403 65887 6437
rect 65677 6387 65887 6403
rect 65407 6370 65558 6386
rect 65407 6336 65508 6370
rect 65542 6336 65558 6370
rect 65407 6320 65558 6336
rect 65407 6281 65467 6320
rect 65827 6281 65887 6387
rect 66181 6446 66241 6613
rect 66299 6587 66359 6613
rect 66324 6446 66391 6453
rect 66181 6437 66391 6446
rect 66181 6403 66341 6437
rect 66375 6403 66391 6437
rect 66181 6387 66391 6403
rect 65943 6353 66009 6369
rect 65943 6319 65959 6353
rect 65993 6319 66009 6353
rect 65943 6303 66009 6319
rect 66061 6354 66127 6369
rect 66061 6320 66077 6354
rect 66111 6320 66127 6354
rect 66061 6304 66127 6320
rect 65945 6281 66005 6303
rect 66063 6281 66123 6304
rect 66181 6281 66241 6387
rect 66705 6385 66765 7086
rect 67312 7066 67372 7092
rect 67430 7066 67490 7277
rect 67783 7271 67843 7303
rect 67901 7277 67961 7303
rect 68019 7277 68079 7303
rect 67780 7255 67846 7271
rect 67780 7221 67796 7255
rect 67830 7221 67846 7255
rect 67780 7205 67846 7221
rect 67662 7138 67728 7154
rect 67662 7104 67678 7138
rect 67712 7104 67728 7138
rect 67662 7088 67728 7104
rect 70658 7125 70713 7185
rect 70913 7125 70939 7185
rect 67665 7066 67725 7088
rect 70658 7067 70697 7125
rect 70658 7007 70713 7067
rect 70913 7007 70939 7067
rect 71059 7043 71125 7059
rect 71059 7009 71075 7043
rect 71109 7009 71125 7043
rect 70658 6949 70697 7007
rect 71059 6993 71125 7009
rect 71062 6949 71122 6993
rect 71598 6949 71643 7757
rect 70658 6889 70713 6949
rect 70913 6889 71643 6949
rect 67665 6840 67725 6866
rect 67312 6644 67372 6666
rect 67430 6644 67490 6666
rect 67309 6628 67375 6644
rect 67309 6594 67325 6628
rect 67359 6594 67375 6628
rect 67309 6578 67375 6594
rect 67427 6628 67493 6644
rect 67427 6594 67443 6628
rect 67477 6594 67493 6628
rect 67427 6578 67493 6594
rect 66615 6369 66765 6385
rect 66615 6335 66631 6369
rect 66665 6335 66765 6369
rect 66615 6319 66765 6335
rect 66705 6281 66765 6319
rect 59693 6152 59753 6178
rect 59811 6152 59871 6178
rect 59929 6152 59989 6178
rect 60047 6152 60107 6178
rect 61591 6152 61651 6178
rect 61709 6152 61769 6178
rect 61827 6152 61887 6178
rect 61945 6152 62005 6178
rect 63467 6172 63527 6198
rect 63585 6172 63645 6198
rect 63703 6172 63763 6198
rect 63821 6178 63881 6198
rect 63821 6172 63882 6178
rect 63939 6172 63999 6198
rect 64057 6172 64117 6198
rect 51291 5889 51351 5911
rect 51409 5889 51469 5911
rect 38203 5803 38269 5819
rect 51288 5873 51354 5889
rect 51288 5839 51304 5873
rect 51338 5839 51354 5873
rect 51288 5823 51354 5839
rect 51406 5873 51472 5889
rect 51406 5839 51422 5873
rect 51456 5839 51472 5873
rect 57916 5957 57976 5979
rect 58034 5957 58094 5979
rect 57913 5941 57979 5957
rect 57913 5907 57929 5941
rect 57963 5907 57979 5941
rect 57913 5891 57979 5907
rect 58031 5941 58097 5957
rect 58031 5907 58047 5941
rect 58081 5907 58097 5941
rect 63704 5987 63762 6172
rect 63704 5961 63764 5987
rect 63822 5961 63882 6172
rect 64175 6166 64235 6198
rect 64293 6172 64353 6198
rect 64411 6172 64471 6198
rect 64172 6150 64238 6166
rect 64172 6116 64188 6150
rect 64222 6116 64238 6150
rect 64172 6100 64238 6116
rect 65407 6055 65467 6081
rect 64054 6033 64120 6049
rect 64054 5999 64070 6033
rect 64104 5999 64120 6033
rect 64054 5983 64120 5999
rect 64057 5961 64117 5983
rect 58031 5891 58097 5907
rect 51406 5823 51472 5839
rect 30084 5536 30152 5596
rect 30352 5536 30422 5596
rect 31273 5568 31339 5584
rect 30509 5546 30563 5562
rect 30084 5478 30135 5536
rect 30509 5512 30519 5546
rect 30553 5512 30563 5546
rect 30509 5494 30563 5512
rect 31273 5534 31289 5568
rect 31323 5534 31339 5568
rect 70658 6189 70713 6249
rect 70913 6190 71643 6249
rect 70913 6189 71216 6190
rect 70658 6131 70697 6189
rect 71199 6132 71216 6189
rect 71271 6189 71643 6190
rect 71271 6132 71286 6189
rect 66705 6055 66765 6081
rect 70658 6071 70713 6131
rect 70913 6071 70939 6131
rect 71199 6113 71286 6132
rect 70658 6013 70697 6071
rect 70658 5953 70713 6013
rect 70913 5953 70939 6013
rect 65827 5855 65887 5881
rect 65945 5855 66005 5881
rect 66063 5855 66123 5881
rect 66181 5855 66241 5881
rect 64057 5735 64117 5761
rect 70459 5748 70513 5808
rect 70913 5748 70939 5808
rect 70459 5690 70498 5748
rect 70459 5630 70513 5690
rect 70913 5630 71388 5690
rect 70459 5572 70498 5630
rect 31273 5494 31339 5534
rect 63704 5539 63764 5561
rect 63822 5539 63882 5561
rect 63701 5523 63767 5539
rect 30371 5478 31377 5494
rect 30084 5418 30152 5478
rect 30352 5434 31377 5478
rect 31577 5434 31603 5494
rect 63701 5489 63717 5523
rect 63751 5489 63767 5523
rect 63701 5473 63767 5489
rect 63819 5523 63885 5539
rect 63819 5489 63835 5523
rect 63869 5489 63885 5523
rect 70459 5512 70513 5572
rect 70913 5512 70939 5572
rect 63819 5473 63885 5489
rect 30352 5419 30422 5434
rect 30352 5418 30378 5419
rect 30084 5360 30135 5418
rect 30084 5300 30152 5360
rect 30352 5300 30378 5360
rect 70459 5281 70513 5341
rect 70913 5281 70939 5341
rect 70459 5223 70498 5281
rect 70459 5163 70513 5223
rect 70913 5222 70939 5223
rect 71100 5222 71166 5225
rect 70913 5209 71166 5222
rect 70913 5175 71116 5209
rect 71150 5175 71166 5209
rect 70913 5163 71166 5175
rect 71331 5223 71388 5630
rect 71598 5415 71643 6189
rect 71598 5355 71846 5415
rect 72046 5355 72072 5415
rect 71487 5223 71566 5234
rect 71331 5221 71846 5223
rect 71331 5163 71500 5221
rect 71555 5163 71846 5221
rect 72246 5163 72272 5223
rect 25099 5107 25250 5123
rect 25099 5073 25115 5107
rect 25149 5073 25250 5107
rect 25099 5057 25250 5073
rect 25190 5018 25250 5057
rect 23122 4794 23182 4820
rect 23892 4792 23952 4818
rect 20279 4592 20339 4618
rect 20397 4592 20457 4618
rect 20515 4592 20575 4618
rect 20633 4592 20693 4618
rect 22348 4594 22408 4620
rect 22466 4594 22526 4620
rect 22584 4594 22644 4620
rect 22702 4594 22762 4620
rect 70459 5105 70498 5163
rect 71099 5159 71166 5163
rect 71487 5153 71566 5163
rect 71200 5105 71287 5122
rect 70459 5045 70513 5105
rect 70913 5045 70939 5105
rect 71200 5103 71846 5105
rect 71200 5045 71215 5103
rect 71270 5045 71846 5103
rect 72246 5045 72272 5105
rect 71200 5027 71287 5045
rect 30699 4871 30759 4887
rect 25190 4792 25250 4818
rect 30126 4788 30152 4848
rect 30352 4788 30420 4848
rect 30369 4730 30420 4788
rect 30126 4670 30152 4730
rect 30352 4723 30420 4730
rect 30699 4837 30713 4871
rect 30747 4837 30759 4871
rect 70459 4927 70513 4987
rect 70913 4927 70939 4987
rect 70459 4869 70498 4927
rect 71238 4869 71287 5027
rect 71720 4987 71786 4990
rect 72319 5032 72385 5048
rect 72319 4998 72335 5032
rect 72369 4998 72385 5032
rect 71720 4974 71846 4987
rect 71720 4940 71736 4974
rect 71770 4940 71846 4974
rect 71720 4927 71846 4940
rect 72246 4927 72272 4987
rect 72319 4982 72385 4998
rect 71720 4924 71786 4927
rect 30699 4723 30759 4837
rect 70459 4809 70513 4869
rect 70913 4809 71287 4869
rect 71329 4869 71398 4874
rect 71329 4855 71846 4869
rect 71329 4821 71346 4855
rect 71380 4821 71846 4855
rect 71329 4809 71846 4821
rect 72246 4809 72272 4869
rect 70459 4751 70498 4809
rect 71329 4805 71396 4809
rect 30352 4670 31377 4723
rect 24416 4592 24476 4618
rect 24534 4592 24594 4618
rect 24652 4592 24712 4618
rect 24770 4592 24830 4618
rect 30369 4663 31377 4670
rect 31577 4663 31603 4723
rect 30369 4612 30420 4663
rect 30126 4552 30152 4612
rect 30352 4552 30420 4612
rect 31272 4622 31338 4663
rect 31272 4588 31288 4622
rect 31322 4588 31338 4622
rect 31272 4572 31338 4588
rect 30369 4364 30420 4552
rect 31205 4437 31271 4453
rect 29886 4304 29952 4364
rect 30352 4304 30420 4364
rect 30562 4361 30645 4421
rect 31045 4361 31071 4421
rect 31205 4403 31221 4437
rect 31255 4403 31271 4437
rect 31205 4386 31271 4403
rect 34925 4407 35221 4443
rect 34925 4386 34985 4407
rect 35043 4386 35103 4407
rect 35161 4386 35221 4407
rect 35279 4406 35575 4442
rect 35279 4386 35339 4406
rect 35397 4386 35457 4406
rect 35515 4386 35575 4406
rect 35633 4406 35929 4442
rect 35633 4386 35693 4406
rect 35751 4386 35811 4406
rect 35869 4386 35929 4406
rect 39982 4438 40048 4454
rect 41112 4444 41178 4460
rect 39982 4404 39998 4438
rect 40032 4431 40048 4438
rect 40032 4404 40557 4431
rect 39982 4388 40557 4404
rect 41112 4410 41128 4444
rect 41162 4435 41178 4444
rect 41162 4410 41699 4435
rect 41112 4392 41699 4410
rect 29886 4246 29937 4304
rect 30562 4303 30622 4361
rect 31212 4303 31271 4386
rect 29886 4186 29952 4246
rect 30352 4186 30378 4246
rect 30562 4243 30645 4303
rect 31045 4243 31377 4303
rect 31777 4243 31803 4303
rect 29886 4128 29937 4186
rect 30562 4185 30622 4243
rect 31289 4185 31355 4187
rect 29886 4068 29952 4128
rect 30352 4068 30378 4128
rect 30562 4125 30645 4185
rect 31045 4125 31071 4185
rect 31289 4171 31377 4185
rect 31289 4137 31305 4171
rect 31339 4137 31377 4171
rect 31289 4125 31377 4137
rect 31777 4125 31803 4185
rect 40513 4336 40557 4388
rect 41655 4340 41699 4392
rect 46533 4436 46599 4452
rect 47663 4442 47729 4458
rect 46533 4402 46549 4436
rect 46583 4429 46599 4436
rect 46583 4402 47108 4429
rect 46533 4386 47108 4402
rect 47663 4408 47679 4442
rect 47713 4433 47729 4442
rect 47713 4408 48250 4433
rect 47663 4390 48250 4408
rect 39982 4320 40455 4336
rect 39982 4286 39998 4320
rect 40032 4295 40455 4320
rect 40032 4294 40219 4295
rect 40032 4286 40048 4294
rect 39982 4270 40048 4286
rect 40159 4274 40219 4294
rect 40277 4274 40337 4295
rect 40395 4274 40455 4295
rect 40513 4295 40809 4336
rect 40513 4274 40573 4295
rect 40631 4274 40691 4295
rect 40749 4274 40809 4295
rect 41112 4324 41597 4340
rect 41112 4290 41128 4324
rect 41162 4299 41597 4324
rect 41162 4298 41361 4299
rect 41162 4290 41178 4298
rect 41112 4274 41178 4290
rect 41301 4278 41361 4298
rect 41419 4278 41479 4299
rect 41537 4278 41597 4299
rect 41655 4299 41951 4340
rect 47064 4334 47108 4386
rect 48206 4338 48250 4390
rect 53188 4437 53254 4453
rect 54318 4443 54384 4459
rect 53188 4403 53204 4437
rect 53238 4430 53254 4437
rect 53238 4403 53763 4430
rect 53188 4387 53763 4403
rect 54318 4409 54334 4443
rect 54368 4434 54384 4443
rect 54368 4409 54905 4434
rect 54318 4391 54905 4409
rect 41655 4278 41715 4299
rect 41773 4278 41833 4299
rect 41891 4278 41951 4299
rect 46533 4318 47006 4334
rect 46533 4284 46549 4318
rect 46583 4293 47006 4318
rect 46583 4292 46770 4293
rect 46583 4284 46599 4292
rect 37834 4223 38130 4259
rect 37834 4202 37894 4223
rect 37952 4202 38012 4223
rect 38070 4202 38130 4223
rect 38188 4222 38484 4258
rect 38188 4202 38248 4222
rect 38306 4202 38366 4222
rect 38424 4202 38484 4222
rect 38542 4222 38838 4258
rect 38542 4202 38602 4222
rect 38660 4202 38720 4222
rect 38778 4202 38838 4222
rect 34925 4160 34985 4186
rect 35043 4160 35103 4186
rect 35161 4160 35221 4186
rect 35279 4166 35339 4186
rect 35279 4160 35340 4166
rect 35397 4160 35457 4186
rect 35515 4160 35575 4186
rect 31289 4121 31355 4125
rect 31289 4067 31354 4069
rect 29926 3950 29952 4010
rect 30352 3950 30422 4010
rect 30371 3892 30422 3950
rect 29926 3832 29952 3892
rect 30352 3832 30422 3892
rect 30371 3774 30422 3832
rect 29926 3714 29952 3774
rect 30352 3714 30422 3774
rect 30561 4007 30645 4067
rect 31045 4007 31071 4067
rect 31289 4053 31377 4067
rect 31289 4019 31304 4053
rect 31338 4019 31377 4053
rect 31289 4007 31377 4019
rect 31777 4007 31803 4067
rect 30561 3949 30621 4007
rect 31289 4003 31354 4007
rect 35162 3975 35220 4160
rect 35162 3949 35222 3975
rect 35280 3949 35340 4160
rect 35633 4154 35693 4186
rect 35751 4160 35811 4186
rect 35869 4160 35929 4186
rect 35630 4138 35696 4154
rect 35630 4104 35646 4138
rect 35680 4104 35696 4138
rect 35630 4088 35696 4104
rect 35512 4021 35578 4037
rect 35512 3987 35528 4021
rect 35562 3987 35578 4021
rect 35512 3971 35578 3987
rect 37834 3976 37894 4002
rect 37952 3976 38012 4002
rect 38070 3976 38130 4002
rect 38188 3982 38248 4002
rect 38188 3976 38249 3982
rect 38306 3976 38366 4002
rect 38424 3976 38484 4002
rect 35515 3949 35575 3971
rect 30561 3889 30645 3949
rect 31045 3889 31377 3949
rect 31777 3889 31803 3949
rect 30561 3831 30621 3889
rect 30561 3771 30645 3831
rect 31045 3771 31071 3831
rect 31212 3806 31271 3889
rect 31205 3789 31271 3806
rect 30371 3527 30422 3714
rect 31205 3755 31221 3789
rect 31255 3755 31271 3789
rect 31205 3739 31271 3755
rect 38071 3791 38129 3976
rect 38071 3765 38131 3791
rect 38189 3765 38249 3976
rect 38542 3970 38602 4002
rect 38660 3976 38720 4002
rect 38778 3976 38838 4002
rect 38539 3954 38605 3970
rect 38539 3920 38555 3954
rect 38589 3920 38605 3954
rect 38539 3904 38605 3920
rect 46533 4268 46599 4284
rect 46710 4272 46770 4292
rect 46828 4272 46888 4293
rect 46946 4272 47006 4293
rect 47064 4293 47360 4334
rect 47064 4272 47124 4293
rect 47182 4272 47242 4293
rect 47300 4272 47360 4293
rect 47663 4322 48148 4338
rect 47663 4288 47679 4322
rect 47713 4297 48148 4322
rect 47713 4296 47912 4297
rect 47713 4288 47729 4296
rect 47663 4272 47729 4288
rect 47852 4276 47912 4296
rect 47970 4276 48030 4297
rect 48088 4276 48148 4297
rect 48206 4297 48502 4338
rect 53719 4335 53763 4387
rect 54861 4339 54905 4391
rect 59810 4438 59876 4454
rect 70459 4691 70513 4751
rect 70913 4691 70939 4751
rect 60940 4444 61006 4460
rect 59810 4404 59826 4438
rect 59860 4431 59876 4438
rect 59860 4404 60385 4431
rect 59810 4388 60385 4404
rect 60940 4410 60956 4444
rect 60990 4435 61006 4444
rect 63538 4499 63834 4535
rect 63538 4478 63598 4499
rect 63656 4478 63716 4499
rect 63774 4478 63834 4499
rect 63892 4498 64188 4534
rect 63892 4478 63952 4498
rect 64010 4478 64070 4498
rect 64128 4478 64188 4498
rect 64246 4498 64542 4534
rect 64246 4478 64306 4498
rect 64364 4478 64424 4498
rect 64482 4478 64542 4498
rect 60990 4410 61527 4435
rect 60940 4392 61527 4410
rect 48206 4276 48266 4297
rect 48324 4276 48384 4297
rect 48442 4276 48502 4297
rect 53188 4319 53661 4335
rect 53188 4285 53204 4319
rect 53238 4294 53661 4319
rect 53238 4293 53425 4294
rect 53238 4285 53254 4293
rect 44385 4221 44681 4257
rect 44385 4200 44445 4221
rect 44503 4200 44563 4221
rect 44621 4200 44681 4221
rect 44739 4220 45035 4256
rect 44739 4200 44799 4220
rect 44857 4200 44917 4220
rect 44975 4200 45035 4220
rect 45093 4220 45389 4256
rect 45093 4200 45153 4220
rect 45211 4200 45271 4220
rect 45329 4200 45389 4220
rect 44385 3974 44445 4000
rect 44503 3974 44563 4000
rect 44621 3974 44681 4000
rect 44739 3980 44799 4000
rect 44739 3974 44800 3980
rect 44857 3974 44917 4000
rect 44975 3974 45035 4000
rect 40159 3857 40219 3874
rect 38421 3837 38487 3853
rect 38421 3803 38437 3837
rect 38471 3803 38487 3837
rect 38421 3787 38487 3803
rect 38424 3765 38484 3787
rect 40159 3768 40220 3857
rect 40277 3848 40337 3874
rect 40395 3848 40455 3874
rect 35515 3723 35575 3749
rect 35162 3527 35222 3549
rect 35280 3527 35340 3549
rect 30084 3467 30152 3527
rect 30352 3467 30422 3527
rect 31273 3499 31339 3515
rect 30509 3477 30563 3493
rect 30084 3409 30135 3467
rect 30509 3443 30519 3477
rect 30553 3443 30563 3477
rect 30509 3425 30563 3443
rect 31273 3465 31289 3499
rect 31323 3465 31339 3499
rect 35159 3511 35225 3527
rect 31273 3425 31339 3465
rect 35159 3477 35175 3511
rect 35209 3477 35225 3511
rect 35159 3461 35225 3477
rect 35277 3511 35343 3527
rect 35277 3477 35293 3511
rect 35327 3477 35343 3511
rect 35277 3461 35343 3477
rect 30371 3409 31377 3425
rect 30084 3349 30152 3409
rect 30352 3365 31377 3409
rect 31577 3365 31603 3425
rect 30352 3350 30422 3365
rect 30352 3349 30378 3350
rect 30084 3291 30135 3349
rect 40069 3715 40220 3768
rect 38424 3539 38484 3565
rect 40069 3491 40129 3715
rect 40513 3673 40573 3874
rect 40631 3848 40691 3874
rect 40749 3848 40809 3874
rect 41301 3861 41361 3878
rect 41301 3772 41362 3861
rect 41419 3852 41479 3878
rect 41537 3852 41597 3878
rect 40187 3622 40573 3673
rect 41211 3719 41362 3772
rect 40187 3491 40247 3622
rect 40302 3564 40368 3580
rect 40302 3530 40318 3564
rect 40352 3530 40368 3564
rect 40302 3514 40368 3530
rect 40305 3491 40365 3514
rect 40588 3491 40648 3517
rect 40706 3491 40766 3517
rect 40824 3491 40884 3517
rect 41211 3495 41271 3719
rect 41655 3677 41715 3878
rect 41773 3852 41833 3878
rect 41891 3852 41951 3878
rect 44622 3789 44680 3974
rect 44622 3763 44682 3789
rect 44740 3763 44800 3974
rect 45093 3968 45153 4000
rect 45211 3974 45271 4000
rect 45329 3974 45389 4000
rect 45090 3952 45156 3968
rect 45090 3918 45106 3952
rect 45140 3918 45156 3952
rect 45090 3902 45156 3918
rect 53188 4269 53254 4285
rect 53365 4273 53425 4293
rect 53483 4273 53543 4294
rect 53601 4273 53661 4294
rect 53719 4294 54015 4335
rect 53719 4273 53779 4294
rect 53837 4273 53897 4294
rect 53955 4273 54015 4294
rect 54318 4323 54803 4339
rect 54318 4289 54334 4323
rect 54368 4298 54803 4323
rect 54368 4297 54567 4298
rect 54368 4289 54384 4297
rect 54318 4273 54384 4289
rect 54507 4277 54567 4297
rect 54625 4277 54685 4298
rect 54743 4277 54803 4298
rect 54861 4298 55157 4339
rect 60341 4336 60385 4388
rect 61483 4340 61527 4392
rect 54861 4277 54921 4298
rect 54979 4277 55039 4298
rect 55097 4277 55157 4298
rect 59810 4320 60283 4336
rect 59810 4286 59826 4320
rect 59860 4295 60283 4320
rect 59860 4294 60047 4295
rect 59860 4286 59876 4294
rect 51040 4222 51336 4258
rect 51040 4201 51100 4222
rect 51158 4201 51218 4222
rect 51276 4201 51336 4222
rect 51394 4221 51690 4257
rect 51394 4201 51454 4221
rect 51512 4201 51572 4221
rect 51630 4201 51690 4221
rect 51748 4221 52044 4257
rect 51748 4201 51808 4221
rect 51866 4201 51926 4221
rect 51984 4201 52044 4221
rect 51040 3975 51100 4001
rect 51158 3975 51218 4001
rect 51276 3975 51336 4001
rect 51394 3981 51454 4001
rect 51394 3975 51455 3981
rect 51512 3975 51572 4001
rect 51630 3975 51690 4001
rect 46710 3855 46770 3872
rect 44972 3835 45038 3851
rect 44972 3801 44988 3835
rect 45022 3801 45038 3835
rect 44972 3785 45038 3801
rect 44975 3763 45035 3785
rect 46710 3766 46771 3855
rect 46828 3846 46888 3872
rect 46946 3846 47006 3872
rect 41329 3626 41715 3677
rect 41329 3495 41389 3626
rect 41444 3568 41510 3584
rect 41444 3534 41460 3568
rect 41494 3534 41510 3568
rect 41444 3518 41510 3534
rect 41447 3495 41507 3518
rect 41730 3495 41790 3521
rect 41848 3495 41908 3521
rect 41966 3495 42026 3521
rect 38071 3343 38131 3365
rect 38189 3343 38249 3365
rect 38068 3327 38134 3343
rect 38068 3293 38084 3327
rect 38118 3293 38134 3327
rect 30084 3231 30152 3291
rect 30352 3231 30378 3291
rect 38068 3277 38134 3293
rect 38186 3327 38252 3343
rect 38186 3293 38202 3327
rect 38236 3293 38252 3327
rect 38186 3277 38252 3293
rect 46620 3713 46771 3766
rect 44975 3537 45035 3563
rect 46620 3489 46680 3713
rect 47064 3671 47124 3872
rect 47182 3846 47242 3872
rect 47300 3846 47360 3872
rect 47852 3859 47912 3876
rect 47852 3770 47913 3859
rect 47970 3850 48030 3876
rect 48088 3850 48148 3876
rect 46738 3620 47124 3671
rect 47762 3717 47913 3770
rect 46738 3489 46798 3620
rect 46853 3562 46919 3578
rect 46853 3528 46869 3562
rect 46903 3528 46919 3562
rect 46853 3512 46919 3528
rect 46856 3489 46916 3512
rect 47139 3489 47199 3515
rect 47257 3489 47317 3515
rect 47375 3489 47435 3515
rect 47762 3493 47822 3717
rect 48206 3675 48266 3876
rect 48324 3850 48384 3876
rect 48442 3850 48502 3876
rect 51277 3790 51335 3975
rect 51277 3764 51337 3790
rect 51395 3764 51455 3975
rect 51748 3969 51808 4001
rect 51866 3975 51926 4001
rect 51984 3975 52044 4001
rect 51745 3953 51811 3969
rect 51745 3919 51761 3953
rect 51795 3919 51811 3953
rect 51745 3903 51811 3919
rect 59810 4270 59876 4286
rect 59987 4274 60047 4294
rect 60105 4274 60165 4295
rect 60223 4274 60283 4295
rect 60341 4295 60637 4336
rect 60341 4274 60401 4295
rect 60459 4274 60519 4295
rect 60577 4274 60637 4295
rect 60940 4324 61425 4340
rect 60940 4290 60956 4324
rect 60990 4299 61425 4324
rect 60990 4298 61189 4299
rect 60990 4290 61006 4298
rect 60940 4274 61006 4290
rect 61129 4278 61189 4298
rect 61247 4278 61307 4299
rect 61365 4278 61425 4299
rect 61483 4299 61779 4340
rect 61483 4278 61543 4299
rect 61601 4278 61661 4299
rect 61719 4278 61779 4299
rect 70459 4454 70513 4514
rect 70913 4454 70939 4514
rect 70459 4396 70498 4454
rect 71329 4396 71386 4805
rect 72327 4673 72378 4982
rect 70459 4336 70513 4396
rect 70913 4336 71386 4396
rect 71598 4613 71846 4673
rect 72046 4613 72378 4673
rect 70459 4278 70498 4336
rect 57662 4223 57958 4259
rect 57662 4202 57722 4223
rect 57780 4202 57840 4223
rect 57898 4202 57958 4223
rect 58016 4222 58312 4258
rect 58016 4202 58076 4222
rect 58134 4202 58194 4222
rect 58252 4202 58312 4222
rect 58370 4222 58666 4258
rect 58370 4202 58430 4222
rect 58488 4202 58548 4222
rect 58606 4202 58666 4222
rect 57662 3976 57722 4002
rect 57780 3976 57840 4002
rect 57898 3976 57958 4002
rect 58016 3982 58076 4002
rect 58016 3976 58077 3982
rect 58134 3976 58194 4002
rect 58252 3976 58312 4002
rect 53365 3856 53425 3873
rect 51627 3836 51693 3852
rect 51627 3802 51643 3836
rect 51677 3802 51693 3836
rect 51627 3786 51693 3802
rect 51630 3764 51690 3786
rect 53365 3767 53426 3856
rect 53483 3847 53543 3873
rect 53601 3847 53661 3873
rect 47880 3624 48266 3675
rect 47880 3493 47940 3624
rect 47995 3566 48061 3582
rect 47995 3532 48011 3566
rect 48045 3532 48061 3566
rect 47995 3516 48061 3532
rect 47998 3493 48058 3516
rect 48281 3493 48341 3519
rect 48399 3493 48459 3519
rect 48517 3493 48577 3519
rect 44622 3341 44682 3363
rect 44740 3341 44800 3363
rect 44619 3325 44685 3341
rect 40069 3265 40129 3291
rect 40187 3265 40247 3291
rect 40305 3259 40365 3291
rect 40588 3259 40648 3291
rect 40706 3259 40766 3291
rect 40824 3259 40884 3291
rect 41211 3269 41271 3295
rect 41329 3269 41389 3295
rect 40305 3218 40884 3259
rect 41447 3263 41507 3295
rect 41730 3263 41790 3295
rect 41848 3263 41908 3295
rect 41966 3263 42026 3295
rect 44619 3291 44635 3325
rect 44669 3291 44685 3325
rect 44619 3275 44685 3291
rect 44737 3325 44803 3341
rect 44737 3291 44753 3325
rect 44787 3291 44803 3325
rect 44737 3275 44803 3291
rect 53275 3714 53426 3767
rect 51630 3538 51690 3564
rect 53275 3490 53335 3714
rect 53719 3672 53779 3873
rect 53837 3847 53897 3873
rect 53955 3847 54015 3873
rect 54507 3860 54567 3877
rect 54507 3771 54568 3860
rect 54625 3851 54685 3877
rect 54743 3851 54803 3877
rect 53393 3621 53779 3672
rect 54417 3718 54568 3771
rect 53393 3490 53453 3621
rect 53508 3563 53574 3579
rect 53508 3529 53524 3563
rect 53558 3529 53574 3563
rect 53508 3513 53574 3529
rect 53511 3490 53571 3513
rect 53794 3490 53854 3516
rect 53912 3490 53972 3516
rect 54030 3490 54090 3516
rect 54417 3494 54477 3718
rect 54861 3676 54921 3877
rect 54979 3851 55039 3877
rect 55097 3851 55157 3877
rect 57899 3791 57957 3976
rect 57899 3765 57959 3791
rect 58017 3765 58077 3976
rect 58370 3970 58430 4002
rect 58488 3976 58548 4002
rect 58606 3976 58666 4002
rect 58367 3954 58433 3970
rect 58367 3920 58383 3954
rect 58417 3920 58433 3954
rect 58367 3904 58433 3920
rect 63538 4252 63598 4278
rect 63656 4252 63716 4278
rect 63774 4252 63834 4278
rect 63892 4258 63952 4278
rect 63892 4252 63953 4258
rect 64010 4252 64070 4278
rect 64128 4252 64188 4278
rect 63775 4067 63833 4252
rect 63775 4041 63835 4067
rect 63893 4041 63953 4252
rect 64246 4246 64306 4278
rect 64364 4252 64424 4278
rect 64482 4252 64542 4278
rect 64243 4230 64309 4246
rect 64243 4196 64259 4230
rect 64293 4196 64309 4230
rect 65766 4226 66062 4277
rect 65766 4211 65826 4226
rect 65884 4211 65944 4226
rect 66002 4211 66062 4226
rect 66120 4211 66180 4237
rect 66238 4211 66298 4237
rect 66356 4211 66416 4237
rect 64243 4180 64309 4196
rect 64125 4113 64191 4129
rect 64125 4079 64141 4113
rect 64175 4079 64191 4113
rect 64125 4063 64191 4079
rect 64128 4041 64188 4063
rect 59987 3857 60047 3874
rect 58249 3837 58315 3853
rect 58249 3803 58265 3837
rect 58299 3803 58315 3837
rect 58249 3787 58315 3803
rect 58252 3765 58312 3787
rect 59987 3768 60048 3857
rect 60105 3848 60165 3874
rect 60223 3848 60283 3874
rect 54535 3625 54921 3676
rect 54535 3494 54595 3625
rect 54650 3567 54716 3583
rect 54650 3533 54666 3567
rect 54700 3533 54716 3567
rect 54650 3517 54716 3533
rect 54653 3494 54713 3517
rect 54936 3494 54996 3520
rect 55054 3494 55114 3520
rect 55172 3494 55232 3520
rect 51277 3342 51337 3364
rect 51395 3342 51455 3364
rect 51274 3326 51340 3342
rect 46620 3263 46680 3289
rect 46738 3263 46798 3289
rect 41447 3222 42026 3263
rect 46856 3257 46916 3289
rect 47139 3257 47199 3289
rect 47257 3257 47317 3289
rect 47375 3257 47435 3289
rect 47762 3267 47822 3293
rect 47880 3267 47940 3293
rect 46856 3216 47435 3257
rect 47998 3261 48058 3293
rect 48281 3261 48341 3293
rect 48399 3261 48459 3293
rect 48517 3261 48577 3293
rect 51274 3292 51290 3326
rect 51324 3292 51340 3326
rect 51274 3276 51340 3292
rect 51392 3326 51458 3342
rect 51392 3292 51408 3326
rect 51442 3292 51458 3326
rect 51392 3276 51458 3292
rect 59897 3715 60048 3768
rect 58252 3539 58312 3565
rect 59897 3491 59957 3715
rect 60341 3673 60401 3874
rect 60459 3848 60519 3874
rect 60577 3848 60637 3874
rect 61129 3861 61189 3878
rect 61129 3772 61190 3861
rect 61247 3852 61307 3878
rect 61365 3852 61425 3878
rect 60015 3622 60401 3673
rect 61039 3719 61190 3772
rect 60015 3491 60075 3622
rect 60130 3564 60196 3580
rect 60130 3530 60146 3564
rect 60180 3530 60196 3564
rect 60130 3514 60196 3530
rect 60133 3491 60193 3514
rect 60416 3491 60476 3517
rect 60534 3491 60594 3517
rect 60652 3491 60712 3517
rect 61039 3495 61099 3719
rect 61483 3677 61543 3878
rect 61601 3852 61661 3878
rect 61719 3852 61779 3878
rect 61157 3626 61543 3677
rect 65282 4011 65342 4037
rect 65400 4011 65460 4037
rect 65518 4011 65578 4037
rect 64128 3815 64188 3841
rect 70459 4218 70513 4278
rect 70913 4218 70939 4278
rect 66603 4028 66899 4079
rect 66603 4011 66663 4028
rect 66721 4011 66781 4028
rect 66839 4011 66899 4028
rect 67075 4029 67371 4065
rect 67075 4008 67135 4029
rect 67193 4008 67253 4029
rect 67311 4008 67371 4029
rect 67429 4028 67725 4064
rect 67429 4008 67489 4028
rect 67547 4008 67607 4028
rect 67665 4008 67725 4028
rect 67783 4028 68079 4064
rect 67783 4008 67843 4028
rect 67901 4008 67961 4028
rect 68019 4008 68079 4028
rect 65282 3794 65342 3811
rect 65400 3794 65460 3811
rect 65518 3794 65578 3811
rect 65766 3794 65826 3811
rect 65282 3743 65826 3794
rect 65884 3785 65944 3811
rect 66002 3785 66062 3811
rect 66120 3792 66180 3811
rect 66238 3792 66298 3811
rect 66356 3792 66416 3811
rect 66603 3792 66663 3811
rect 66721 3792 66781 3811
rect 61157 3495 61217 3626
rect 63775 3619 63835 3641
rect 63893 3619 63953 3641
rect 63772 3603 63838 3619
rect 61272 3568 61338 3584
rect 61272 3534 61288 3568
rect 61322 3534 61338 3568
rect 63772 3569 63788 3603
rect 63822 3569 63838 3603
rect 63772 3553 63838 3569
rect 63890 3603 63956 3619
rect 63890 3569 63906 3603
rect 63940 3569 63956 3603
rect 63890 3553 63956 3569
rect 61272 3518 61338 3534
rect 65407 3539 65467 3743
rect 66120 3741 66663 3792
rect 66705 3785 66781 3792
rect 66839 3785 66899 3811
rect 70658 3981 70713 4041
rect 70913 3981 70939 4041
rect 70658 3923 70697 3981
rect 70658 3863 70713 3923
rect 70913 3863 70939 3923
rect 71059 3899 71125 3915
rect 71059 3865 71075 3899
rect 71109 3865 71125 3899
rect 66705 3741 66780 3785
rect 67075 3782 67135 3808
rect 67193 3782 67253 3808
rect 67311 3782 67371 3808
rect 67429 3788 67489 3808
rect 67429 3782 67490 3788
rect 67547 3782 67607 3808
rect 67665 3782 67725 3808
rect 66705 3659 66765 3741
rect 66705 3641 66939 3659
rect 66705 3607 66888 3641
rect 66922 3607 66939 3641
rect 65709 3541 66005 3601
rect 61275 3495 61335 3518
rect 61558 3495 61618 3521
rect 61676 3495 61736 3521
rect 61794 3495 61854 3521
rect 57899 3343 57959 3365
rect 58017 3343 58077 3365
rect 57896 3327 57962 3343
rect 53275 3264 53335 3290
rect 53393 3264 53453 3290
rect 47998 3220 48577 3261
rect 53511 3258 53571 3290
rect 53794 3258 53854 3290
rect 53912 3258 53972 3290
rect 54030 3258 54090 3290
rect 54417 3268 54477 3294
rect 54535 3268 54595 3294
rect 53511 3217 54090 3258
rect 54653 3262 54713 3294
rect 54936 3262 54996 3294
rect 55054 3262 55114 3294
rect 55172 3262 55232 3294
rect 57896 3293 57912 3327
rect 57946 3293 57962 3327
rect 57896 3277 57962 3293
rect 58014 3327 58080 3343
rect 58014 3293 58030 3327
rect 58064 3293 58080 3327
rect 58014 3277 58080 3293
rect 65407 3522 65538 3539
rect 65407 3488 65488 3522
rect 65522 3488 65538 3522
rect 65709 3518 65769 3541
rect 65827 3518 65887 3541
rect 65945 3518 66005 3541
rect 66063 3542 66359 3602
rect 66063 3518 66123 3542
rect 66181 3518 66241 3542
rect 66299 3518 66359 3542
rect 66705 3591 66939 3607
rect 67312 3597 67370 3782
rect 65407 3471 65538 3488
rect 59897 3265 59957 3291
rect 60015 3265 60075 3291
rect 54653 3221 55232 3262
rect 60133 3259 60193 3291
rect 60416 3259 60476 3291
rect 60534 3259 60594 3291
rect 60652 3259 60712 3291
rect 61039 3269 61099 3295
rect 61157 3269 61217 3295
rect 60133 3218 60712 3259
rect 61275 3263 61335 3295
rect 61558 3263 61618 3295
rect 61676 3263 61736 3295
rect 61794 3263 61854 3295
rect 61275 3222 61854 3263
rect 30697 2803 30757 2819
rect 30124 2720 30150 2780
rect 30350 2720 30418 2780
rect 30367 2662 30418 2720
rect 30124 2602 30150 2662
rect 30350 2655 30418 2662
rect 30697 2769 30711 2803
rect 30745 2769 30757 2803
rect 30697 2655 30757 2769
rect 65407 2891 65467 3471
rect 65709 3092 65769 3118
rect 65677 2951 65744 2958
rect 65827 2951 65887 3118
rect 65945 3092 66005 3118
rect 66063 3092 66123 3118
rect 65677 2942 65887 2951
rect 65677 2908 65693 2942
rect 65727 2908 65887 2942
rect 65677 2892 65887 2908
rect 65407 2875 65558 2891
rect 65407 2841 65508 2875
rect 65542 2841 65558 2875
rect 65407 2825 65558 2841
rect 65407 2786 65467 2825
rect 65827 2786 65887 2892
rect 66181 2951 66241 3118
rect 66299 3092 66359 3118
rect 66324 2951 66391 2958
rect 66181 2942 66391 2951
rect 66181 2908 66341 2942
rect 66375 2908 66391 2942
rect 66181 2892 66391 2908
rect 65943 2858 66009 2874
rect 65943 2824 65959 2858
rect 65993 2824 66009 2858
rect 65943 2808 66009 2824
rect 66061 2859 66127 2874
rect 66061 2825 66077 2859
rect 66111 2825 66127 2859
rect 66061 2809 66127 2825
rect 65945 2786 66005 2808
rect 66063 2786 66123 2809
rect 66181 2786 66241 2892
rect 66705 2890 66765 3591
rect 67312 3571 67372 3597
rect 67430 3571 67490 3782
rect 67783 3776 67843 3808
rect 67901 3782 67961 3808
rect 68019 3782 68079 3808
rect 70658 3805 70697 3863
rect 71059 3849 71125 3865
rect 71062 3805 71122 3849
rect 71598 3805 71643 4613
rect 67780 3760 67846 3776
rect 67780 3726 67796 3760
rect 67830 3726 67846 3760
rect 70658 3745 70713 3805
rect 70913 3745 71643 3805
rect 67780 3710 67846 3726
rect 67662 3643 67728 3659
rect 67662 3609 67678 3643
rect 67712 3609 67728 3643
rect 67662 3593 67728 3609
rect 67665 3571 67725 3593
rect 67665 3345 67725 3371
rect 67312 3149 67372 3171
rect 67430 3149 67490 3171
rect 67309 3133 67375 3149
rect 67309 3099 67325 3133
rect 67359 3099 67375 3133
rect 67309 3083 67375 3099
rect 67427 3133 67493 3149
rect 67427 3099 67443 3133
rect 67477 3099 67493 3133
rect 67427 3083 67493 3099
rect 70654 3057 70709 3117
rect 70909 3058 71639 3117
rect 70909 3057 71212 3058
rect 70654 2999 70693 3057
rect 71195 3000 71212 3057
rect 71267 3057 71639 3058
rect 71267 3000 71282 3057
rect 66615 2874 66765 2890
rect 66615 2840 66631 2874
rect 66665 2840 66765 2874
rect 66615 2824 66765 2840
rect 66705 2786 66765 2824
rect 70654 2939 70709 2999
rect 70909 2939 70935 2999
rect 71195 2981 71282 3000
rect 70654 2881 70693 2939
rect 70654 2821 70709 2881
rect 70909 2821 70935 2881
rect 30350 2602 31375 2655
rect 30367 2595 31375 2602
rect 31575 2595 31601 2655
rect 30367 2544 30418 2595
rect 30124 2484 30150 2544
rect 30350 2484 30418 2544
rect 31270 2554 31336 2595
rect 31270 2520 31286 2554
rect 31320 2520 31336 2554
rect 37848 2573 38144 2609
rect 37848 2552 37908 2573
rect 37966 2552 38026 2573
rect 38084 2552 38144 2573
rect 38202 2572 38498 2608
rect 38202 2552 38262 2572
rect 38320 2552 38380 2572
rect 38438 2552 38498 2572
rect 38556 2572 38852 2608
rect 38556 2552 38616 2572
rect 38674 2552 38734 2572
rect 38792 2552 38852 2572
rect 31270 2504 31336 2520
rect 30367 2296 30418 2484
rect 31203 2369 31269 2385
rect 29884 2236 29950 2296
rect 30350 2236 30418 2296
rect 30560 2293 30643 2353
rect 31043 2293 31069 2353
rect 31203 2335 31219 2369
rect 31253 2335 31269 2369
rect 44399 2571 44695 2607
rect 44399 2550 44459 2571
rect 44517 2550 44577 2571
rect 44635 2550 44695 2571
rect 44753 2570 45049 2606
rect 44753 2550 44813 2570
rect 44871 2550 44931 2570
rect 44989 2550 45049 2570
rect 45107 2570 45403 2606
rect 45107 2550 45167 2570
rect 45225 2550 45285 2570
rect 45343 2550 45403 2570
rect 31203 2318 31269 2335
rect 37848 2326 37908 2352
rect 37966 2326 38026 2352
rect 38084 2326 38144 2352
rect 38202 2332 38262 2352
rect 38202 2326 38263 2332
rect 38320 2326 38380 2352
rect 38438 2326 38498 2352
rect 747 2155 1043 2194
rect 747 2140 807 2155
rect 865 2140 925 2155
rect 983 2140 1043 2155
rect 1214 2155 1510 2194
rect 1214 2140 1274 2155
rect 1332 2140 1392 2155
rect 1450 2140 1510 2155
rect 1568 2155 1864 2194
rect 1568 2140 1628 2155
rect 1686 2140 1746 2155
rect 1804 2140 1864 2155
rect 2041 2155 2337 2194
rect 2041 2140 2101 2155
rect 2159 2140 2219 2155
rect 2277 2140 2337 2155
rect 3891 2155 4187 2194
rect 3891 2140 3951 2155
rect 4009 2140 4069 2155
rect 4127 2140 4187 2155
rect 4358 2155 4654 2194
rect 4358 2140 4418 2155
rect 4476 2140 4536 2155
rect 4594 2140 4654 2155
rect 4712 2155 5008 2194
rect 4712 2140 4772 2155
rect 4830 2140 4890 2155
rect 4948 2140 5008 2155
rect 5185 2155 5481 2194
rect 5185 2140 5245 2155
rect 5303 2140 5363 2155
rect 5421 2140 5481 2155
rect 7023 2159 7319 2198
rect 7023 2144 7083 2159
rect 7141 2144 7201 2159
rect 7259 2144 7319 2159
rect 7490 2159 7786 2198
rect 7490 2144 7550 2159
rect 7608 2144 7668 2159
rect 7726 2144 7786 2159
rect 7844 2159 8140 2198
rect 7844 2144 7904 2159
rect 7962 2144 8022 2159
rect 8080 2144 8140 2159
rect 8317 2159 8613 2198
rect 8317 2144 8377 2159
rect 8435 2144 8495 2159
rect 8553 2144 8613 2159
rect 10167 2159 10463 2198
rect 10167 2144 10227 2159
rect 10285 2144 10345 2159
rect 10403 2144 10463 2159
rect 10634 2159 10930 2198
rect 10634 2144 10694 2159
rect 10752 2144 10812 2159
rect 10870 2144 10930 2159
rect 10988 2159 11284 2198
rect 10988 2144 11048 2159
rect 11106 2144 11166 2159
rect 11224 2144 11284 2159
rect 11461 2159 11757 2198
rect 11461 2144 11521 2159
rect 11579 2144 11639 2159
rect 11697 2144 11757 2159
rect 13369 2155 13665 2194
rect 306 1956 602 1995
rect 306 1940 366 1956
rect 424 1940 484 1956
rect 542 1940 602 1956
rect 2514 1956 2810 1995
rect 2514 1940 2574 1956
rect 2632 1940 2692 1956
rect 2750 1940 2810 1956
rect 3450 1956 3746 1995
rect 3450 1940 3510 1956
rect 3568 1940 3628 1956
rect 3686 1940 3746 1956
rect 5658 1956 5954 1995
rect 5658 1940 5718 1956
rect 5776 1940 5836 1956
rect 5894 1940 5954 1956
rect 6582 1960 6878 1999
rect 6582 1944 6642 1960
rect 6700 1944 6760 1960
rect 6818 1944 6878 1960
rect 8790 1960 9086 1999
rect 8790 1944 8850 1960
rect 8908 1944 8968 1960
rect 9026 1944 9086 1960
rect 9726 1960 10022 1999
rect 9726 1944 9786 1960
rect 9844 1944 9904 1960
rect 9962 1944 10022 1960
rect 13369 2140 13429 2155
rect 13487 2140 13547 2155
rect 13605 2140 13665 2155
rect 13836 2155 14132 2194
rect 13836 2140 13896 2155
rect 13954 2140 14014 2155
rect 14072 2140 14132 2155
rect 14190 2155 14486 2194
rect 14190 2140 14250 2155
rect 14308 2140 14368 2155
rect 14426 2140 14486 2155
rect 14663 2155 14959 2194
rect 14663 2140 14723 2155
rect 14781 2140 14841 2155
rect 14899 2140 14959 2155
rect 16513 2155 16809 2194
rect 16513 2140 16573 2155
rect 16631 2140 16691 2155
rect 16749 2140 16809 2155
rect 16980 2155 17276 2194
rect 16980 2140 17040 2155
rect 17098 2140 17158 2155
rect 17216 2140 17276 2155
rect 17334 2155 17630 2194
rect 17334 2140 17394 2155
rect 17452 2140 17512 2155
rect 17570 2140 17630 2155
rect 17807 2155 18103 2194
rect 17807 2140 17867 2155
rect 17925 2140 17985 2155
rect 18043 2140 18103 2155
rect 19645 2159 19941 2198
rect 19645 2144 19705 2159
rect 19763 2144 19823 2159
rect 19881 2144 19941 2159
rect 20112 2159 20408 2198
rect 20112 2144 20172 2159
rect 20230 2144 20290 2159
rect 20348 2144 20408 2159
rect 20466 2159 20762 2198
rect 20466 2144 20526 2159
rect 20584 2144 20644 2159
rect 20702 2144 20762 2159
rect 20939 2159 21235 2198
rect 20939 2144 20999 2159
rect 21057 2144 21117 2159
rect 21175 2144 21235 2159
rect 22789 2159 23085 2198
rect 22789 2144 22849 2159
rect 22907 2144 22967 2159
rect 23025 2144 23085 2159
rect 23256 2159 23552 2198
rect 23256 2144 23316 2159
rect 23374 2144 23434 2159
rect 23492 2144 23552 2159
rect 23610 2159 23906 2198
rect 23610 2144 23670 2159
rect 23728 2144 23788 2159
rect 23846 2144 23906 2159
rect 24083 2159 24379 2198
rect 29884 2178 29935 2236
rect 30560 2235 30620 2293
rect 31210 2235 31269 2318
rect 24083 2144 24143 2159
rect 24201 2144 24261 2159
rect 24319 2144 24379 2159
rect 11934 1960 12230 1999
rect 11934 1944 11994 1960
rect 12052 1944 12112 1960
rect 12170 1944 12230 1960
rect 12928 1956 13224 1995
rect 12928 1940 12988 1956
rect 13046 1940 13106 1956
rect 13164 1940 13224 1956
rect 306 1454 366 1740
rect 424 1714 484 1740
rect 542 1714 602 1740
rect 747 1714 807 1740
rect 306 1437 442 1454
rect 306 1382 365 1437
rect 423 1382 442 1437
rect 306 1367 442 1382
rect 306 1055 366 1367
rect 865 1322 925 1740
rect 983 1714 1043 1740
rect 1214 1714 1274 1740
rect 1332 1714 1392 1740
rect 1450 1714 1510 1740
rect 1568 1714 1628 1740
rect 1333 1554 1392 1714
rect 1333 1553 1396 1554
rect 1330 1537 1396 1553
rect 1330 1503 1346 1537
rect 1380 1503 1396 1537
rect 1330 1487 1396 1503
rect 1433 1438 1528 1453
rect 1433 1383 1452 1438
rect 1510 1415 1528 1438
rect 1686 1415 1746 1740
rect 1804 1714 1864 1740
rect 2041 1714 2101 1740
rect 1510 1383 1746 1415
rect 1433 1366 1746 1383
rect 865 1265 1392 1322
rect 1332 1166 1392 1265
rect 1321 1153 1402 1166
rect 1321 1098 1334 1153
rect 1392 1098 1402 1153
rect 1321 1087 1402 1098
rect 306 1010 1200 1055
rect 1140 807 1200 1010
rect 1332 807 1392 1087
rect 1450 807 1510 1366
rect 2159 1324 2219 1740
rect 2277 1714 2337 1740
rect 2514 1714 2574 1740
rect 2632 1714 2692 1740
rect 2640 1591 2706 1594
rect 2750 1591 2810 1740
rect 2640 1578 2810 1591
rect 2640 1544 2656 1578
rect 2690 1544 2810 1578
rect 2640 1531 2810 1544
rect 2640 1528 2706 1531
rect 1681 1307 2219 1324
rect 1681 1273 1700 1307
rect 1734 1273 2219 1307
rect 1681 1267 2219 1273
rect 1681 1257 1750 1267
rect 1681 1255 1746 1257
rect 1565 917 1631 933
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1568 807 1628 867
rect 1686 807 1746 1255
rect 2750 1055 2810 1531
rect 1882 1010 2810 1055
rect 3450 1454 3510 1740
rect 3568 1714 3628 1740
rect 3686 1714 3746 1740
rect 3891 1714 3951 1740
rect 3450 1437 3586 1454
rect 3450 1382 3509 1437
rect 3567 1382 3586 1437
rect 3450 1367 3586 1382
rect 3450 1055 3510 1367
rect 4009 1322 4069 1740
rect 4127 1714 4187 1740
rect 4358 1714 4418 1740
rect 4476 1714 4536 1740
rect 4594 1714 4654 1740
rect 4712 1714 4772 1740
rect 4477 1554 4536 1714
rect 4477 1553 4540 1554
rect 4474 1537 4540 1553
rect 4474 1503 4490 1537
rect 4524 1503 4540 1537
rect 4474 1487 4540 1503
rect 4577 1438 4672 1453
rect 4577 1383 4596 1438
rect 4654 1415 4672 1438
rect 4830 1415 4890 1740
rect 4948 1714 5008 1740
rect 5185 1714 5245 1740
rect 4654 1383 4890 1415
rect 4577 1366 4890 1383
rect 4009 1265 4536 1322
rect 4476 1166 4536 1265
rect 4465 1153 4546 1166
rect 4465 1098 4478 1153
rect 4536 1098 4546 1153
rect 4465 1087 4546 1098
rect 3450 1010 4344 1055
rect 1882 807 1942 1010
rect 4284 807 4344 1010
rect 4476 807 4536 1087
rect 4594 807 4654 1366
rect 5303 1324 5363 1740
rect 5421 1714 5481 1740
rect 5658 1714 5718 1740
rect 5776 1714 5836 1740
rect 5784 1591 5850 1594
rect 5894 1591 5954 1740
rect 5784 1578 5954 1591
rect 5784 1544 5800 1578
rect 5834 1544 5954 1578
rect 5784 1531 5954 1544
rect 5784 1528 5850 1531
rect 4825 1307 5363 1324
rect 4825 1273 4844 1307
rect 4878 1273 5363 1307
rect 4825 1267 5363 1273
rect 4825 1257 4894 1267
rect 4825 1255 4890 1257
rect 4709 917 4775 933
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 4712 807 4772 867
rect 4830 807 4890 1255
rect 5894 1055 5954 1531
rect 5026 1010 5954 1055
rect 6582 1458 6642 1744
rect 6700 1718 6760 1744
rect 6818 1718 6878 1744
rect 7023 1718 7083 1744
rect 6582 1441 6718 1458
rect 6582 1386 6641 1441
rect 6699 1386 6718 1441
rect 6582 1371 6718 1386
rect 6582 1059 6642 1371
rect 7141 1326 7201 1744
rect 7259 1718 7319 1744
rect 7490 1718 7550 1744
rect 7608 1718 7668 1744
rect 7726 1718 7786 1744
rect 7844 1718 7904 1744
rect 7609 1558 7668 1718
rect 7609 1557 7672 1558
rect 7606 1541 7672 1557
rect 7606 1507 7622 1541
rect 7656 1507 7672 1541
rect 7606 1491 7672 1507
rect 7709 1442 7804 1457
rect 7709 1387 7728 1442
rect 7786 1419 7804 1442
rect 7962 1419 8022 1744
rect 8080 1718 8140 1744
rect 8317 1718 8377 1744
rect 7786 1387 8022 1419
rect 7709 1370 8022 1387
rect 7141 1269 7668 1326
rect 7608 1170 7668 1269
rect 7597 1157 7678 1170
rect 7597 1102 7610 1157
rect 7668 1102 7678 1157
rect 7597 1091 7678 1102
rect 6582 1014 7476 1059
rect 5026 807 5086 1010
rect 7416 811 7476 1014
rect 7608 811 7668 1091
rect 7726 811 7786 1370
rect 8435 1328 8495 1744
rect 8553 1718 8613 1744
rect 8790 1718 8850 1744
rect 8908 1718 8968 1744
rect 8916 1595 8982 1598
rect 9026 1595 9086 1744
rect 8916 1582 9086 1595
rect 8916 1548 8932 1582
rect 8966 1548 9086 1582
rect 8916 1535 9086 1548
rect 8916 1532 8982 1535
rect 7957 1311 8495 1328
rect 7957 1277 7976 1311
rect 8010 1277 8495 1311
rect 7957 1271 8495 1277
rect 7957 1261 8026 1271
rect 7957 1259 8022 1261
rect 7841 921 7907 937
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 7844 811 7904 871
rect 7962 811 8022 1259
rect 9026 1059 9086 1535
rect 8158 1014 9086 1059
rect 9726 1458 9786 1744
rect 9844 1718 9904 1744
rect 9962 1718 10022 1744
rect 10167 1718 10227 1744
rect 9726 1441 9862 1458
rect 9726 1386 9785 1441
rect 9843 1386 9862 1441
rect 9726 1371 9862 1386
rect 9726 1059 9786 1371
rect 10285 1326 10345 1744
rect 10403 1718 10463 1744
rect 10634 1718 10694 1744
rect 10752 1718 10812 1744
rect 10870 1718 10930 1744
rect 10988 1718 11048 1744
rect 10753 1558 10812 1718
rect 10753 1557 10816 1558
rect 10750 1541 10816 1557
rect 10750 1507 10766 1541
rect 10800 1507 10816 1541
rect 10750 1491 10816 1507
rect 10853 1442 10948 1457
rect 10853 1387 10872 1442
rect 10930 1419 10948 1442
rect 11106 1419 11166 1744
rect 11224 1718 11284 1744
rect 11461 1718 11521 1744
rect 10930 1387 11166 1419
rect 10853 1370 11166 1387
rect 10285 1269 10812 1326
rect 10752 1170 10812 1269
rect 10741 1157 10822 1170
rect 10741 1102 10754 1157
rect 10812 1102 10822 1157
rect 10741 1091 10822 1102
rect 9726 1014 10620 1059
rect 8158 811 8218 1014
rect 10560 811 10620 1014
rect 10752 811 10812 1091
rect 10870 811 10930 1370
rect 11579 1328 11639 1744
rect 11697 1718 11757 1744
rect 11934 1718 11994 1744
rect 12052 1718 12112 1744
rect 12060 1595 12126 1598
rect 12170 1595 12230 1744
rect 15136 1956 15432 1995
rect 15136 1940 15196 1956
rect 15254 1940 15314 1956
rect 15372 1940 15432 1956
rect 16072 1956 16368 1995
rect 16072 1940 16132 1956
rect 16190 1940 16250 1956
rect 16308 1940 16368 1956
rect 18280 1956 18576 1995
rect 18280 1940 18340 1956
rect 18398 1940 18458 1956
rect 18516 1940 18576 1956
rect 19204 1960 19500 1999
rect 19204 1944 19264 1960
rect 19322 1944 19382 1960
rect 19440 1944 19500 1960
rect 21412 1960 21708 1999
rect 21412 1944 21472 1960
rect 21530 1944 21590 1960
rect 21648 1944 21708 1960
rect 22348 1960 22644 1999
rect 22348 1944 22408 1960
rect 22466 1944 22526 1960
rect 22584 1944 22644 1960
rect 24556 1960 24852 1999
rect 24556 1944 24616 1960
rect 24674 1944 24734 1960
rect 24792 1944 24852 1960
rect 29884 2118 29950 2178
rect 30350 2118 30376 2178
rect 30560 2175 30643 2235
rect 31043 2175 31375 2235
rect 31775 2175 31801 2235
rect 29884 2060 29935 2118
rect 30560 2117 30620 2175
rect 31287 2117 31353 2119
rect 29884 2000 29950 2060
rect 30350 2000 30376 2060
rect 30560 2057 30643 2117
rect 31043 2057 31069 2117
rect 31287 2103 31375 2117
rect 31287 2069 31303 2103
rect 31337 2069 31375 2103
rect 31287 2057 31375 2069
rect 31775 2057 31801 2117
rect 38085 2141 38143 2326
rect 38085 2115 38145 2141
rect 38203 2115 38263 2326
rect 38556 2320 38616 2352
rect 38674 2326 38734 2352
rect 38792 2326 38852 2352
rect 51054 2572 51350 2608
rect 51054 2551 51114 2572
rect 51172 2551 51232 2572
rect 51290 2551 51350 2572
rect 51408 2571 51704 2607
rect 51408 2551 51468 2571
rect 51526 2551 51586 2571
rect 51644 2551 51704 2571
rect 51762 2571 52058 2607
rect 51762 2551 51822 2571
rect 51880 2551 51940 2571
rect 51998 2551 52058 2571
rect 57676 2573 57972 2609
rect 57676 2552 57736 2573
rect 57794 2552 57854 2573
rect 57912 2552 57972 2573
rect 58030 2572 58326 2608
rect 58030 2552 58090 2572
rect 58148 2552 58208 2572
rect 58266 2552 58326 2572
rect 58384 2572 58680 2608
rect 58384 2552 58444 2572
rect 58502 2552 58562 2572
rect 58620 2552 58680 2572
rect 65407 2560 65467 2586
rect 70455 2616 70509 2676
rect 70909 2616 70935 2676
rect 66705 2560 66765 2586
rect 70455 2558 70494 2616
rect 70455 2498 70509 2558
rect 70909 2498 71384 2558
rect 70455 2440 70494 2498
rect 65827 2360 65887 2386
rect 65945 2360 66005 2386
rect 66063 2360 66123 2386
rect 66181 2360 66241 2386
rect 70455 2380 70509 2440
rect 70909 2380 70935 2440
rect 44399 2324 44459 2350
rect 44517 2324 44577 2350
rect 44635 2324 44695 2350
rect 44753 2330 44813 2350
rect 44753 2324 44814 2330
rect 44871 2324 44931 2350
rect 44989 2324 45049 2350
rect 38553 2304 38619 2320
rect 38553 2270 38569 2304
rect 38603 2270 38619 2304
rect 38553 2254 38619 2270
rect 38435 2187 38501 2203
rect 38435 2153 38451 2187
rect 38485 2153 38501 2187
rect 38435 2137 38501 2153
rect 39796 2150 40092 2201
rect 38438 2115 38498 2137
rect 39796 2135 39856 2150
rect 39914 2135 39974 2150
rect 40032 2135 40092 2150
rect 40150 2135 40210 2161
rect 40268 2135 40328 2161
rect 40386 2135 40446 2161
rect 41694 2150 41990 2201
rect 41694 2135 41754 2150
rect 41812 2135 41872 2150
rect 41930 2135 41990 2150
rect 42048 2135 42108 2161
rect 42166 2135 42226 2161
rect 42284 2135 42344 2161
rect 44636 2139 44694 2324
rect 31287 2053 31353 2057
rect 31287 1999 31352 2001
rect 29924 1882 29950 1942
rect 30350 1882 30420 1942
rect 30369 1824 30420 1882
rect 29924 1764 29950 1824
rect 30350 1764 30420 1824
rect 12060 1582 12230 1595
rect 12060 1548 12076 1582
rect 12110 1548 12230 1582
rect 12060 1535 12230 1548
rect 12060 1532 12126 1535
rect 11101 1311 11639 1328
rect 11101 1277 11120 1311
rect 11154 1277 11639 1311
rect 11101 1271 11639 1277
rect 11101 1261 11170 1271
rect 11101 1259 11166 1261
rect 10985 921 11051 937
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 10988 811 11048 871
rect 11106 811 11166 1259
rect 12170 1059 12230 1535
rect 11302 1014 12230 1059
rect 12928 1454 12988 1740
rect 13046 1714 13106 1740
rect 13164 1714 13224 1740
rect 13369 1714 13429 1740
rect 12928 1437 13064 1454
rect 12928 1382 12987 1437
rect 13045 1382 13064 1437
rect 12928 1367 13064 1382
rect 12928 1055 12988 1367
rect 13487 1322 13547 1740
rect 13605 1714 13665 1740
rect 13836 1714 13896 1740
rect 13954 1714 14014 1740
rect 14072 1714 14132 1740
rect 14190 1714 14250 1740
rect 13955 1554 14014 1714
rect 13955 1553 14018 1554
rect 13952 1537 14018 1553
rect 13952 1503 13968 1537
rect 14002 1503 14018 1537
rect 13952 1487 14018 1503
rect 14055 1438 14150 1453
rect 14055 1383 14074 1438
rect 14132 1415 14150 1438
rect 14308 1415 14368 1740
rect 14426 1714 14486 1740
rect 14663 1714 14723 1740
rect 14132 1383 14368 1415
rect 14055 1366 14368 1383
rect 13487 1265 14014 1322
rect 13954 1166 14014 1265
rect 13943 1153 14024 1166
rect 13943 1098 13956 1153
rect 14014 1098 14024 1153
rect 13943 1087 14024 1098
rect 11302 811 11362 1014
rect 12928 1010 13822 1055
rect 1140 581 1200 607
rect 1332 381 1392 407
rect 1450 381 1510 407
rect 1568 381 1628 407
rect 1686 381 1746 407
rect 1507 326 1573 334
rect 1882 326 1942 607
rect 4284 581 4344 607
rect 4476 381 4536 407
rect 4594 381 4654 407
rect 4712 381 4772 407
rect 4830 381 4890 407
rect 1507 318 1942 326
rect 1507 284 1523 318
rect 1557 284 1942 318
rect 1507 275 1942 284
rect 4651 326 4717 334
rect 5026 326 5086 607
rect 7416 585 7476 611
rect 7608 385 7668 411
rect 7726 385 7786 411
rect 7844 385 7904 411
rect 7962 385 8022 411
rect 4651 318 5086 326
rect 4651 284 4667 318
rect 4701 284 5086 318
rect 4651 275 5086 284
rect 7783 330 7849 338
rect 8158 330 8218 611
rect 10560 585 10620 611
rect 13762 807 13822 1010
rect 13954 807 14014 1087
rect 14072 807 14132 1366
rect 14781 1324 14841 1740
rect 14899 1714 14959 1740
rect 15136 1714 15196 1740
rect 15254 1714 15314 1740
rect 15262 1591 15328 1594
rect 15372 1591 15432 1740
rect 15262 1578 15432 1591
rect 15262 1544 15278 1578
rect 15312 1544 15432 1578
rect 15262 1531 15432 1544
rect 15262 1528 15328 1531
rect 14303 1307 14841 1324
rect 14303 1273 14322 1307
rect 14356 1273 14841 1307
rect 14303 1267 14841 1273
rect 14303 1257 14372 1267
rect 14303 1255 14368 1257
rect 14187 917 14253 933
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14190 807 14250 867
rect 14308 807 14368 1255
rect 15372 1055 15432 1531
rect 14504 1010 15432 1055
rect 16072 1454 16132 1740
rect 16190 1714 16250 1740
rect 16308 1714 16368 1740
rect 16513 1714 16573 1740
rect 16072 1437 16208 1454
rect 16072 1382 16131 1437
rect 16189 1382 16208 1437
rect 16072 1367 16208 1382
rect 16072 1055 16132 1367
rect 16631 1322 16691 1740
rect 16749 1714 16809 1740
rect 16980 1714 17040 1740
rect 17098 1714 17158 1740
rect 17216 1714 17276 1740
rect 17334 1714 17394 1740
rect 17099 1554 17158 1714
rect 17099 1553 17162 1554
rect 17096 1537 17162 1553
rect 17096 1503 17112 1537
rect 17146 1503 17162 1537
rect 17096 1487 17162 1503
rect 17199 1438 17294 1453
rect 17199 1383 17218 1438
rect 17276 1415 17294 1438
rect 17452 1415 17512 1740
rect 17570 1714 17630 1740
rect 17807 1714 17867 1740
rect 17276 1383 17512 1415
rect 17199 1366 17512 1383
rect 16631 1265 17158 1322
rect 17098 1166 17158 1265
rect 17087 1153 17168 1166
rect 17087 1098 17100 1153
rect 17158 1098 17168 1153
rect 17087 1087 17168 1098
rect 16072 1010 16966 1055
rect 14504 807 14564 1010
rect 16906 807 16966 1010
rect 17098 807 17158 1087
rect 17216 807 17276 1366
rect 17925 1324 17985 1740
rect 18043 1714 18103 1740
rect 18280 1714 18340 1740
rect 18398 1714 18458 1740
rect 18406 1591 18472 1594
rect 18516 1591 18576 1740
rect 18406 1578 18576 1591
rect 18406 1544 18422 1578
rect 18456 1544 18576 1578
rect 18406 1531 18576 1544
rect 18406 1528 18472 1531
rect 17447 1307 17985 1324
rect 17447 1273 17466 1307
rect 17500 1273 17985 1307
rect 17447 1267 17985 1273
rect 17447 1257 17516 1267
rect 17447 1255 17512 1257
rect 17331 917 17397 933
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17334 807 17394 867
rect 17452 807 17512 1255
rect 18516 1055 18576 1531
rect 17648 1010 18576 1055
rect 19204 1458 19264 1744
rect 19322 1718 19382 1744
rect 19440 1718 19500 1744
rect 19645 1718 19705 1744
rect 19204 1441 19340 1458
rect 19204 1386 19263 1441
rect 19321 1386 19340 1441
rect 19204 1371 19340 1386
rect 19204 1059 19264 1371
rect 19763 1326 19823 1744
rect 19881 1718 19941 1744
rect 20112 1718 20172 1744
rect 20230 1718 20290 1744
rect 20348 1718 20408 1744
rect 20466 1718 20526 1744
rect 20231 1558 20290 1718
rect 20231 1557 20294 1558
rect 20228 1541 20294 1557
rect 20228 1507 20244 1541
rect 20278 1507 20294 1541
rect 20228 1491 20294 1507
rect 20331 1442 20426 1457
rect 20331 1387 20350 1442
rect 20408 1419 20426 1442
rect 20584 1419 20644 1744
rect 20702 1718 20762 1744
rect 20939 1718 20999 1744
rect 20408 1387 20644 1419
rect 20331 1370 20644 1387
rect 19763 1269 20290 1326
rect 20230 1170 20290 1269
rect 20219 1157 20300 1170
rect 20219 1102 20232 1157
rect 20290 1102 20300 1157
rect 20219 1091 20300 1102
rect 19204 1014 20098 1059
rect 17648 807 17708 1010
rect 20038 811 20098 1014
rect 20230 811 20290 1091
rect 20348 811 20408 1370
rect 21057 1328 21117 1744
rect 21175 1718 21235 1744
rect 21412 1718 21472 1744
rect 21530 1718 21590 1744
rect 21538 1595 21604 1598
rect 21648 1595 21708 1744
rect 21538 1582 21708 1595
rect 21538 1548 21554 1582
rect 21588 1548 21708 1582
rect 21538 1535 21708 1548
rect 21538 1532 21604 1535
rect 20579 1311 21117 1328
rect 20579 1277 20598 1311
rect 20632 1277 21117 1311
rect 20579 1271 21117 1277
rect 20579 1261 20648 1271
rect 20579 1259 20644 1261
rect 20463 921 20529 937
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20466 811 20526 871
rect 20584 811 20644 1259
rect 21648 1059 21708 1535
rect 20780 1014 21708 1059
rect 22348 1458 22408 1744
rect 22466 1718 22526 1744
rect 22584 1718 22644 1744
rect 22789 1718 22849 1744
rect 22348 1441 22484 1458
rect 22348 1386 22407 1441
rect 22465 1386 22484 1441
rect 22348 1371 22484 1386
rect 22348 1059 22408 1371
rect 22907 1326 22967 1744
rect 23025 1718 23085 1744
rect 23256 1718 23316 1744
rect 23374 1718 23434 1744
rect 23492 1718 23552 1744
rect 23610 1718 23670 1744
rect 23375 1558 23434 1718
rect 23375 1557 23438 1558
rect 23372 1541 23438 1557
rect 23372 1507 23388 1541
rect 23422 1507 23438 1541
rect 23372 1491 23438 1507
rect 23475 1442 23570 1457
rect 23475 1387 23494 1442
rect 23552 1419 23570 1442
rect 23728 1419 23788 1744
rect 23846 1718 23906 1744
rect 24083 1718 24143 1744
rect 23552 1387 23788 1419
rect 23475 1370 23788 1387
rect 22907 1269 23434 1326
rect 23374 1170 23434 1269
rect 23363 1157 23444 1170
rect 23363 1102 23376 1157
rect 23434 1102 23444 1157
rect 23363 1091 23444 1102
rect 22348 1014 23242 1059
rect 20780 811 20840 1014
rect 23182 811 23242 1014
rect 23374 811 23434 1091
rect 23492 811 23552 1370
rect 24201 1328 24261 1744
rect 24319 1718 24379 1744
rect 24556 1718 24616 1744
rect 24674 1718 24734 1744
rect 24682 1595 24748 1598
rect 24792 1595 24852 1744
rect 30369 1706 30420 1764
rect 29924 1646 29950 1706
rect 30350 1646 30420 1706
rect 30559 1939 30643 1999
rect 31043 1939 31069 1999
rect 31287 1985 31375 1999
rect 31287 1951 31302 1985
rect 31336 1951 31375 1985
rect 31287 1939 31375 1951
rect 31775 1939 31801 1999
rect 30559 1881 30619 1939
rect 31287 1935 31352 1939
rect 30559 1821 30643 1881
rect 31043 1821 31375 1881
rect 31775 1821 31801 1881
rect 30559 1763 30619 1821
rect 30559 1703 30643 1763
rect 31043 1703 31069 1763
rect 31210 1738 31269 1821
rect 31203 1721 31269 1738
rect 24682 1582 24852 1595
rect 24682 1548 24698 1582
rect 24732 1548 24852 1582
rect 24682 1535 24852 1548
rect 24682 1532 24748 1535
rect 23723 1311 24261 1328
rect 23723 1277 23742 1311
rect 23776 1277 24261 1311
rect 23723 1271 24261 1277
rect 23723 1261 23792 1271
rect 23723 1259 23788 1261
rect 23607 921 23673 937
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23610 811 23670 871
rect 23728 811 23788 1259
rect 24792 1059 24852 1535
rect 30369 1459 30420 1646
rect 31203 1687 31219 1721
rect 31253 1687 31269 1721
rect 39312 1935 39372 1961
rect 39430 1935 39490 1961
rect 39548 1935 39608 1961
rect 38438 1889 38498 1915
rect 38085 1693 38145 1715
rect 38203 1699 38263 1715
rect 31203 1671 31269 1687
rect 34941 1647 35237 1683
rect 34941 1626 35001 1647
rect 35059 1626 35119 1647
rect 35177 1626 35237 1647
rect 35295 1646 35591 1682
rect 35295 1626 35355 1646
rect 35413 1626 35473 1646
rect 35531 1626 35591 1646
rect 35649 1646 35945 1682
rect 35649 1626 35709 1646
rect 35767 1626 35827 1646
rect 35885 1626 35945 1646
rect 38082 1677 38148 1693
rect 38082 1643 38098 1677
rect 38132 1643 38148 1677
rect 38082 1627 38148 1643
rect 38197 1677 38271 1699
rect 38197 1643 38216 1677
rect 38250 1643 38271 1677
rect 40633 1952 40929 2003
rect 40633 1935 40693 1952
rect 40751 1935 40811 1952
rect 40869 1935 40929 1952
rect 41210 1935 41270 1961
rect 41328 1935 41388 1961
rect 41446 1935 41506 1961
rect 44636 2113 44696 2139
rect 44754 2113 44814 2324
rect 45107 2318 45167 2350
rect 45225 2324 45285 2350
rect 45343 2324 45403 2350
rect 51054 2325 51114 2351
rect 51172 2325 51232 2351
rect 51290 2325 51350 2351
rect 51408 2331 51468 2351
rect 51408 2325 51469 2331
rect 51526 2325 51586 2351
rect 51644 2325 51704 2351
rect 45104 2302 45170 2318
rect 45104 2268 45120 2302
rect 45154 2268 45170 2302
rect 45104 2252 45170 2268
rect 44986 2185 45052 2201
rect 44986 2151 45002 2185
rect 45036 2151 45052 2185
rect 44986 2135 45052 2151
rect 46347 2148 46643 2199
rect 44989 2113 45049 2135
rect 46347 2133 46407 2148
rect 46465 2133 46525 2148
rect 46583 2133 46643 2148
rect 46701 2133 46761 2159
rect 46819 2133 46879 2159
rect 46937 2133 46997 2159
rect 48245 2148 48541 2199
rect 48245 2133 48305 2148
rect 48363 2133 48423 2148
rect 48481 2133 48541 2148
rect 48599 2133 48659 2159
rect 48717 2133 48777 2159
rect 48835 2133 48895 2159
rect 51291 2140 51349 2325
rect 42531 1952 42827 2003
rect 42531 1935 42591 1952
rect 42649 1935 42709 1952
rect 42767 1935 42827 1952
rect 39312 1718 39372 1735
rect 39430 1718 39490 1735
rect 39548 1718 39608 1735
rect 39796 1718 39856 1735
rect 39312 1667 39856 1718
rect 39914 1709 39974 1735
rect 40032 1709 40092 1735
rect 40150 1716 40210 1735
rect 40268 1716 40328 1735
rect 40386 1716 40446 1735
rect 40633 1716 40693 1735
rect 40751 1716 40811 1735
rect 30082 1399 30150 1459
rect 30350 1399 30420 1459
rect 31271 1431 31337 1447
rect 30507 1409 30561 1425
rect 30082 1341 30133 1399
rect 30507 1375 30517 1409
rect 30551 1375 30561 1409
rect 30507 1357 30561 1375
rect 31271 1397 31287 1431
rect 31321 1397 31337 1431
rect 38197 1586 38271 1643
rect 39437 1586 39497 1667
rect 40150 1665 40693 1716
rect 40735 1709 40811 1716
rect 40869 1709 40929 1735
rect 41210 1718 41270 1735
rect 41328 1718 41388 1735
rect 41446 1718 41506 1735
rect 41694 1718 41754 1735
rect 40735 1665 40810 1709
rect 41210 1667 41754 1718
rect 41812 1709 41872 1735
rect 41930 1709 41990 1735
rect 42048 1716 42108 1735
rect 42166 1716 42226 1735
rect 42284 1716 42344 1735
rect 42531 1716 42591 1735
rect 42649 1716 42709 1735
rect 38197 1561 39497 1586
rect 38196 1513 39497 1561
rect 40735 1545 40795 1665
rect 31271 1357 31337 1397
rect 34941 1400 35001 1426
rect 35059 1400 35119 1426
rect 35177 1400 35237 1426
rect 35295 1406 35355 1426
rect 35295 1400 35356 1406
rect 35413 1400 35473 1426
rect 35531 1400 35591 1426
rect 30369 1341 31375 1357
rect 30082 1281 30150 1341
rect 30350 1297 31375 1341
rect 31575 1297 31601 1357
rect 30350 1282 30420 1297
rect 30350 1281 30376 1282
rect 30082 1223 30133 1281
rect 30082 1163 30150 1223
rect 30350 1163 30376 1223
rect 35178 1215 35236 1400
rect 35178 1189 35238 1215
rect 35296 1189 35356 1400
rect 35649 1394 35709 1426
rect 35767 1400 35827 1426
rect 35885 1400 35945 1426
rect 35646 1378 35712 1394
rect 35646 1344 35662 1378
rect 35696 1344 35712 1378
rect 35646 1328 35712 1344
rect 35528 1261 35594 1277
rect 35528 1227 35544 1261
rect 35578 1227 35594 1261
rect 35528 1211 35594 1227
rect 35531 1189 35591 1211
rect 23924 1014 24852 1059
rect 23924 811 23984 1014
rect 10752 385 10812 411
rect 10870 385 10930 411
rect 10988 385 11048 411
rect 11106 385 11166 411
rect 7783 322 8218 330
rect 7783 288 7799 322
rect 7833 288 8218 322
rect 7783 279 8218 288
rect 10927 330 10993 338
rect 11302 330 11362 611
rect 13762 581 13822 607
rect 13954 381 14014 407
rect 14072 381 14132 407
rect 14190 381 14250 407
rect 14308 381 14368 407
rect 10927 322 11362 330
rect 10927 288 10943 322
rect 10977 288 11362 322
rect 10927 279 11362 288
rect 14129 326 14195 334
rect 14504 326 14564 607
rect 16906 581 16966 607
rect 17098 381 17158 407
rect 17216 381 17276 407
rect 17334 381 17394 407
rect 17452 381 17512 407
rect 14129 318 14564 326
rect 14129 284 14145 318
rect 14179 284 14564 318
rect 1507 268 1573 275
rect 4651 268 4717 275
rect 7783 272 7849 279
rect 10927 272 10993 279
rect 14129 275 14564 284
rect 17273 326 17339 334
rect 17648 326 17708 607
rect 20038 585 20098 611
rect 20230 385 20290 411
rect 20348 385 20408 411
rect 20466 385 20526 411
rect 20584 385 20644 411
rect 17273 318 17708 326
rect 17273 284 17289 318
rect 17323 284 17708 318
rect 17273 275 17708 284
rect 20405 330 20471 338
rect 20780 330 20840 611
rect 23182 585 23242 611
rect 35531 963 35591 989
rect 37843 969 38139 1005
rect 37843 948 37903 969
rect 37961 948 38021 969
rect 38079 948 38139 969
rect 38197 968 38493 1004
rect 38197 948 38257 968
rect 38315 948 38375 968
rect 38433 948 38493 968
rect 38551 968 38847 1004
rect 38551 948 38611 968
rect 38669 948 38729 968
rect 38787 948 38847 968
rect 35178 767 35238 789
rect 35296 767 35356 789
rect 35175 751 35241 767
rect 30699 734 30759 750
rect 30126 651 30152 711
rect 30352 651 30420 711
rect 23374 385 23434 411
rect 23492 385 23552 411
rect 23610 385 23670 411
rect 23728 385 23788 411
rect 20405 322 20840 330
rect 20405 288 20421 322
rect 20455 288 20840 322
rect 20405 279 20840 288
rect 23549 330 23615 338
rect 23924 330 23984 611
rect 30369 593 30420 651
rect 30126 533 30152 593
rect 30352 586 30420 593
rect 30699 700 30713 734
rect 30747 700 30759 734
rect 35175 717 35191 751
rect 35225 717 35241 751
rect 35175 701 35241 717
rect 35293 751 35359 767
rect 35293 717 35309 751
rect 35343 717 35359 751
rect 39437 815 39497 1513
rect 39739 1465 40035 1525
rect 39739 1442 39799 1465
rect 39857 1442 39917 1465
rect 39975 1442 40035 1465
rect 40093 1466 40389 1526
rect 40734 1525 40795 1545
rect 40093 1442 40153 1466
rect 40211 1442 40271 1466
rect 40329 1442 40389 1466
rect 40715 1509 40795 1525
rect 40715 1475 40730 1509
rect 40764 1475 40795 1509
rect 40715 1459 40795 1475
rect 40734 1436 40795 1459
rect 40735 1290 40795 1436
rect 40734 1117 40795 1290
rect 39739 1016 39799 1042
rect 39707 875 39774 882
rect 39857 875 39917 1042
rect 39975 1016 40035 1042
rect 40093 1016 40153 1042
rect 39707 866 39917 875
rect 39707 832 39723 866
rect 39757 832 39917 866
rect 39707 816 39917 832
rect 39437 799 39588 815
rect 39437 765 39538 799
rect 39572 765 39588 799
rect 39437 749 39588 765
rect 37843 722 37903 748
rect 37961 722 38021 748
rect 38079 722 38139 748
rect 38197 728 38257 748
rect 38197 722 38258 728
rect 38315 722 38375 748
rect 38433 722 38493 748
rect 35293 701 35359 717
rect 30699 586 30759 700
rect 30352 533 31377 586
rect 30369 526 31377 533
rect 31577 526 31603 586
rect 38080 537 38138 722
rect 30369 475 30420 526
rect 30126 415 30152 475
rect 30352 415 30420 475
rect 31272 485 31338 526
rect 31272 451 31288 485
rect 31322 451 31338 485
rect 38080 511 38140 537
rect 38198 511 38258 722
rect 38551 716 38611 748
rect 38669 722 38729 748
rect 38787 722 38847 748
rect 38548 700 38614 716
rect 39437 710 39497 749
rect 39857 710 39917 816
rect 40211 875 40271 1042
rect 40329 1016 40389 1042
rect 40354 875 40421 882
rect 40211 866 40421 875
rect 40211 832 40371 866
rect 40405 832 40421 866
rect 40211 816 40421 832
rect 39973 782 40039 798
rect 39973 748 39989 782
rect 40023 748 40039 782
rect 39973 732 40039 748
rect 40091 783 40157 798
rect 40091 749 40107 783
rect 40141 749 40157 783
rect 40091 733 40157 749
rect 39975 710 40035 732
rect 40093 710 40153 733
rect 40211 710 40271 816
rect 40735 814 40795 1117
rect 40645 798 40795 814
rect 40645 764 40661 798
rect 40695 764 40795 798
rect 40645 748 40795 764
rect 40735 710 40795 748
rect 41335 1009 41395 1667
rect 42048 1665 42591 1716
rect 42633 1709 42709 1716
rect 42767 1709 42827 1735
rect 45863 1933 45923 1959
rect 45981 1933 46041 1959
rect 46099 1933 46159 1959
rect 44989 1887 45049 1913
rect 42633 1665 42708 1709
rect 44636 1691 44696 1713
rect 44754 1697 44814 1713
rect 44633 1675 44699 1691
rect 41637 1465 41933 1525
rect 41637 1442 41697 1465
rect 41755 1442 41815 1465
rect 41873 1442 41933 1465
rect 41991 1466 42287 1526
rect 41991 1442 42051 1466
rect 42109 1442 42169 1466
rect 42227 1442 42287 1466
rect 42633 1512 42693 1665
rect 44633 1641 44649 1675
rect 44683 1641 44699 1675
rect 44633 1625 44699 1641
rect 44748 1675 44822 1697
rect 44748 1641 44767 1675
rect 44801 1641 44822 1675
rect 47184 1950 47480 2001
rect 47184 1933 47244 1950
rect 47302 1933 47362 1950
rect 47420 1933 47480 1950
rect 47761 1933 47821 1959
rect 47879 1933 47939 1959
rect 47997 1933 48057 1959
rect 51291 2114 51351 2140
rect 51409 2114 51469 2325
rect 51762 2319 51822 2351
rect 51880 2325 51940 2351
rect 51998 2325 52058 2351
rect 57676 2326 57736 2352
rect 57794 2326 57854 2352
rect 57912 2326 57972 2352
rect 58030 2332 58090 2352
rect 58030 2326 58091 2332
rect 58148 2326 58208 2352
rect 58266 2326 58326 2352
rect 51759 2303 51825 2319
rect 51759 2269 51775 2303
rect 51809 2269 51825 2303
rect 51759 2253 51825 2269
rect 51641 2186 51707 2202
rect 51641 2152 51657 2186
rect 51691 2152 51707 2186
rect 51641 2136 51707 2152
rect 53002 2149 53298 2200
rect 51644 2114 51704 2136
rect 53002 2134 53062 2149
rect 53120 2134 53180 2149
rect 53238 2134 53298 2149
rect 53356 2134 53416 2160
rect 53474 2134 53534 2160
rect 53592 2134 53652 2160
rect 54900 2149 55196 2200
rect 54900 2134 54960 2149
rect 55018 2134 55078 2149
rect 55136 2134 55196 2149
rect 55254 2134 55314 2160
rect 55372 2134 55432 2160
rect 55490 2134 55550 2160
rect 57913 2141 57971 2326
rect 49082 1950 49378 2001
rect 49082 1933 49142 1950
rect 49200 1933 49260 1950
rect 49318 1933 49378 1950
rect 45863 1716 45923 1733
rect 45981 1716 46041 1733
rect 46099 1716 46159 1733
rect 46347 1716 46407 1733
rect 45863 1665 46407 1716
rect 46465 1707 46525 1733
rect 46583 1707 46643 1733
rect 46701 1714 46761 1733
rect 46819 1714 46879 1733
rect 46937 1714 46997 1733
rect 47184 1714 47244 1733
rect 47302 1714 47362 1733
rect 44748 1584 44822 1641
rect 45988 1584 46048 1665
rect 46701 1663 47244 1714
rect 47286 1707 47362 1714
rect 47420 1707 47480 1733
rect 47761 1716 47821 1733
rect 47879 1716 47939 1733
rect 47997 1716 48057 1733
rect 48245 1716 48305 1733
rect 47286 1663 47361 1707
rect 47761 1665 48305 1716
rect 48363 1707 48423 1733
rect 48481 1707 48541 1733
rect 48599 1714 48659 1733
rect 48717 1714 48777 1733
rect 48835 1714 48895 1733
rect 49082 1714 49142 1733
rect 49200 1714 49260 1733
rect 44748 1559 46048 1584
rect 42633 1488 42887 1512
rect 44747 1511 46048 1559
rect 47286 1543 47346 1663
rect 42633 1454 42837 1488
rect 42871 1454 42887 1488
rect 42633 1438 42887 1454
rect 41637 1016 41697 1042
rect 41335 993 41402 1009
rect 41335 959 41351 993
rect 41385 959 41402 993
rect 41335 943 41402 959
rect 41335 815 41395 943
rect 41605 875 41672 882
rect 41755 875 41815 1042
rect 41873 1016 41933 1042
rect 41991 1016 42051 1042
rect 41605 866 41815 875
rect 41605 832 41621 866
rect 41655 832 41815 866
rect 41605 816 41815 832
rect 41335 799 41486 815
rect 41335 765 41436 799
rect 41470 765 41486 799
rect 41335 749 41486 765
rect 41335 710 41395 749
rect 41755 710 41815 816
rect 42109 875 42169 1042
rect 42227 1016 42287 1042
rect 42250 876 42317 883
rect 42244 875 42317 876
rect 42109 867 42317 875
rect 42109 833 42267 867
rect 42301 833 42317 867
rect 42109 817 42317 833
rect 42109 816 42306 817
rect 41871 782 41937 798
rect 41871 748 41887 782
rect 41921 748 41937 782
rect 41871 732 41937 748
rect 41989 783 42055 798
rect 41989 749 42005 783
rect 42039 749 42055 783
rect 41989 733 42055 749
rect 41873 710 41933 732
rect 41991 710 42051 733
rect 42109 710 42169 816
rect 42633 814 42693 1438
rect 44394 967 44690 1003
rect 44394 946 44454 967
rect 44512 946 44572 967
rect 44630 946 44690 967
rect 44748 966 45044 1002
rect 44748 946 44808 966
rect 44866 946 44926 966
rect 44984 946 45044 966
rect 45102 966 45398 1002
rect 45102 946 45162 966
rect 45220 946 45280 966
rect 45338 946 45398 966
rect 42543 798 42693 814
rect 42543 764 42559 798
rect 42593 764 42693 798
rect 42543 748 42693 764
rect 42633 710 42693 748
rect 45988 813 46048 1511
rect 46290 1463 46586 1523
rect 46290 1440 46350 1463
rect 46408 1440 46468 1463
rect 46526 1440 46586 1463
rect 46644 1464 46940 1524
rect 47285 1523 47346 1543
rect 46644 1440 46704 1464
rect 46762 1440 46822 1464
rect 46880 1440 46940 1464
rect 47266 1507 47346 1523
rect 47266 1473 47281 1507
rect 47315 1473 47346 1507
rect 47266 1457 47346 1473
rect 47285 1434 47346 1457
rect 47286 1288 47346 1434
rect 47285 1115 47346 1288
rect 46290 1014 46350 1040
rect 46258 873 46325 880
rect 46408 873 46468 1040
rect 46526 1014 46586 1040
rect 46644 1014 46704 1040
rect 46258 864 46468 873
rect 46258 830 46274 864
rect 46308 830 46468 864
rect 46258 814 46468 830
rect 45988 797 46139 813
rect 45988 763 46089 797
rect 46123 763 46139 797
rect 45988 747 46139 763
rect 44394 720 44454 746
rect 44512 720 44572 746
rect 44630 720 44690 746
rect 44748 726 44808 746
rect 44748 720 44809 726
rect 44866 720 44926 746
rect 44984 720 45044 746
rect 38548 666 38564 700
rect 38598 666 38614 700
rect 38548 650 38614 666
rect 38430 583 38496 599
rect 38430 549 38446 583
rect 38480 549 38496 583
rect 38430 533 38496 549
rect 38433 511 38493 533
rect 31272 435 31338 451
rect 23549 322 23984 330
rect 23549 288 23565 322
rect 23599 288 23984 322
rect 23549 279 23984 288
rect 14129 268 14195 275
rect 17273 268 17339 275
rect 20405 272 20471 279
rect 23549 272 23615 279
rect 30369 227 30420 415
rect 31205 300 31271 316
rect 29886 167 29952 227
rect 30352 167 30420 227
rect 30562 224 30645 284
rect 31045 224 31071 284
rect 31205 266 31221 300
rect 31255 266 31271 300
rect 31205 249 31271 266
rect 29886 109 29937 167
rect 30562 166 30622 224
rect 31212 166 31271 249
rect 29886 49 29952 109
rect 30352 49 30378 109
rect 30562 106 30645 166
rect 31045 106 31377 166
rect 31777 106 31803 166
rect 39437 484 39497 510
rect 38433 285 38493 311
rect 40735 484 40795 510
rect 41335 484 41395 510
rect 44631 535 44689 720
rect 42633 484 42693 510
rect 44631 509 44691 535
rect 44749 509 44809 720
rect 45102 714 45162 746
rect 45220 720 45280 746
rect 45338 720 45398 746
rect 45099 698 45165 714
rect 45988 708 46048 747
rect 46408 708 46468 814
rect 46762 873 46822 1040
rect 46880 1014 46940 1040
rect 46905 873 46972 880
rect 46762 864 46972 873
rect 46762 830 46922 864
rect 46956 830 46972 864
rect 46762 814 46972 830
rect 46524 780 46590 796
rect 46524 746 46540 780
rect 46574 746 46590 780
rect 46524 730 46590 746
rect 46642 781 46708 796
rect 46642 747 46658 781
rect 46692 747 46708 781
rect 46642 731 46708 747
rect 46526 708 46586 730
rect 46644 708 46704 731
rect 46762 708 46822 814
rect 47286 812 47346 1115
rect 47196 796 47346 812
rect 47196 762 47212 796
rect 47246 762 47346 796
rect 47196 746 47346 762
rect 47286 708 47346 746
rect 47886 1007 47946 1665
rect 48599 1663 49142 1714
rect 49184 1707 49260 1714
rect 49318 1707 49378 1733
rect 52518 1934 52578 1960
rect 52636 1934 52696 1960
rect 52754 1934 52814 1960
rect 51644 1888 51704 1914
rect 49184 1663 49259 1707
rect 51291 1692 51351 1714
rect 51409 1698 51469 1714
rect 51288 1676 51354 1692
rect 48188 1463 48484 1523
rect 48188 1440 48248 1463
rect 48306 1440 48366 1463
rect 48424 1440 48484 1463
rect 48542 1464 48838 1524
rect 48542 1440 48602 1464
rect 48660 1440 48720 1464
rect 48778 1440 48838 1464
rect 49184 1510 49244 1663
rect 51288 1642 51304 1676
rect 51338 1642 51354 1676
rect 51288 1626 51354 1642
rect 51403 1676 51477 1698
rect 51403 1642 51422 1676
rect 51456 1642 51477 1676
rect 53839 1951 54135 2002
rect 53839 1934 53899 1951
rect 53957 1934 54017 1951
rect 54075 1934 54135 1951
rect 54416 1934 54476 1960
rect 54534 1934 54594 1960
rect 54652 1934 54712 1960
rect 57913 2115 57973 2141
rect 58031 2115 58091 2326
rect 58384 2320 58444 2352
rect 58502 2326 58562 2352
rect 58620 2326 58680 2352
rect 58381 2304 58447 2320
rect 58381 2270 58397 2304
rect 58431 2270 58447 2304
rect 58381 2254 58447 2270
rect 58263 2187 58329 2203
rect 58263 2153 58279 2187
rect 58313 2153 58329 2187
rect 58263 2137 58329 2153
rect 59624 2150 59920 2201
rect 58266 2115 58326 2137
rect 59624 2135 59684 2150
rect 59742 2135 59802 2150
rect 59860 2135 59920 2150
rect 59978 2135 60038 2161
rect 60096 2135 60156 2161
rect 60214 2135 60274 2161
rect 61522 2150 61818 2201
rect 61522 2135 61582 2150
rect 61640 2135 61700 2150
rect 61758 2135 61818 2150
rect 61876 2135 61936 2161
rect 61994 2135 62054 2161
rect 62112 2135 62172 2161
rect 55737 1951 56033 2002
rect 55737 1934 55797 1951
rect 55855 1934 55915 1951
rect 55973 1934 56033 1951
rect 52518 1717 52578 1734
rect 52636 1717 52696 1734
rect 52754 1717 52814 1734
rect 53002 1717 53062 1734
rect 52518 1666 53062 1717
rect 53120 1708 53180 1734
rect 53238 1708 53298 1734
rect 53356 1715 53416 1734
rect 53474 1715 53534 1734
rect 53592 1715 53652 1734
rect 53839 1715 53899 1734
rect 53957 1715 54017 1734
rect 51403 1585 51477 1642
rect 52643 1585 52703 1666
rect 53356 1664 53899 1715
rect 53941 1708 54017 1715
rect 54075 1708 54135 1734
rect 54416 1717 54476 1734
rect 54534 1717 54594 1734
rect 54652 1717 54712 1734
rect 54900 1717 54960 1734
rect 53941 1664 54016 1708
rect 54416 1666 54960 1717
rect 55018 1708 55078 1734
rect 55136 1708 55196 1734
rect 55254 1715 55314 1734
rect 55372 1715 55432 1734
rect 55490 1715 55550 1734
rect 55737 1715 55797 1734
rect 55855 1715 55915 1734
rect 51403 1560 52703 1585
rect 51402 1512 52703 1560
rect 53941 1544 54001 1664
rect 49184 1486 49438 1510
rect 49184 1452 49388 1486
rect 49422 1452 49438 1486
rect 49184 1436 49438 1452
rect 48188 1014 48248 1040
rect 47886 991 47953 1007
rect 47886 957 47902 991
rect 47936 957 47953 991
rect 47886 941 47953 957
rect 47886 813 47946 941
rect 48156 873 48223 880
rect 48306 873 48366 1040
rect 48424 1014 48484 1040
rect 48542 1014 48602 1040
rect 48156 864 48366 873
rect 48156 830 48172 864
rect 48206 830 48366 864
rect 48156 814 48366 830
rect 47886 797 48037 813
rect 47886 763 47987 797
rect 48021 763 48037 797
rect 47886 747 48037 763
rect 47886 708 47946 747
rect 48306 708 48366 814
rect 48660 873 48720 1040
rect 48778 1014 48838 1040
rect 48801 874 48868 881
rect 48795 873 48868 874
rect 48660 865 48868 873
rect 48660 831 48818 865
rect 48852 831 48868 865
rect 48660 815 48868 831
rect 48660 814 48857 815
rect 48422 780 48488 796
rect 48422 746 48438 780
rect 48472 746 48488 780
rect 48422 730 48488 746
rect 48540 781 48606 796
rect 48540 747 48556 781
rect 48590 747 48606 781
rect 48540 731 48606 747
rect 48424 708 48484 730
rect 48542 708 48602 731
rect 48660 708 48720 814
rect 49184 812 49244 1436
rect 51049 968 51345 1004
rect 51049 947 51109 968
rect 51167 947 51227 968
rect 51285 947 51345 968
rect 51403 967 51699 1003
rect 51403 947 51463 967
rect 51521 947 51581 967
rect 51639 947 51699 967
rect 51757 967 52053 1003
rect 51757 947 51817 967
rect 51875 947 51935 967
rect 51993 947 52053 967
rect 49094 796 49244 812
rect 49094 762 49110 796
rect 49144 762 49244 796
rect 49094 746 49244 762
rect 52643 814 52703 1512
rect 52945 1464 53241 1524
rect 52945 1441 53005 1464
rect 53063 1441 53123 1464
rect 53181 1441 53241 1464
rect 53299 1465 53595 1525
rect 53940 1524 54001 1544
rect 53299 1441 53359 1465
rect 53417 1441 53477 1465
rect 53535 1441 53595 1465
rect 53921 1508 54001 1524
rect 53921 1474 53936 1508
rect 53970 1474 54001 1508
rect 53921 1458 54001 1474
rect 53940 1435 54001 1458
rect 53941 1289 54001 1435
rect 53940 1116 54001 1289
rect 52945 1015 53005 1041
rect 52913 874 52980 881
rect 53063 874 53123 1041
rect 53181 1015 53241 1041
rect 53299 1015 53359 1041
rect 52913 865 53123 874
rect 52913 831 52929 865
rect 52963 831 53123 865
rect 52913 815 53123 831
rect 52643 798 52794 814
rect 52643 764 52744 798
rect 52778 764 52794 798
rect 52643 748 52794 764
rect 49184 708 49244 746
rect 51049 721 51109 747
rect 51167 721 51227 747
rect 51285 721 51345 747
rect 51403 727 51463 747
rect 51403 721 51464 727
rect 51521 721 51581 747
rect 51639 721 51699 747
rect 45099 664 45115 698
rect 45149 664 45165 698
rect 45099 648 45165 664
rect 44981 581 45047 597
rect 44981 547 44997 581
rect 45031 547 45047 581
rect 44981 531 45047 547
rect 44984 509 45044 531
rect 39857 284 39917 310
rect 39975 284 40035 310
rect 40093 284 40153 310
rect 40211 284 40271 310
rect 41755 284 41815 310
rect 41873 284 41933 310
rect 41991 284 42051 310
rect 42109 284 42169 310
rect 29886 -9 29937 49
rect 30562 48 30622 106
rect 38080 89 38140 111
rect 38198 89 38258 111
rect 31289 48 31355 50
rect 29886 -69 29952 -9
rect 30352 -69 30378 -9
rect 30562 -12 30645 48
rect 31045 -12 31071 48
rect 31289 34 31377 48
rect 31289 0 31305 34
rect 31339 0 31377 34
rect 31289 -12 31377 0
rect 31777 -12 31803 48
rect 38077 73 38143 89
rect 38077 39 38093 73
rect 38127 39 38143 73
rect 38077 23 38143 39
rect 38195 73 38261 89
rect 38195 39 38211 73
rect 38245 39 38261 73
rect 45988 482 46048 508
rect 44984 283 45044 309
rect 47286 482 47346 508
rect 47886 482 47946 508
rect 51286 536 51344 721
rect 51286 510 51346 536
rect 51404 510 51464 721
rect 51757 715 51817 747
rect 51875 721 51935 747
rect 51993 721 52053 747
rect 51754 699 51820 715
rect 52643 709 52703 748
rect 53063 709 53123 815
rect 53417 874 53477 1041
rect 53535 1015 53595 1041
rect 53560 874 53627 881
rect 53417 865 53627 874
rect 53417 831 53577 865
rect 53611 831 53627 865
rect 53417 815 53627 831
rect 53179 781 53245 797
rect 53179 747 53195 781
rect 53229 747 53245 781
rect 53179 731 53245 747
rect 53297 782 53363 797
rect 53297 748 53313 782
rect 53347 748 53363 782
rect 53297 732 53363 748
rect 53181 709 53241 731
rect 53299 709 53359 732
rect 53417 709 53477 815
rect 53941 813 54001 1116
rect 53851 797 54001 813
rect 53851 763 53867 797
rect 53901 763 54001 797
rect 53851 747 54001 763
rect 53941 709 54001 747
rect 54541 1008 54601 1666
rect 55254 1664 55797 1715
rect 55839 1708 55915 1715
rect 55973 1708 56033 1734
rect 59140 1935 59200 1961
rect 59258 1935 59318 1961
rect 59376 1935 59436 1961
rect 58266 1889 58326 1915
rect 55839 1664 55914 1708
rect 57913 1693 57973 1715
rect 58031 1699 58091 1715
rect 57910 1677 57976 1693
rect 54843 1464 55139 1524
rect 54843 1441 54903 1464
rect 54961 1441 55021 1464
rect 55079 1441 55139 1464
rect 55197 1465 55493 1525
rect 55197 1441 55257 1465
rect 55315 1441 55375 1465
rect 55433 1441 55493 1465
rect 55839 1511 55899 1664
rect 57910 1643 57926 1677
rect 57960 1643 57976 1677
rect 57910 1627 57976 1643
rect 58025 1677 58099 1699
rect 58025 1643 58044 1677
rect 58078 1643 58099 1677
rect 60461 1952 60757 2003
rect 60461 1935 60521 1952
rect 60579 1935 60639 1952
rect 60697 1935 60757 1952
rect 61038 1935 61098 1961
rect 61156 1935 61216 1961
rect 61274 1935 61334 1961
rect 70455 2149 70509 2209
rect 70909 2149 70935 2209
rect 70455 2091 70494 2149
rect 70455 2031 70509 2091
rect 70909 2090 70935 2091
rect 71096 2090 71162 2093
rect 70909 2077 71162 2090
rect 70909 2043 71112 2077
rect 71146 2043 71162 2077
rect 70909 2031 71162 2043
rect 71327 2091 71384 2498
rect 71594 2283 71639 3057
rect 71594 2223 71842 2283
rect 72042 2223 72068 2283
rect 71483 2091 71562 2102
rect 71327 2089 71842 2091
rect 71327 2031 71496 2089
rect 71551 2031 71842 2089
rect 72242 2031 72268 2091
rect 62359 1952 62655 2003
rect 62359 1935 62419 1952
rect 62477 1935 62537 1952
rect 62595 1935 62655 1952
rect 70455 1973 70494 2031
rect 71095 2027 71162 2031
rect 71483 2021 71562 2031
rect 71196 1973 71283 1990
rect 70455 1913 70509 1973
rect 70909 1913 70935 1973
rect 71196 1971 71842 1973
rect 71196 1913 71211 1971
rect 71266 1913 71842 1971
rect 72242 1913 72268 1973
rect 71196 1895 71283 1913
rect 59140 1718 59200 1735
rect 59258 1718 59318 1735
rect 59376 1718 59436 1735
rect 59624 1718 59684 1735
rect 59140 1667 59684 1718
rect 59742 1709 59802 1735
rect 59860 1709 59920 1735
rect 59978 1716 60038 1735
rect 60096 1716 60156 1735
rect 60214 1716 60274 1735
rect 60461 1716 60521 1735
rect 60579 1716 60639 1735
rect 58025 1586 58099 1643
rect 59265 1586 59325 1667
rect 59978 1665 60521 1716
rect 60563 1709 60639 1716
rect 60697 1709 60757 1735
rect 61038 1718 61098 1735
rect 61156 1718 61216 1735
rect 61274 1718 61334 1735
rect 61522 1718 61582 1735
rect 60563 1665 60638 1709
rect 61038 1667 61582 1718
rect 61640 1709 61700 1735
rect 61758 1709 61818 1735
rect 61876 1716 61936 1735
rect 61994 1716 62054 1735
rect 62112 1716 62172 1735
rect 62359 1716 62419 1735
rect 62477 1716 62537 1735
rect 58025 1561 59325 1586
rect 58024 1513 59325 1561
rect 60563 1545 60623 1665
rect 55839 1487 56093 1511
rect 55839 1453 56043 1487
rect 56077 1453 56093 1487
rect 55839 1437 56093 1453
rect 54843 1015 54903 1041
rect 54541 992 54608 1008
rect 54541 958 54557 992
rect 54591 958 54608 992
rect 54541 942 54608 958
rect 54541 814 54601 942
rect 54811 874 54878 881
rect 54961 874 55021 1041
rect 55079 1015 55139 1041
rect 55197 1015 55257 1041
rect 54811 865 55021 874
rect 54811 831 54827 865
rect 54861 831 55021 865
rect 54811 815 55021 831
rect 54541 798 54692 814
rect 54541 764 54642 798
rect 54676 764 54692 798
rect 54541 748 54692 764
rect 54541 709 54601 748
rect 54961 709 55021 815
rect 55315 874 55375 1041
rect 55433 1015 55493 1041
rect 55456 875 55523 882
rect 55450 874 55523 875
rect 55315 866 55523 874
rect 55315 832 55473 866
rect 55507 832 55523 866
rect 55315 816 55523 832
rect 55315 815 55512 816
rect 55077 781 55143 797
rect 55077 747 55093 781
rect 55127 747 55143 781
rect 55077 731 55143 747
rect 55195 782 55261 797
rect 55195 748 55211 782
rect 55245 748 55261 782
rect 55195 732 55261 748
rect 55079 709 55139 731
rect 55197 709 55257 732
rect 55315 709 55375 815
rect 55839 813 55899 1437
rect 57671 969 57967 1005
rect 57671 948 57731 969
rect 57789 948 57849 969
rect 57907 948 57967 969
rect 58025 968 58321 1004
rect 58025 948 58085 968
rect 58143 948 58203 968
rect 58261 948 58321 968
rect 58379 968 58675 1004
rect 58379 948 58439 968
rect 58497 948 58557 968
rect 58615 948 58675 968
rect 55749 797 55899 813
rect 55749 763 55765 797
rect 55799 763 55899 797
rect 55749 747 55899 763
rect 59265 815 59325 1513
rect 59567 1465 59863 1525
rect 59567 1442 59627 1465
rect 59685 1442 59745 1465
rect 59803 1442 59863 1465
rect 59921 1466 60217 1526
rect 60562 1525 60623 1545
rect 59921 1442 59981 1466
rect 60039 1442 60099 1466
rect 60157 1442 60217 1466
rect 60543 1509 60623 1525
rect 60543 1475 60558 1509
rect 60592 1475 60623 1509
rect 60543 1459 60623 1475
rect 60562 1436 60623 1459
rect 60563 1290 60623 1436
rect 60562 1117 60623 1290
rect 59567 1016 59627 1042
rect 59535 875 59602 882
rect 59685 875 59745 1042
rect 59803 1016 59863 1042
rect 59921 1016 59981 1042
rect 59535 866 59745 875
rect 59535 832 59551 866
rect 59585 832 59745 866
rect 59535 816 59745 832
rect 59265 799 59416 815
rect 59265 765 59366 799
rect 59400 765 59416 799
rect 59265 749 59416 765
rect 55839 709 55899 747
rect 57671 722 57731 748
rect 57789 722 57849 748
rect 57907 722 57967 748
rect 58025 728 58085 748
rect 58025 722 58086 728
rect 58143 722 58203 748
rect 58261 722 58321 748
rect 51754 665 51770 699
rect 51804 665 51820 699
rect 51754 649 51820 665
rect 51636 582 51702 598
rect 51636 548 51652 582
rect 51686 548 51702 582
rect 51636 532 51702 548
rect 51639 510 51699 532
rect 49184 482 49244 508
rect 46408 282 46468 308
rect 46526 282 46586 308
rect 46644 282 46704 308
rect 46762 282 46822 308
rect 48306 282 48366 308
rect 48424 282 48484 308
rect 48542 282 48602 308
rect 48660 282 48720 308
rect 44631 87 44691 109
rect 44749 87 44809 109
rect 44628 71 44694 87
rect 38195 23 38261 39
rect 31289 -16 31355 -12
rect 31289 -70 31354 -68
rect 29926 -187 29952 -127
rect 30352 -187 30422 -127
rect 30371 -245 30422 -187
rect 29926 -305 29952 -245
rect 30352 -305 30422 -245
rect 30371 -363 30422 -305
rect 29926 -423 29952 -363
rect 30352 -423 30422 -363
rect 30561 -130 30645 -70
rect 31045 -130 31071 -70
rect 31289 -84 31377 -70
rect 31289 -118 31304 -84
rect 31338 -118 31377 -84
rect 31289 -130 31377 -118
rect 31777 -130 31803 -70
rect 30561 -188 30621 -130
rect 31289 -134 31354 -130
rect 44628 37 44644 71
rect 44678 37 44694 71
rect 44628 21 44694 37
rect 44746 71 44812 87
rect 44746 37 44762 71
rect 44796 37 44812 71
rect 52643 483 52703 509
rect 51639 284 51699 310
rect 53941 483 54001 509
rect 54541 483 54601 509
rect 57908 537 57966 722
rect 57908 511 57968 537
rect 58026 511 58086 722
rect 58379 716 58439 748
rect 58497 722 58557 748
rect 58615 722 58675 748
rect 58376 700 58442 716
rect 59265 710 59325 749
rect 59685 710 59745 816
rect 60039 875 60099 1042
rect 60157 1016 60217 1042
rect 60182 875 60249 882
rect 60039 866 60249 875
rect 60039 832 60199 866
rect 60233 832 60249 866
rect 60039 816 60249 832
rect 59801 782 59867 798
rect 59801 748 59817 782
rect 59851 748 59867 782
rect 59801 732 59867 748
rect 59919 783 59985 798
rect 59919 749 59935 783
rect 59969 749 59985 783
rect 59919 733 59985 749
rect 59803 710 59863 732
rect 59921 710 59981 733
rect 60039 710 60099 816
rect 60563 814 60623 1117
rect 60473 798 60623 814
rect 60473 764 60489 798
rect 60523 764 60623 798
rect 60473 748 60623 764
rect 60563 710 60623 748
rect 61163 1009 61223 1667
rect 61876 1665 62419 1716
rect 62461 1709 62537 1716
rect 62595 1709 62655 1735
rect 70455 1795 70509 1855
rect 70909 1795 70935 1855
rect 70455 1737 70494 1795
rect 71234 1737 71283 1895
rect 71716 1855 71782 1858
rect 72315 1900 72381 1916
rect 72315 1866 72331 1900
rect 72365 1866 72381 1900
rect 71716 1842 71842 1855
rect 71716 1808 71732 1842
rect 71766 1808 71842 1842
rect 71716 1795 71842 1808
rect 72242 1795 72268 1855
rect 72315 1850 72381 1866
rect 71716 1792 71782 1795
rect 62461 1665 62536 1709
rect 70455 1677 70509 1737
rect 70909 1677 71283 1737
rect 71325 1737 71394 1742
rect 71325 1723 71842 1737
rect 71325 1689 71342 1723
rect 71376 1689 71842 1723
rect 71325 1677 71842 1689
rect 72242 1677 72268 1737
rect 61465 1465 61761 1525
rect 61465 1442 61525 1465
rect 61583 1442 61643 1465
rect 61701 1442 61761 1465
rect 61819 1466 62115 1526
rect 61819 1442 61879 1466
rect 61937 1442 61997 1466
rect 62055 1442 62115 1466
rect 62461 1512 62521 1665
rect 70455 1619 70494 1677
rect 71325 1673 71392 1677
rect 70455 1559 70509 1619
rect 70909 1559 70935 1619
rect 62461 1488 62715 1512
rect 62461 1454 62665 1488
rect 62699 1454 62715 1488
rect 62461 1438 62715 1454
rect 61465 1016 61525 1042
rect 61163 993 61230 1009
rect 61163 959 61179 993
rect 61213 959 61230 993
rect 61163 943 61230 959
rect 61163 815 61223 943
rect 61433 875 61500 882
rect 61583 875 61643 1042
rect 61701 1016 61761 1042
rect 61819 1016 61879 1042
rect 61433 866 61643 875
rect 61433 832 61449 866
rect 61483 832 61643 866
rect 61433 816 61643 832
rect 61163 799 61314 815
rect 61163 765 61264 799
rect 61298 765 61314 799
rect 61163 749 61314 765
rect 61163 710 61223 749
rect 61583 710 61643 816
rect 61937 875 61997 1042
rect 62055 1016 62115 1042
rect 62078 876 62145 883
rect 62072 875 62145 876
rect 61937 867 62145 875
rect 61937 833 62095 867
rect 62129 833 62145 867
rect 61937 817 62145 833
rect 61937 816 62134 817
rect 61699 782 61765 798
rect 61699 748 61715 782
rect 61749 748 61765 782
rect 61699 732 61765 748
rect 61817 783 61883 798
rect 61817 749 61833 783
rect 61867 749 61883 783
rect 61817 733 61883 749
rect 61701 710 61761 732
rect 61819 710 61879 733
rect 61937 710 61997 816
rect 62461 814 62521 1438
rect 63535 1429 63831 1465
rect 63535 1408 63595 1429
rect 63653 1408 63713 1429
rect 63771 1408 63831 1429
rect 63889 1428 64185 1464
rect 63889 1408 63949 1428
rect 64007 1408 64067 1428
rect 64125 1408 64185 1428
rect 64243 1428 64539 1464
rect 64243 1408 64303 1428
rect 64361 1408 64421 1428
rect 64479 1408 64539 1428
rect 70455 1322 70509 1382
rect 70909 1322 70935 1382
rect 70455 1264 70494 1322
rect 71325 1264 71382 1673
rect 72323 1541 72374 1850
rect 63535 1182 63595 1208
rect 63653 1182 63713 1208
rect 63771 1182 63831 1208
rect 63889 1188 63949 1208
rect 63889 1182 63950 1188
rect 64007 1182 64067 1208
rect 64125 1182 64185 1208
rect 63772 997 63830 1182
rect 63772 971 63832 997
rect 63890 971 63950 1182
rect 64243 1176 64303 1208
rect 64361 1182 64421 1208
rect 64479 1182 64539 1208
rect 70455 1204 70509 1264
rect 70909 1204 71382 1264
rect 71594 1481 71842 1541
rect 72042 1481 72374 1541
rect 64240 1160 64306 1176
rect 64240 1126 64256 1160
rect 64290 1126 64306 1160
rect 64240 1110 64306 1126
rect 70455 1146 70494 1204
rect 70455 1086 70509 1146
rect 70909 1086 70935 1146
rect 64122 1043 64188 1059
rect 64122 1009 64138 1043
rect 64172 1009 64188 1043
rect 64122 993 64188 1009
rect 64125 971 64185 993
rect 62371 798 62521 814
rect 62371 764 62387 798
rect 62421 764 62521 798
rect 62371 748 62521 764
rect 62461 710 62521 748
rect 58376 666 58392 700
rect 58426 666 58442 700
rect 58376 650 58442 666
rect 58258 583 58324 599
rect 58258 549 58274 583
rect 58308 549 58324 583
rect 58258 533 58324 549
rect 58261 511 58321 533
rect 55839 483 55899 509
rect 53063 283 53123 309
rect 53181 283 53241 309
rect 53299 283 53359 309
rect 53417 283 53477 309
rect 54961 283 55021 309
rect 55079 283 55139 309
rect 55197 283 55257 309
rect 55315 283 55375 309
rect 51286 88 51346 110
rect 51404 88 51464 110
rect 51283 72 51349 88
rect 44746 21 44812 37
rect 51283 38 51299 72
rect 51333 38 51349 72
rect 51283 22 51349 38
rect 51401 72 51467 88
rect 51401 38 51417 72
rect 51451 38 51467 72
rect 59265 484 59325 510
rect 58261 285 58321 311
rect 60563 484 60623 510
rect 61163 484 61223 510
rect 70654 849 70709 909
rect 70909 849 70935 909
rect 70654 791 70693 849
rect 64125 745 64185 771
rect 70654 731 70709 791
rect 70909 731 70935 791
rect 71055 767 71121 783
rect 71055 733 71071 767
rect 71105 733 71121 767
rect 70654 673 70693 731
rect 71055 717 71121 733
rect 71058 673 71118 717
rect 71594 673 71639 1481
rect 70654 613 70709 673
rect 70909 613 71639 673
rect 63772 549 63832 571
rect 63890 549 63950 571
rect 63769 533 63835 549
rect 62461 484 62521 510
rect 63769 499 63785 533
rect 63819 499 63835 533
rect 63769 483 63835 499
rect 63887 533 63953 549
rect 63887 499 63903 533
rect 63937 499 63953 533
rect 63887 483 63953 499
rect 59685 284 59745 310
rect 59803 284 59863 310
rect 59921 284 59981 310
rect 60039 284 60099 310
rect 61583 284 61643 310
rect 61701 284 61761 310
rect 61819 284 61879 310
rect 61937 284 61997 310
rect 57908 89 57968 111
rect 58026 89 58086 111
rect 57905 73 57971 89
rect 51401 22 51467 38
rect 57905 39 57921 73
rect 57955 39 57971 73
rect 57905 23 57971 39
rect 58023 73 58089 89
rect 58023 39 58039 73
rect 58073 39 58089 73
rect 58023 23 58089 39
rect 65766 -122 66062 -71
rect 65766 -137 65826 -122
rect 65884 -137 65944 -122
rect 66002 -137 66062 -122
rect 66120 -137 66180 -111
rect 66238 -137 66298 -111
rect 66356 -137 66416 -111
rect 30561 -248 30645 -188
rect 31045 -248 31377 -188
rect 31777 -248 31803 -188
rect 30561 -306 30621 -248
rect 30561 -366 30645 -306
rect 31045 -366 31071 -306
rect 31212 -331 31271 -248
rect 31205 -348 31271 -331
rect 65282 -337 65342 -311
rect 65400 -337 65460 -311
rect 65518 -337 65578 -311
rect 30371 -610 30422 -423
rect 31205 -382 31221 -348
rect 31255 -382 31271 -348
rect 31205 -398 31271 -382
rect 70654 -87 70709 -27
rect 70909 -86 71639 -27
rect 70909 -87 71212 -86
rect 70654 -145 70693 -87
rect 71195 -144 71212 -87
rect 71267 -87 71639 -86
rect 71267 -144 71282 -87
rect 70654 -205 70709 -145
rect 70909 -205 70935 -145
rect 71195 -163 71282 -144
rect 70654 -263 70693 -205
rect 66603 -320 66899 -269
rect 66603 -337 66663 -320
rect 66721 -337 66781 -320
rect 66839 -337 66899 -320
rect 67075 -319 67371 -283
rect 67075 -340 67135 -319
rect 67193 -340 67253 -319
rect 67311 -340 67371 -319
rect 67429 -320 67725 -284
rect 67429 -340 67489 -320
rect 67547 -340 67607 -320
rect 67665 -340 67725 -320
rect 67783 -320 68079 -284
rect 67783 -340 67843 -320
rect 67901 -340 67961 -320
rect 68019 -340 68079 -320
rect 70654 -323 70709 -263
rect 70909 -323 70935 -263
rect 65282 -554 65342 -537
rect 65400 -554 65460 -537
rect 65518 -554 65578 -537
rect 65766 -554 65826 -537
rect 65282 -605 65826 -554
rect 65884 -563 65944 -537
rect 66002 -563 66062 -537
rect 66120 -556 66180 -537
rect 66238 -556 66298 -537
rect 66356 -556 66416 -537
rect 66603 -556 66663 -537
rect 66721 -556 66781 -537
rect 30084 -670 30152 -610
rect 30352 -670 30422 -610
rect 31273 -638 31339 -622
rect 30509 -660 30563 -644
rect 30084 -728 30135 -670
rect 30509 -694 30519 -660
rect 30553 -694 30563 -660
rect 30509 -712 30563 -694
rect 31273 -672 31289 -638
rect 31323 -672 31339 -638
rect 31273 -712 31339 -672
rect 30371 -728 31377 -712
rect 30084 -788 30152 -728
rect 30352 -772 31377 -728
rect 31577 -772 31603 -712
rect 30352 -787 30422 -772
rect 30352 -788 30378 -787
rect 30084 -846 30135 -788
rect 65407 -809 65467 -605
rect 66120 -607 66663 -556
rect 66705 -563 66781 -556
rect 66839 -563 66899 -537
rect 70455 -528 70509 -468
rect 70909 -528 70935 -468
rect 66705 -607 66780 -563
rect 67075 -566 67135 -540
rect 67193 -566 67253 -540
rect 67311 -566 67371 -540
rect 67429 -560 67489 -540
rect 67429 -566 67490 -560
rect 67547 -566 67607 -540
rect 67665 -566 67725 -540
rect 66705 -689 66765 -607
rect 66705 -707 66939 -689
rect 66705 -741 66888 -707
rect 66922 -741 66939 -707
rect 65709 -807 66005 -747
rect 41885 -846 41951 -830
rect 30084 -906 30152 -846
rect 30352 -906 30378 -846
rect 41885 -880 41901 -846
rect 41935 -880 41951 -846
rect 41885 -896 41951 -880
rect 42003 -846 42069 -830
rect 42003 -880 42019 -846
rect 42053 -880 42069 -846
rect 42003 -896 42069 -880
rect 48439 -841 48505 -825
rect 48439 -875 48455 -841
rect 48489 -875 48505 -841
rect 48439 -891 48505 -875
rect 48557 -841 48623 -825
rect 65407 -826 65538 -809
rect 48557 -875 48573 -841
rect 48607 -875 48623 -841
rect 48557 -891 48623 -875
rect 55088 -853 55154 -837
rect 55088 -887 55104 -853
rect 55138 -887 55154 -853
rect 41888 -918 41948 -896
rect 42006 -918 42066 -896
rect 48442 -913 48502 -891
rect 48560 -913 48620 -891
rect 55088 -903 55154 -887
rect 55206 -853 55272 -837
rect 55206 -887 55222 -853
rect 55256 -887 55272 -853
rect 55206 -903 55272 -887
rect 65407 -860 65488 -826
rect 65522 -860 65538 -826
rect 65709 -830 65769 -807
rect 65827 -830 65887 -807
rect 65945 -830 66005 -807
rect 66063 -806 66359 -746
rect 66063 -830 66123 -806
rect 66181 -830 66241 -806
rect 66299 -830 66359 -806
rect 66705 -757 66939 -741
rect 67312 -751 67370 -566
rect 65407 -877 65538 -860
rect 42241 -1118 42301 -1092
rect 55091 -925 55151 -903
rect 55209 -925 55269 -903
rect 48795 -1113 48855 -1087
rect 30697 -1334 30757 -1318
rect 30124 -1417 30150 -1357
rect 30350 -1417 30418 -1357
rect 30367 -1475 30418 -1417
rect 30124 -1535 30150 -1475
rect 30350 -1482 30418 -1475
rect 30697 -1368 30711 -1334
rect 30745 -1368 30757 -1334
rect 30697 -1482 30757 -1368
rect 41888 -1344 41948 -1318
rect 30350 -1535 31375 -1482
rect 30367 -1542 31375 -1535
rect 31575 -1542 31601 -1482
rect 41888 -1529 41946 -1344
rect 42006 -1529 42066 -1318
rect 42241 -1340 42301 -1318
rect 48442 -1339 48502 -1313
rect 42238 -1356 42304 -1340
rect 42238 -1390 42254 -1356
rect 42288 -1390 42304 -1356
rect 42238 -1406 42304 -1390
rect 42356 -1473 42422 -1457
rect 42356 -1507 42372 -1473
rect 42406 -1507 42422 -1473
rect 42356 -1523 42422 -1507
rect 30367 -1593 30418 -1542
rect 30124 -1653 30150 -1593
rect 30350 -1653 30418 -1593
rect 31270 -1583 31336 -1542
rect 31270 -1617 31286 -1583
rect 31320 -1617 31336 -1583
rect 41651 -1555 41711 -1529
rect 41769 -1555 41829 -1529
rect 41887 -1555 41947 -1529
rect 42005 -1535 42066 -1529
rect 42005 -1555 42065 -1535
rect 42123 -1555 42183 -1529
rect 42241 -1555 42301 -1529
rect 42359 -1555 42419 -1523
rect 48442 -1524 48500 -1339
rect 48560 -1524 48620 -1313
rect 48795 -1335 48855 -1313
rect 55444 -1125 55504 -1099
rect 48792 -1351 48858 -1335
rect 48792 -1385 48808 -1351
rect 48842 -1385 48858 -1351
rect 48792 -1401 48858 -1385
rect 55091 -1351 55151 -1325
rect 48910 -1468 48976 -1452
rect 48910 -1502 48926 -1468
rect 48960 -1502 48976 -1468
rect 48910 -1518 48976 -1502
rect 42477 -1555 42537 -1529
rect 42595 -1555 42655 -1529
rect 48205 -1550 48265 -1524
rect 48323 -1550 48383 -1524
rect 48441 -1550 48501 -1524
rect 48559 -1530 48620 -1524
rect 48559 -1550 48619 -1530
rect 48677 -1550 48737 -1524
rect 48795 -1550 48855 -1524
rect 48913 -1550 48973 -1518
rect 49031 -1550 49091 -1524
rect 49149 -1550 49209 -1524
rect 55091 -1536 55149 -1351
rect 55209 -1536 55269 -1325
rect 55444 -1347 55504 -1325
rect 55441 -1363 55507 -1347
rect 55441 -1397 55457 -1363
rect 55491 -1397 55507 -1363
rect 55441 -1413 55507 -1397
rect 63542 -1416 63838 -1380
rect 63542 -1437 63602 -1416
rect 63660 -1437 63720 -1416
rect 63778 -1437 63838 -1416
rect 63896 -1417 64192 -1381
rect 63896 -1437 63956 -1417
rect 64014 -1437 64074 -1417
rect 64132 -1437 64192 -1417
rect 64250 -1417 64546 -1381
rect 64250 -1437 64310 -1417
rect 64368 -1437 64428 -1417
rect 64486 -1437 64546 -1417
rect 55559 -1480 55625 -1464
rect 55559 -1514 55575 -1480
rect 55609 -1514 55625 -1480
rect 55559 -1530 55625 -1514
rect 31270 -1633 31336 -1617
rect 779 -1737 1075 -1698
rect 779 -1752 839 -1737
rect 897 -1752 957 -1737
rect 1015 -1752 1075 -1737
rect 1246 -1737 1542 -1698
rect 1246 -1752 1306 -1737
rect 1364 -1752 1424 -1737
rect 1482 -1752 1542 -1737
rect 1600 -1737 1896 -1698
rect 1600 -1752 1660 -1737
rect 1718 -1752 1778 -1737
rect 1836 -1752 1896 -1737
rect 2073 -1737 2369 -1698
rect 2073 -1752 2133 -1737
rect 2191 -1752 2251 -1737
rect 2309 -1752 2369 -1737
rect 3923 -1737 4219 -1698
rect 3923 -1752 3983 -1737
rect 4041 -1752 4101 -1737
rect 4159 -1752 4219 -1737
rect 4390 -1737 4686 -1698
rect 4390 -1752 4450 -1737
rect 4508 -1752 4568 -1737
rect 4626 -1752 4686 -1737
rect 4744 -1737 5040 -1698
rect 4744 -1752 4804 -1737
rect 4862 -1752 4922 -1737
rect 4980 -1752 5040 -1737
rect 5217 -1737 5513 -1698
rect 5217 -1752 5277 -1737
rect 5335 -1752 5395 -1737
rect 5453 -1752 5513 -1737
rect 7055 -1733 7351 -1694
rect 7055 -1748 7115 -1733
rect 7173 -1748 7233 -1733
rect 7291 -1748 7351 -1733
rect 7522 -1733 7818 -1694
rect 7522 -1748 7582 -1733
rect 7640 -1748 7700 -1733
rect 7758 -1748 7818 -1733
rect 7876 -1733 8172 -1694
rect 7876 -1748 7936 -1733
rect 7994 -1748 8054 -1733
rect 8112 -1748 8172 -1733
rect 8349 -1733 8645 -1694
rect 8349 -1748 8409 -1733
rect 8467 -1748 8527 -1733
rect 8585 -1748 8645 -1733
rect 10199 -1733 10495 -1694
rect 10199 -1748 10259 -1733
rect 10317 -1748 10377 -1733
rect 10435 -1748 10495 -1733
rect 10666 -1733 10962 -1694
rect 10666 -1748 10726 -1733
rect 10784 -1748 10844 -1733
rect 10902 -1748 10962 -1733
rect 11020 -1733 11316 -1694
rect 11020 -1748 11080 -1733
rect 11138 -1748 11198 -1733
rect 11256 -1748 11316 -1733
rect 11493 -1733 11789 -1694
rect 11493 -1748 11553 -1733
rect 11611 -1748 11671 -1733
rect 11729 -1748 11789 -1733
rect 13401 -1737 13697 -1698
rect 338 -1936 634 -1897
rect 338 -1952 398 -1936
rect 456 -1952 516 -1936
rect 574 -1952 634 -1936
rect 2546 -1936 2842 -1897
rect 2546 -1952 2606 -1936
rect 2664 -1952 2724 -1936
rect 2782 -1952 2842 -1936
rect 3482 -1936 3778 -1897
rect 3482 -1952 3542 -1936
rect 3600 -1952 3660 -1936
rect 3718 -1952 3778 -1936
rect 5690 -1936 5986 -1897
rect 5690 -1952 5750 -1936
rect 5808 -1952 5868 -1936
rect 5926 -1952 5986 -1936
rect 6614 -1932 6910 -1893
rect 6614 -1948 6674 -1932
rect 6732 -1948 6792 -1932
rect 6850 -1948 6910 -1932
rect 8822 -1932 9118 -1893
rect 8822 -1948 8882 -1932
rect 8940 -1948 9000 -1932
rect 9058 -1948 9118 -1932
rect 9758 -1932 10054 -1893
rect 9758 -1948 9818 -1932
rect 9876 -1948 9936 -1932
rect 9994 -1948 10054 -1932
rect 13401 -1752 13461 -1737
rect 13519 -1752 13579 -1737
rect 13637 -1752 13697 -1737
rect 13868 -1737 14164 -1698
rect 13868 -1752 13928 -1737
rect 13986 -1752 14046 -1737
rect 14104 -1752 14164 -1737
rect 14222 -1737 14518 -1698
rect 14222 -1752 14282 -1737
rect 14340 -1752 14400 -1737
rect 14458 -1752 14518 -1737
rect 14695 -1737 14991 -1698
rect 14695 -1752 14755 -1737
rect 14813 -1752 14873 -1737
rect 14931 -1752 14991 -1737
rect 16545 -1737 16841 -1698
rect 16545 -1752 16605 -1737
rect 16663 -1752 16723 -1737
rect 16781 -1752 16841 -1737
rect 17012 -1737 17308 -1698
rect 17012 -1752 17072 -1737
rect 17130 -1752 17190 -1737
rect 17248 -1752 17308 -1737
rect 17366 -1737 17662 -1698
rect 17366 -1752 17426 -1737
rect 17484 -1752 17544 -1737
rect 17602 -1752 17662 -1737
rect 17839 -1737 18135 -1698
rect 17839 -1752 17899 -1737
rect 17957 -1752 18017 -1737
rect 18075 -1752 18135 -1737
rect 19677 -1733 19973 -1694
rect 19677 -1748 19737 -1733
rect 19795 -1748 19855 -1733
rect 19913 -1748 19973 -1733
rect 20144 -1733 20440 -1694
rect 20144 -1748 20204 -1733
rect 20262 -1748 20322 -1733
rect 20380 -1748 20440 -1733
rect 20498 -1733 20794 -1694
rect 20498 -1748 20558 -1733
rect 20616 -1748 20676 -1733
rect 20734 -1748 20794 -1733
rect 20971 -1733 21267 -1694
rect 20971 -1748 21031 -1733
rect 21089 -1748 21149 -1733
rect 21207 -1748 21267 -1733
rect 22821 -1733 23117 -1694
rect 22821 -1748 22881 -1733
rect 22939 -1748 22999 -1733
rect 23057 -1748 23117 -1733
rect 23288 -1733 23584 -1694
rect 23288 -1748 23348 -1733
rect 23406 -1748 23466 -1733
rect 23524 -1748 23584 -1733
rect 23642 -1733 23938 -1694
rect 23642 -1748 23702 -1733
rect 23760 -1748 23820 -1733
rect 23878 -1748 23938 -1733
rect 24115 -1733 24411 -1694
rect 24115 -1748 24175 -1733
rect 24233 -1748 24293 -1733
rect 24351 -1748 24411 -1733
rect 11966 -1932 12262 -1893
rect 11966 -1948 12026 -1932
rect 12084 -1948 12144 -1932
rect 12202 -1948 12262 -1932
rect 12960 -1936 13256 -1897
rect 12960 -1952 13020 -1936
rect 13078 -1952 13138 -1936
rect 13196 -1952 13256 -1936
rect 338 -2438 398 -2152
rect 456 -2178 516 -2152
rect 574 -2178 634 -2152
rect 779 -2178 839 -2152
rect 338 -2455 474 -2438
rect 338 -2510 397 -2455
rect 455 -2510 474 -2455
rect 338 -2525 474 -2510
rect 338 -2837 398 -2525
rect 897 -2570 957 -2152
rect 1015 -2178 1075 -2152
rect 1246 -2178 1306 -2152
rect 1364 -2178 1424 -2152
rect 1482 -2178 1542 -2152
rect 1600 -2178 1660 -2152
rect 1365 -2338 1424 -2178
rect 1365 -2339 1428 -2338
rect 1362 -2355 1428 -2339
rect 1362 -2389 1378 -2355
rect 1412 -2389 1428 -2355
rect 1362 -2405 1428 -2389
rect 1465 -2454 1560 -2439
rect 1465 -2509 1484 -2454
rect 1542 -2477 1560 -2454
rect 1718 -2477 1778 -2152
rect 1836 -2178 1896 -2152
rect 2073 -2178 2133 -2152
rect 1542 -2509 1778 -2477
rect 1465 -2526 1778 -2509
rect 897 -2627 1424 -2570
rect 1364 -2726 1424 -2627
rect 1353 -2739 1434 -2726
rect 1353 -2794 1366 -2739
rect 1424 -2794 1434 -2739
rect 1353 -2805 1434 -2794
rect 338 -2882 1232 -2837
rect 1172 -3085 1232 -2882
rect 1364 -3085 1424 -2805
rect 1482 -3085 1542 -2526
rect 2191 -2568 2251 -2152
rect 2309 -2178 2369 -2152
rect 2546 -2178 2606 -2152
rect 2664 -2178 2724 -2152
rect 2672 -2301 2738 -2298
rect 2782 -2301 2842 -2152
rect 2672 -2314 2842 -2301
rect 2672 -2348 2688 -2314
rect 2722 -2348 2842 -2314
rect 2672 -2361 2842 -2348
rect 2672 -2364 2738 -2361
rect 1713 -2585 2251 -2568
rect 1713 -2619 1732 -2585
rect 1766 -2619 2251 -2585
rect 1713 -2625 2251 -2619
rect 1713 -2635 1782 -2625
rect 1713 -2637 1778 -2635
rect 1597 -2975 1663 -2959
rect 1597 -3009 1613 -2975
rect 1647 -3009 1663 -2975
rect 1597 -3025 1663 -3009
rect 1600 -3085 1660 -3025
rect 1718 -3085 1778 -2637
rect 2782 -2837 2842 -2361
rect 1914 -2882 2842 -2837
rect 3482 -2438 3542 -2152
rect 3600 -2178 3660 -2152
rect 3718 -2178 3778 -2152
rect 3923 -2178 3983 -2152
rect 3482 -2455 3618 -2438
rect 3482 -2510 3541 -2455
rect 3599 -2510 3618 -2455
rect 3482 -2525 3618 -2510
rect 3482 -2837 3542 -2525
rect 4041 -2570 4101 -2152
rect 4159 -2178 4219 -2152
rect 4390 -2178 4450 -2152
rect 4508 -2178 4568 -2152
rect 4626 -2178 4686 -2152
rect 4744 -2178 4804 -2152
rect 4509 -2338 4568 -2178
rect 4509 -2339 4572 -2338
rect 4506 -2355 4572 -2339
rect 4506 -2389 4522 -2355
rect 4556 -2389 4572 -2355
rect 4506 -2405 4572 -2389
rect 4609 -2454 4704 -2439
rect 4609 -2509 4628 -2454
rect 4686 -2477 4704 -2454
rect 4862 -2477 4922 -2152
rect 4980 -2178 5040 -2152
rect 5217 -2178 5277 -2152
rect 4686 -2509 4922 -2477
rect 4609 -2526 4922 -2509
rect 4041 -2627 4568 -2570
rect 4508 -2726 4568 -2627
rect 4497 -2739 4578 -2726
rect 4497 -2794 4510 -2739
rect 4568 -2794 4578 -2739
rect 4497 -2805 4578 -2794
rect 3482 -2882 4376 -2837
rect 1914 -3085 1974 -2882
rect 4316 -3085 4376 -2882
rect 4508 -3085 4568 -2805
rect 4626 -3085 4686 -2526
rect 5335 -2568 5395 -2152
rect 5453 -2178 5513 -2152
rect 5690 -2178 5750 -2152
rect 5808 -2178 5868 -2152
rect 5816 -2301 5882 -2298
rect 5926 -2301 5986 -2152
rect 5816 -2314 5986 -2301
rect 5816 -2348 5832 -2314
rect 5866 -2348 5986 -2314
rect 5816 -2361 5986 -2348
rect 5816 -2364 5882 -2361
rect 4857 -2585 5395 -2568
rect 4857 -2619 4876 -2585
rect 4910 -2619 5395 -2585
rect 4857 -2625 5395 -2619
rect 4857 -2635 4926 -2625
rect 4857 -2637 4922 -2635
rect 4741 -2975 4807 -2959
rect 4741 -3009 4757 -2975
rect 4791 -3009 4807 -2975
rect 4741 -3025 4807 -3009
rect 4744 -3085 4804 -3025
rect 4862 -3085 4922 -2637
rect 5926 -2837 5986 -2361
rect 5058 -2882 5986 -2837
rect 6614 -2434 6674 -2148
rect 6732 -2174 6792 -2148
rect 6850 -2174 6910 -2148
rect 7055 -2174 7115 -2148
rect 6614 -2451 6750 -2434
rect 6614 -2506 6673 -2451
rect 6731 -2506 6750 -2451
rect 6614 -2521 6750 -2506
rect 6614 -2833 6674 -2521
rect 7173 -2566 7233 -2148
rect 7291 -2174 7351 -2148
rect 7522 -2174 7582 -2148
rect 7640 -2174 7700 -2148
rect 7758 -2174 7818 -2148
rect 7876 -2174 7936 -2148
rect 7641 -2334 7700 -2174
rect 7641 -2335 7704 -2334
rect 7638 -2351 7704 -2335
rect 7638 -2385 7654 -2351
rect 7688 -2385 7704 -2351
rect 7638 -2401 7704 -2385
rect 7741 -2450 7836 -2435
rect 7741 -2505 7760 -2450
rect 7818 -2473 7836 -2450
rect 7994 -2473 8054 -2148
rect 8112 -2174 8172 -2148
rect 8349 -2174 8409 -2148
rect 7818 -2505 8054 -2473
rect 7741 -2522 8054 -2505
rect 7173 -2623 7700 -2566
rect 7640 -2722 7700 -2623
rect 7629 -2735 7710 -2722
rect 7629 -2790 7642 -2735
rect 7700 -2790 7710 -2735
rect 7629 -2801 7710 -2790
rect 6614 -2878 7508 -2833
rect 5058 -3085 5118 -2882
rect 7448 -3081 7508 -2878
rect 7640 -3081 7700 -2801
rect 7758 -3081 7818 -2522
rect 8467 -2564 8527 -2148
rect 8585 -2174 8645 -2148
rect 8822 -2174 8882 -2148
rect 8940 -2174 9000 -2148
rect 8948 -2297 9014 -2294
rect 9058 -2297 9118 -2148
rect 8948 -2310 9118 -2297
rect 8948 -2344 8964 -2310
rect 8998 -2344 9118 -2310
rect 8948 -2357 9118 -2344
rect 8948 -2360 9014 -2357
rect 7989 -2581 8527 -2564
rect 7989 -2615 8008 -2581
rect 8042 -2615 8527 -2581
rect 7989 -2621 8527 -2615
rect 7989 -2631 8058 -2621
rect 7989 -2633 8054 -2631
rect 7873 -2971 7939 -2955
rect 7873 -3005 7889 -2971
rect 7923 -3005 7939 -2971
rect 7873 -3021 7939 -3005
rect 7876 -3081 7936 -3021
rect 7994 -3081 8054 -2633
rect 9058 -2833 9118 -2357
rect 8190 -2878 9118 -2833
rect 9758 -2434 9818 -2148
rect 9876 -2174 9936 -2148
rect 9994 -2174 10054 -2148
rect 10199 -2174 10259 -2148
rect 9758 -2451 9894 -2434
rect 9758 -2506 9817 -2451
rect 9875 -2506 9894 -2451
rect 9758 -2521 9894 -2506
rect 9758 -2833 9818 -2521
rect 10317 -2566 10377 -2148
rect 10435 -2174 10495 -2148
rect 10666 -2174 10726 -2148
rect 10784 -2174 10844 -2148
rect 10902 -2174 10962 -2148
rect 11020 -2174 11080 -2148
rect 10785 -2334 10844 -2174
rect 10785 -2335 10848 -2334
rect 10782 -2351 10848 -2335
rect 10782 -2385 10798 -2351
rect 10832 -2385 10848 -2351
rect 10782 -2401 10848 -2385
rect 10885 -2450 10980 -2435
rect 10885 -2505 10904 -2450
rect 10962 -2473 10980 -2450
rect 11138 -2473 11198 -2148
rect 11256 -2174 11316 -2148
rect 11493 -2174 11553 -2148
rect 10962 -2505 11198 -2473
rect 10885 -2522 11198 -2505
rect 10317 -2623 10844 -2566
rect 10784 -2722 10844 -2623
rect 10773 -2735 10854 -2722
rect 10773 -2790 10786 -2735
rect 10844 -2790 10854 -2735
rect 10773 -2801 10854 -2790
rect 9758 -2878 10652 -2833
rect 8190 -3081 8250 -2878
rect 10592 -3081 10652 -2878
rect 10784 -3081 10844 -2801
rect 10902 -3081 10962 -2522
rect 11611 -2564 11671 -2148
rect 11729 -2174 11789 -2148
rect 11966 -2174 12026 -2148
rect 12084 -2174 12144 -2148
rect 12092 -2297 12158 -2294
rect 12202 -2297 12262 -2148
rect 15168 -1936 15464 -1897
rect 15168 -1952 15228 -1936
rect 15286 -1952 15346 -1936
rect 15404 -1952 15464 -1936
rect 16104 -1936 16400 -1897
rect 16104 -1952 16164 -1936
rect 16222 -1952 16282 -1936
rect 16340 -1952 16400 -1936
rect 18312 -1936 18608 -1897
rect 18312 -1952 18372 -1936
rect 18430 -1952 18490 -1936
rect 18548 -1952 18608 -1936
rect 19236 -1932 19532 -1893
rect 19236 -1948 19296 -1932
rect 19354 -1948 19414 -1932
rect 19472 -1948 19532 -1932
rect 21444 -1932 21740 -1893
rect 21444 -1948 21504 -1932
rect 21562 -1948 21622 -1932
rect 21680 -1948 21740 -1932
rect 22380 -1932 22676 -1893
rect 22380 -1948 22440 -1932
rect 22498 -1948 22558 -1932
rect 22616 -1948 22676 -1932
rect 30367 -1841 30418 -1653
rect 31203 -1768 31269 -1752
rect 54854 -1562 54914 -1536
rect 54972 -1562 55032 -1536
rect 55090 -1562 55150 -1536
rect 55208 -1542 55269 -1536
rect 55208 -1562 55268 -1542
rect 55326 -1562 55386 -1536
rect 55444 -1562 55504 -1536
rect 55562 -1562 55622 -1530
rect 55680 -1562 55740 -1536
rect 55798 -1562 55858 -1536
rect 24588 -1932 24884 -1893
rect 24588 -1948 24648 -1932
rect 24706 -1948 24766 -1932
rect 24824 -1948 24884 -1932
rect 29884 -1901 29950 -1841
rect 30350 -1901 30418 -1841
rect 30560 -1844 30643 -1784
rect 31043 -1844 31069 -1784
rect 31203 -1802 31219 -1768
rect 31253 -1802 31269 -1768
rect 31203 -1819 31269 -1802
rect 41651 -1776 41711 -1755
rect 41769 -1776 41829 -1755
rect 41887 -1776 41947 -1755
rect 41651 -1812 41947 -1776
rect 42005 -1775 42065 -1755
rect 42123 -1775 42183 -1755
rect 42241 -1775 42301 -1755
rect 42005 -1811 42301 -1775
rect 42359 -1775 42419 -1755
rect 42477 -1775 42537 -1755
rect 42595 -1775 42655 -1755
rect 42359 -1811 42655 -1775
rect 48205 -1771 48265 -1750
rect 48323 -1771 48383 -1750
rect 48441 -1771 48501 -1750
rect 48205 -1807 48501 -1771
rect 48559 -1770 48619 -1750
rect 48677 -1770 48737 -1750
rect 48795 -1770 48855 -1750
rect 48559 -1806 48855 -1770
rect 48913 -1770 48973 -1750
rect 49031 -1770 49091 -1750
rect 49149 -1770 49209 -1750
rect 65407 -1457 65467 -877
rect 65709 -1256 65769 -1230
rect 65677 -1397 65744 -1390
rect 65827 -1397 65887 -1230
rect 65945 -1256 66005 -1230
rect 66063 -1256 66123 -1230
rect 65677 -1406 65887 -1397
rect 65677 -1440 65693 -1406
rect 65727 -1440 65887 -1406
rect 65677 -1456 65887 -1440
rect 65407 -1473 65558 -1457
rect 65407 -1507 65508 -1473
rect 65542 -1507 65558 -1473
rect 65407 -1523 65558 -1507
rect 65407 -1562 65467 -1523
rect 65827 -1562 65887 -1456
rect 66181 -1397 66241 -1230
rect 66299 -1256 66359 -1230
rect 66324 -1397 66391 -1390
rect 66181 -1406 66391 -1397
rect 66181 -1440 66341 -1406
rect 66375 -1440 66391 -1406
rect 66181 -1456 66391 -1440
rect 65943 -1490 66009 -1474
rect 65943 -1524 65959 -1490
rect 65993 -1524 66009 -1490
rect 65943 -1540 66009 -1524
rect 66061 -1489 66127 -1474
rect 66061 -1523 66077 -1489
rect 66111 -1523 66127 -1489
rect 66061 -1539 66127 -1523
rect 65945 -1562 66005 -1540
rect 66063 -1562 66123 -1539
rect 66181 -1562 66241 -1456
rect 66705 -1458 66765 -757
rect 67312 -777 67372 -751
rect 67430 -777 67490 -566
rect 67783 -572 67843 -540
rect 67901 -566 67961 -540
rect 68019 -566 68079 -540
rect 67780 -588 67846 -572
rect 67780 -622 67796 -588
rect 67830 -622 67846 -588
rect 67780 -638 67846 -622
rect 70455 -586 70494 -528
rect 70455 -646 70509 -586
rect 70909 -646 71384 -586
rect 67662 -705 67728 -689
rect 67662 -739 67678 -705
rect 67712 -739 67728 -705
rect 67662 -755 67728 -739
rect 70455 -704 70494 -646
rect 67665 -777 67725 -755
rect 70455 -764 70509 -704
rect 70909 -764 70935 -704
rect 67665 -1003 67725 -977
rect 70455 -995 70509 -935
rect 70909 -995 70935 -935
rect 70455 -1053 70494 -995
rect 70455 -1113 70509 -1053
rect 70909 -1054 70935 -1053
rect 71096 -1054 71162 -1051
rect 70909 -1067 71162 -1054
rect 70909 -1101 71112 -1067
rect 71146 -1101 71162 -1067
rect 70909 -1113 71162 -1101
rect 71327 -1053 71384 -646
rect 71594 -861 71639 -87
rect 71594 -921 71842 -861
rect 72042 -921 72068 -861
rect 71483 -1053 71562 -1042
rect 71327 -1055 71842 -1053
rect 71327 -1113 71496 -1055
rect 71551 -1113 71842 -1055
rect 72242 -1113 72268 -1053
rect 67312 -1199 67372 -1177
rect 67430 -1199 67490 -1177
rect 67309 -1215 67375 -1199
rect 67309 -1249 67325 -1215
rect 67359 -1249 67375 -1215
rect 67309 -1265 67375 -1249
rect 67427 -1215 67493 -1199
rect 67427 -1249 67443 -1215
rect 67477 -1249 67493 -1215
rect 67427 -1265 67493 -1249
rect 70455 -1171 70494 -1113
rect 71095 -1117 71162 -1113
rect 71483 -1123 71562 -1113
rect 71196 -1171 71283 -1154
rect 70455 -1231 70509 -1171
rect 70909 -1231 70935 -1171
rect 71196 -1173 71842 -1171
rect 71196 -1231 71211 -1173
rect 71266 -1231 71842 -1173
rect 72242 -1231 72268 -1171
rect 71196 -1249 71283 -1231
rect 70455 -1349 70509 -1289
rect 70909 -1349 70935 -1289
rect 70455 -1407 70494 -1349
rect 71234 -1407 71283 -1249
rect 71716 -1289 71782 -1286
rect 72315 -1244 72381 -1228
rect 72315 -1278 72331 -1244
rect 72365 -1278 72381 -1244
rect 71716 -1302 71842 -1289
rect 71716 -1336 71732 -1302
rect 71766 -1336 71842 -1302
rect 71716 -1349 71842 -1336
rect 72242 -1349 72268 -1289
rect 72315 -1294 72381 -1278
rect 71716 -1352 71782 -1349
rect 66615 -1474 66765 -1458
rect 66615 -1508 66631 -1474
rect 66665 -1508 66765 -1474
rect 66615 -1524 66765 -1508
rect 66705 -1562 66765 -1524
rect 70455 -1467 70509 -1407
rect 70909 -1467 71283 -1407
rect 71325 -1407 71394 -1402
rect 71325 -1421 71842 -1407
rect 71325 -1455 71342 -1421
rect 71376 -1455 71842 -1421
rect 71325 -1467 71842 -1455
rect 72242 -1467 72268 -1407
rect 70455 -1525 70494 -1467
rect 71325 -1471 71392 -1467
rect 63542 -1663 63602 -1637
rect 63660 -1663 63720 -1637
rect 63778 -1663 63838 -1637
rect 63896 -1657 63956 -1637
rect 63896 -1663 63957 -1657
rect 64014 -1663 64074 -1637
rect 64132 -1663 64192 -1637
rect 48913 -1806 49209 -1770
rect 54854 -1783 54914 -1762
rect 54972 -1783 55032 -1762
rect 55090 -1783 55150 -1762
rect 54854 -1819 55150 -1783
rect 55208 -1782 55268 -1762
rect 55326 -1782 55386 -1762
rect 55444 -1782 55504 -1762
rect 55208 -1818 55504 -1782
rect 55562 -1782 55622 -1762
rect 55680 -1782 55740 -1762
rect 55798 -1782 55858 -1762
rect 55562 -1818 55858 -1782
rect 29884 -1959 29935 -1901
rect 30560 -1902 30620 -1844
rect 31210 -1902 31269 -1819
rect 63779 -1848 63837 -1663
rect 63779 -1874 63839 -1848
rect 63897 -1874 63957 -1663
rect 64250 -1669 64310 -1637
rect 64368 -1663 64428 -1637
rect 64486 -1663 64546 -1637
rect 64247 -1685 64313 -1669
rect 64247 -1719 64263 -1685
rect 64297 -1719 64313 -1685
rect 64247 -1735 64313 -1719
rect 64129 -1802 64195 -1786
rect 65407 -1788 65467 -1762
rect 64129 -1836 64145 -1802
rect 64179 -1836 64195 -1802
rect 64129 -1852 64195 -1836
rect 64132 -1874 64192 -1852
rect 12092 -2310 12262 -2297
rect 12092 -2344 12108 -2310
rect 12142 -2344 12262 -2310
rect 12092 -2357 12262 -2344
rect 12092 -2360 12158 -2357
rect 11133 -2581 11671 -2564
rect 11133 -2615 11152 -2581
rect 11186 -2615 11671 -2581
rect 11133 -2621 11671 -2615
rect 11133 -2631 11202 -2621
rect 11133 -2633 11198 -2631
rect 11017 -2971 11083 -2955
rect 11017 -3005 11033 -2971
rect 11067 -3005 11083 -2971
rect 11017 -3021 11083 -3005
rect 11020 -3081 11080 -3021
rect 11138 -3081 11198 -2633
rect 12202 -2833 12262 -2357
rect 11334 -2878 12262 -2833
rect 12960 -2438 13020 -2152
rect 13078 -2178 13138 -2152
rect 13196 -2178 13256 -2152
rect 13401 -2178 13461 -2152
rect 12960 -2455 13096 -2438
rect 12960 -2510 13019 -2455
rect 13077 -2510 13096 -2455
rect 12960 -2525 13096 -2510
rect 12960 -2837 13020 -2525
rect 13519 -2570 13579 -2152
rect 13637 -2178 13697 -2152
rect 13868 -2178 13928 -2152
rect 13986 -2178 14046 -2152
rect 14104 -2178 14164 -2152
rect 14222 -2178 14282 -2152
rect 13987 -2338 14046 -2178
rect 13987 -2339 14050 -2338
rect 13984 -2355 14050 -2339
rect 13984 -2389 14000 -2355
rect 14034 -2389 14050 -2355
rect 13984 -2405 14050 -2389
rect 14087 -2454 14182 -2439
rect 14087 -2509 14106 -2454
rect 14164 -2477 14182 -2454
rect 14340 -2477 14400 -2152
rect 14458 -2178 14518 -2152
rect 14695 -2178 14755 -2152
rect 14164 -2509 14400 -2477
rect 14087 -2526 14400 -2509
rect 13519 -2627 14046 -2570
rect 13986 -2726 14046 -2627
rect 13975 -2739 14056 -2726
rect 13975 -2794 13988 -2739
rect 14046 -2794 14056 -2739
rect 13975 -2805 14056 -2794
rect 11334 -3081 11394 -2878
rect 12960 -2882 13854 -2837
rect 1172 -3311 1232 -3285
rect 1364 -3511 1424 -3485
rect 1482 -3511 1542 -3485
rect 1600 -3511 1660 -3485
rect 1718 -3511 1778 -3485
rect 1539 -3566 1605 -3558
rect 1914 -3566 1974 -3285
rect 4316 -3311 4376 -3285
rect 4508 -3511 4568 -3485
rect 4626 -3511 4686 -3485
rect 4744 -3511 4804 -3485
rect 4862 -3511 4922 -3485
rect 1539 -3574 1974 -3566
rect 1539 -3608 1555 -3574
rect 1589 -3608 1974 -3574
rect 1539 -3617 1974 -3608
rect 4683 -3566 4749 -3558
rect 5058 -3566 5118 -3285
rect 7448 -3307 7508 -3281
rect 7640 -3507 7700 -3481
rect 7758 -3507 7818 -3481
rect 7876 -3507 7936 -3481
rect 7994 -3507 8054 -3481
rect 4683 -3574 5118 -3566
rect 4683 -3608 4699 -3574
rect 4733 -3608 5118 -3574
rect 4683 -3617 5118 -3608
rect 7815 -3562 7881 -3554
rect 8190 -3562 8250 -3281
rect 10592 -3307 10652 -3281
rect 13794 -3085 13854 -2882
rect 13986 -3085 14046 -2805
rect 14104 -3085 14164 -2526
rect 14813 -2568 14873 -2152
rect 14931 -2178 14991 -2152
rect 15168 -2178 15228 -2152
rect 15286 -2178 15346 -2152
rect 15294 -2301 15360 -2298
rect 15404 -2301 15464 -2152
rect 15294 -2314 15464 -2301
rect 15294 -2348 15310 -2314
rect 15344 -2348 15464 -2314
rect 15294 -2361 15464 -2348
rect 15294 -2364 15360 -2361
rect 14335 -2585 14873 -2568
rect 14335 -2619 14354 -2585
rect 14388 -2619 14873 -2585
rect 14335 -2625 14873 -2619
rect 14335 -2635 14404 -2625
rect 14335 -2637 14400 -2635
rect 14219 -2975 14285 -2959
rect 14219 -3009 14235 -2975
rect 14269 -3009 14285 -2975
rect 14219 -3025 14285 -3009
rect 14222 -3085 14282 -3025
rect 14340 -3085 14400 -2637
rect 15404 -2837 15464 -2361
rect 14536 -2882 15464 -2837
rect 16104 -2438 16164 -2152
rect 16222 -2178 16282 -2152
rect 16340 -2178 16400 -2152
rect 16545 -2178 16605 -2152
rect 16104 -2455 16240 -2438
rect 16104 -2510 16163 -2455
rect 16221 -2510 16240 -2455
rect 16104 -2525 16240 -2510
rect 16104 -2837 16164 -2525
rect 16663 -2570 16723 -2152
rect 16781 -2178 16841 -2152
rect 17012 -2178 17072 -2152
rect 17130 -2178 17190 -2152
rect 17248 -2178 17308 -2152
rect 17366 -2178 17426 -2152
rect 17131 -2338 17190 -2178
rect 17131 -2339 17194 -2338
rect 17128 -2355 17194 -2339
rect 17128 -2389 17144 -2355
rect 17178 -2389 17194 -2355
rect 17128 -2405 17194 -2389
rect 17231 -2454 17326 -2439
rect 17231 -2509 17250 -2454
rect 17308 -2477 17326 -2454
rect 17484 -2477 17544 -2152
rect 17602 -2178 17662 -2152
rect 17839 -2178 17899 -2152
rect 17308 -2509 17544 -2477
rect 17231 -2526 17544 -2509
rect 16663 -2627 17190 -2570
rect 17130 -2726 17190 -2627
rect 17119 -2739 17200 -2726
rect 17119 -2794 17132 -2739
rect 17190 -2794 17200 -2739
rect 17119 -2805 17200 -2794
rect 16104 -2882 16998 -2837
rect 14536 -3085 14596 -2882
rect 16938 -3085 16998 -2882
rect 17130 -3085 17190 -2805
rect 17248 -3085 17308 -2526
rect 17957 -2568 18017 -2152
rect 18075 -2178 18135 -2152
rect 18312 -2178 18372 -2152
rect 18430 -2178 18490 -2152
rect 18438 -2301 18504 -2298
rect 18548 -2301 18608 -2152
rect 18438 -2314 18608 -2301
rect 18438 -2348 18454 -2314
rect 18488 -2348 18608 -2314
rect 18438 -2361 18608 -2348
rect 18438 -2364 18504 -2361
rect 17479 -2585 18017 -2568
rect 17479 -2619 17498 -2585
rect 17532 -2619 18017 -2585
rect 17479 -2625 18017 -2619
rect 17479 -2635 17548 -2625
rect 17479 -2637 17544 -2635
rect 17363 -2975 17429 -2959
rect 17363 -3009 17379 -2975
rect 17413 -3009 17429 -2975
rect 17363 -3025 17429 -3009
rect 17366 -3085 17426 -3025
rect 17484 -3085 17544 -2637
rect 18548 -2837 18608 -2361
rect 17680 -2882 18608 -2837
rect 19236 -2434 19296 -2148
rect 19354 -2174 19414 -2148
rect 19472 -2174 19532 -2148
rect 19677 -2174 19737 -2148
rect 19236 -2451 19372 -2434
rect 19236 -2506 19295 -2451
rect 19353 -2506 19372 -2451
rect 19236 -2521 19372 -2506
rect 19236 -2833 19296 -2521
rect 19795 -2566 19855 -2148
rect 19913 -2174 19973 -2148
rect 20144 -2174 20204 -2148
rect 20262 -2174 20322 -2148
rect 20380 -2174 20440 -2148
rect 20498 -2174 20558 -2148
rect 20263 -2334 20322 -2174
rect 20263 -2335 20326 -2334
rect 20260 -2351 20326 -2335
rect 20260 -2385 20276 -2351
rect 20310 -2385 20326 -2351
rect 20260 -2401 20326 -2385
rect 20363 -2450 20458 -2435
rect 20363 -2505 20382 -2450
rect 20440 -2473 20458 -2450
rect 20616 -2473 20676 -2148
rect 20734 -2174 20794 -2148
rect 20971 -2174 21031 -2148
rect 20440 -2505 20676 -2473
rect 20363 -2522 20676 -2505
rect 19795 -2623 20322 -2566
rect 20262 -2722 20322 -2623
rect 20251 -2735 20332 -2722
rect 20251 -2790 20264 -2735
rect 20322 -2790 20332 -2735
rect 20251 -2801 20332 -2790
rect 19236 -2878 20130 -2833
rect 17680 -3085 17740 -2882
rect 20070 -3081 20130 -2878
rect 20262 -3081 20322 -2801
rect 20380 -3081 20440 -2522
rect 21089 -2564 21149 -2148
rect 21207 -2174 21267 -2148
rect 21444 -2174 21504 -2148
rect 21562 -2174 21622 -2148
rect 21570 -2297 21636 -2294
rect 21680 -2297 21740 -2148
rect 21570 -2310 21740 -2297
rect 21570 -2344 21586 -2310
rect 21620 -2344 21740 -2310
rect 21570 -2357 21740 -2344
rect 21570 -2360 21636 -2357
rect 20611 -2581 21149 -2564
rect 20611 -2615 20630 -2581
rect 20664 -2615 21149 -2581
rect 20611 -2621 21149 -2615
rect 20611 -2631 20680 -2621
rect 20611 -2633 20676 -2631
rect 20495 -2971 20561 -2955
rect 20495 -3005 20511 -2971
rect 20545 -3005 20561 -2971
rect 20495 -3021 20561 -3005
rect 20498 -3081 20558 -3021
rect 20616 -3081 20676 -2633
rect 21680 -2833 21740 -2357
rect 20812 -2878 21740 -2833
rect 22380 -2434 22440 -2148
rect 22498 -2174 22558 -2148
rect 22616 -2174 22676 -2148
rect 22821 -2174 22881 -2148
rect 22380 -2451 22516 -2434
rect 22380 -2506 22439 -2451
rect 22497 -2506 22516 -2451
rect 22380 -2521 22516 -2506
rect 22380 -2833 22440 -2521
rect 22939 -2566 22999 -2148
rect 23057 -2174 23117 -2148
rect 23288 -2174 23348 -2148
rect 23406 -2174 23466 -2148
rect 23524 -2174 23584 -2148
rect 23642 -2174 23702 -2148
rect 23407 -2334 23466 -2174
rect 23407 -2335 23470 -2334
rect 23404 -2351 23470 -2335
rect 23404 -2385 23420 -2351
rect 23454 -2385 23470 -2351
rect 23404 -2401 23470 -2385
rect 23507 -2450 23602 -2435
rect 23507 -2505 23526 -2450
rect 23584 -2473 23602 -2450
rect 23760 -2473 23820 -2148
rect 23878 -2174 23938 -2148
rect 24115 -2174 24175 -2148
rect 23584 -2505 23820 -2473
rect 23507 -2522 23820 -2505
rect 22939 -2623 23466 -2566
rect 23406 -2722 23466 -2623
rect 23395 -2735 23476 -2722
rect 23395 -2790 23408 -2735
rect 23466 -2790 23476 -2735
rect 23395 -2801 23476 -2790
rect 22380 -2878 23274 -2833
rect 20812 -3081 20872 -2878
rect 23214 -3081 23274 -2878
rect 23406 -3081 23466 -2801
rect 23524 -3081 23584 -2522
rect 24233 -2564 24293 -2148
rect 24351 -2174 24411 -2148
rect 24588 -2174 24648 -2148
rect 24706 -2174 24766 -2148
rect 24714 -2297 24780 -2294
rect 24824 -2297 24884 -2148
rect 24714 -2310 24884 -2297
rect 24714 -2344 24730 -2310
rect 24764 -2344 24884 -2310
rect 24714 -2357 24884 -2344
rect 24714 -2360 24780 -2357
rect 23755 -2581 24293 -2564
rect 23755 -2615 23774 -2581
rect 23808 -2615 24293 -2581
rect 23755 -2621 24293 -2615
rect 23755 -2631 23824 -2621
rect 23755 -2633 23820 -2631
rect 23639 -2971 23705 -2955
rect 23639 -3005 23655 -2971
rect 23689 -3005 23705 -2971
rect 23639 -3021 23705 -3005
rect 23642 -3081 23702 -3021
rect 23760 -3081 23820 -2633
rect 24824 -2833 24884 -2357
rect 29884 -2019 29950 -1959
rect 30350 -2019 30376 -1959
rect 30560 -1962 30643 -1902
rect 31043 -1962 31375 -1902
rect 31775 -1962 31801 -1902
rect 29884 -2077 29935 -2019
rect 30560 -2020 30620 -1962
rect 31287 -2020 31353 -2018
rect 29884 -2137 29950 -2077
rect 30350 -2137 30376 -2077
rect 30560 -2080 30643 -2020
rect 31043 -2080 31069 -2020
rect 31287 -2034 31375 -2020
rect 31287 -2068 31303 -2034
rect 31337 -2068 31375 -2034
rect 31287 -2080 31375 -2068
rect 31775 -2080 31801 -2020
rect 31287 -2084 31353 -2080
rect 31287 -2138 31352 -2136
rect 29924 -2255 29950 -2195
rect 30350 -2255 30420 -2195
rect 30369 -2313 30420 -2255
rect 29924 -2373 29950 -2313
rect 30350 -2373 30420 -2313
rect 30369 -2431 30420 -2373
rect 29924 -2491 29950 -2431
rect 30350 -2491 30420 -2431
rect 30559 -2198 30643 -2138
rect 31043 -2198 31069 -2138
rect 31287 -2152 31375 -2138
rect 31287 -2186 31302 -2152
rect 31336 -2186 31375 -2152
rect 31287 -2198 31375 -2186
rect 31775 -2198 31801 -2138
rect 30559 -2256 30619 -2198
rect 31287 -2202 31352 -2198
rect 30559 -2316 30643 -2256
rect 31043 -2316 31375 -2256
rect 31775 -2316 31801 -2256
rect 70455 -1585 70509 -1525
rect 70909 -1585 70935 -1525
rect 66705 -1788 66765 -1762
rect 70455 -1822 70509 -1762
rect 70909 -1822 70935 -1762
rect 70455 -1880 70494 -1822
rect 71325 -1880 71382 -1471
rect 72323 -1603 72374 -1294
rect 70455 -1940 70509 -1880
rect 70909 -1940 71382 -1880
rect 71594 -1663 71842 -1603
rect 72042 -1663 72374 -1603
rect 65827 -1988 65887 -1962
rect 65945 -1988 66005 -1962
rect 66063 -1988 66123 -1962
rect 66181 -1988 66241 -1962
rect 70455 -1998 70494 -1940
rect 70455 -2058 70509 -1998
rect 70909 -2058 70935 -1998
rect 64132 -2100 64192 -2074
rect 63779 -2296 63839 -2274
rect 63897 -2296 63957 -2274
rect 70654 -2295 70709 -2235
rect 70909 -2295 70935 -2235
rect 63776 -2312 63842 -2296
rect 30559 -2374 30619 -2316
rect 30559 -2434 30643 -2374
rect 31043 -2434 31069 -2374
rect 31210 -2399 31269 -2316
rect 63776 -2346 63792 -2312
rect 63826 -2346 63842 -2312
rect 63776 -2362 63842 -2346
rect 63894 -2312 63960 -2296
rect 63894 -2346 63910 -2312
rect 63944 -2346 63960 -2312
rect 63894 -2362 63960 -2346
rect 70654 -2353 70693 -2295
rect 31203 -2416 31269 -2399
rect 30369 -2678 30420 -2491
rect 31203 -2450 31219 -2416
rect 31253 -2450 31269 -2416
rect 31203 -2466 31269 -2450
rect 70654 -2413 70709 -2353
rect 70909 -2413 70935 -2353
rect 71055 -2377 71121 -2361
rect 71055 -2411 71071 -2377
rect 71105 -2411 71121 -2377
rect 70654 -2471 70693 -2413
rect 71055 -2427 71121 -2411
rect 71058 -2471 71118 -2427
rect 71594 -2471 71639 -1663
rect 70654 -2531 70709 -2471
rect 70909 -2531 71639 -2471
rect 23956 -2878 24884 -2833
rect 30082 -2738 30150 -2678
rect 30350 -2738 30420 -2678
rect 31271 -2706 31337 -2690
rect 30507 -2728 30561 -2712
rect 30082 -2796 30133 -2738
rect 30507 -2762 30517 -2728
rect 30551 -2762 30561 -2728
rect 30507 -2780 30561 -2762
rect 31271 -2740 31287 -2706
rect 31321 -2740 31337 -2706
rect 31271 -2780 31337 -2740
rect 30369 -2796 31375 -2780
rect 30082 -2856 30150 -2796
rect 30350 -2840 31375 -2796
rect 31575 -2840 31601 -2780
rect 30350 -2855 30420 -2840
rect 30350 -2856 30376 -2855
rect 23956 -3081 24016 -2878
rect 30082 -2914 30133 -2856
rect 30082 -2974 30150 -2914
rect 30350 -2974 30376 -2914
rect 10784 -3507 10844 -3481
rect 10902 -3507 10962 -3481
rect 11020 -3507 11080 -3481
rect 11138 -3507 11198 -3481
rect 7815 -3570 8250 -3562
rect 7815 -3604 7831 -3570
rect 7865 -3604 8250 -3570
rect 7815 -3613 8250 -3604
rect 10959 -3562 11025 -3554
rect 11334 -3562 11394 -3281
rect 13794 -3311 13854 -3285
rect 13986 -3511 14046 -3485
rect 14104 -3511 14164 -3485
rect 14222 -3511 14282 -3485
rect 14340 -3511 14400 -3485
rect 10959 -3570 11394 -3562
rect 10959 -3604 10975 -3570
rect 11009 -3604 11394 -3570
rect 10959 -3613 11394 -3604
rect 14161 -3566 14227 -3558
rect 14536 -3566 14596 -3285
rect 16938 -3311 16998 -3285
rect 17130 -3511 17190 -3485
rect 17248 -3511 17308 -3485
rect 17366 -3511 17426 -3485
rect 17484 -3511 17544 -3485
rect 14161 -3574 14596 -3566
rect 14161 -3608 14177 -3574
rect 14211 -3608 14596 -3574
rect 1539 -3624 1605 -3617
rect 4683 -3624 4749 -3617
rect 7815 -3620 7881 -3613
rect 10959 -3620 11025 -3613
rect 14161 -3617 14596 -3608
rect 17305 -3566 17371 -3558
rect 17680 -3566 17740 -3285
rect 20070 -3307 20130 -3281
rect 20262 -3507 20322 -3481
rect 20380 -3507 20440 -3481
rect 20498 -3507 20558 -3481
rect 20616 -3507 20676 -3481
rect 17305 -3574 17740 -3566
rect 17305 -3608 17321 -3574
rect 17355 -3608 17740 -3574
rect 17305 -3617 17740 -3608
rect 20437 -3562 20503 -3554
rect 20812 -3562 20872 -3281
rect 23214 -3307 23274 -3281
rect 23406 -3507 23466 -3481
rect 23524 -3507 23584 -3481
rect 23642 -3507 23702 -3481
rect 23760 -3507 23820 -3481
rect 20437 -3570 20872 -3562
rect 20437 -3604 20453 -3570
rect 20487 -3604 20872 -3570
rect 20437 -3613 20872 -3604
rect 23581 -3562 23647 -3554
rect 23956 -3562 24016 -3281
rect 23581 -3570 24016 -3562
rect 23581 -3604 23597 -3570
rect 23631 -3604 24016 -3570
rect 23581 -3613 24016 -3604
rect 14161 -3624 14227 -3617
rect 17305 -3624 17371 -3617
rect 20437 -3620 20503 -3613
rect 23581 -3620 23647 -3613
<< polycont >>
rect 41810 24735 41844 24769
rect 42940 24741 42974 24775
rect 48323 24732 48357 24766
rect 49453 24738 49487 24772
rect 41810 24617 41844 24651
rect 42940 24621 42974 24655
rect 54857 24727 54891 24761
rect 55987 24733 56021 24767
rect 48323 24614 48357 24648
rect 40367 24251 40401 24285
rect 49453 24618 49487 24652
rect 61415 24731 61449 24765
rect 62545 24737 62579 24771
rect 54857 24609 54891 24643
rect 40249 24134 40283 24168
rect 42130 23861 42164 23895
rect 46880 24248 46914 24282
rect 55987 24613 56021 24647
rect 61415 24613 61449 24647
rect 46762 24131 46796 24165
rect 43272 23865 43306 23899
rect 39896 23624 39930 23658
rect 40014 23624 40048 23658
rect 48643 23858 48677 23892
rect 53414 24243 53448 24277
rect 62545 24617 62579 24651
rect 53296 24126 53330 24160
rect 49785 23862 49819 23896
rect 46409 23621 46443 23655
rect 46527 23621 46561 23655
rect 55177 23853 55211 23887
rect 59972 24247 60006 24281
rect 59854 24130 59888 24164
rect 56319 23857 56353 23891
rect 52943 23616 52977 23650
rect 53061 23616 53095 23650
rect 61735 23857 61769 23891
rect 62877 23861 62911 23895
rect 59501 23620 59535 23654
rect 59619 23620 59653 23654
rect 40381 22601 40415 22635
rect 40263 22484 40297 22518
rect 3178 21400 3212 21434
rect 4488 21359 4522 21393
rect 4358 21239 4416 21294
rect 4134 21129 4168 21163
rect 4253 20739 4287 20773
rect 5445 21238 5503 21293
rect 4476 20954 4534 21009
rect 6322 21400 6356 21434
rect 7632 21359 7666 21393
rect 7502 21239 7560 21294
rect 7278 21129 7312 21163
rect 7397 20739 7431 20773
rect 8589 21238 8647 21293
rect 7620 20954 7678 21009
rect 9454 21396 9488 21430
rect 10764 21355 10798 21389
rect 10634 21235 10692 21290
rect 10410 21125 10444 21159
rect 4311 20140 4345 20174
rect 10529 20735 10563 20769
rect 11721 21234 11779 21289
rect 10752 20950 10810 21005
rect 12598 21396 12632 21430
rect 13908 21355 13942 21389
rect 13778 21235 13836 21290
rect 13554 21125 13588 21159
rect 13673 20735 13707 20769
rect 14865 21234 14923 21289
rect 13896 20950 13954 21005
rect 15800 21400 15834 21434
rect 17110 21359 17144 21393
rect 16980 21239 17038 21294
rect 16756 21129 16790 21163
rect 16875 20739 16909 20773
rect 18067 21238 18125 21293
rect 17098 20954 17156 21009
rect 18944 21400 18978 21434
rect 20254 21359 20288 21393
rect 20124 21239 20182 21294
rect 19900 21129 19934 21163
rect 20019 20739 20053 20773
rect 39910 21974 39944 22008
rect 40028 21974 40062 22008
rect 46894 22598 46928 22632
rect 46776 22481 46810 22515
rect 21211 21238 21269 21293
rect 20242 20954 20300 21009
rect 22076 21396 22110 21430
rect 23386 21355 23420 21389
rect 23256 21235 23314 21290
rect 23032 21125 23066 21159
rect 7455 20140 7489 20174
rect 10587 20136 10621 20170
rect 13731 20136 13765 20170
rect 16933 20140 16967 20174
rect 23151 20735 23185 20769
rect 24343 21234 24401 21289
rect 23374 20950 23432 21005
rect 25220 21396 25254 21430
rect 26530 21355 26564 21389
rect 26400 21235 26458 21290
rect 26176 21125 26210 21159
rect 26295 20735 26329 20769
rect 27487 21234 27545 21289
rect 26518 20950 26576 21005
rect 42542 21806 42576 21840
rect 41535 21163 41569 21197
rect 41350 21096 41384 21130
rect 42183 21163 42217 21197
rect 41801 21079 41835 21113
rect 41919 21080 41953 21114
rect 42473 21095 42507 21129
rect 46423 21971 46457 22005
rect 46541 21971 46575 22005
rect 53428 22593 53462 22627
rect 53310 22476 53344 22510
rect 44649 21785 44683 21819
rect 43163 21290 43197 21324
rect 43433 21163 43467 21197
rect 43248 21096 43282 21130
rect 44079 21164 44113 21198
rect 43699 21079 43733 21113
rect 43817 21080 43851 21114
rect 44371 21095 44405 21129
rect 49055 21803 49089 21837
rect 48048 21160 48082 21194
rect 47863 21093 47897 21127
rect 40376 20997 40410 21031
rect 40258 20880 40292 20914
rect 20077 20140 20111 20174
rect 23209 20136 23243 20170
rect 48696 21160 48730 21194
rect 48314 21076 48348 21110
rect 48432 21077 48466 21111
rect 48986 21092 49020 21126
rect 52957 21966 52991 22000
rect 53075 21966 53109 22000
rect 59986 22597 60020 22631
rect 59868 22480 59902 22514
rect 51162 21782 51196 21816
rect 49676 21287 49710 21321
rect 49946 21160 49980 21194
rect 49761 21093 49795 21127
rect 50592 21161 50626 21195
rect 50212 21076 50246 21110
rect 50330 21077 50364 21111
rect 50884 21092 50918 21126
rect 55589 21798 55623 21832
rect 54582 21155 54616 21189
rect 54397 21088 54431 21122
rect 46889 20994 46923 21028
rect 46771 20877 46805 20911
rect 39905 20370 39939 20404
rect 40023 20370 40057 20404
rect 55230 21155 55264 21189
rect 54848 21071 54882 21105
rect 54966 21072 55000 21106
rect 55520 21087 55554 21121
rect 59515 21970 59549 22004
rect 59633 21970 59667 22004
rect 57696 21777 57730 21811
rect 56210 21282 56244 21316
rect 56480 21155 56514 21189
rect 56295 21088 56329 21122
rect 57126 21156 57160 21190
rect 56746 21071 56780 21105
rect 56864 21072 56898 21106
rect 57418 21087 57452 21121
rect 62147 21802 62181 21836
rect 61140 21159 61174 21193
rect 60955 21092 60989 21126
rect 53423 20989 53457 21023
rect 53305 20872 53339 20906
rect 46418 20367 46452 20401
rect 46536 20367 46570 20401
rect 61788 21159 61822 21193
rect 61406 21075 61440 21109
rect 61524 21076 61558 21110
rect 62078 21091 62112 21125
rect 71216 21898 71271 21956
rect 64254 21781 64288 21815
rect 62768 21286 62802 21320
rect 63038 21159 63072 21193
rect 62853 21092 62887 21126
rect 63684 21160 63718 21194
rect 63304 21075 63338 21109
rect 63422 21076 63456 21110
rect 63976 21091 64010 21125
rect 59981 20993 60015 21027
rect 59863 20876 59897 20910
rect 26353 20136 26387 20170
rect 52952 20362 52986 20396
rect 53070 20362 53104 20396
rect 71116 20941 71150 20975
rect 71500 20929 71555 20987
rect 71215 20811 71270 20869
rect 72335 20764 72369 20798
rect 71736 20706 71770 20740
rect 71346 20587 71380 20621
rect 59510 20366 59544 20400
rect 59628 20366 59662 20400
rect 71075 19631 71109 19665
rect 40446 19133 40480 19167
rect 41576 19127 41610 19161
rect 47004 19129 47038 19163
rect 48134 19123 48168 19157
rect 40446 19013 40480 19047
rect 41576 19009 41610 19043
rect 53538 19134 53572 19168
rect 54668 19128 54702 19162
rect 47004 19009 47038 19043
rect 43019 18643 43053 18677
rect 40114 18257 40148 18291
rect 43137 18526 43171 18560
rect 48134 19005 48168 19039
rect 41256 18253 41290 18287
rect 60051 19137 60085 19171
rect 61181 19131 61215 19165
rect 53538 19014 53572 19048
rect 49577 18639 49611 18673
rect 46672 18253 46706 18287
rect 49695 18522 49729 18556
rect 54668 19010 54702 19044
rect 47814 18249 47848 18283
rect 43372 18016 43406 18050
rect 43490 18016 43524 18050
rect 60051 19017 60085 19051
rect 56111 18644 56145 18678
rect 53206 18258 53240 18292
rect 56229 18527 56263 18561
rect 61181 19013 61215 19047
rect 54348 18254 54382 18288
rect 49930 18012 49964 18046
rect 50048 18012 50082 18046
rect 71216 18754 71271 18812
rect 62624 18647 62658 18681
rect 59719 18261 59753 18295
rect 62742 18530 62776 18564
rect 60861 18257 60895 18291
rect 56464 18017 56498 18051
rect 56582 18017 56616 18051
rect 62977 18020 63011 18054
rect 63095 18020 63129 18054
rect 71116 17797 71150 17831
rect 71500 17785 71555 17843
rect 71215 17667 71270 17725
rect 72335 17620 72369 17654
rect 71736 17562 71770 17596
rect 71346 17443 71380 17477
rect 5318 16936 5352 16970
rect 6486 16936 6520 16970
rect 7654 16936 7688 16970
rect 8822 16936 8856 16970
rect 9996 16934 10030 16968
rect 5318 16828 5352 16862
rect 6486 16828 6520 16862
rect 7654 16828 7688 16862
rect 11164 16934 11198 16968
rect 12332 16934 12366 16968
rect 43005 16993 43039 17027
rect 13500 16934 13534 16968
rect 8822 16828 8856 16862
rect 5023 16065 5057 16099
rect 9996 16826 10030 16860
rect 6191 16065 6225 16099
rect 7359 16065 7393 16099
rect 11164 16826 11198 16860
rect 12332 16826 12366 16860
rect 13500 16826 13534 16860
rect 8527 16065 8561 16099
rect 43123 16876 43157 16910
rect 9701 16063 9735 16097
rect 10869 16063 10903 16097
rect 12037 16063 12071 16097
rect 14098 16331 14132 16365
rect 13205 16063 13239 16097
rect 14216 16214 14250 16248
rect 15546 16331 15580 16365
rect 15664 16214 15698 16248
rect 17044 16329 17078 16363
rect 17162 16212 17196 16246
rect 18492 16329 18526 16363
rect 18610 16212 18644 16246
rect 20012 16331 20046 16365
rect 20130 16214 20164 16248
rect 49563 16989 49597 17023
rect 49681 16872 49715 16906
rect 21460 16331 21494 16365
rect 21578 16214 21612 16248
rect 22958 16329 22992 16363
rect 23076 16212 23110 16246
rect 24406 16329 24440 16363
rect 24524 16212 24558 16246
rect 38737 16177 38771 16211
rect 14451 15704 14485 15738
rect 14569 15704 14603 15738
rect 15899 15704 15933 15738
rect 16017 15704 16051 15738
rect 17397 15702 17431 15736
rect 17515 15702 17549 15736
rect 18845 15702 18879 15736
rect 18963 15702 18997 15736
rect 20365 15704 20399 15738
rect 20483 15704 20517 15738
rect 21813 15704 21847 15738
rect 21931 15704 21965 15738
rect 23311 15702 23345 15736
rect 23429 15702 23463 15736
rect 24759 15702 24793 15736
rect 24877 15702 24911 15736
rect 39307 15556 39341 15590
rect 39015 15487 39049 15521
rect 56097 16994 56131 17028
rect 56215 16877 56249 16911
rect 40223 15682 40257 15716
rect 39953 15555 39987 15589
rect 39569 15472 39603 15506
rect 39687 15471 39721 15505
rect 40138 15488 40172 15522
rect 43358 16366 43392 16400
rect 43476 16366 43510 16400
rect 40844 16198 40878 16232
rect 41203 15555 41237 15589
rect 40913 15487 40947 15521
rect 41851 15555 41885 15589
rect 41467 15472 41501 15506
rect 41585 15471 41619 15505
rect 45295 16173 45329 16207
rect 42036 15488 42070 15522
rect 45865 15552 45899 15586
rect 45573 15483 45607 15517
rect 43010 15389 43044 15423
rect 43128 15272 43162 15306
rect 62610 16997 62644 17031
rect 62728 16880 62762 16914
rect 46781 15678 46815 15712
rect 46511 15551 46545 15585
rect 46127 15468 46161 15502
rect 46245 15467 46279 15501
rect 46696 15484 46730 15518
rect 49916 16362 49950 16396
rect 50034 16362 50068 16396
rect 47402 16194 47436 16228
rect 47761 15551 47795 15585
rect 47471 15483 47505 15517
rect 48409 15551 48443 15585
rect 48025 15468 48059 15502
rect 48143 15467 48177 15501
rect 51829 16178 51863 16212
rect 48594 15484 48628 15518
rect 52399 15557 52433 15591
rect 52107 15488 52141 15522
rect 676 14262 710 14296
rect 1986 14221 2020 14255
rect 1856 14101 1914 14156
rect 1632 13991 1666 14025
rect 1751 13601 1785 13635
rect 2943 14100 3001 14155
rect 1974 13816 2032 13871
rect 3820 14262 3854 14296
rect 5130 14221 5164 14255
rect 5000 14101 5058 14156
rect 4776 13991 4810 14025
rect 4895 13601 4929 13635
rect 6087 14100 6145 14155
rect 5118 13816 5176 13871
rect 6952 14258 6986 14292
rect 8262 14217 8296 14251
rect 8132 14097 8190 14152
rect 7908 13987 7942 14021
rect 1809 13002 1843 13036
rect 8027 13597 8061 13631
rect 9219 14096 9277 14151
rect 8250 13812 8308 13867
rect 10096 14258 10130 14292
rect 11406 14217 11440 14251
rect 11276 14097 11334 14152
rect 11052 13987 11086 14021
rect 11171 13597 11205 13631
rect 12363 14096 12421 14151
rect 11394 13812 11452 13867
rect 13298 14262 13332 14296
rect 14608 14221 14642 14255
rect 14478 14101 14536 14156
rect 14254 13991 14288 14025
rect 14373 13601 14407 13635
rect 15565 14100 15623 14155
rect 14596 13816 14654 13871
rect 16442 14262 16476 14296
rect 17752 14221 17786 14255
rect 17622 14101 17680 14156
rect 17398 13991 17432 14025
rect 17517 13601 17551 13635
rect 49568 15385 49602 15419
rect 49686 15268 49720 15302
rect 53315 15683 53349 15717
rect 53045 15556 53079 15590
rect 52661 15473 52695 15507
rect 52779 15472 52813 15506
rect 53230 15489 53264 15523
rect 56450 16367 56484 16401
rect 56568 16367 56602 16401
rect 53936 16199 53970 16233
rect 54295 15556 54329 15590
rect 54005 15488 54039 15522
rect 54943 15556 54977 15590
rect 54559 15473 54593 15507
rect 54677 15472 54711 15506
rect 58342 16181 58376 16215
rect 55128 15489 55162 15523
rect 58912 15560 58946 15594
rect 58620 15491 58654 15525
rect 43363 14762 43397 14796
rect 43481 14762 43515 14796
rect 56102 15390 56136 15424
rect 56220 15273 56254 15307
rect 71075 16487 71109 16521
rect 59828 15686 59862 15720
rect 59558 15559 59592 15593
rect 59174 15476 59208 15510
rect 59292 15475 59326 15509
rect 59743 15492 59777 15526
rect 62963 16370 62997 16404
rect 63081 16370 63115 16404
rect 60449 16202 60483 16236
rect 60808 15559 60842 15593
rect 60518 15491 60552 15525
rect 61456 15559 61490 15593
rect 61072 15476 61106 15510
rect 61190 15475 61224 15509
rect 61641 15492 61675 15526
rect 71212 15622 71267 15680
rect 49921 14758 49955 14792
rect 50039 14758 50073 14792
rect 62615 15393 62649 15427
rect 62733 15276 62767 15310
rect 56455 14763 56489 14797
rect 56573 14763 56607 14797
rect 62968 14766 63002 14800
rect 63086 14766 63120 14800
rect 71112 14665 71146 14699
rect 71496 14653 71551 14711
rect 18709 14100 18767 14155
rect 17740 13816 17798 13871
rect 19574 14258 19608 14292
rect 20884 14217 20918 14251
rect 20754 14097 20812 14152
rect 20530 13987 20564 14021
rect 4953 13002 4987 13036
rect 8085 12998 8119 13032
rect 11229 12998 11263 13032
rect 14431 13002 14465 13036
rect 20649 13597 20683 13631
rect 21841 14096 21899 14151
rect 20872 13812 20930 13867
rect 22718 14258 22752 14292
rect 24028 14217 24062 14251
rect 23898 14097 23956 14152
rect 23674 13987 23708 14021
rect 23793 13597 23827 13631
rect 71211 14535 71266 14593
rect 72331 14488 72365 14522
rect 71732 14430 71766 14464
rect 71342 14311 71376 14345
rect 24985 14096 25043 14151
rect 24016 13812 24074 13867
rect 17575 13002 17609 13036
rect 20707 12998 20741 13032
rect 71071 13355 71105 13389
rect 23851 12998 23885 13032
rect 30715 13111 30749 13145
rect 31290 12862 31324 12896
rect 31223 12677 31257 12711
rect 31307 12411 31341 12445
rect 71212 12478 71267 12536
rect 676 11528 710 11562
rect 1986 11487 2020 11521
rect 1856 11367 1914 11422
rect 1632 11257 1666 11291
rect 1751 10867 1785 10901
rect 2943 11366 3001 11421
rect 1974 11082 2032 11137
rect 3820 11528 3854 11562
rect 5130 11487 5164 11521
rect 5000 11367 5058 11422
rect 4776 11257 4810 11291
rect 4895 10867 4929 10901
rect 6087 11366 6145 11421
rect 5118 11082 5176 11137
rect 6952 11524 6986 11558
rect 8262 11483 8296 11517
rect 8132 11363 8190 11418
rect 7908 11253 7942 11287
rect 1809 10268 1843 10302
rect 8027 10863 8061 10897
rect 9219 11362 9277 11417
rect 8250 11078 8308 11133
rect 10096 11524 10130 11558
rect 11406 11483 11440 11517
rect 11276 11363 11334 11418
rect 11052 11253 11086 11287
rect 11171 10863 11205 10897
rect 12363 11362 12421 11417
rect 11394 11078 11452 11133
rect 13298 11528 13332 11562
rect 14608 11487 14642 11521
rect 14478 11367 14536 11422
rect 14254 11257 14288 11291
rect 14373 10867 14407 10901
rect 15565 11366 15623 11421
rect 14596 11082 14654 11137
rect 16442 11528 16476 11562
rect 17752 11487 17786 11521
rect 17622 11367 17680 11422
rect 17398 11257 17432 11291
rect 17517 10867 17551 10901
rect 31306 12293 31340 12327
rect 31223 12029 31257 12063
rect 18709 11366 18767 11421
rect 17740 11082 17798 11137
rect 19574 11524 19608 11558
rect 20884 11483 20918 11517
rect 20754 11363 20812 11418
rect 20530 11253 20564 11287
rect 4953 10268 4987 10302
rect 8085 10264 8119 10298
rect 11229 10264 11263 10298
rect 14431 10268 14465 10302
rect 20649 10863 20683 10897
rect 21841 11362 21899 11417
rect 20872 11078 20930 11133
rect 22718 11524 22752 11558
rect 24028 11483 24062 11517
rect 23898 11363 23956 11418
rect 23674 11253 23708 11287
rect 23793 10863 23827 10897
rect 30521 11717 30555 11751
rect 31291 11739 31325 11773
rect 42337 11867 42371 11901
rect 42219 11750 42253 11784
rect 24985 11362 25043 11417
rect 24016 11078 24074 11133
rect 48886 11866 48920 11900
rect 48768 11749 48802 11783
rect 55540 11887 55574 11921
rect 55422 11770 55456 11804
rect 64193 11720 64227 11754
rect 64075 11603 64109 11637
rect 41866 11240 41900 11274
rect 41984 11240 42018 11274
rect 48415 11239 48449 11273
rect 48533 11239 48567 11273
rect 55069 11260 55103 11294
rect 55187 11260 55221 11294
rect 63722 11093 63756 11127
rect 63840 11093 63874 11127
rect 71112 11521 71146 11555
rect 71496 11509 71551 11567
rect 66886 11193 66920 11227
rect 30713 11043 30747 11077
rect 65486 11074 65520 11108
rect 17575 10268 17609 10302
rect 20707 10264 20741 10298
rect 31288 10794 31322 10828
rect 31221 10609 31255 10643
rect 23851 10264 23885 10298
rect 31305 10343 31339 10377
rect 31304 10225 31338 10259
rect 40006 10184 40040 10218
rect 41136 10190 41170 10224
rect 46555 10272 46589 10306
rect 47685 10278 47719 10312
rect 46555 10154 46589 10188
rect 47685 10158 47719 10192
rect 53209 10204 53243 10238
rect 54339 10210 54373 10244
rect 59834 10272 59868 10306
rect 60964 10278 60998 10312
rect 65691 10494 65725 10528
rect 65506 10427 65540 10461
rect 66339 10494 66373 10528
rect 65957 10410 65991 10444
rect 66075 10411 66109 10445
rect 67794 11312 67828 11346
rect 71211 11391 71266 11449
rect 67676 11195 67710 11229
rect 72331 11344 72365 11378
rect 71732 11286 71766 11320
rect 71342 11167 71376 11201
rect 67323 10685 67357 10719
rect 67441 10685 67475 10719
rect 66629 10426 66663 10460
rect 40006 10066 40040 10100
rect 41136 10070 41170 10104
rect 31221 9961 31255 9995
rect 35673 9967 35707 10001
rect 35555 9850 35589 9884
rect 30519 9649 30553 9683
rect 31289 9671 31323 9705
rect 686 8796 720 8830
rect 1996 8755 2030 8789
rect 1866 8635 1924 8690
rect 1642 8525 1676 8559
rect 1761 8135 1795 8169
rect 2953 8634 3011 8689
rect 1984 8350 2042 8405
rect 3830 8796 3864 8830
rect 5140 8755 5174 8789
rect 5010 8635 5068 8690
rect 4786 8525 4820 8559
rect 4905 8135 4939 8169
rect 38563 9700 38597 9734
rect 38445 9583 38479 9617
rect 6097 8634 6155 8689
rect 5128 8350 5186 8405
rect 6962 8792 6996 8826
rect 8272 8751 8306 8785
rect 8142 8631 8200 8686
rect 7918 8521 7952 8555
rect 1819 7536 1853 7570
rect 8037 8131 8071 8165
rect 9229 8630 9287 8685
rect 8260 8346 8318 8401
rect 10106 8792 10140 8826
rect 11416 8751 11450 8785
rect 11286 8631 11344 8686
rect 11062 8521 11096 8555
rect 11181 8131 11215 8165
rect 12373 8630 12431 8685
rect 11404 8346 11462 8401
rect 13308 8796 13342 8830
rect 14618 8755 14652 8789
rect 14488 8635 14546 8690
rect 14264 8525 14298 8559
rect 14383 8135 14417 8169
rect 15575 8634 15633 8689
rect 14606 8350 14664 8405
rect 16452 8796 16486 8830
rect 17762 8755 17796 8789
rect 17632 8635 17690 8690
rect 17408 8525 17442 8559
rect 17527 8135 17561 8169
rect 35202 9340 35236 9374
rect 35320 9340 35354 9374
rect 40326 9310 40360 9344
rect 45112 9788 45146 9822
rect 59834 10154 59868 10188
rect 53209 10086 53243 10120
rect 54339 10090 54373 10124
rect 60964 10158 60998 10192
rect 44994 9671 45028 9705
rect 41468 9314 41502 9348
rect 38092 9073 38126 9107
rect 38210 9073 38244 9107
rect 46875 9398 46909 9432
rect 51766 9720 51800 9754
rect 51648 9603 51682 9637
rect 48017 9402 48051 9436
rect 44641 9161 44675 9195
rect 44759 9161 44793 9195
rect 53529 9330 53563 9364
rect 58391 9788 58425 9822
rect 71071 10211 71105 10245
rect 58273 9671 58307 9705
rect 54671 9334 54705 9368
rect 51295 9093 51329 9127
rect 51413 9093 51447 9127
rect 60154 9398 60188 9432
rect 61296 9402 61330 9436
rect 57920 9161 57954 9195
rect 58038 9161 58072 9195
rect 71216 9276 71271 9334
rect 18719 8634 18777 8689
rect 17750 8350 17808 8405
rect 19584 8792 19618 8826
rect 20894 8751 20928 8785
rect 20764 8631 20822 8686
rect 20540 8521 20574 8555
rect 4963 7536 4997 7570
rect 8095 7532 8129 7566
rect 11239 7532 11273 7566
rect 14441 7536 14475 7570
rect 20659 8131 20693 8165
rect 21851 8630 21909 8685
rect 20882 8346 20940 8401
rect 22728 8792 22762 8826
rect 24038 8751 24072 8785
rect 23908 8631 23966 8686
rect 23684 8521 23718 8555
rect 23803 8131 23837 8165
rect 30715 8974 30749 9008
rect 64188 9149 64222 9183
rect 64070 9032 64104 9066
rect 31290 8725 31324 8759
rect 24995 8630 25053 8685
rect 24026 8346 24084 8401
rect 31223 8540 31257 8574
rect 63717 8522 63751 8556
rect 31307 8274 31341 8308
rect 17585 7536 17619 7570
rect 20717 7532 20751 7566
rect 31306 8156 31340 8190
rect 63835 8522 63869 8556
rect 31223 7892 31257 7926
rect 38577 8050 38611 8084
rect 45126 8138 45160 8172
rect 71116 8319 71150 8353
rect 71500 8307 71555 8365
rect 45008 8021 45042 8055
rect 38459 7933 38493 7967
rect 23861 7532 23895 7566
rect 30521 7580 30555 7614
rect 31291 7602 31325 7636
rect 35665 7382 35699 7416
rect 38106 7423 38140 7457
rect 38224 7423 38258 7457
rect 35547 7265 35581 7299
rect 30713 6906 30747 6940
rect 35194 6755 35228 6789
rect 35312 6755 35346 6789
rect 31288 6657 31322 6691
rect 3307 6229 3341 6263
rect 4045 6229 4079 6263
rect 4783 6229 4817 6263
rect 5521 6229 5555 6263
rect 6261 6229 6295 6263
rect 7003 6229 7037 6263
rect 7741 6229 7775 6263
rect 8479 6231 8513 6265
rect 9491 5846 9525 5880
rect 11559 5844 11593 5878
rect 10885 5652 10919 5686
rect 9803 5144 9837 5178
rect 9513 5076 9547 5110
rect 10451 5144 10485 5178
rect 10067 5061 10101 5095
rect 10185 5060 10219 5094
rect 10636 5077 10670 5111
rect 13628 5846 13662 5880
rect 12953 5650 12987 5684
rect 11871 5142 11905 5176
rect 11581 5074 11615 5108
rect 12519 5142 12553 5176
rect 12135 5059 12169 5093
rect 12253 5058 12287 5092
rect 12704 5075 12738 5109
rect 15696 5844 15730 5878
rect 15022 5652 15056 5686
rect 13940 5144 13974 5178
rect 13650 5076 13684 5110
rect 14588 5144 14622 5178
rect 14204 5061 14238 5095
rect 14322 5060 14356 5094
rect 14773 5077 14807 5111
rect 17765 5844 17799 5878
rect 17090 5650 17124 5684
rect 16008 5142 16042 5176
rect 15718 5074 15752 5108
rect 16656 5142 16690 5176
rect 16272 5059 16306 5093
rect 16390 5058 16424 5092
rect 16841 5075 16875 5109
rect 40738 7255 40772 7289
rect 39731 6612 39765 6646
rect 39546 6545 39580 6579
rect 31221 6472 31255 6506
rect 40379 6612 40413 6646
rect 39997 6528 40031 6562
rect 40115 6529 40149 6563
rect 40669 6544 40703 6578
rect 44655 7511 44689 7545
rect 44773 7511 44807 7545
rect 51780 8070 51814 8104
rect 51662 7953 51696 7987
rect 58405 8138 58439 8172
rect 58287 8021 58321 8055
rect 71215 8189 71270 8247
rect 72335 8142 72369 8176
rect 71736 8084 71770 8118
rect 42845 7234 42879 7268
rect 41359 6739 41393 6773
rect 41629 6612 41663 6646
rect 41444 6545 41478 6579
rect 42275 6613 42309 6647
rect 41895 6528 41929 6562
rect 42013 6529 42047 6563
rect 47287 7343 47321 7377
rect 46280 6700 46314 6734
rect 46095 6633 46129 6667
rect 42567 6544 42601 6578
rect 38572 6446 38606 6480
rect 38454 6329 38488 6363
rect 31305 6206 31339 6240
rect 19833 5842 19867 5876
rect 19159 5650 19193 5684
rect 18077 5142 18111 5176
rect 17787 5074 17821 5108
rect 18725 5142 18759 5176
rect 18341 5059 18375 5093
rect 18459 5058 18493 5092
rect 18910 5075 18944 5109
rect 21902 5844 21936 5878
rect 21227 5648 21261 5682
rect 20145 5140 20179 5174
rect 19855 5072 19889 5106
rect 20793 5140 20827 5174
rect 20409 5057 20443 5091
rect 20527 5056 20561 5090
rect 20978 5073 21012 5107
rect 23970 5842 24004 5876
rect 23296 5650 23330 5684
rect 22214 5142 22248 5176
rect 21924 5074 21958 5108
rect 22862 5142 22896 5176
rect 22478 5059 22512 5093
rect 22596 5058 22630 5092
rect 23047 5075 23081 5109
rect 31304 6088 31338 6122
rect 46928 6700 46962 6734
rect 46546 6616 46580 6650
rect 46664 6617 46698 6651
rect 47218 6632 47252 6666
rect 51309 7443 51343 7477
rect 51427 7443 51461 7477
rect 49394 7322 49428 7356
rect 47908 6827 47942 6861
rect 48178 6700 48212 6734
rect 47993 6633 48027 6667
rect 48824 6701 48858 6735
rect 48444 6616 48478 6650
rect 48562 6617 48596 6651
rect 49116 6632 49150 6666
rect 45121 6534 45155 6568
rect 45003 6417 45037 6451
rect 53941 7275 53975 7309
rect 52934 6632 52968 6666
rect 52749 6565 52783 6599
rect 53582 6632 53616 6666
rect 53200 6548 53234 6582
rect 53318 6549 53352 6583
rect 53872 6564 53906 6598
rect 57934 7511 57968 7545
rect 58052 7511 58086 7545
rect 71346 7965 71380 7999
rect 56048 7254 56082 7288
rect 54562 6759 54596 6793
rect 54832 6632 54866 6666
rect 54647 6565 54681 6599
rect 55478 6633 55512 6667
rect 55098 6548 55132 6582
rect 55216 6549 55250 6583
rect 60566 7343 60600 7377
rect 59559 6700 59593 6734
rect 59374 6633 59408 6667
rect 55770 6564 55804 6598
rect 51775 6466 51809 6500
rect 51657 6349 51691 6383
rect 25364 5648 25398 5682
rect 24282 5140 24316 5174
rect 23992 5072 24026 5106
rect 24930 5140 24964 5174
rect 24546 5057 24580 5091
rect 24664 5056 24698 5090
rect 31221 5824 31255 5858
rect 38101 5819 38135 5853
rect 38219 5819 38253 5853
rect 44650 5907 44684 5941
rect 44768 5907 44802 5941
rect 60207 6700 60241 6734
rect 59825 6616 59859 6650
rect 59943 6617 59977 6651
rect 60497 6632 60531 6666
rect 62673 7322 62707 7356
rect 61187 6827 61221 6861
rect 61457 6700 61491 6734
rect 61272 6633 61306 6667
rect 62103 6701 62137 6735
rect 61723 6616 61757 6650
rect 61841 6617 61875 6651
rect 62395 6632 62429 6666
rect 66888 7102 66922 7136
rect 65488 6983 65522 7017
rect 58400 6534 58434 6568
rect 58282 6417 58316 6451
rect 65693 6403 65727 6437
rect 65508 6336 65542 6370
rect 66341 6403 66375 6437
rect 65959 6319 65993 6353
rect 66077 6320 66111 6354
rect 67796 7221 67830 7255
rect 67678 7104 67712 7138
rect 71075 7009 71109 7043
rect 67325 6594 67359 6628
rect 67443 6594 67477 6628
rect 66631 6335 66665 6369
rect 51304 5839 51338 5873
rect 51422 5839 51456 5873
rect 57929 5907 57963 5941
rect 58047 5907 58081 5941
rect 64188 6116 64222 6150
rect 64070 5999 64104 6033
rect 30519 5512 30553 5546
rect 31289 5534 31323 5568
rect 71216 6132 71271 6190
rect 63717 5489 63751 5523
rect 63835 5489 63869 5523
rect 71116 5175 71150 5209
rect 71500 5163 71555 5221
rect 25115 5073 25149 5107
rect 71215 5045 71270 5103
rect 30713 4837 30747 4871
rect 72335 4998 72369 5032
rect 71736 4940 71770 4974
rect 71346 4821 71380 4855
rect 31288 4588 31322 4622
rect 31221 4403 31255 4437
rect 39998 4404 40032 4438
rect 41128 4410 41162 4444
rect 31305 4137 31339 4171
rect 46549 4402 46583 4436
rect 47679 4408 47713 4442
rect 39998 4286 40032 4320
rect 41128 4290 41162 4324
rect 53204 4403 53238 4437
rect 54334 4409 54368 4443
rect 46549 4284 46583 4318
rect 31304 4019 31338 4053
rect 35646 4104 35680 4138
rect 35528 3987 35562 4021
rect 31221 3755 31255 3789
rect 38555 3920 38589 3954
rect 47679 4288 47713 4322
rect 59826 4404 59860 4438
rect 60956 4410 60990 4444
rect 53204 4285 53238 4319
rect 38437 3803 38471 3837
rect 30519 3443 30553 3477
rect 31289 3465 31323 3499
rect 35175 3477 35209 3511
rect 35293 3477 35327 3511
rect 40318 3530 40352 3564
rect 45106 3918 45140 3952
rect 54334 4289 54368 4323
rect 59826 4286 59860 4320
rect 44988 3801 45022 3835
rect 41460 3534 41494 3568
rect 38084 3293 38118 3327
rect 38202 3293 38236 3327
rect 46869 3528 46903 3562
rect 51761 3919 51795 3953
rect 60956 4290 60990 4324
rect 51643 3802 51677 3836
rect 48011 3532 48045 3566
rect 44635 3291 44669 3325
rect 44753 3291 44787 3325
rect 53524 3529 53558 3563
rect 58383 3920 58417 3954
rect 64259 4196 64293 4230
rect 64141 4079 64175 4113
rect 58265 3803 58299 3837
rect 54666 3533 54700 3567
rect 51290 3292 51324 3326
rect 51408 3292 51442 3326
rect 60146 3530 60180 3564
rect 61288 3534 61322 3568
rect 63788 3569 63822 3603
rect 63906 3569 63940 3603
rect 71075 3865 71109 3899
rect 66888 3607 66922 3641
rect 57912 3293 57946 3327
rect 58030 3293 58064 3327
rect 65488 3488 65522 3522
rect 30711 2769 30745 2803
rect 65693 2908 65727 2942
rect 65508 2841 65542 2875
rect 66341 2908 66375 2942
rect 65959 2824 65993 2858
rect 66077 2825 66111 2859
rect 67796 3726 67830 3760
rect 67678 3609 67712 3643
rect 67325 3099 67359 3133
rect 67443 3099 67477 3133
rect 71212 3000 71267 3058
rect 66631 2840 66665 2874
rect 31286 2520 31320 2554
rect 31219 2335 31253 2369
rect 365 1382 423 1437
rect 1346 1503 1380 1537
rect 1452 1383 1510 1438
rect 1334 1098 1392 1153
rect 2656 1544 2690 1578
rect 1700 1273 1734 1307
rect 1581 883 1615 917
rect 3509 1382 3567 1437
rect 4490 1503 4524 1537
rect 4596 1383 4654 1438
rect 4478 1098 4536 1153
rect 5800 1544 5834 1578
rect 4844 1273 4878 1307
rect 4725 883 4759 917
rect 6641 1386 6699 1441
rect 7622 1507 7656 1541
rect 7728 1387 7786 1442
rect 7610 1102 7668 1157
rect 8932 1548 8966 1582
rect 7976 1277 8010 1311
rect 7857 887 7891 921
rect 9785 1386 9843 1441
rect 10766 1507 10800 1541
rect 10872 1387 10930 1442
rect 10754 1102 10812 1157
rect 31303 2069 31337 2103
rect 38569 2270 38603 2304
rect 38451 2153 38485 2187
rect 12076 1548 12110 1582
rect 11120 1277 11154 1311
rect 11001 887 11035 921
rect 12987 1382 13045 1437
rect 13968 1503 14002 1537
rect 14074 1383 14132 1438
rect 13956 1098 14014 1153
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 15278 1544 15312 1578
rect 14322 1273 14356 1307
rect 14203 883 14237 917
rect 16131 1382 16189 1437
rect 17112 1503 17146 1537
rect 17218 1383 17276 1438
rect 17100 1098 17158 1153
rect 18422 1544 18456 1578
rect 17466 1273 17500 1307
rect 17347 883 17381 917
rect 19263 1386 19321 1441
rect 20244 1507 20278 1541
rect 20350 1387 20408 1442
rect 20232 1102 20290 1157
rect 21554 1548 21588 1582
rect 20598 1277 20632 1311
rect 20479 887 20513 921
rect 22407 1386 22465 1441
rect 23388 1507 23422 1541
rect 23494 1387 23552 1442
rect 23376 1102 23434 1157
rect 31302 1951 31336 1985
rect 24698 1548 24732 1582
rect 23742 1277 23776 1311
rect 23623 887 23657 921
rect 31219 1687 31253 1721
rect 38098 1643 38132 1677
rect 38216 1643 38250 1677
rect 45120 2268 45154 2302
rect 45002 2151 45036 2185
rect 30517 1375 30551 1409
rect 31287 1397 31321 1431
rect 35662 1344 35696 1378
rect 35544 1227 35578 1261
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 30713 700 30747 734
rect 35191 717 35225 751
rect 35309 717 35343 751
rect 40730 1475 40764 1509
rect 39723 832 39757 866
rect 39538 765 39572 799
rect 31288 451 31322 485
rect 40371 832 40405 866
rect 39989 748 40023 782
rect 40107 749 40141 783
rect 40661 764 40695 798
rect 44649 1641 44683 1675
rect 44767 1641 44801 1675
rect 51775 2269 51809 2303
rect 51657 2152 51691 2186
rect 42837 1454 42871 1488
rect 41351 959 41385 993
rect 41621 832 41655 866
rect 41436 765 41470 799
rect 42267 833 42301 867
rect 41887 748 41921 782
rect 42005 749 42039 783
rect 42559 764 42593 798
rect 47281 1473 47315 1507
rect 46274 830 46308 864
rect 46089 763 46123 797
rect 38564 666 38598 700
rect 38446 549 38480 583
rect 23565 288 23599 322
rect 31221 266 31255 300
rect 46922 830 46956 864
rect 46540 746 46574 780
rect 46658 747 46692 781
rect 47212 762 47246 796
rect 51304 1642 51338 1676
rect 51422 1642 51456 1676
rect 58397 2270 58431 2304
rect 58279 2153 58313 2187
rect 49388 1452 49422 1486
rect 47902 957 47936 991
rect 48172 830 48206 864
rect 47987 763 48021 797
rect 48818 831 48852 865
rect 48438 746 48472 780
rect 48556 747 48590 781
rect 49110 762 49144 796
rect 53936 1474 53970 1508
rect 52929 831 52963 865
rect 52744 764 52778 798
rect 45115 664 45149 698
rect 44997 547 45031 581
rect 31305 0 31339 34
rect 38093 39 38127 73
rect 38211 39 38245 73
rect 53577 831 53611 865
rect 53195 747 53229 781
rect 53313 748 53347 782
rect 53867 763 53901 797
rect 57926 1643 57960 1677
rect 58044 1643 58078 1677
rect 71112 2043 71146 2077
rect 71496 2031 71551 2089
rect 71211 1913 71266 1971
rect 56043 1453 56077 1487
rect 54557 958 54591 992
rect 54827 831 54861 865
rect 54642 764 54676 798
rect 55473 832 55507 866
rect 55093 747 55127 781
rect 55211 748 55245 782
rect 55765 763 55799 797
rect 60558 1475 60592 1509
rect 59551 832 59585 866
rect 59366 765 59400 799
rect 51770 665 51804 699
rect 51652 548 51686 582
rect 31304 -118 31338 -84
rect 44644 37 44678 71
rect 44762 37 44796 71
rect 60199 832 60233 866
rect 59817 748 59851 782
rect 59935 749 59969 783
rect 60489 764 60523 798
rect 72331 1866 72365 1900
rect 71732 1808 71766 1842
rect 71342 1689 71376 1723
rect 62665 1454 62699 1488
rect 61179 959 61213 993
rect 61449 832 61483 866
rect 61264 765 61298 799
rect 62095 833 62129 867
rect 61715 748 61749 782
rect 61833 749 61867 783
rect 64256 1126 64290 1160
rect 64138 1009 64172 1043
rect 62387 764 62421 798
rect 58392 666 58426 700
rect 58274 549 58308 583
rect 51299 38 51333 72
rect 51417 38 51451 72
rect 71071 733 71105 767
rect 63785 499 63819 533
rect 63903 499 63937 533
rect 57921 39 57955 73
rect 58039 39 58073 73
rect 31221 -382 31255 -348
rect 71212 -144 71267 -86
rect 30519 -694 30553 -660
rect 31289 -672 31323 -638
rect 66888 -741 66922 -707
rect 41901 -880 41935 -846
rect 42019 -880 42053 -846
rect 48455 -875 48489 -841
rect 48573 -875 48607 -841
rect 55104 -887 55138 -853
rect 55222 -887 55256 -853
rect 65488 -860 65522 -826
rect 30711 -1368 30745 -1334
rect 42254 -1390 42288 -1356
rect 42372 -1507 42406 -1473
rect 31286 -1617 31320 -1583
rect 48808 -1385 48842 -1351
rect 48926 -1502 48960 -1468
rect 55457 -1397 55491 -1363
rect 55575 -1514 55609 -1480
rect 397 -2510 455 -2455
rect 1378 -2389 1412 -2355
rect 1484 -2509 1542 -2454
rect 1366 -2794 1424 -2739
rect 2688 -2348 2722 -2314
rect 1732 -2619 1766 -2585
rect 1613 -3009 1647 -2975
rect 3541 -2510 3599 -2455
rect 4522 -2389 4556 -2355
rect 4628 -2509 4686 -2454
rect 4510 -2794 4568 -2739
rect 5832 -2348 5866 -2314
rect 4876 -2619 4910 -2585
rect 4757 -3009 4791 -2975
rect 6673 -2506 6731 -2451
rect 7654 -2385 7688 -2351
rect 7760 -2505 7818 -2450
rect 7642 -2790 7700 -2735
rect 8964 -2344 8998 -2310
rect 8008 -2615 8042 -2581
rect 7889 -3005 7923 -2971
rect 9817 -2506 9875 -2451
rect 10798 -2385 10832 -2351
rect 10904 -2505 10962 -2450
rect 10786 -2790 10844 -2735
rect 31219 -1802 31253 -1768
rect 65693 -1440 65727 -1406
rect 65508 -1507 65542 -1473
rect 66341 -1440 66375 -1406
rect 65959 -1524 65993 -1490
rect 66077 -1523 66111 -1489
rect 67796 -622 67830 -588
rect 67678 -739 67712 -705
rect 71112 -1101 71146 -1067
rect 71496 -1113 71551 -1055
rect 67325 -1249 67359 -1215
rect 67443 -1249 67477 -1215
rect 71211 -1231 71266 -1173
rect 72331 -1278 72365 -1244
rect 71732 -1336 71766 -1302
rect 66631 -1508 66665 -1474
rect 71342 -1455 71376 -1421
rect 64263 -1719 64297 -1685
rect 64145 -1836 64179 -1802
rect 12108 -2344 12142 -2310
rect 11152 -2615 11186 -2581
rect 11033 -3005 11067 -2971
rect 13019 -2510 13077 -2455
rect 14000 -2389 14034 -2355
rect 14106 -2509 14164 -2454
rect 13988 -2794 14046 -2739
rect 1555 -3608 1589 -3574
rect 4699 -3608 4733 -3574
rect 15310 -2348 15344 -2314
rect 14354 -2619 14388 -2585
rect 14235 -3009 14269 -2975
rect 16163 -2510 16221 -2455
rect 17144 -2389 17178 -2355
rect 17250 -2509 17308 -2454
rect 17132 -2794 17190 -2739
rect 18454 -2348 18488 -2314
rect 17498 -2619 17532 -2585
rect 17379 -3009 17413 -2975
rect 19295 -2506 19353 -2451
rect 20276 -2385 20310 -2351
rect 20382 -2505 20440 -2450
rect 20264 -2790 20322 -2735
rect 21586 -2344 21620 -2310
rect 20630 -2615 20664 -2581
rect 20511 -3005 20545 -2971
rect 22439 -2506 22497 -2451
rect 23420 -2385 23454 -2351
rect 23526 -2505 23584 -2450
rect 23408 -2790 23466 -2735
rect 24730 -2344 24764 -2310
rect 23774 -2615 23808 -2581
rect 23655 -3005 23689 -2971
rect 31303 -2068 31337 -2034
rect 31302 -2186 31336 -2152
rect 63792 -2346 63826 -2312
rect 63910 -2346 63944 -2312
rect 31219 -2450 31253 -2416
rect 71071 -2411 71105 -2377
rect 30517 -2762 30551 -2728
rect 31287 -2740 31321 -2706
rect 7831 -3604 7865 -3570
rect 10975 -3604 11009 -3570
rect 14177 -3608 14211 -3574
rect 17321 -3608 17355 -3574
rect 20453 -3604 20487 -3570
rect 23597 -3604 23631 -3570
<< locali >>
rect 39995 24935 40218 25011
rect 39995 24786 40074 24935
rect 40141 24786 40218 24935
rect 39995 24680 40218 24786
rect 42477 24989 42700 25065
rect 42477 24840 42556 24989
rect 42623 24840 42700 24989
rect 41810 24769 41844 24785
rect 41810 24719 41844 24735
rect 42477 24734 42700 24840
rect 43624 24989 43847 25065
rect 43624 24840 43703 24989
rect 43770 24840 43847 24989
rect 42940 24775 42974 24791
rect 42940 24725 42974 24741
rect 43624 24734 43847 24840
rect 46508 24932 46731 25008
rect 46508 24783 46587 24932
rect 46654 24783 46731 24932
rect 46508 24677 46731 24783
rect 48990 24986 49213 25062
rect 48990 24837 49069 24986
rect 49136 24837 49213 24986
rect 48323 24766 48357 24782
rect 48323 24716 48357 24732
rect 48990 24731 49213 24837
rect 50137 24986 50360 25062
rect 50137 24837 50216 24986
rect 50283 24837 50360 24986
rect 49453 24772 49487 24788
rect 49453 24722 49487 24738
rect 50137 24731 50360 24837
rect 53042 24927 53265 25003
rect 53042 24778 53121 24927
rect 53188 24778 53265 24927
rect 53042 24672 53265 24778
rect 55524 24981 55747 25057
rect 55524 24832 55603 24981
rect 55670 24832 55747 24981
rect 54857 24761 54891 24777
rect 54857 24711 54891 24727
rect 55524 24726 55747 24832
rect 56671 24981 56894 25057
rect 56671 24832 56750 24981
rect 56817 24832 56894 24981
rect 55987 24767 56021 24783
rect 55987 24717 56021 24733
rect 56671 24726 56894 24832
rect 59600 24931 59823 25007
rect 59600 24782 59679 24931
rect 59746 24782 59823 24931
rect 59600 24676 59823 24782
rect 62082 24985 62305 25061
rect 62082 24836 62161 24985
rect 62228 24836 62305 24985
rect 61415 24765 61449 24781
rect 61415 24715 61449 24731
rect 62082 24730 62305 24836
rect 63229 24985 63452 25061
rect 63229 24836 63308 24985
rect 63375 24836 63452 24985
rect 62545 24771 62579 24787
rect 62545 24721 62579 24737
rect 63229 24730 63452 24836
rect 41810 24651 41844 24667
rect 40426 24571 40696 24605
rect 41810 24601 41844 24617
rect 42940 24655 42974 24671
rect 39600 24521 39634 24537
rect 39600 24329 39634 24345
rect 39718 24521 39752 24537
rect 39718 24329 39752 24345
rect 39836 24521 39870 24537
rect 39836 24329 39870 24345
rect 39954 24521 39988 24537
rect 39954 24329 39988 24345
rect 40072 24521 40106 24537
rect 40072 24329 40106 24345
rect 40190 24521 40224 24537
rect 40190 24329 40224 24345
rect 40308 24521 40342 24537
rect 40308 24329 40342 24345
rect 40426 24521 40460 24571
rect 40426 24329 40460 24345
rect 40544 24521 40578 24537
rect 40544 24329 40578 24345
rect 40662 24521 40696 24571
rect 40662 24329 40696 24345
rect 41925 24593 41959 24609
rect 40351 24251 40367 24285
rect 40401 24251 40417 24285
rect 41925 24201 41959 24217
rect 42043 24593 42077 24609
rect 42043 24201 42077 24217
rect 42161 24593 42195 24609
rect 42161 24201 42195 24217
rect 42279 24593 42313 24609
rect 42279 24201 42313 24217
rect 42397 24593 42431 24609
rect 42397 24201 42431 24217
rect 42515 24593 42549 24609
rect 42515 24201 42549 24217
rect 42633 24593 42667 24609
rect 42940 24605 42974 24621
rect 48323 24648 48357 24664
rect 42633 24201 42667 24217
rect 43067 24597 43101 24613
rect 43067 24205 43101 24221
rect 43185 24597 43219 24613
rect 43185 24205 43219 24221
rect 43303 24597 43337 24613
rect 43303 24205 43337 24221
rect 43421 24597 43455 24613
rect 43421 24205 43455 24221
rect 43539 24597 43573 24613
rect 43539 24205 43573 24221
rect 43657 24597 43691 24613
rect 43657 24205 43691 24221
rect 43775 24597 43809 24613
rect 46939 24568 47209 24602
rect 48323 24598 48357 24614
rect 49453 24652 49487 24668
rect 46113 24518 46147 24534
rect 46113 24326 46147 24342
rect 46231 24518 46265 24534
rect 46231 24326 46265 24342
rect 46349 24518 46383 24534
rect 46349 24326 46383 24342
rect 46467 24518 46501 24534
rect 46467 24326 46501 24342
rect 46585 24518 46619 24534
rect 46585 24326 46619 24342
rect 46703 24518 46737 24534
rect 46703 24326 46737 24342
rect 46821 24518 46855 24534
rect 46821 24326 46855 24342
rect 46939 24518 46973 24568
rect 46939 24326 46973 24342
rect 47057 24518 47091 24534
rect 47057 24326 47091 24342
rect 47175 24518 47209 24568
rect 47175 24326 47209 24342
rect 48438 24590 48472 24606
rect 46864 24248 46880 24282
rect 46914 24248 46930 24282
rect 43775 24205 43809 24221
rect 48438 24198 48472 24214
rect 48556 24590 48590 24606
rect 48556 24198 48590 24214
rect 48674 24590 48708 24606
rect 48674 24198 48708 24214
rect 48792 24590 48826 24606
rect 48792 24198 48826 24214
rect 48910 24590 48944 24606
rect 48910 24198 48944 24214
rect 49028 24590 49062 24606
rect 49028 24198 49062 24214
rect 49146 24590 49180 24606
rect 49453 24602 49487 24618
rect 54857 24643 54891 24659
rect 49146 24198 49180 24214
rect 49580 24594 49614 24610
rect 49580 24202 49614 24218
rect 49698 24594 49732 24610
rect 49698 24202 49732 24218
rect 49816 24594 49850 24610
rect 49816 24202 49850 24218
rect 49934 24594 49968 24610
rect 49934 24202 49968 24218
rect 50052 24594 50086 24610
rect 50052 24202 50086 24218
rect 50170 24594 50204 24610
rect 50170 24202 50204 24218
rect 50288 24594 50322 24610
rect 53473 24563 53743 24597
rect 54857 24593 54891 24609
rect 55987 24647 56021 24663
rect 52647 24513 52681 24529
rect 52647 24321 52681 24337
rect 52765 24513 52799 24529
rect 52765 24321 52799 24337
rect 52883 24513 52917 24529
rect 52883 24321 52917 24337
rect 53001 24513 53035 24529
rect 53001 24321 53035 24337
rect 53119 24513 53153 24529
rect 53119 24321 53153 24337
rect 53237 24513 53271 24529
rect 53237 24321 53271 24337
rect 53355 24513 53389 24529
rect 53355 24321 53389 24337
rect 53473 24513 53507 24563
rect 53473 24321 53507 24337
rect 53591 24513 53625 24529
rect 53591 24321 53625 24337
rect 53709 24513 53743 24563
rect 53709 24321 53743 24337
rect 54972 24585 55006 24601
rect 53398 24243 53414 24277
rect 53448 24243 53464 24277
rect 50288 24202 50322 24218
rect 54972 24193 55006 24209
rect 55090 24585 55124 24601
rect 55090 24193 55124 24209
rect 55208 24585 55242 24601
rect 55208 24193 55242 24209
rect 55326 24585 55360 24601
rect 55326 24193 55360 24209
rect 55444 24585 55478 24601
rect 55444 24193 55478 24209
rect 55562 24585 55596 24601
rect 55562 24193 55596 24209
rect 55680 24585 55714 24601
rect 55987 24597 56021 24613
rect 61415 24647 61449 24663
rect 55680 24193 55714 24209
rect 56114 24589 56148 24605
rect 56114 24197 56148 24213
rect 56232 24589 56266 24605
rect 56232 24197 56266 24213
rect 56350 24589 56384 24605
rect 56350 24197 56384 24213
rect 56468 24589 56502 24605
rect 56468 24197 56502 24213
rect 56586 24589 56620 24605
rect 56586 24197 56620 24213
rect 56704 24589 56738 24605
rect 56704 24197 56738 24213
rect 56822 24589 56856 24605
rect 60031 24567 60301 24601
rect 61415 24597 61449 24613
rect 62545 24651 62579 24667
rect 59205 24517 59239 24533
rect 59205 24325 59239 24341
rect 59323 24517 59357 24533
rect 59323 24325 59357 24341
rect 59441 24517 59475 24533
rect 59441 24325 59475 24341
rect 59559 24517 59593 24533
rect 59559 24325 59593 24341
rect 59677 24517 59711 24533
rect 59677 24325 59711 24341
rect 59795 24517 59829 24533
rect 59795 24325 59829 24341
rect 59913 24517 59947 24533
rect 59913 24325 59947 24341
rect 60031 24517 60065 24567
rect 60031 24325 60065 24341
rect 60149 24517 60183 24533
rect 60149 24325 60183 24341
rect 60267 24517 60301 24567
rect 60267 24325 60301 24341
rect 61530 24589 61564 24605
rect 59956 24247 59972 24281
rect 60006 24247 60022 24281
rect 56822 24197 56856 24213
rect 61530 24197 61564 24213
rect 61648 24589 61682 24605
rect 61648 24197 61682 24213
rect 61766 24589 61800 24605
rect 61766 24197 61800 24213
rect 61884 24589 61918 24605
rect 61884 24197 61918 24213
rect 62002 24589 62036 24605
rect 62002 24197 62036 24213
rect 62120 24589 62154 24605
rect 62120 24197 62154 24213
rect 62238 24589 62272 24605
rect 62545 24601 62579 24617
rect 62238 24197 62272 24213
rect 62672 24593 62706 24609
rect 62672 24201 62706 24217
rect 62790 24593 62824 24609
rect 62790 24201 62824 24217
rect 62908 24593 62942 24609
rect 62908 24201 62942 24217
rect 63026 24593 63060 24609
rect 63026 24201 63060 24217
rect 63144 24593 63178 24609
rect 63144 24201 63178 24217
rect 63262 24593 63296 24609
rect 63262 24201 63296 24217
rect 63380 24593 63414 24609
rect 63380 24201 63414 24217
rect 28274 24163 28352 24172
rect 28274 24096 28285 24163
rect 28342 24096 28352 24163
rect 40233 24134 40249 24168
rect 40283 24134 40299 24168
rect 46746 24131 46762 24165
rect 46796 24131 46812 24165
rect 53280 24126 53296 24160
rect 53330 24126 53346 24160
rect 59838 24130 59854 24164
rect 59888 24130 59904 24164
rect 4210 22254 4438 22272
rect 4210 22178 4226 22254
rect 4422 22178 4438 22254
rect 4210 22162 4438 22178
rect 7354 22254 7582 22272
rect 7354 22178 7370 22254
rect 7566 22178 7582 22254
rect 7354 22162 7582 22178
rect 10486 22250 10714 22268
rect 10486 22174 10502 22250
rect 10698 22174 10714 22250
rect 10486 22158 10714 22174
rect 13630 22250 13858 22268
rect 13630 22174 13646 22250
rect 13842 22174 13858 22250
rect 13630 22158 13858 22174
rect 16832 22254 17060 22272
rect 16832 22178 16848 22254
rect 17044 22178 17060 22254
rect 16832 22162 17060 22178
rect 19976 22254 20204 22272
rect 19976 22178 19992 22254
rect 20188 22178 20204 22254
rect 19976 22162 20204 22178
rect 23108 22250 23336 22268
rect 23108 22174 23124 22250
rect 23320 22174 23336 22250
rect 23108 22158 23336 22174
rect 26252 22250 26480 22268
rect 26252 22174 26268 22250
rect 26464 22174 26480 22250
rect 26252 22158 26480 22174
rect 3485 22036 3755 22075
rect 3485 21984 3519 22036
rect 3012 21834 3282 21871
rect 3012 21784 3046 21834
rect 3012 21592 3046 21608
rect 3130 21784 3164 21800
rect 3130 21554 3164 21608
rect 3248 21784 3282 21834
rect 3248 21592 3282 21608
rect 3366 21784 3400 21800
rect 3366 21554 3400 21608
rect 3485 21592 3519 21608
rect 3603 21984 3637 22000
rect 3130 21515 3400 21554
rect 3603 21557 3637 21608
rect 3721 21984 3755 22036
rect 3958 22036 4228 22075
rect 3721 21592 3755 21608
rect 3839 21984 3873 22000
rect 3839 21557 3873 21608
rect 3958 21984 3992 22036
rect 3958 21592 3992 21608
rect 4076 21984 4110 22000
rect 4076 21557 4110 21608
rect 4194 21984 4228 22036
rect 4430 22036 4700 22075
rect 4194 21592 4228 21608
rect 4312 21984 4346 22000
rect 4312 21557 4346 21608
rect 4430 21984 4464 22036
rect 4430 21592 4464 21608
rect 4548 21984 4582 22000
rect 4548 21557 4582 21608
rect 4666 21984 4700 22036
rect 4897 22037 5167 22076
rect 4666 21592 4700 21608
rect 4779 21984 4813 22000
rect 4779 21557 4813 21608
rect 4897 21984 4931 22037
rect 4897 21592 4931 21608
rect 5015 21984 5049 22000
rect 5015 21557 5049 21608
rect 5133 21984 5167 22037
rect 6629 22036 6899 22075
rect 6629 21984 6663 22036
rect 5338 21835 5608 21874
rect 5133 21592 5167 21608
rect 5220 21784 5254 21800
rect 3603 21518 5049 21557
rect 5220 21557 5254 21608
rect 5338 21784 5372 21835
rect 5338 21592 5372 21608
rect 5456 21784 5490 21800
rect 5456 21557 5490 21608
rect 5574 21784 5608 21835
rect 5574 21592 5608 21608
rect 6156 21834 6426 21871
rect 6156 21784 6190 21834
rect 6156 21592 6190 21608
rect 6274 21784 6308 21800
rect 5220 21518 5490 21557
rect 6274 21554 6308 21608
rect 6392 21784 6426 21834
rect 6392 21592 6426 21608
rect 6510 21784 6544 21800
rect 6510 21554 6544 21608
rect 6629 21592 6663 21608
rect 6747 21984 6781 22000
rect 6274 21515 6544 21554
rect 6747 21557 6781 21608
rect 6865 21984 6899 22036
rect 7102 22036 7372 22075
rect 6865 21592 6899 21608
rect 6983 21984 7017 22000
rect 6983 21557 7017 21608
rect 7102 21984 7136 22036
rect 7102 21592 7136 21608
rect 7220 21984 7254 22000
rect 7220 21557 7254 21608
rect 7338 21984 7372 22036
rect 7574 22036 7844 22075
rect 7338 21592 7372 21608
rect 7456 21984 7490 22000
rect 7456 21557 7490 21608
rect 7574 21984 7608 22036
rect 7574 21592 7608 21608
rect 7692 21984 7726 22000
rect 7692 21557 7726 21608
rect 7810 21984 7844 22036
rect 8041 22037 8311 22076
rect 7810 21592 7844 21608
rect 7923 21984 7957 22000
rect 7923 21557 7957 21608
rect 8041 21984 8075 22037
rect 8041 21592 8075 21608
rect 8159 21984 8193 22000
rect 8159 21557 8193 21608
rect 8277 21984 8311 22037
rect 9761 22032 10031 22071
rect 9761 21980 9795 22032
rect 8482 21835 8752 21874
rect 8277 21592 8311 21608
rect 8364 21784 8398 21800
rect 6747 21518 8193 21557
rect 8364 21557 8398 21608
rect 8482 21784 8516 21835
rect 8482 21592 8516 21608
rect 8600 21784 8634 21800
rect 8600 21557 8634 21608
rect 8718 21784 8752 21835
rect 8718 21592 8752 21608
rect 9288 21830 9558 21867
rect 9288 21780 9322 21830
rect 9288 21588 9322 21604
rect 9406 21780 9440 21796
rect 8364 21518 8634 21557
rect 9406 21550 9440 21604
rect 9524 21780 9558 21830
rect 9524 21588 9558 21604
rect 9642 21780 9676 21796
rect 9642 21550 9676 21604
rect 9761 21588 9795 21604
rect 9879 21980 9913 21996
rect 9406 21511 9676 21550
rect 9879 21553 9913 21604
rect 9997 21980 10031 22032
rect 10234 22032 10504 22071
rect 9997 21588 10031 21604
rect 10115 21980 10149 21996
rect 10115 21553 10149 21604
rect 10234 21980 10268 22032
rect 10234 21588 10268 21604
rect 10352 21980 10386 21996
rect 10352 21553 10386 21604
rect 10470 21980 10504 22032
rect 10706 22032 10976 22071
rect 10470 21588 10504 21604
rect 10588 21980 10622 21996
rect 10588 21553 10622 21604
rect 10706 21980 10740 22032
rect 10706 21588 10740 21604
rect 10824 21980 10858 21996
rect 10824 21553 10858 21604
rect 10942 21980 10976 22032
rect 11173 22033 11443 22072
rect 10942 21588 10976 21604
rect 11055 21980 11089 21996
rect 11055 21553 11089 21604
rect 11173 21980 11207 22033
rect 11173 21588 11207 21604
rect 11291 21980 11325 21996
rect 11291 21553 11325 21604
rect 11409 21980 11443 22033
rect 12905 22032 13175 22071
rect 12905 21980 12939 22032
rect 11614 21831 11884 21870
rect 11409 21588 11443 21604
rect 11496 21780 11530 21796
rect 9879 21514 11325 21553
rect 11496 21553 11530 21604
rect 11614 21780 11648 21831
rect 11614 21588 11648 21604
rect 11732 21780 11766 21796
rect 11732 21553 11766 21604
rect 11850 21780 11884 21831
rect 11850 21588 11884 21604
rect 12432 21830 12702 21867
rect 12432 21780 12466 21830
rect 12432 21588 12466 21604
rect 12550 21780 12584 21796
rect 11496 21514 11766 21553
rect 12550 21550 12584 21604
rect 12668 21780 12702 21830
rect 12668 21588 12702 21604
rect 12786 21780 12820 21796
rect 12786 21550 12820 21604
rect 12905 21588 12939 21604
rect 13023 21980 13057 21996
rect 12550 21511 12820 21550
rect 13023 21553 13057 21604
rect 13141 21980 13175 22032
rect 13378 22032 13648 22071
rect 13141 21588 13175 21604
rect 13259 21980 13293 21996
rect 13259 21553 13293 21604
rect 13378 21980 13412 22032
rect 13378 21588 13412 21604
rect 13496 21980 13530 21996
rect 13496 21553 13530 21604
rect 13614 21980 13648 22032
rect 13850 22032 14120 22071
rect 13614 21588 13648 21604
rect 13732 21980 13766 21996
rect 13732 21553 13766 21604
rect 13850 21980 13884 22032
rect 13850 21588 13884 21604
rect 13968 21980 14002 21996
rect 13968 21553 14002 21604
rect 14086 21980 14120 22032
rect 14317 22033 14587 22072
rect 14086 21588 14120 21604
rect 14199 21980 14233 21996
rect 14199 21553 14233 21604
rect 14317 21980 14351 22033
rect 14317 21588 14351 21604
rect 14435 21980 14469 21996
rect 14435 21553 14469 21604
rect 14553 21980 14587 22033
rect 16107 22036 16377 22075
rect 16107 21984 16141 22036
rect 14758 21831 15028 21870
rect 14553 21588 14587 21604
rect 14640 21780 14674 21796
rect 13023 21514 14469 21553
rect 14640 21553 14674 21604
rect 14758 21780 14792 21831
rect 14758 21588 14792 21604
rect 14876 21780 14910 21796
rect 14876 21553 14910 21604
rect 14994 21780 15028 21831
rect 14994 21588 15028 21604
rect 15634 21834 15904 21871
rect 15634 21784 15668 21834
rect 15634 21592 15668 21608
rect 15752 21784 15786 21800
rect 14640 21514 14910 21553
rect 15752 21554 15786 21608
rect 15870 21784 15904 21834
rect 15870 21592 15904 21608
rect 15988 21784 16022 21800
rect 15988 21554 16022 21608
rect 16107 21592 16141 21608
rect 16225 21984 16259 22000
rect 15752 21515 16022 21554
rect 16225 21557 16259 21608
rect 16343 21984 16377 22036
rect 16580 22036 16850 22075
rect 16343 21592 16377 21608
rect 16461 21984 16495 22000
rect 16461 21557 16495 21608
rect 16580 21984 16614 22036
rect 16580 21592 16614 21608
rect 16698 21984 16732 22000
rect 16698 21557 16732 21608
rect 16816 21984 16850 22036
rect 17052 22036 17322 22075
rect 16816 21592 16850 21608
rect 16934 21984 16968 22000
rect 16934 21557 16968 21608
rect 17052 21984 17086 22036
rect 17052 21592 17086 21608
rect 17170 21984 17204 22000
rect 17170 21557 17204 21608
rect 17288 21984 17322 22036
rect 17519 22037 17789 22076
rect 17288 21592 17322 21608
rect 17401 21984 17435 22000
rect 17401 21557 17435 21608
rect 17519 21984 17553 22037
rect 17519 21592 17553 21608
rect 17637 21984 17671 22000
rect 17637 21557 17671 21608
rect 17755 21984 17789 22037
rect 19251 22036 19521 22075
rect 19251 21984 19285 22036
rect 17960 21835 18230 21874
rect 17755 21592 17789 21608
rect 17842 21784 17876 21800
rect 16225 21518 17671 21557
rect 17842 21557 17876 21608
rect 17960 21784 17994 21835
rect 17960 21592 17994 21608
rect 18078 21784 18112 21800
rect 18078 21557 18112 21608
rect 18196 21784 18230 21835
rect 18196 21592 18230 21608
rect 18778 21834 19048 21871
rect 18778 21784 18812 21834
rect 18778 21592 18812 21608
rect 18896 21784 18930 21800
rect 17842 21518 18112 21557
rect 18896 21554 18930 21608
rect 19014 21784 19048 21834
rect 19014 21592 19048 21608
rect 19132 21784 19166 21800
rect 19132 21554 19166 21608
rect 19251 21592 19285 21608
rect 19369 21984 19403 22000
rect 18896 21515 19166 21554
rect 19369 21557 19403 21608
rect 19487 21984 19521 22036
rect 19724 22036 19994 22075
rect 19487 21592 19521 21608
rect 19605 21984 19639 22000
rect 19605 21557 19639 21608
rect 19724 21984 19758 22036
rect 19724 21592 19758 21608
rect 19842 21984 19876 22000
rect 19842 21557 19876 21608
rect 19960 21984 19994 22036
rect 20196 22036 20466 22075
rect 19960 21592 19994 21608
rect 20078 21984 20112 22000
rect 20078 21557 20112 21608
rect 20196 21984 20230 22036
rect 20196 21592 20230 21608
rect 20314 21984 20348 22000
rect 20314 21557 20348 21608
rect 20432 21984 20466 22036
rect 20663 22037 20933 22076
rect 20432 21592 20466 21608
rect 20545 21984 20579 22000
rect 20545 21557 20579 21608
rect 20663 21984 20697 22037
rect 20663 21592 20697 21608
rect 20781 21984 20815 22000
rect 20781 21557 20815 21608
rect 20899 21984 20933 22037
rect 22383 22032 22653 22071
rect 22383 21980 22417 22032
rect 21104 21835 21374 21874
rect 20899 21592 20933 21608
rect 20986 21784 21020 21800
rect 19369 21518 20815 21557
rect 20986 21557 21020 21608
rect 21104 21784 21138 21835
rect 21104 21592 21138 21608
rect 21222 21784 21256 21800
rect 21222 21557 21256 21608
rect 21340 21784 21374 21835
rect 21340 21592 21374 21608
rect 21910 21830 22180 21867
rect 21910 21780 21944 21830
rect 21910 21588 21944 21604
rect 22028 21780 22062 21796
rect 20986 21518 21256 21557
rect 22028 21550 22062 21604
rect 22146 21780 22180 21830
rect 22146 21588 22180 21604
rect 22264 21780 22298 21796
rect 22264 21550 22298 21604
rect 22383 21588 22417 21604
rect 22501 21980 22535 21996
rect 22028 21511 22298 21550
rect 22501 21553 22535 21604
rect 22619 21980 22653 22032
rect 22856 22032 23126 22071
rect 22619 21588 22653 21604
rect 22737 21980 22771 21996
rect 22737 21553 22771 21604
rect 22856 21980 22890 22032
rect 22856 21588 22890 21604
rect 22974 21980 23008 21996
rect 22974 21553 23008 21604
rect 23092 21980 23126 22032
rect 23328 22032 23598 22071
rect 23092 21588 23126 21604
rect 23210 21980 23244 21996
rect 23210 21553 23244 21604
rect 23328 21980 23362 22032
rect 23328 21588 23362 21604
rect 23446 21980 23480 21996
rect 23446 21553 23480 21604
rect 23564 21980 23598 22032
rect 23795 22033 24065 22072
rect 23564 21588 23598 21604
rect 23677 21980 23711 21996
rect 23677 21553 23711 21604
rect 23795 21980 23829 22033
rect 23795 21588 23829 21604
rect 23913 21980 23947 21996
rect 23913 21553 23947 21604
rect 24031 21980 24065 22033
rect 25527 22032 25797 22071
rect 25527 21980 25561 22032
rect 24236 21831 24506 21870
rect 24031 21588 24065 21604
rect 24118 21780 24152 21796
rect 22501 21514 23947 21553
rect 24118 21553 24152 21604
rect 24236 21780 24270 21831
rect 24236 21588 24270 21604
rect 24354 21780 24388 21796
rect 24354 21553 24388 21604
rect 24472 21780 24506 21831
rect 24472 21588 24506 21604
rect 25054 21830 25324 21867
rect 25054 21780 25088 21830
rect 25054 21588 25088 21604
rect 25172 21780 25206 21796
rect 24118 21514 24388 21553
rect 25172 21550 25206 21604
rect 25290 21780 25324 21830
rect 25290 21588 25324 21604
rect 25408 21780 25442 21796
rect 25408 21550 25442 21604
rect 25527 21588 25561 21604
rect 25645 21980 25679 21996
rect 25172 21511 25442 21550
rect 25645 21553 25679 21604
rect 25763 21980 25797 22032
rect 26000 22032 26270 22071
rect 25763 21588 25797 21604
rect 25881 21980 25915 21996
rect 25881 21553 25915 21604
rect 26000 21980 26034 22032
rect 26000 21588 26034 21604
rect 26118 21980 26152 21996
rect 26118 21553 26152 21604
rect 26236 21980 26270 22032
rect 26472 22032 26742 22071
rect 26236 21588 26270 21604
rect 26354 21980 26388 21996
rect 26354 21553 26388 21604
rect 26472 21980 26506 22032
rect 26472 21588 26506 21604
rect 26590 21980 26624 21996
rect 26590 21553 26624 21604
rect 26708 21980 26742 22032
rect 26939 22033 27209 22072
rect 26708 21588 26742 21604
rect 26821 21980 26855 21996
rect 26821 21553 26855 21604
rect 26939 21980 26973 22033
rect 26939 21588 26973 21604
rect 27057 21980 27091 21996
rect 27057 21553 27091 21604
rect 27175 21980 27209 22033
rect 27380 21831 27650 21870
rect 27175 21588 27209 21604
rect 27262 21780 27296 21796
rect 25645 21514 27091 21553
rect 27262 21553 27296 21604
rect 27380 21780 27414 21831
rect 27380 21588 27414 21604
rect 27498 21780 27532 21796
rect 27498 21553 27532 21604
rect 27616 21780 27650 21831
rect 27616 21588 27650 21604
rect 27262 21514 27532 21553
rect 28274 21445 28352 24096
rect 39837 24084 39871 24100
rect 27937 21436 28352 21445
rect 3162 21400 3178 21434
rect 3212 21400 3228 21434
rect 4488 21393 4522 21409
rect 6306 21400 6322 21434
rect 6356 21400 6372 21434
rect 4488 21343 4522 21359
rect 7632 21393 7666 21409
rect 9438 21396 9454 21430
rect 9488 21396 9504 21430
rect 7632 21343 7666 21359
rect 10764 21389 10798 21405
rect 12582 21396 12598 21430
rect 12632 21396 12648 21430
rect 10764 21339 10798 21355
rect 13908 21389 13942 21405
rect 15784 21400 15800 21434
rect 15834 21400 15850 21434
rect 13908 21339 13942 21355
rect 17110 21393 17144 21409
rect 18928 21400 18944 21434
rect 18978 21400 18994 21434
rect 17110 21343 17144 21359
rect 20254 21393 20288 21409
rect 22060 21396 22076 21430
rect 22110 21396 22126 21430
rect 20254 21343 20288 21359
rect 23386 21389 23420 21405
rect 25204 21396 25220 21430
rect 25254 21396 25270 21430
rect 23386 21339 23420 21355
rect 26530 21389 26564 21405
rect 27937 21392 27950 21436
rect 28042 21392 28352 21436
rect 27937 21381 28352 21392
rect 28402 24042 28480 24053
rect 28402 23975 28412 24042
rect 28469 23975 28480 24042
rect 26530 21339 26564 21355
rect 4342 21294 4434 21307
rect 4342 21239 4358 21294
rect 4418 21239 4434 21294
rect 4342 21222 4434 21239
rect 5427 21293 5519 21310
rect 5427 21238 5443 21293
rect 5503 21238 5519 21293
rect 5427 21225 5519 21238
rect 7486 21294 7578 21307
rect 7486 21239 7502 21294
rect 7562 21239 7578 21294
rect 7486 21222 7578 21239
rect 8571 21293 8663 21310
rect 8571 21238 8587 21293
rect 8647 21238 8663 21293
rect 8571 21225 8663 21238
rect 10618 21290 10710 21303
rect 10618 21235 10634 21290
rect 10694 21235 10710 21290
rect 10618 21218 10710 21235
rect 11703 21289 11795 21306
rect 11703 21234 11719 21289
rect 11779 21234 11795 21289
rect 11703 21221 11795 21234
rect 13762 21290 13854 21303
rect 13762 21235 13778 21290
rect 13838 21235 13854 21290
rect 13762 21218 13854 21235
rect 14847 21289 14939 21306
rect 14847 21234 14863 21289
rect 14923 21234 14939 21289
rect 14847 21221 14939 21234
rect 16964 21294 17056 21307
rect 16964 21239 16980 21294
rect 17040 21239 17056 21294
rect 16964 21222 17056 21239
rect 18049 21293 18141 21310
rect 18049 21238 18065 21293
rect 18125 21238 18141 21293
rect 18049 21225 18141 21238
rect 20108 21294 20200 21307
rect 20108 21239 20124 21294
rect 20184 21239 20200 21294
rect 20108 21222 20200 21239
rect 21193 21293 21285 21310
rect 21193 21238 21209 21293
rect 21269 21238 21285 21293
rect 21193 21225 21285 21238
rect 23240 21290 23332 21303
rect 23240 21235 23256 21290
rect 23316 21235 23332 21290
rect 23240 21218 23332 21235
rect 24325 21289 24417 21306
rect 24325 21234 24341 21289
rect 24401 21234 24417 21289
rect 24325 21221 24417 21234
rect 26384 21290 26476 21303
rect 26384 21235 26400 21290
rect 26460 21235 26476 21290
rect 26384 21218 26476 21235
rect 27469 21289 27561 21306
rect 27469 21234 27485 21289
rect 27545 21234 27561 21289
rect 27469 21221 27561 21234
rect 27736 21290 27793 21294
rect 27736 21230 27740 21290
rect 27789 21230 27793 21290
rect 27736 21226 27793 21230
rect 4134 21163 4168 21179
rect 4134 21113 4168 21129
rect 5694 21178 5945 21182
rect 5694 21118 5698 21178
rect 5747 21118 5945 21178
rect 5694 21114 5945 21118
rect 4460 21009 4552 21022
rect 4460 20954 4476 21009
rect 4536 20954 4552 21009
rect 4460 20937 4552 20954
rect 5888 20888 5945 21114
rect 7278 21163 7312 21179
rect 7278 21113 7312 21129
rect 8838 21178 8895 21182
rect 11994 21178 12248 21179
rect 8838 21118 8842 21178
rect 8891 21118 8895 21178
rect 8838 21114 8895 21118
rect 10410 21159 10444 21175
rect 10410 21109 10444 21125
rect 11970 21174 12248 21178
rect 11970 21114 11974 21174
rect 12023 21114 12248 21174
rect 11970 21110 12248 21114
rect 7604 21009 7696 21022
rect 7604 20954 7620 21009
rect 7680 20954 7696 21009
rect 7604 20937 7696 20954
rect 8838 21010 8895 21014
rect 8838 20950 8842 21010
rect 8891 20950 8895 21010
rect 8838 20946 8895 20950
rect 9891 21005 10828 21018
rect 9891 20950 10752 21005
rect 10812 20950 10828 21005
rect 9891 20933 10828 20950
rect 11970 21006 12027 21010
rect 11970 20946 11974 21006
rect 12023 20946 12027 21006
rect 11970 20942 12027 20946
rect 9891 20888 9966 20933
rect 5888 20823 9966 20888
rect 12180 20882 12248 21110
rect 13554 21159 13588 21175
rect 13554 21109 13588 21125
rect 16756 21163 16790 21179
rect 16756 21113 16790 21129
rect 18304 21178 18499 21182
rect 18304 21118 18320 21178
rect 18369 21118 18499 21178
rect 18304 21110 18499 21118
rect 19900 21163 19934 21179
rect 19900 21113 19934 21129
rect 23032 21159 23066 21175
rect 18441 21107 18499 21110
rect 23032 21109 23066 21125
rect 24592 21174 24649 21178
rect 24592 21114 24596 21174
rect 24645 21114 24649 21174
rect 24592 21110 24649 21114
rect 26176 21159 26210 21175
rect 26176 21109 26210 21125
rect 18441 21050 18672 21107
rect 13880 21005 13972 21018
rect 13880 20950 13896 21005
rect 13956 20950 13972 21005
rect 13880 20933 13972 20950
rect 15114 21006 15171 21010
rect 15114 20946 15118 21006
rect 15167 20946 15171 21006
rect 15114 20942 15171 20946
rect 16302 21009 17174 21022
rect 16302 20954 17098 21009
rect 17158 20954 17174 21009
rect 16302 20937 17174 20954
rect 18316 21010 18373 21014
rect 18316 20950 18320 21010
rect 18369 20950 18373 21010
rect 18316 20946 18373 20950
rect 16302 20882 16379 20937
rect 12180 20820 16379 20882
rect 18595 20876 18672 21050
rect 20226 21009 20318 21022
rect 28402 21019 28480 23975
rect 20226 20954 20242 21009
rect 20302 20954 20318 21009
rect 20226 20937 20318 20954
rect 21460 21010 21517 21014
rect 21460 20950 21464 21010
rect 21513 20950 21517 21010
rect 21460 20946 21517 20950
rect 22043 21005 23450 21018
rect 22043 20950 23374 21005
rect 23434 20950 23450 21005
rect 22043 20933 23450 20950
rect 24592 21006 24649 21010
rect 24592 20946 24596 21006
rect 24645 20946 24649 21006
rect 24592 20942 24649 20946
rect 26502 21005 26594 21018
rect 26502 20950 26518 21005
rect 26578 20950 26594 21005
rect 26502 20933 26594 20950
rect 27736 21006 27793 21010
rect 27736 20946 27740 21006
rect 27789 20946 27793 21006
rect 27736 20942 27793 20946
rect 27938 20998 28480 21019
rect 27938 20954 27950 20998
rect 28042 20954 28480 20998
rect 22043 20876 22123 20933
rect 27938 20932 28480 20954
rect 28524 23924 28602 23935
rect 28524 23857 28534 23924
rect 28591 23857 28602 23924
rect 18595 20823 22123 20876
rect 28524 20861 28602 23857
rect 28524 20820 28541 20861
rect 28591 20820 28602 20861
rect 4253 20773 4287 20789
rect 4253 20723 4287 20739
rect 7397 20773 7431 20789
rect 7397 20723 7431 20739
rect 10529 20769 10563 20785
rect 10529 20719 10563 20735
rect 13673 20769 13707 20785
rect 13673 20719 13707 20735
rect 16875 20773 16909 20789
rect 16875 20723 16909 20739
rect 20019 20773 20053 20789
rect 20019 20723 20053 20739
rect 23151 20769 23185 20785
rect 23151 20719 23185 20735
rect 26295 20769 26329 20785
rect 28524 20777 28602 20820
rect 28647 23802 28725 23813
rect 28647 23735 28658 23802
rect 28715 23735 28725 23802
rect 28524 20770 28603 20777
rect 26295 20719 26329 20735
rect 27936 20758 28603 20770
rect 27936 20714 27950 20758
rect 28042 20714 28603 20758
rect 27936 20705 28603 20714
rect 3880 20651 3914 20667
rect 3880 20459 3914 20475
rect 3998 20663 4032 20667
rect 4076 20663 4110 20667
rect 3998 20651 4110 20663
rect 4032 20475 4076 20651
rect 3998 20463 4076 20475
rect 3998 20459 4032 20463
rect 4076 20259 4110 20275
rect 4194 20651 4228 20667
rect 4194 20259 4228 20275
rect 4312 20651 4346 20667
rect 4312 20259 4346 20275
rect 4430 20651 4464 20667
rect 4430 20259 4464 20275
rect 4548 20663 4582 20667
rect 4622 20663 4656 20667
rect 4548 20651 4656 20663
rect 4582 20475 4622 20651
rect 4582 20463 4656 20475
rect 4622 20459 4656 20463
rect 4740 20651 4774 20667
rect 4740 20459 4774 20475
rect 7024 20651 7058 20667
rect 7024 20459 7058 20475
rect 7142 20663 7176 20667
rect 7220 20663 7254 20667
rect 7142 20651 7254 20663
rect 7176 20475 7220 20651
rect 7142 20463 7220 20475
rect 7142 20459 7176 20463
rect 4548 20259 4582 20275
rect 7220 20259 7254 20275
rect 7338 20651 7372 20667
rect 7338 20259 7372 20275
rect 7456 20651 7490 20667
rect 7456 20259 7490 20275
rect 7574 20651 7608 20667
rect 7574 20259 7608 20275
rect 7692 20663 7726 20667
rect 7766 20663 7800 20667
rect 7692 20651 7800 20663
rect 7726 20475 7766 20651
rect 7726 20463 7800 20475
rect 7766 20459 7800 20463
rect 7884 20651 7918 20667
rect 7884 20459 7918 20475
rect 10156 20647 10190 20663
rect 10156 20455 10190 20471
rect 10274 20659 10308 20663
rect 10352 20659 10386 20663
rect 10274 20647 10386 20659
rect 10308 20471 10352 20647
rect 10274 20459 10352 20471
rect 10274 20455 10308 20459
rect 7692 20259 7726 20275
rect 10352 20255 10386 20271
rect 10470 20647 10504 20663
rect 10470 20255 10504 20271
rect 10588 20647 10622 20663
rect 10588 20255 10622 20271
rect 10706 20647 10740 20663
rect 10706 20255 10740 20271
rect 10824 20659 10858 20663
rect 10898 20659 10932 20663
rect 10824 20647 10932 20659
rect 10858 20471 10898 20647
rect 10858 20459 10932 20471
rect 10898 20455 10932 20459
rect 11016 20647 11050 20663
rect 11016 20455 11050 20471
rect 13300 20647 13334 20663
rect 13300 20455 13334 20471
rect 13418 20659 13452 20663
rect 13496 20659 13530 20663
rect 13418 20647 13530 20659
rect 13452 20471 13496 20647
rect 13418 20459 13496 20471
rect 13418 20455 13452 20459
rect 10824 20255 10858 20271
rect 13496 20255 13530 20271
rect 13614 20647 13648 20663
rect 13614 20255 13648 20271
rect 13732 20647 13766 20663
rect 13732 20255 13766 20271
rect 13850 20647 13884 20663
rect 13850 20255 13884 20271
rect 13968 20659 14002 20663
rect 14042 20659 14076 20663
rect 13968 20647 14076 20659
rect 14002 20471 14042 20647
rect 14002 20459 14076 20471
rect 14042 20455 14076 20459
rect 14160 20647 14194 20663
rect 14160 20455 14194 20471
rect 16502 20651 16536 20667
rect 16502 20459 16536 20475
rect 16620 20663 16654 20667
rect 16698 20663 16732 20667
rect 16620 20651 16732 20663
rect 16654 20475 16698 20651
rect 16620 20463 16698 20475
rect 16620 20459 16654 20463
rect 13968 20255 14002 20271
rect 16698 20259 16732 20275
rect 16816 20651 16850 20667
rect 16816 20259 16850 20275
rect 16934 20651 16968 20667
rect 16934 20259 16968 20275
rect 17052 20651 17086 20667
rect 17052 20259 17086 20275
rect 17170 20663 17204 20667
rect 17244 20663 17278 20667
rect 17170 20651 17278 20663
rect 17204 20475 17244 20651
rect 17204 20463 17278 20475
rect 17244 20459 17278 20463
rect 17362 20651 17396 20667
rect 17362 20459 17396 20475
rect 19646 20651 19680 20667
rect 19646 20459 19680 20475
rect 19764 20663 19798 20667
rect 19842 20663 19876 20667
rect 19764 20651 19876 20663
rect 19798 20475 19842 20651
rect 19764 20463 19842 20475
rect 19764 20459 19798 20463
rect 17170 20259 17204 20275
rect 19842 20259 19876 20275
rect 19960 20651 19994 20667
rect 19960 20259 19994 20275
rect 20078 20651 20112 20667
rect 20078 20259 20112 20275
rect 20196 20651 20230 20667
rect 20196 20259 20230 20275
rect 20314 20663 20348 20667
rect 20388 20663 20422 20667
rect 20314 20651 20422 20663
rect 20348 20475 20388 20651
rect 20348 20463 20422 20475
rect 20388 20459 20422 20463
rect 20506 20651 20540 20667
rect 20506 20459 20540 20475
rect 22778 20647 22812 20663
rect 22778 20455 22812 20471
rect 22896 20659 22930 20663
rect 22974 20659 23008 20663
rect 22896 20647 23008 20659
rect 22930 20471 22974 20647
rect 22896 20459 22974 20471
rect 22896 20455 22930 20459
rect 20314 20259 20348 20275
rect 22974 20255 23008 20271
rect 23092 20647 23126 20663
rect 23092 20255 23126 20271
rect 23210 20647 23244 20663
rect 23210 20255 23244 20271
rect 23328 20647 23362 20663
rect 23328 20255 23362 20271
rect 23446 20659 23480 20663
rect 23520 20659 23554 20663
rect 23446 20647 23554 20659
rect 23480 20471 23520 20647
rect 23480 20459 23554 20471
rect 23520 20455 23554 20459
rect 23638 20647 23672 20663
rect 23638 20455 23672 20471
rect 25922 20647 25956 20663
rect 25922 20455 25956 20471
rect 26040 20659 26074 20663
rect 26118 20659 26152 20663
rect 26040 20647 26152 20659
rect 26074 20471 26118 20647
rect 26040 20459 26118 20471
rect 26040 20455 26074 20459
rect 23446 20255 23480 20271
rect 26118 20255 26152 20271
rect 26236 20647 26270 20663
rect 26236 20255 26270 20271
rect 26354 20647 26388 20663
rect 26354 20255 26388 20271
rect 26472 20647 26506 20663
rect 26472 20255 26506 20271
rect 26590 20659 26624 20663
rect 26664 20659 26698 20663
rect 26590 20647 26698 20659
rect 26624 20471 26664 20647
rect 26624 20459 26698 20471
rect 26664 20455 26698 20459
rect 26782 20647 26816 20663
rect 28647 20634 28725 23735
rect 28772 23683 28850 23694
rect 39837 23692 39871 23708
rect 39955 24084 39989 24100
rect 39955 23692 39989 23708
rect 40073 24084 40107 24100
rect 40190 24084 40224 24100
rect 40190 23892 40224 23908
rect 40308 24084 40342 24100
rect 40308 23892 40342 23908
rect 46350 24081 46384 24097
rect 42114 23861 42130 23895
rect 42164 23861 42180 23895
rect 43256 23865 43272 23899
rect 43306 23865 43322 23899
rect 41835 23810 41869 23826
rect 40073 23692 40107 23708
rect 40360 23758 40609 23801
rect 28772 23616 28780 23683
rect 28837 23616 28850 23683
rect 40360 23668 40407 23758
rect 40570 23668 40609 23758
rect 39880 23624 39896 23658
rect 39930 23624 39946 23658
rect 39998 23624 40014 23658
rect 40048 23624 40064 23658
rect 40360 23629 40609 23668
rect 41835 23618 41869 23634
rect 41953 23810 41987 23826
rect 41953 23618 41987 23634
rect 42071 23810 42105 23826
rect 42071 23618 42105 23634
rect 42189 23810 42223 23826
rect 42189 23618 42223 23634
rect 42354 23810 42388 23826
rect 42354 23618 42388 23634
rect 42472 23810 42506 23826
rect 42472 23618 42506 23634
rect 42590 23810 42624 23826
rect 42590 23618 42624 23634
rect 42708 23810 42742 23826
rect 42708 23618 42742 23634
rect 42977 23814 43011 23830
rect 42977 23622 43011 23638
rect 43095 23814 43129 23830
rect 43095 23622 43129 23638
rect 43213 23814 43247 23830
rect 43213 23622 43247 23638
rect 43331 23814 43365 23830
rect 43331 23622 43365 23638
rect 43496 23814 43530 23830
rect 43496 23622 43530 23638
rect 43614 23814 43648 23830
rect 43614 23622 43648 23638
rect 43732 23814 43766 23830
rect 43732 23622 43766 23638
rect 43850 23814 43884 23830
rect 46350 23689 46384 23705
rect 46468 24081 46502 24097
rect 46468 23689 46502 23705
rect 46586 24081 46620 24097
rect 46703 24081 46737 24097
rect 46703 23889 46737 23905
rect 46821 24081 46855 24097
rect 46821 23889 46855 23905
rect 52884 24076 52918 24092
rect 48627 23858 48643 23892
rect 48677 23858 48693 23892
rect 49769 23862 49785 23896
rect 49819 23862 49835 23896
rect 48348 23807 48382 23823
rect 46586 23689 46620 23705
rect 46873 23755 47122 23798
rect 46873 23665 46920 23755
rect 47083 23665 47122 23755
rect 43850 23622 43884 23638
rect 46393 23621 46409 23655
rect 46443 23621 46459 23655
rect 46511 23621 46527 23655
rect 46561 23621 46577 23655
rect 46873 23626 47122 23665
rect 28772 23285 28850 23616
rect 48348 23615 48382 23631
rect 48466 23807 48500 23823
rect 48466 23615 48500 23631
rect 48584 23807 48618 23823
rect 48584 23615 48618 23631
rect 48702 23807 48736 23823
rect 48702 23615 48736 23631
rect 48867 23807 48901 23823
rect 48867 23615 48901 23631
rect 48985 23807 49019 23823
rect 48985 23615 49019 23631
rect 49103 23807 49137 23823
rect 49103 23615 49137 23631
rect 49221 23807 49255 23823
rect 49221 23615 49255 23631
rect 49490 23811 49524 23827
rect 49490 23619 49524 23635
rect 49608 23811 49642 23827
rect 49608 23619 49642 23635
rect 49726 23811 49760 23827
rect 49726 23619 49760 23635
rect 49844 23811 49878 23827
rect 49844 23619 49878 23635
rect 50009 23811 50043 23827
rect 50009 23619 50043 23635
rect 50127 23811 50161 23827
rect 50127 23619 50161 23635
rect 50245 23811 50279 23827
rect 50245 23619 50279 23635
rect 50363 23811 50397 23827
rect 52884 23684 52918 23700
rect 53002 24076 53036 24092
rect 53002 23684 53036 23700
rect 53120 24076 53154 24092
rect 53237 24076 53271 24092
rect 53237 23884 53271 23900
rect 53355 24076 53389 24092
rect 53355 23884 53389 23900
rect 59442 24080 59476 24096
rect 55161 23853 55177 23887
rect 55211 23853 55227 23887
rect 56303 23857 56319 23891
rect 56353 23857 56369 23891
rect 54882 23802 54916 23818
rect 53120 23684 53154 23700
rect 53407 23750 53656 23793
rect 53407 23660 53454 23750
rect 53617 23660 53656 23750
rect 50363 23619 50397 23635
rect 52927 23616 52943 23650
rect 52977 23616 52993 23650
rect 53045 23616 53061 23650
rect 53095 23616 53111 23650
rect 53407 23621 53656 23660
rect 54882 23610 54916 23626
rect 55000 23802 55034 23818
rect 55000 23610 55034 23626
rect 55118 23802 55152 23818
rect 55118 23610 55152 23626
rect 55236 23802 55270 23818
rect 55236 23610 55270 23626
rect 55401 23802 55435 23818
rect 55401 23610 55435 23626
rect 55519 23802 55553 23818
rect 55519 23610 55553 23626
rect 55637 23802 55671 23818
rect 55637 23610 55671 23626
rect 55755 23802 55789 23818
rect 55755 23610 55789 23626
rect 56024 23806 56058 23822
rect 56024 23614 56058 23630
rect 56142 23806 56176 23822
rect 56142 23614 56176 23630
rect 56260 23806 56294 23822
rect 56260 23614 56294 23630
rect 56378 23806 56412 23822
rect 56378 23614 56412 23630
rect 56543 23806 56577 23822
rect 56543 23614 56577 23630
rect 56661 23806 56695 23822
rect 56661 23614 56695 23630
rect 56779 23806 56813 23822
rect 56779 23614 56813 23630
rect 56897 23806 56931 23822
rect 59442 23688 59476 23704
rect 59560 24080 59594 24096
rect 59560 23688 59594 23704
rect 59678 24080 59712 24096
rect 59795 24080 59829 24096
rect 59795 23888 59829 23904
rect 59913 24080 59947 24096
rect 59913 23888 59947 23904
rect 61719 23857 61735 23891
rect 61769 23857 61785 23891
rect 62861 23861 62877 23895
rect 62911 23861 62927 23895
rect 61440 23806 61474 23822
rect 59678 23688 59712 23704
rect 59965 23754 60214 23797
rect 59965 23664 60012 23754
rect 60175 23664 60214 23754
rect 56897 23614 56931 23630
rect 59485 23620 59501 23654
rect 59535 23620 59551 23654
rect 59603 23620 59619 23654
rect 59653 23620 59669 23654
rect 59965 23625 60214 23664
rect 61440 23614 61474 23630
rect 61558 23806 61592 23822
rect 61558 23614 61592 23630
rect 61676 23806 61710 23822
rect 61676 23614 61710 23630
rect 61794 23806 61828 23822
rect 61794 23614 61828 23630
rect 61959 23806 61993 23822
rect 61959 23614 61993 23630
rect 62077 23806 62111 23822
rect 62077 23614 62111 23630
rect 62195 23806 62229 23822
rect 62195 23614 62229 23630
rect 62313 23806 62347 23822
rect 62313 23614 62347 23630
rect 62582 23810 62616 23826
rect 62582 23618 62616 23634
rect 62700 23810 62734 23826
rect 62700 23618 62734 23634
rect 62818 23810 62852 23826
rect 62818 23618 62852 23634
rect 62936 23810 62970 23826
rect 62936 23618 62970 23634
rect 63101 23810 63135 23826
rect 63101 23618 63135 23634
rect 63219 23810 63253 23826
rect 63219 23618 63253 23634
rect 63337 23810 63371 23826
rect 63337 23618 63371 23634
rect 63455 23810 63489 23826
rect 63455 23618 63489 23634
rect 41850 23387 42022 23434
rect 27936 20622 28725 20634
rect 27936 20578 27951 20622
rect 28043 20578 28725 20622
rect 27936 20571 28725 20578
rect 28770 21302 28850 23285
rect 40009 23285 40232 23361
rect 40009 23136 40088 23285
rect 40155 23136 40232 23285
rect 41850 23224 41889 23387
rect 41979 23224 42022 23387
rect 41850 23185 42022 23224
rect 42992 23385 43164 23432
rect 42992 23222 43031 23385
rect 43121 23222 43164 23385
rect 48363 23384 48535 23431
rect 42992 23183 43164 23222
rect 46522 23282 46745 23358
rect 40009 23030 40232 23136
rect 46522 23133 46601 23282
rect 46668 23133 46745 23282
rect 48363 23221 48402 23384
rect 48492 23221 48535 23384
rect 48363 23182 48535 23221
rect 49505 23382 49677 23429
rect 49505 23219 49544 23382
rect 49634 23219 49677 23382
rect 54897 23379 55069 23426
rect 49505 23180 49677 23219
rect 53056 23277 53279 23353
rect 46522 23027 46745 23133
rect 53056 23128 53135 23277
rect 53202 23128 53279 23277
rect 54897 23216 54936 23379
rect 55026 23216 55069 23379
rect 54897 23177 55069 23216
rect 56039 23377 56211 23424
rect 56039 23214 56078 23377
rect 56168 23214 56211 23377
rect 61455 23383 61627 23430
rect 56039 23175 56211 23214
rect 59614 23281 59837 23357
rect 53056 23022 53279 23128
rect 59614 23132 59693 23281
rect 59760 23132 59837 23281
rect 61455 23220 61494 23383
rect 61584 23220 61627 23383
rect 61455 23181 61627 23220
rect 62597 23381 62769 23428
rect 62597 23218 62636 23381
rect 62726 23218 62769 23381
rect 62597 23179 62769 23218
rect 59614 23026 59837 23132
rect 40440 22921 40710 22955
rect 39614 22871 39648 22887
rect 33812 22852 33883 22859
rect 33812 22803 33822 22852
rect 33876 22803 33883 22852
rect 33658 22431 33743 22440
rect 33658 22360 33666 22431
rect 33735 22360 33743 22431
rect 28899 22039 28980 22049
rect 28899 21963 28910 22039
rect 28970 21988 28980 22039
rect 33511 22007 33601 22016
rect 28970 21963 28979 21988
rect 28770 20523 28848 21302
rect 26782 20455 26816 20471
rect 27936 20512 28848 20523
rect 27936 20468 27950 20512
rect 28042 20468 28848 20512
rect 27936 20459 28848 20468
rect 28899 20397 28979 21963
rect 33511 21936 33519 22007
rect 33590 21936 33601 22007
rect 27937 20385 28979 20397
rect 27937 20341 27949 20385
rect 28042 20341 28979 20385
rect 27937 20334 28979 20341
rect 29036 21584 29116 21604
rect 29036 21508 29049 21584
rect 29109 21508 29116 21584
rect 26590 20255 26624 20271
rect 4295 20140 4311 20174
rect 4345 20140 4361 20174
rect 7439 20140 7455 20174
rect 7489 20140 7505 20174
rect 10571 20136 10587 20170
rect 10621 20136 10637 20170
rect 13715 20136 13731 20170
rect 13765 20136 13781 20170
rect 16917 20140 16933 20174
rect 16967 20140 16983 20174
rect 20061 20140 20077 20174
rect 20111 20140 20127 20174
rect 23193 20136 23209 20170
rect 23243 20136 23259 20170
rect 26337 20136 26353 20170
rect 26387 20136 26403 20170
rect 29036 20156 29116 21508
rect 33364 21547 33458 21560
rect 33364 21486 33376 21547
rect 33447 21486 33458 21547
rect 27937 20147 29116 20156
rect 27937 20103 27949 20147
rect 28042 20103 29116 20147
rect 27937 20092 29116 20103
rect 29183 21165 29263 21177
rect 29183 21089 29192 21165
rect 29252 21089 29263 21165
rect 4244 20022 4380 20026
rect 4244 20008 4284 20022
rect 4342 20008 4380 20022
rect 4244 19962 4260 20008
rect 4364 19962 4380 20008
rect 4244 19940 4380 19962
rect 7388 20022 7524 20026
rect 16866 20022 17002 20026
rect 7388 20008 7428 20022
rect 7486 20008 7524 20022
rect 7388 19962 7404 20008
rect 7508 19962 7524 20008
rect 7388 19940 7524 19962
rect 10520 20018 10656 20022
rect 10520 20004 10560 20018
rect 10618 20004 10656 20018
rect 10520 19958 10536 20004
rect 10640 19958 10656 20004
rect 10520 19936 10656 19958
rect 13664 20018 13800 20022
rect 13664 20004 13704 20018
rect 13762 20004 13800 20018
rect 13664 19958 13680 20004
rect 13784 19958 13800 20004
rect 13664 19936 13800 19958
rect 16866 20008 16906 20022
rect 16964 20008 17002 20022
rect 16866 19962 16882 20008
rect 16986 19962 17002 20008
rect 16866 19940 17002 19962
rect 20010 20022 20146 20026
rect 20010 20008 20050 20022
rect 20108 20008 20146 20022
rect 20010 19962 20026 20008
rect 20130 19962 20146 20008
rect 20010 19940 20146 19962
rect 23142 20018 23278 20022
rect 23142 20004 23182 20018
rect 23240 20004 23278 20018
rect 23142 19958 23158 20004
rect 23262 19958 23278 20004
rect 23142 19936 23278 19958
rect 26286 20018 26422 20022
rect 26286 20004 26326 20018
rect 26384 20004 26422 20018
rect 26286 19958 26302 20004
rect 26406 19958 26422 20004
rect 26286 19936 26422 19958
rect 29183 19935 29263 21089
rect 27937 19923 29263 19935
rect 27937 19879 27948 19923
rect 28041 19879 29263 19923
rect 27937 19871 29263 19879
rect 4562 17048 4766 17060
rect 4562 16976 4590 17048
rect 4734 16976 4766 17048
rect 4562 16974 4624 16976
rect 4704 16974 4766 16976
rect 4562 16958 4766 16974
rect 5730 17048 5934 17060
rect 5730 16976 5758 17048
rect 5902 16976 5934 17048
rect 5730 16974 5792 16976
rect 5872 16974 5934 16976
rect 5302 16936 5318 16970
rect 5352 16936 5368 16970
rect 5730 16958 5934 16974
rect 6898 17048 7102 17060
rect 6898 16976 6926 17048
rect 7070 16976 7102 17048
rect 6898 16974 6960 16976
rect 7040 16974 7102 16976
rect 6470 16936 6486 16970
rect 6520 16936 6536 16970
rect 6898 16958 7102 16974
rect 8066 17048 8270 17060
rect 8066 16976 8094 17048
rect 8238 16976 8270 17048
rect 8066 16974 8128 16976
rect 8208 16974 8270 16976
rect 7638 16936 7654 16970
rect 7688 16936 7704 16970
rect 8066 16958 8270 16974
rect 9240 17046 9444 17058
rect 9240 16974 9268 17046
rect 9412 16974 9444 17046
rect 9240 16972 9302 16974
rect 9382 16972 9444 16974
rect 8806 16936 8822 16970
rect 8856 16936 8872 16970
rect 9240 16956 9444 16972
rect 10408 17046 10612 17058
rect 10408 16974 10436 17046
rect 10580 16974 10612 17046
rect 10408 16972 10470 16974
rect 10550 16972 10612 16974
rect 9980 16934 9996 16968
rect 10030 16934 10046 16968
rect 10408 16956 10612 16972
rect 11576 17046 11780 17058
rect 11576 16974 11604 17046
rect 11748 16974 11780 17046
rect 11576 16972 11638 16974
rect 11718 16972 11780 16974
rect 11148 16934 11164 16968
rect 11198 16934 11214 16968
rect 11576 16956 11780 16972
rect 12744 17046 12948 17058
rect 12744 16974 12772 17046
rect 12916 16974 12948 17046
rect 12744 16972 12806 16974
rect 12886 16972 12948 16974
rect 12316 16934 12332 16968
rect 12366 16934 12382 16968
rect 12744 16956 12948 16972
rect 13484 16934 13500 16968
rect 13534 16934 13550 16968
rect 5302 16828 5318 16862
rect 5352 16828 5368 16862
rect 6470 16828 6486 16862
rect 6520 16828 6536 16862
rect 7638 16828 7654 16862
rect 7688 16828 7704 16862
rect 8806 16828 8822 16862
rect 8856 16828 8872 16862
rect 9980 16826 9996 16860
rect 10030 16826 10046 16860
rect 11148 16826 11164 16860
rect 11198 16826 11214 16860
rect 12316 16826 12332 16860
rect 12366 16826 12382 16860
rect 13484 16826 13500 16860
rect 13534 16826 13550 16860
rect 14442 16841 14610 16857
rect 4520 16796 4554 16812
rect 4520 16404 4554 16420
rect 4638 16796 4672 16812
rect 4638 16404 4672 16420
rect 4756 16796 4790 16812
rect 4756 16404 4790 16420
rect 4874 16796 4908 16812
rect 4874 16404 4908 16420
rect 4992 16796 5026 16812
rect 4992 16404 5026 16420
rect 5110 16796 5144 16812
rect 5110 16404 5144 16420
rect 5228 16796 5262 16812
rect 5228 16404 5262 16420
rect 5688 16798 5722 16814
rect 5688 16406 5722 16422
rect 5806 16798 5840 16814
rect 5806 16406 5840 16422
rect 5924 16798 5958 16814
rect 5924 16406 5958 16422
rect 6042 16798 6076 16814
rect 6042 16406 6076 16422
rect 6160 16798 6194 16814
rect 6160 16406 6194 16422
rect 6278 16798 6312 16814
rect 6278 16406 6312 16422
rect 6396 16798 6430 16814
rect 6396 16406 6430 16422
rect 6856 16796 6890 16812
rect 6856 16404 6890 16420
rect 6974 16796 7008 16812
rect 6974 16404 7008 16420
rect 7092 16796 7126 16812
rect 7092 16404 7126 16420
rect 7210 16796 7244 16812
rect 7210 16404 7244 16420
rect 7328 16796 7362 16812
rect 7328 16404 7362 16420
rect 7446 16796 7480 16812
rect 7446 16404 7480 16420
rect 7564 16796 7598 16812
rect 7564 16404 7598 16420
rect 8024 16798 8058 16814
rect 8024 16406 8058 16422
rect 8142 16798 8176 16814
rect 8142 16406 8176 16422
rect 8260 16798 8294 16814
rect 8260 16406 8294 16422
rect 8378 16798 8412 16814
rect 8378 16406 8412 16422
rect 8496 16798 8530 16814
rect 8496 16406 8530 16422
rect 8614 16798 8648 16814
rect 8614 16406 8648 16422
rect 8732 16798 8766 16814
rect 8732 16406 8766 16422
rect 9198 16796 9232 16812
rect 9198 16404 9232 16420
rect 9316 16796 9350 16812
rect 9316 16404 9350 16420
rect 9434 16796 9468 16812
rect 9434 16404 9468 16420
rect 9552 16796 9586 16812
rect 9552 16404 9586 16420
rect 9670 16796 9704 16812
rect 9670 16404 9704 16420
rect 9788 16796 9822 16812
rect 9788 16404 9822 16420
rect 9906 16796 9940 16812
rect 9906 16404 9940 16420
rect 10366 16794 10400 16810
rect 10366 16402 10400 16418
rect 10484 16794 10518 16810
rect 10484 16402 10518 16418
rect 10602 16794 10636 16810
rect 10602 16402 10636 16418
rect 10720 16794 10754 16810
rect 10720 16402 10754 16418
rect 10838 16794 10872 16810
rect 10838 16402 10872 16418
rect 10956 16794 10990 16810
rect 10956 16402 10990 16418
rect 11074 16794 11108 16810
rect 11074 16402 11108 16418
rect 11534 16796 11568 16812
rect 11534 16404 11568 16420
rect 11652 16796 11686 16812
rect 11652 16404 11686 16420
rect 11770 16796 11804 16812
rect 11770 16404 11804 16420
rect 11888 16796 11922 16812
rect 11888 16404 11922 16420
rect 12006 16796 12040 16812
rect 12006 16404 12040 16420
rect 12124 16796 12158 16812
rect 12124 16404 12158 16420
rect 12242 16796 12276 16812
rect 12242 16404 12276 16420
rect 12702 16796 12736 16812
rect 12702 16404 12736 16420
rect 12820 16796 12854 16812
rect 12820 16404 12854 16420
rect 12938 16796 12972 16812
rect 12938 16404 12972 16420
rect 13056 16796 13090 16812
rect 13056 16404 13090 16420
rect 13174 16796 13208 16812
rect 13174 16404 13208 16420
rect 13292 16796 13326 16812
rect 13292 16404 13326 16420
rect 13410 16796 13444 16812
rect 14442 16771 14458 16841
rect 14594 16771 14610 16841
rect 14442 16755 14610 16771
rect 15890 16841 16058 16857
rect 15890 16771 15906 16841
rect 16042 16771 16058 16841
rect 15890 16755 16058 16771
rect 17388 16839 17556 16855
rect 17388 16769 17404 16839
rect 17540 16769 17556 16839
rect 17388 16753 17556 16769
rect 18836 16839 19004 16855
rect 18836 16769 18852 16839
rect 18988 16769 19004 16839
rect 18836 16753 19004 16769
rect 20356 16841 20524 16857
rect 20356 16771 20372 16841
rect 20508 16771 20524 16841
rect 20356 16755 20524 16771
rect 21804 16841 21972 16857
rect 21804 16771 21820 16841
rect 21956 16771 21972 16841
rect 21804 16755 21972 16771
rect 23302 16839 23470 16855
rect 23302 16769 23318 16839
rect 23454 16769 23470 16839
rect 23302 16753 23470 16769
rect 24750 16839 24918 16855
rect 24750 16769 24766 16839
rect 24902 16769 24918 16839
rect 24750 16753 24918 16769
rect 13410 16404 13444 16420
rect 13803 16651 14073 16685
rect 13803 16601 13837 16651
rect 13803 16409 13837 16425
rect 13921 16601 13955 16617
rect 13921 16409 13955 16425
rect 14039 16601 14073 16651
rect 15251 16651 15521 16685
rect 14039 16409 14073 16425
rect 14157 16601 14191 16617
rect 14157 16409 14191 16425
rect 14275 16601 14309 16617
rect 14275 16409 14309 16425
rect 14393 16601 14427 16617
rect 14393 16409 14427 16425
rect 14511 16601 14545 16617
rect 14511 16409 14545 16425
rect 14629 16601 14663 16617
rect 14629 16409 14663 16425
rect 14747 16601 14781 16617
rect 14747 16409 14781 16425
rect 14865 16601 14899 16617
rect 14865 16409 14899 16425
rect 15251 16601 15285 16651
rect 15251 16409 15285 16425
rect 15369 16601 15403 16617
rect 15369 16409 15403 16425
rect 15487 16601 15521 16651
rect 16749 16649 17019 16683
rect 15487 16409 15521 16425
rect 15605 16601 15639 16617
rect 15605 16409 15639 16425
rect 15723 16601 15757 16617
rect 15723 16409 15757 16425
rect 15841 16601 15875 16617
rect 15841 16409 15875 16425
rect 15959 16601 15993 16617
rect 15959 16409 15993 16425
rect 16077 16601 16111 16617
rect 16077 16409 16111 16425
rect 16195 16601 16229 16617
rect 16195 16409 16229 16425
rect 16313 16601 16347 16617
rect 16313 16409 16347 16425
rect 16749 16599 16783 16649
rect 16749 16407 16783 16423
rect 16867 16599 16901 16615
rect 16867 16407 16901 16423
rect 16985 16599 17019 16649
rect 18197 16649 18467 16683
rect 16985 16407 17019 16423
rect 17103 16599 17137 16615
rect 17103 16407 17137 16423
rect 17221 16599 17255 16615
rect 17221 16407 17255 16423
rect 17339 16599 17373 16615
rect 17339 16407 17373 16423
rect 17457 16599 17491 16615
rect 17457 16407 17491 16423
rect 17575 16599 17609 16615
rect 17575 16407 17609 16423
rect 17693 16599 17727 16615
rect 17693 16407 17727 16423
rect 17811 16599 17845 16615
rect 17811 16407 17845 16423
rect 18197 16599 18231 16649
rect 18197 16407 18231 16423
rect 18315 16599 18349 16615
rect 18315 16407 18349 16423
rect 18433 16599 18467 16649
rect 19717 16651 19987 16685
rect 18433 16407 18467 16423
rect 18551 16599 18585 16615
rect 18551 16407 18585 16423
rect 18669 16599 18703 16615
rect 18669 16407 18703 16423
rect 18787 16599 18821 16615
rect 18787 16407 18821 16423
rect 18905 16599 18939 16615
rect 18905 16407 18939 16423
rect 19023 16599 19057 16615
rect 19023 16407 19057 16423
rect 19141 16599 19175 16615
rect 19141 16407 19175 16423
rect 19259 16599 19293 16615
rect 19259 16407 19293 16423
rect 19717 16601 19751 16651
rect 19717 16409 19751 16425
rect 19835 16601 19869 16617
rect 19835 16409 19869 16425
rect 19953 16601 19987 16651
rect 21165 16651 21435 16685
rect 19953 16409 19987 16425
rect 20071 16601 20105 16617
rect 20071 16409 20105 16425
rect 20189 16601 20223 16617
rect 20189 16409 20223 16425
rect 20307 16601 20341 16617
rect 20307 16409 20341 16425
rect 20425 16601 20459 16617
rect 20425 16409 20459 16425
rect 20543 16601 20577 16617
rect 20543 16409 20577 16425
rect 20661 16601 20695 16617
rect 20661 16409 20695 16425
rect 20779 16601 20813 16617
rect 20779 16409 20813 16425
rect 21165 16601 21199 16651
rect 21165 16409 21199 16425
rect 21283 16601 21317 16617
rect 21283 16409 21317 16425
rect 21401 16601 21435 16651
rect 22663 16649 22933 16683
rect 21401 16409 21435 16425
rect 21519 16601 21553 16617
rect 21519 16409 21553 16425
rect 21637 16601 21671 16617
rect 21637 16409 21671 16425
rect 21755 16601 21789 16617
rect 21755 16409 21789 16425
rect 21873 16601 21907 16617
rect 21873 16409 21907 16425
rect 21991 16601 22025 16617
rect 21991 16409 22025 16425
rect 22109 16601 22143 16617
rect 22109 16409 22143 16425
rect 22227 16601 22261 16617
rect 22227 16409 22261 16425
rect 22663 16599 22697 16649
rect 22663 16407 22697 16423
rect 22781 16599 22815 16615
rect 22781 16407 22815 16423
rect 22899 16599 22933 16649
rect 24111 16649 24381 16683
rect 22899 16407 22933 16423
rect 23017 16599 23051 16615
rect 23017 16407 23051 16423
rect 23135 16599 23169 16615
rect 23135 16407 23169 16423
rect 23253 16599 23287 16615
rect 23253 16407 23287 16423
rect 23371 16599 23405 16615
rect 23371 16407 23405 16423
rect 23489 16599 23523 16615
rect 23489 16407 23523 16423
rect 23607 16599 23641 16615
rect 23607 16407 23641 16423
rect 23725 16599 23759 16615
rect 23725 16407 23759 16423
rect 24111 16599 24145 16649
rect 24111 16407 24145 16423
rect 24229 16599 24263 16615
rect 24229 16407 24263 16423
rect 24347 16599 24381 16649
rect 24347 16407 24381 16423
rect 24465 16599 24499 16615
rect 24465 16407 24499 16423
rect 24583 16599 24617 16615
rect 24583 16407 24617 16423
rect 24701 16599 24735 16615
rect 24701 16407 24735 16423
rect 24819 16599 24853 16615
rect 24819 16407 24853 16423
rect 24937 16599 24971 16615
rect 24937 16407 24971 16423
rect 25055 16599 25089 16615
rect 25055 16407 25089 16423
rect 25173 16599 25207 16615
rect 25173 16407 25207 16423
rect 14082 16331 14098 16365
rect 14132 16331 14148 16365
rect 15530 16331 15546 16365
rect 15580 16331 15596 16365
rect 17028 16329 17044 16363
rect 17078 16329 17094 16363
rect 18476 16329 18492 16363
rect 18526 16329 18542 16363
rect 19996 16331 20012 16365
rect 20046 16331 20062 16365
rect 21444 16331 21460 16365
rect 21494 16331 21510 16365
rect 22942 16329 22958 16363
rect 22992 16329 23008 16363
rect 24390 16329 24406 16363
rect 24440 16329 24456 16363
rect 14200 16214 14216 16248
rect 14250 16214 14266 16248
rect 15648 16214 15664 16248
rect 15698 16214 15714 16248
rect 17146 16212 17162 16246
rect 17196 16212 17212 16246
rect 18594 16212 18610 16246
rect 18644 16212 18660 16246
rect 20114 16214 20130 16248
rect 20164 16214 20180 16248
rect 21562 16214 21578 16248
rect 21612 16214 21628 16248
rect 23060 16212 23076 16246
rect 23110 16212 23126 16246
rect 24508 16212 24524 16246
rect 24558 16212 24574 16246
rect 9360 16134 10160 16168
rect 5007 16065 5023 16099
rect 5057 16065 5073 16099
rect 6175 16065 6191 16099
rect 6225 16065 6241 16099
rect 7343 16065 7359 16099
rect 7393 16065 7409 16099
rect 8511 16065 8527 16099
rect 8561 16065 8577 16099
rect 9360 16096 9394 16134
rect 9240 16062 9510 16096
rect 9685 16063 9701 16097
rect 9735 16063 9751 16097
rect 4445 16008 4479 16024
rect 4445 15816 4479 15832
rect 4563 16008 4597 16024
rect 4563 15741 4597 15832
rect 4681 16008 4715 16024
rect 4681 15816 4715 15832
rect 4799 16008 4833 16024
rect 4799 15741 4833 15832
rect 4964 16014 4998 16030
rect 4964 15822 4998 15838
rect 5082 16014 5116 16030
rect 5082 15822 5116 15838
rect 5200 16014 5234 16030
rect 5200 15822 5234 15838
rect 5318 16014 5352 16030
rect 5318 15822 5352 15838
rect 5613 16007 5647 16023
rect 5613 15815 5647 15831
rect 5731 16007 5765 16023
rect 3399 15704 4833 15741
rect 5731 15746 5765 15831
rect 5849 16007 5883 16023
rect 5849 15815 5883 15831
rect 5967 16007 6001 16023
rect 5967 15746 6001 15831
rect 6132 16014 6166 16030
rect 6132 15822 6166 15838
rect 6250 16014 6284 16030
rect 6250 15822 6284 15838
rect 6368 16014 6402 16030
rect 6368 15822 6402 15838
rect 6486 16014 6520 16030
rect 6486 15822 6520 15838
rect 6781 16007 6815 16023
rect 6781 15815 6815 15831
rect 6899 16007 6933 16023
rect 5066 15708 5208 15720
rect 5731 15711 6001 15746
rect 6899 15746 6933 15831
rect 7017 16007 7051 16023
rect 7017 15815 7051 15831
rect 7135 16007 7169 16023
rect 7135 15746 7169 15831
rect 7300 16012 7334 16028
rect 7300 15820 7334 15836
rect 7418 16012 7452 16028
rect 7418 15820 7452 15836
rect 7536 16012 7570 16028
rect 7536 15820 7570 15836
rect 7654 16012 7688 16028
rect 7654 15820 7688 15836
rect 7950 16008 7984 16024
rect 7950 15816 7984 15832
rect 8068 16008 8102 16024
rect 5066 15704 5102 15708
rect 5168 15704 5208 15708
rect 1708 15116 1936 15134
rect 1708 15040 1724 15116
rect 1920 15040 1936 15116
rect 1708 15024 1936 15040
rect 983 14898 1253 14937
rect 983 14846 1017 14898
rect 510 14696 780 14733
rect 510 14646 544 14696
rect 510 14454 544 14470
rect 628 14646 662 14662
rect 628 14416 662 14470
rect 746 14646 780 14696
rect 746 14454 780 14470
rect 864 14646 898 14662
rect 864 14416 898 14470
rect 983 14454 1017 14470
rect 1101 14846 1135 14862
rect 628 14377 898 14416
rect 1101 14419 1135 14470
rect 1219 14846 1253 14898
rect 1456 14898 1726 14937
rect 1219 14454 1253 14470
rect 1337 14846 1371 14862
rect 1337 14419 1371 14470
rect 1456 14846 1490 14898
rect 1456 14454 1490 14470
rect 1574 14846 1608 14862
rect 1574 14419 1608 14470
rect 1692 14846 1726 14898
rect 1928 14898 2198 14937
rect 1692 14454 1726 14470
rect 1810 14846 1844 14862
rect 1810 14419 1844 14470
rect 1928 14846 1962 14898
rect 1928 14454 1962 14470
rect 2046 14846 2080 14862
rect 2046 14419 2080 14470
rect 2164 14846 2198 14898
rect 2395 14899 2665 14938
rect 2164 14454 2198 14470
rect 2277 14846 2311 14862
rect 2277 14419 2311 14470
rect 2395 14846 2429 14899
rect 2395 14454 2429 14470
rect 2513 14846 2547 14862
rect 2513 14419 2547 14470
rect 2631 14846 2665 14899
rect 2836 14697 3106 14736
rect 2631 14454 2665 14470
rect 2718 14646 2752 14662
rect 1101 14380 2547 14419
rect 2718 14419 2752 14470
rect 2836 14646 2870 14697
rect 2836 14454 2870 14470
rect 2954 14646 2988 14662
rect 2954 14419 2988 14470
rect 3072 14646 3106 14697
rect 3072 14454 3106 14470
rect 2718 14380 2988 14419
rect 660 14262 676 14296
rect 710 14262 726 14296
rect 1986 14255 2020 14271
rect 1986 14205 2020 14221
rect 1840 14156 1932 14169
rect 1840 14101 1856 14156
rect 1916 14101 1932 14156
rect 1840 14084 1932 14101
rect 2925 14155 3017 14172
rect 2925 14100 2941 14155
rect 3001 14100 3017 14155
rect 2925 14087 3017 14100
rect 1632 14025 1666 14041
rect 1632 13975 1666 13991
rect 3192 14040 3249 14044
rect 3192 13980 3196 14040
rect 3245 13980 3249 14040
rect 3192 13976 3249 13980
rect 1958 13871 2050 13884
rect 3399 13876 3437 15704
rect 5066 15638 5072 15704
rect 5190 15638 5208 15704
rect 5066 15612 5208 15638
rect 5844 15346 5887 15711
rect 6234 15708 6376 15720
rect 6899 15711 7169 15746
rect 8068 15732 8102 15832
rect 8186 16008 8220 16024
rect 8186 15816 8220 15832
rect 8304 16008 8338 16024
rect 8304 15732 8338 15832
rect 8468 16012 8502 16028
rect 8468 15820 8502 15836
rect 8586 16012 8620 16028
rect 8586 15820 8620 15836
rect 8704 16012 8738 16028
rect 8704 15820 8738 15836
rect 8822 16012 8856 16028
rect 8822 15820 8856 15836
rect 9122 16012 9156 16028
rect 9122 15820 9156 15836
rect 9240 16012 9274 16062
rect 9240 15820 9274 15836
rect 9358 16012 9392 16028
rect 9358 15820 9392 15836
rect 9476 16012 9510 16062
rect 9476 15820 9510 15836
rect 9642 16012 9676 16028
rect 9642 15820 9676 15836
rect 9760 16012 9794 16028
rect 9760 15820 9794 15836
rect 9878 16012 9912 16028
rect 9878 15820 9912 15836
rect 9996 16012 10030 16028
rect 9996 15820 10030 15836
rect 6234 15704 6270 15708
rect 6336 15704 6376 15708
rect 6234 15638 6240 15704
rect 6358 15638 6376 15704
rect 6234 15612 6376 15638
rect 6997 15369 7064 15711
rect 7402 15708 7544 15720
rect 7402 15704 7438 15708
rect 7504 15704 7544 15708
rect 7402 15638 7408 15704
rect 7526 15638 7544 15704
rect 8068 15697 8338 15732
rect 8570 15708 8712 15720
rect 8570 15704 8606 15708
rect 8672 15704 8712 15708
rect 7402 15612 7544 15638
rect 8158 15464 8216 15697
rect 8570 15638 8576 15704
rect 8694 15638 8712 15704
rect 8570 15612 8712 15638
rect 9744 15706 9886 15718
rect 9744 15702 9780 15706
rect 9846 15702 9886 15706
rect 9744 15636 9750 15702
rect 9868 15636 9886 15702
rect 9744 15610 9886 15636
rect 8158 15405 9867 15464
rect 5844 15287 6585 15346
rect 6997 15305 9714 15369
rect 4852 15116 5080 15134
rect 4852 15040 4868 15116
rect 5064 15040 5080 15116
rect 4852 15024 5080 15040
rect 4127 14898 4397 14937
rect 4127 14846 4161 14898
rect 3654 14696 3924 14733
rect 3654 14646 3688 14696
rect 3654 14454 3688 14470
rect 3772 14646 3806 14662
rect 3772 14416 3806 14470
rect 3890 14646 3924 14696
rect 3890 14454 3924 14470
rect 4008 14646 4042 14662
rect 4008 14416 4042 14470
rect 4127 14454 4161 14470
rect 4245 14846 4279 14862
rect 3772 14377 4042 14416
rect 4245 14419 4279 14470
rect 4363 14846 4397 14898
rect 4600 14898 4870 14937
rect 4363 14454 4397 14470
rect 4481 14846 4515 14862
rect 4481 14419 4515 14470
rect 4600 14846 4634 14898
rect 4600 14454 4634 14470
rect 4718 14846 4752 14862
rect 4718 14419 4752 14470
rect 4836 14846 4870 14898
rect 5072 14898 5342 14937
rect 4836 14454 4870 14470
rect 4954 14846 4988 14862
rect 4954 14419 4988 14470
rect 5072 14846 5106 14898
rect 5072 14454 5106 14470
rect 5190 14846 5224 14862
rect 5190 14419 5224 14470
rect 5308 14846 5342 14898
rect 5539 14899 5809 14938
rect 5308 14454 5342 14470
rect 5421 14846 5455 14862
rect 5421 14419 5455 14470
rect 5539 14846 5573 14899
rect 5539 14454 5573 14470
rect 5657 14846 5691 14862
rect 5657 14419 5691 14470
rect 5775 14846 5809 14899
rect 5980 14697 6250 14736
rect 5775 14454 5809 14470
rect 5862 14646 5896 14662
rect 4245 14380 5691 14419
rect 5862 14419 5896 14470
rect 5980 14646 6014 14697
rect 5980 14454 6014 14470
rect 6098 14646 6132 14662
rect 6098 14419 6132 14470
rect 6216 14646 6250 14697
rect 6216 14454 6250 14470
rect 5862 14380 6132 14419
rect 3804 14262 3820 14296
rect 3854 14262 3870 14296
rect 5130 14255 5164 14271
rect 6518 14234 6585 15287
rect 7984 15112 8212 15130
rect 7984 15036 8000 15112
rect 8196 15036 8212 15112
rect 7984 15020 8212 15036
rect 7259 14894 7529 14933
rect 7259 14842 7293 14894
rect 6786 14692 7056 14729
rect 6786 14642 6820 14692
rect 6786 14450 6820 14466
rect 6904 14642 6938 14658
rect 6904 14412 6938 14466
rect 7022 14642 7056 14692
rect 7022 14450 7056 14466
rect 7140 14642 7174 14658
rect 7140 14412 7174 14466
rect 7259 14450 7293 14466
rect 7377 14842 7411 14858
rect 6904 14373 7174 14412
rect 7377 14415 7411 14466
rect 7495 14842 7529 14894
rect 7732 14894 8002 14933
rect 7495 14450 7529 14466
rect 7613 14842 7647 14858
rect 7613 14415 7647 14466
rect 7732 14842 7766 14894
rect 7732 14450 7766 14466
rect 7850 14842 7884 14858
rect 7850 14415 7884 14466
rect 7968 14842 8002 14894
rect 8204 14894 8474 14933
rect 7968 14450 8002 14466
rect 8086 14842 8120 14858
rect 8086 14415 8120 14466
rect 8204 14842 8238 14894
rect 8204 14450 8238 14466
rect 8322 14842 8356 14858
rect 8322 14415 8356 14466
rect 8440 14842 8474 14894
rect 8671 14895 8941 14934
rect 8440 14450 8474 14466
rect 8553 14842 8587 14858
rect 8553 14415 8587 14466
rect 8671 14842 8705 14895
rect 8671 14450 8705 14466
rect 8789 14842 8823 14858
rect 8789 14415 8823 14466
rect 8907 14842 8941 14895
rect 9112 14693 9382 14732
rect 8907 14450 8941 14466
rect 8994 14642 9028 14658
rect 7377 14376 8823 14415
rect 8994 14415 9028 14466
rect 9112 14642 9146 14693
rect 9112 14450 9146 14466
rect 9230 14642 9264 14658
rect 9230 14415 9264 14466
rect 9348 14642 9382 14693
rect 9348 14450 9382 14466
rect 8994 14376 9264 14415
rect 6936 14258 6952 14292
rect 6986 14258 7002 14292
rect 5130 14205 5164 14221
rect 4984 14156 5076 14169
rect 4984 14101 5000 14156
rect 5060 14101 5076 14156
rect 4984 14084 5076 14101
rect 6069 14155 6161 14172
rect 6069 14100 6085 14155
rect 6145 14100 6161 14155
rect 6069 14087 6161 14100
rect 4776 14025 4810 14041
rect 4776 13975 4810 13991
rect 6336 14040 6393 14044
rect 6336 13980 6340 14040
rect 6389 13980 6393 14040
rect 6336 13976 6393 13980
rect 1958 13816 1974 13871
rect 2034 13816 2050 13871
rect 1958 13799 2050 13816
rect 3183 13872 3437 13876
rect 3183 13812 3196 13872
rect 3245 13812 3437 13872
rect 3183 13808 3437 13812
rect 5102 13871 5194 13884
rect 5102 13816 5118 13871
rect 5178 13816 5194 13871
rect 5102 13799 5194 13816
rect 6336 13875 6393 13876
rect 6517 13875 6585 14234
rect 8262 14251 8296 14267
rect 8262 14201 8296 14217
rect 8116 14152 8208 14165
rect 8116 14097 8132 14152
rect 8192 14097 8208 14152
rect 8116 14080 8208 14097
rect 9201 14151 9293 14168
rect 9201 14096 9217 14151
rect 9277 14096 9293 14151
rect 9201 14083 9293 14096
rect 7908 14021 7942 14037
rect 7908 13971 7942 13987
rect 9468 14036 9525 14040
rect 9468 13976 9472 14036
rect 9521 13976 9525 14036
rect 9468 13972 9525 13976
rect 6336 13872 6585 13875
rect 6336 13812 6340 13872
rect 6389 13812 6585 13872
rect 6336 13808 6585 13812
rect 6339 13807 6585 13808
rect 8234 13867 8326 13880
rect 9646 13872 9714 15305
rect 8234 13812 8250 13867
rect 8310 13812 8326 13867
rect 8234 13795 8326 13812
rect 9468 13868 9714 13872
rect 9468 13808 9472 13868
rect 9521 13808 9714 13868
rect 9468 13804 9714 13808
rect 9788 13872 9867 15405
rect 10087 15265 10160 16134
rect 14157 16164 14191 16180
rect 10853 16063 10869 16097
rect 10903 16063 10919 16097
rect 12021 16063 12037 16097
rect 12071 16063 12087 16097
rect 13189 16063 13205 16097
rect 13239 16063 13255 16097
rect 10291 16012 10325 16028
rect 10291 15820 10325 15836
rect 10409 16012 10443 16028
rect 10409 15725 10443 15836
rect 10527 16012 10561 16028
rect 10527 15820 10561 15836
rect 10645 16012 10679 16028
rect 10645 15725 10679 15836
rect 10810 16012 10844 16028
rect 10810 15820 10844 15836
rect 10928 16012 10962 16028
rect 10928 15820 10962 15836
rect 11046 16012 11080 16028
rect 11046 15820 11080 15836
rect 11164 16012 11198 16028
rect 11164 15820 11198 15836
rect 11459 16012 11493 16028
rect 11459 15820 11493 15836
rect 11577 16012 11611 16028
rect 10409 15689 10679 15725
rect 11577 15742 11611 15836
rect 11695 16012 11729 16028
rect 11695 15820 11729 15836
rect 11813 16012 11847 16028
rect 11813 15742 11847 15836
rect 11978 16012 12012 16028
rect 11978 15820 12012 15836
rect 12096 16012 12130 16028
rect 12096 15820 12130 15836
rect 12214 16012 12248 16028
rect 12214 15820 12248 15836
rect 12332 16012 12366 16028
rect 12332 15820 12366 15836
rect 12626 16006 12660 16022
rect 12626 15814 12660 15830
rect 12744 16006 12778 16022
rect 10912 15706 11054 15718
rect 11577 15708 11847 15742
rect 12744 15730 12778 15830
rect 12862 16006 12896 16022
rect 12862 15814 12896 15830
rect 12980 16006 13014 16022
rect 12980 15730 13014 15830
rect 13146 16010 13180 16026
rect 13146 15818 13180 15834
rect 13264 16010 13298 16026
rect 13264 15818 13298 15834
rect 13382 16010 13416 16026
rect 13382 15818 13416 15834
rect 13500 16010 13534 16026
rect 14157 15972 14191 15988
rect 14275 16164 14309 16180
rect 14275 15972 14309 15988
rect 14392 16164 14426 16180
rect 13500 15818 13534 15834
rect 14392 15772 14426 15788
rect 14510 16164 14544 16180
rect 14510 15772 14544 15788
rect 14628 16164 14662 16180
rect 15605 16164 15639 16180
rect 15605 15972 15639 15988
rect 15723 16164 15757 16180
rect 15723 15972 15757 15988
rect 15840 16164 15874 16180
rect 14628 15772 14662 15788
rect 15840 15772 15874 15788
rect 15958 16164 15992 16180
rect 15958 15772 15992 15788
rect 16076 16164 16110 16180
rect 17103 16162 17137 16178
rect 17103 15970 17137 15986
rect 17221 16162 17255 16178
rect 17221 15970 17255 15986
rect 17338 16162 17372 16178
rect 16076 15772 16110 15788
rect 17338 15770 17372 15786
rect 17456 16162 17490 16178
rect 17456 15770 17490 15786
rect 17574 16162 17608 16178
rect 18551 16162 18585 16178
rect 18551 15970 18585 15986
rect 18669 16162 18703 16178
rect 18669 15970 18703 15986
rect 18786 16162 18820 16178
rect 17574 15770 17608 15786
rect 18786 15770 18820 15786
rect 18904 16162 18938 16178
rect 18904 15770 18938 15786
rect 19022 16162 19056 16178
rect 20071 16164 20105 16180
rect 20071 15972 20105 15988
rect 20189 16164 20223 16180
rect 20189 15972 20223 15988
rect 20306 16164 20340 16180
rect 19022 15770 19056 15786
rect 20306 15772 20340 15788
rect 20424 16164 20458 16180
rect 20424 15772 20458 15788
rect 20542 16164 20576 16180
rect 21519 16164 21553 16180
rect 21519 15972 21553 15988
rect 21637 16164 21671 16180
rect 21637 15972 21671 15988
rect 21754 16164 21788 16180
rect 20542 15772 20576 15788
rect 21754 15772 21788 15788
rect 21872 16164 21906 16180
rect 21872 15772 21906 15788
rect 21990 16164 22024 16180
rect 23017 16162 23051 16178
rect 23017 15970 23051 15986
rect 23135 16162 23169 16178
rect 23135 15970 23169 15986
rect 23252 16162 23286 16178
rect 21990 15772 22024 15788
rect 23252 15770 23286 15786
rect 23370 16162 23404 16178
rect 23370 15770 23404 15786
rect 23488 16162 23522 16178
rect 24465 16162 24499 16178
rect 24465 15970 24499 15986
rect 24583 16162 24617 16178
rect 24583 15970 24617 15986
rect 24700 16162 24734 16178
rect 23488 15770 23522 15786
rect 24700 15770 24734 15786
rect 24818 16162 24852 16178
rect 24818 15770 24852 15786
rect 24936 16162 24970 16178
rect 24936 15770 24970 15786
rect 10912 15702 10948 15706
rect 11014 15702 11054 15706
rect 10544 15347 10593 15689
rect 10912 15636 10918 15702
rect 11036 15636 11054 15702
rect 10912 15610 11054 15636
rect 11695 15435 11729 15708
rect 12080 15706 12222 15718
rect 12080 15702 12116 15706
rect 12182 15702 12222 15706
rect 12080 15636 12086 15702
rect 12204 15636 12222 15702
rect 12744 15696 13014 15730
rect 13248 15706 13390 15718
rect 13248 15702 13284 15706
rect 13350 15702 13390 15706
rect 14435 15704 14451 15738
rect 14485 15704 14501 15738
rect 14553 15704 14569 15738
rect 14603 15704 14619 15738
rect 15883 15704 15899 15738
rect 15933 15704 15949 15738
rect 16001 15704 16017 15738
rect 16051 15704 16067 15738
rect 17381 15702 17397 15736
rect 17431 15702 17447 15736
rect 17499 15702 17515 15736
rect 17549 15702 17565 15736
rect 18829 15702 18845 15736
rect 18879 15702 18895 15736
rect 18947 15702 18963 15736
rect 18997 15702 19013 15736
rect 20349 15704 20365 15738
rect 20399 15704 20415 15738
rect 20467 15704 20483 15738
rect 20517 15704 20533 15738
rect 21797 15704 21813 15738
rect 21847 15704 21863 15738
rect 21915 15704 21931 15738
rect 21965 15704 21981 15738
rect 23295 15702 23311 15736
rect 23345 15702 23361 15736
rect 23413 15702 23429 15736
rect 23463 15702 23479 15736
rect 24743 15702 24759 15736
rect 24793 15702 24809 15736
rect 24861 15702 24877 15736
rect 24911 15702 24927 15736
rect 12080 15610 12222 15636
rect 12877 15523 12922 15696
rect 13248 15636 13254 15702
rect 13372 15636 13390 15702
rect 13248 15610 13390 15636
rect 14218 15633 14386 15651
rect 14218 15577 14236 15633
rect 14370 15577 14386 15633
rect 14218 15561 14386 15577
rect 15666 15633 15834 15651
rect 15666 15577 15684 15633
rect 15818 15577 15834 15633
rect 15666 15561 15834 15577
rect 17164 15631 17332 15649
rect 17164 15575 17182 15631
rect 17316 15575 17332 15631
rect 17164 15559 17332 15575
rect 18612 15631 18780 15649
rect 18612 15575 18630 15631
rect 18764 15575 18780 15631
rect 18612 15559 18780 15575
rect 20132 15633 20300 15651
rect 20132 15577 20150 15633
rect 20284 15577 20300 15633
rect 20132 15561 20300 15577
rect 21580 15633 21748 15651
rect 21580 15577 21598 15633
rect 21732 15577 21748 15633
rect 21580 15561 21748 15577
rect 23078 15631 23246 15649
rect 23078 15575 23096 15631
rect 23230 15575 23246 15631
rect 23078 15559 23246 15575
rect 24526 15631 24694 15649
rect 24526 15575 24544 15631
rect 24678 15575 24694 15631
rect 24526 15559 24694 15575
rect 12877 15469 25542 15523
rect 11695 15381 22319 15435
rect 10544 15299 19195 15347
rect 10087 15211 13079 15265
rect 11128 15112 11356 15130
rect 11128 15036 11144 15112
rect 11340 15036 11356 15112
rect 11128 15020 11356 15036
rect 10403 14894 10673 14933
rect 10403 14842 10437 14894
rect 9930 14692 10200 14729
rect 9930 14642 9964 14692
rect 9930 14450 9964 14466
rect 10048 14642 10082 14658
rect 10048 14412 10082 14466
rect 10166 14642 10200 14692
rect 10166 14450 10200 14466
rect 10284 14642 10318 14658
rect 10284 14412 10318 14466
rect 10403 14450 10437 14466
rect 10521 14842 10555 14858
rect 10048 14373 10318 14412
rect 10521 14415 10555 14466
rect 10639 14842 10673 14894
rect 10876 14894 11146 14933
rect 10639 14450 10673 14466
rect 10757 14842 10791 14858
rect 10757 14415 10791 14466
rect 10876 14842 10910 14894
rect 10876 14450 10910 14466
rect 10994 14842 11028 14858
rect 10994 14415 11028 14466
rect 11112 14842 11146 14894
rect 11348 14894 11618 14933
rect 11112 14450 11146 14466
rect 11230 14842 11264 14858
rect 11230 14415 11264 14466
rect 11348 14842 11382 14894
rect 11348 14450 11382 14466
rect 11466 14842 11500 14858
rect 11466 14415 11500 14466
rect 11584 14842 11618 14894
rect 11815 14895 12085 14934
rect 11584 14450 11618 14466
rect 11697 14842 11731 14858
rect 11697 14415 11731 14466
rect 11815 14842 11849 14895
rect 11815 14450 11849 14466
rect 11933 14842 11967 14858
rect 11933 14415 11967 14466
rect 12051 14842 12085 14895
rect 12256 14693 12526 14732
rect 12051 14450 12085 14466
rect 12138 14642 12172 14658
rect 10521 14376 11967 14415
rect 12138 14415 12172 14466
rect 12256 14642 12290 14693
rect 12256 14450 12290 14466
rect 12374 14642 12408 14658
rect 12374 14415 12408 14466
rect 12492 14642 12526 14693
rect 12492 14450 12526 14466
rect 12138 14376 12408 14415
rect 10080 14258 10096 14292
rect 10130 14258 10146 14292
rect 11406 14251 11440 14267
rect 11406 14201 11440 14217
rect 11260 14152 11352 14165
rect 11260 14097 11276 14152
rect 11336 14097 11352 14152
rect 11260 14080 11352 14097
rect 12345 14151 12437 14168
rect 12345 14096 12361 14151
rect 12421 14096 12437 14151
rect 12345 14083 12437 14096
rect 11052 14021 11086 14037
rect 11052 13971 11086 13987
rect 12612 14036 12669 14040
rect 12612 13976 12616 14036
rect 12665 13976 12669 14036
rect 12612 13972 12669 13976
rect 11378 13872 11470 13880
rect 9788 13867 11470 13872
rect 9788 13812 11394 13867
rect 11452 13812 11470 13867
rect 9788 13801 11470 13812
rect 13007 13877 13079 15211
rect 14330 15116 14558 15134
rect 14330 15040 14346 15116
rect 14542 15040 14558 15116
rect 14330 15024 14558 15040
rect 17474 15116 17702 15134
rect 17474 15040 17490 15116
rect 17686 15040 17702 15116
rect 17474 15024 17702 15040
rect 13605 14898 13875 14937
rect 13605 14846 13639 14898
rect 13132 14696 13402 14733
rect 13132 14646 13166 14696
rect 13132 14454 13166 14470
rect 13250 14646 13284 14662
rect 13250 14416 13284 14470
rect 13368 14646 13402 14696
rect 13368 14454 13402 14470
rect 13486 14646 13520 14662
rect 13486 14416 13520 14470
rect 13605 14454 13639 14470
rect 13723 14846 13757 14862
rect 13250 14377 13520 14416
rect 13723 14419 13757 14470
rect 13841 14846 13875 14898
rect 14078 14898 14348 14937
rect 13841 14454 13875 14470
rect 13959 14846 13993 14862
rect 13959 14419 13993 14470
rect 14078 14846 14112 14898
rect 14078 14454 14112 14470
rect 14196 14846 14230 14862
rect 14196 14419 14230 14470
rect 14314 14846 14348 14898
rect 14550 14898 14820 14937
rect 14314 14454 14348 14470
rect 14432 14846 14466 14862
rect 14432 14419 14466 14470
rect 14550 14846 14584 14898
rect 14550 14454 14584 14470
rect 14668 14846 14702 14862
rect 14668 14419 14702 14470
rect 14786 14846 14820 14898
rect 15017 14899 15287 14938
rect 14786 14454 14820 14470
rect 14899 14846 14933 14862
rect 14899 14419 14933 14470
rect 15017 14846 15051 14899
rect 15017 14454 15051 14470
rect 15135 14846 15169 14862
rect 15135 14419 15169 14470
rect 15253 14846 15287 14899
rect 16749 14898 17019 14937
rect 16749 14846 16783 14898
rect 15458 14697 15728 14736
rect 15253 14454 15287 14470
rect 15340 14646 15374 14662
rect 13723 14380 15169 14419
rect 15340 14419 15374 14470
rect 15458 14646 15492 14697
rect 15458 14454 15492 14470
rect 15576 14646 15610 14662
rect 15576 14419 15610 14470
rect 15694 14646 15728 14697
rect 15694 14454 15728 14470
rect 16276 14696 16546 14733
rect 16276 14646 16310 14696
rect 16276 14454 16310 14470
rect 16394 14646 16428 14662
rect 15340 14380 15610 14419
rect 16394 14416 16428 14470
rect 16512 14646 16546 14696
rect 16512 14454 16546 14470
rect 16630 14646 16664 14662
rect 16630 14416 16664 14470
rect 16749 14454 16783 14470
rect 16867 14846 16901 14862
rect 16394 14377 16664 14416
rect 16867 14419 16901 14470
rect 16985 14846 17019 14898
rect 17222 14898 17492 14937
rect 16985 14454 17019 14470
rect 17103 14846 17137 14862
rect 17103 14419 17137 14470
rect 17222 14846 17256 14898
rect 17222 14454 17256 14470
rect 17340 14846 17374 14862
rect 17340 14419 17374 14470
rect 17458 14846 17492 14898
rect 17694 14898 17964 14937
rect 17458 14454 17492 14470
rect 17576 14846 17610 14862
rect 17576 14419 17610 14470
rect 17694 14846 17728 14898
rect 17694 14454 17728 14470
rect 17812 14846 17846 14862
rect 17812 14419 17846 14470
rect 17930 14846 17964 14898
rect 18161 14899 18431 14938
rect 17930 14454 17964 14470
rect 18043 14846 18077 14862
rect 18043 14419 18077 14470
rect 18161 14846 18195 14899
rect 18161 14454 18195 14470
rect 18279 14846 18313 14862
rect 18279 14419 18313 14470
rect 18397 14846 18431 14899
rect 18602 14697 18872 14736
rect 18397 14454 18431 14470
rect 18484 14646 18518 14662
rect 16867 14380 18313 14419
rect 18484 14419 18518 14470
rect 18602 14646 18636 14697
rect 18602 14454 18636 14470
rect 18720 14646 18754 14662
rect 18720 14419 18754 14470
rect 18838 14646 18872 14697
rect 18838 14454 18872 14470
rect 18484 14380 18754 14419
rect 13282 14262 13298 14296
rect 13332 14262 13348 14296
rect 14608 14255 14642 14271
rect 16426 14262 16442 14296
rect 16476 14262 16492 14296
rect 14608 14205 14642 14221
rect 17752 14255 17786 14271
rect 17752 14205 17786 14221
rect 14462 14156 14554 14169
rect 14462 14101 14478 14156
rect 14538 14101 14554 14156
rect 14462 14084 14554 14101
rect 15547 14155 15639 14172
rect 15547 14100 15563 14155
rect 15623 14100 15639 14155
rect 15547 14087 15639 14100
rect 17606 14156 17698 14169
rect 17606 14101 17622 14156
rect 17682 14101 17698 14156
rect 17606 14084 17698 14101
rect 18691 14155 18783 14172
rect 18691 14100 18707 14155
rect 18767 14100 18783 14155
rect 18691 14087 18783 14100
rect 14254 14025 14288 14041
rect 14254 13975 14288 13991
rect 15814 14040 15871 14044
rect 15814 13980 15818 14040
rect 15867 13980 15871 14040
rect 15814 13976 15871 13980
rect 17398 14025 17432 14041
rect 17398 13975 17432 13991
rect 18958 14040 19015 14044
rect 18958 13980 18962 14040
rect 19011 13980 19015 14040
rect 18958 13976 19015 13980
rect 14580 13877 14672 13884
rect 13007 13871 14672 13877
rect 13007 13816 14596 13871
rect 14654 13816 14672 13871
rect 13007 13806 14672 13816
rect 11378 13795 11470 13801
rect 14580 13799 14672 13806
rect 17724 13871 17816 13884
rect 19127 13876 19195 15299
rect 20606 15112 20834 15130
rect 20606 15036 20622 15112
rect 20818 15036 20834 15112
rect 20606 15020 20834 15036
rect 19881 14894 20151 14933
rect 19881 14842 19915 14894
rect 19408 14692 19678 14729
rect 19408 14642 19442 14692
rect 19408 14450 19442 14466
rect 19526 14642 19560 14658
rect 19526 14412 19560 14466
rect 19644 14642 19678 14692
rect 19644 14450 19678 14466
rect 19762 14642 19796 14658
rect 19762 14412 19796 14466
rect 19881 14450 19915 14466
rect 19999 14842 20033 14858
rect 19526 14373 19796 14412
rect 19999 14415 20033 14466
rect 20117 14842 20151 14894
rect 20354 14894 20624 14933
rect 20117 14450 20151 14466
rect 20235 14842 20269 14858
rect 20235 14415 20269 14466
rect 20354 14842 20388 14894
rect 20354 14450 20388 14466
rect 20472 14842 20506 14858
rect 20472 14415 20506 14466
rect 20590 14842 20624 14894
rect 20826 14894 21096 14933
rect 20590 14450 20624 14466
rect 20708 14842 20742 14858
rect 20708 14415 20742 14466
rect 20826 14842 20860 14894
rect 20826 14450 20860 14466
rect 20944 14842 20978 14858
rect 20944 14415 20978 14466
rect 21062 14842 21096 14894
rect 21293 14895 21563 14934
rect 21062 14450 21096 14466
rect 21175 14842 21209 14858
rect 21175 14415 21209 14466
rect 21293 14842 21327 14895
rect 21293 14450 21327 14466
rect 21411 14842 21445 14858
rect 21411 14415 21445 14466
rect 21529 14842 21563 14895
rect 21734 14693 22004 14732
rect 21529 14450 21563 14466
rect 21616 14642 21650 14658
rect 19999 14376 21445 14415
rect 21616 14415 21650 14466
rect 21734 14642 21768 14693
rect 21734 14450 21768 14466
rect 21852 14642 21886 14658
rect 21852 14415 21886 14466
rect 21970 14642 22004 14693
rect 21970 14450 22004 14466
rect 21616 14376 21886 14415
rect 19558 14258 19574 14292
rect 19608 14258 19624 14292
rect 20884 14251 20918 14267
rect 20884 14201 20918 14217
rect 20738 14152 20830 14165
rect 20738 14097 20754 14152
rect 20814 14097 20830 14152
rect 20738 14080 20830 14097
rect 21823 14151 21915 14168
rect 21823 14096 21839 14151
rect 21899 14096 21915 14151
rect 21823 14083 21915 14096
rect 20530 14021 20564 14037
rect 20530 13971 20564 13987
rect 22090 14036 22147 14040
rect 22090 13976 22094 14036
rect 22143 13976 22147 14036
rect 22090 13972 22147 13976
rect 17724 13816 17740 13871
rect 17800 13816 17816 13871
rect 17724 13799 17816 13816
rect 18957 13872 19195 13876
rect 18957 13812 18962 13872
rect 19011 13812 19195 13872
rect 18957 13807 19195 13812
rect 20856 13867 20948 13880
rect 22241 13872 22319 15381
rect 23750 15112 23978 15130
rect 23750 15036 23766 15112
rect 23962 15036 23978 15112
rect 23750 15020 23978 15036
rect 23025 14894 23295 14933
rect 23025 14842 23059 14894
rect 22552 14692 22822 14729
rect 22552 14642 22586 14692
rect 22552 14450 22586 14466
rect 22670 14642 22704 14658
rect 22670 14412 22704 14466
rect 22788 14642 22822 14692
rect 22788 14450 22822 14466
rect 22906 14642 22940 14658
rect 22906 14412 22940 14466
rect 23025 14450 23059 14466
rect 23143 14842 23177 14858
rect 22670 14373 22940 14412
rect 23143 14415 23177 14466
rect 23261 14842 23295 14894
rect 23498 14894 23768 14933
rect 23261 14450 23295 14466
rect 23379 14842 23413 14858
rect 23379 14415 23413 14466
rect 23498 14842 23532 14894
rect 23498 14450 23532 14466
rect 23616 14842 23650 14858
rect 23616 14415 23650 14466
rect 23734 14842 23768 14894
rect 23970 14894 24240 14933
rect 23734 14450 23768 14466
rect 23852 14842 23886 14858
rect 23852 14415 23886 14466
rect 23970 14842 24004 14894
rect 23970 14450 24004 14466
rect 24088 14842 24122 14858
rect 24088 14415 24122 14466
rect 24206 14842 24240 14894
rect 24437 14895 24707 14934
rect 24206 14450 24240 14466
rect 24319 14842 24353 14858
rect 24319 14415 24353 14466
rect 24437 14842 24471 14895
rect 24437 14450 24471 14466
rect 24555 14842 24589 14858
rect 24555 14415 24589 14466
rect 24673 14842 24707 14895
rect 24878 14693 25148 14732
rect 24673 14450 24707 14466
rect 24760 14642 24794 14658
rect 23143 14376 24589 14415
rect 24760 14415 24794 14466
rect 24878 14642 24912 14693
rect 24878 14450 24912 14466
rect 24996 14642 25030 14658
rect 24996 14415 25030 14466
rect 25114 14642 25148 14693
rect 25114 14450 25148 14466
rect 24760 14376 25030 14415
rect 25450 14322 25542 15469
rect 22702 14258 22718 14292
rect 22752 14258 22768 14292
rect 24028 14251 24062 14267
rect 24028 14201 24062 14217
rect 23882 14152 23974 14165
rect 23882 14097 23898 14152
rect 23958 14097 23974 14152
rect 23882 14080 23974 14097
rect 24967 14151 25059 14168
rect 24967 14096 24983 14151
rect 25043 14096 25059 14151
rect 24967 14083 25059 14096
rect 23674 14021 23708 14037
rect 23674 13971 23708 13987
rect 25234 14036 25291 14040
rect 25234 13976 25238 14036
rect 25287 13976 25291 14036
rect 25234 13972 25291 13976
rect 25449 13881 25542 14322
rect 20856 13812 20872 13867
rect 20932 13812 20948 13867
rect 20856 13795 20948 13812
rect 22090 13868 22319 13872
rect 22090 13808 22094 13868
rect 22143 13808 22319 13868
rect 22090 13804 22319 13808
rect 24000 13867 24092 13880
rect 24000 13812 24016 13867
rect 24076 13812 24092 13867
rect 24000 13795 24092 13812
rect 25231 13868 25542 13881
rect 25231 13808 25238 13868
rect 25287 13808 25542 13868
rect 25231 13795 25542 13808
rect 1751 13635 1785 13651
rect 1751 13585 1785 13601
rect 4895 13635 4929 13651
rect 4895 13585 4929 13601
rect 8027 13631 8061 13647
rect 8027 13581 8061 13597
rect 11171 13631 11205 13647
rect 11171 13581 11205 13597
rect 14373 13635 14407 13651
rect 14373 13585 14407 13601
rect 17517 13635 17551 13651
rect 17517 13585 17551 13601
rect 20649 13631 20683 13647
rect 20649 13581 20683 13597
rect 23793 13631 23827 13647
rect 23793 13581 23827 13597
rect 1378 13513 1412 13529
rect 1378 13321 1412 13337
rect 1496 13525 1530 13529
rect 1574 13525 1608 13529
rect 1496 13513 1608 13525
rect 1530 13337 1574 13513
rect 1496 13325 1574 13337
rect 1496 13321 1530 13325
rect 1574 13121 1608 13137
rect 1692 13513 1726 13529
rect 1692 13121 1726 13137
rect 1810 13513 1844 13529
rect 1810 13121 1844 13137
rect 1928 13513 1962 13529
rect 1928 13121 1962 13137
rect 2046 13525 2080 13529
rect 2120 13525 2154 13529
rect 2046 13513 2154 13525
rect 2080 13337 2120 13513
rect 2080 13325 2154 13337
rect 2120 13321 2154 13325
rect 2238 13513 2272 13529
rect 2238 13321 2272 13337
rect 4522 13513 4556 13529
rect 4522 13321 4556 13337
rect 4640 13525 4674 13529
rect 4718 13525 4752 13529
rect 4640 13513 4752 13525
rect 4674 13337 4718 13513
rect 4640 13325 4718 13337
rect 4640 13321 4674 13325
rect 2046 13121 2080 13137
rect 4718 13121 4752 13137
rect 4836 13513 4870 13529
rect 4836 13121 4870 13137
rect 4954 13513 4988 13529
rect 4954 13121 4988 13137
rect 5072 13513 5106 13529
rect 5072 13121 5106 13137
rect 5190 13525 5224 13529
rect 5264 13525 5298 13529
rect 5190 13513 5298 13525
rect 5224 13337 5264 13513
rect 5224 13325 5298 13337
rect 5264 13321 5298 13325
rect 5382 13513 5416 13529
rect 5382 13321 5416 13337
rect 7654 13509 7688 13525
rect 7654 13317 7688 13333
rect 7772 13521 7806 13525
rect 7850 13521 7884 13525
rect 7772 13509 7884 13521
rect 7806 13333 7850 13509
rect 7772 13321 7850 13333
rect 7772 13317 7806 13321
rect 5190 13121 5224 13137
rect 7850 13117 7884 13133
rect 7968 13509 8002 13525
rect 7968 13117 8002 13133
rect 8086 13509 8120 13525
rect 8086 13117 8120 13133
rect 8204 13509 8238 13525
rect 8204 13117 8238 13133
rect 8322 13521 8356 13525
rect 8396 13521 8430 13525
rect 8322 13509 8430 13521
rect 8356 13333 8396 13509
rect 8356 13321 8430 13333
rect 8396 13317 8430 13321
rect 8514 13509 8548 13525
rect 8514 13317 8548 13333
rect 10798 13509 10832 13525
rect 10798 13317 10832 13333
rect 10916 13521 10950 13525
rect 10994 13521 11028 13525
rect 10916 13509 11028 13521
rect 10950 13333 10994 13509
rect 10916 13321 10994 13333
rect 10916 13317 10950 13321
rect 8322 13117 8356 13133
rect 10994 13117 11028 13133
rect 11112 13509 11146 13525
rect 11112 13117 11146 13133
rect 11230 13509 11264 13525
rect 11230 13117 11264 13133
rect 11348 13509 11382 13525
rect 11348 13117 11382 13133
rect 11466 13521 11500 13525
rect 11540 13521 11574 13525
rect 11466 13509 11574 13521
rect 11500 13333 11540 13509
rect 11500 13321 11574 13333
rect 11540 13317 11574 13321
rect 11658 13509 11692 13525
rect 11658 13317 11692 13333
rect 14000 13513 14034 13529
rect 14000 13321 14034 13337
rect 14118 13525 14152 13529
rect 14196 13525 14230 13529
rect 14118 13513 14230 13525
rect 14152 13337 14196 13513
rect 14118 13325 14196 13337
rect 14118 13321 14152 13325
rect 11466 13117 11500 13133
rect 14196 13121 14230 13137
rect 14314 13513 14348 13529
rect 14314 13121 14348 13137
rect 14432 13513 14466 13529
rect 14432 13121 14466 13137
rect 14550 13513 14584 13529
rect 14550 13121 14584 13137
rect 14668 13525 14702 13529
rect 14742 13525 14776 13529
rect 14668 13513 14776 13525
rect 14702 13337 14742 13513
rect 14702 13325 14776 13337
rect 14742 13321 14776 13325
rect 14860 13513 14894 13529
rect 14860 13321 14894 13337
rect 17144 13513 17178 13529
rect 17144 13321 17178 13337
rect 17262 13525 17296 13529
rect 17340 13525 17374 13529
rect 17262 13513 17374 13525
rect 17296 13337 17340 13513
rect 17262 13325 17340 13337
rect 17262 13321 17296 13325
rect 14668 13121 14702 13137
rect 17340 13121 17374 13137
rect 17458 13513 17492 13529
rect 17458 13121 17492 13137
rect 17576 13513 17610 13529
rect 17576 13121 17610 13137
rect 17694 13513 17728 13529
rect 17694 13121 17728 13137
rect 17812 13525 17846 13529
rect 17886 13525 17920 13529
rect 17812 13513 17920 13525
rect 17846 13337 17886 13513
rect 17846 13325 17920 13337
rect 17886 13321 17920 13325
rect 18004 13513 18038 13529
rect 18004 13321 18038 13337
rect 20276 13509 20310 13525
rect 20276 13317 20310 13333
rect 20394 13521 20428 13525
rect 20472 13521 20506 13525
rect 20394 13509 20506 13521
rect 20428 13333 20472 13509
rect 20394 13321 20472 13333
rect 20394 13317 20428 13321
rect 17812 13121 17846 13137
rect 20472 13117 20506 13133
rect 20590 13509 20624 13525
rect 20590 13117 20624 13133
rect 20708 13509 20742 13525
rect 20708 13117 20742 13133
rect 20826 13509 20860 13525
rect 20826 13117 20860 13133
rect 20944 13521 20978 13525
rect 21018 13521 21052 13525
rect 20944 13509 21052 13521
rect 20978 13333 21018 13509
rect 20978 13321 21052 13333
rect 21018 13317 21052 13321
rect 21136 13509 21170 13525
rect 21136 13317 21170 13333
rect 23420 13509 23454 13525
rect 23420 13317 23454 13333
rect 23538 13521 23572 13525
rect 23616 13521 23650 13525
rect 23538 13509 23650 13521
rect 23572 13333 23616 13509
rect 23538 13321 23616 13333
rect 23538 13317 23572 13321
rect 20944 13117 20978 13133
rect 23616 13117 23650 13133
rect 23734 13509 23768 13525
rect 23734 13117 23768 13133
rect 23852 13509 23886 13525
rect 23852 13117 23886 13133
rect 23970 13509 24004 13525
rect 23970 13117 24004 13133
rect 24088 13521 24122 13525
rect 24162 13521 24196 13525
rect 24088 13509 24196 13521
rect 24122 13333 24162 13509
rect 24122 13321 24196 13333
rect 24162 13317 24196 13321
rect 24280 13509 24314 13525
rect 24280 13317 24314 13333
rect 24088 13117 24122 13133
rect 30077 13134 30166 13168
rect 30342 13134 30358 13168
rect 1793 13002 1809 13036
rect 1843 13002 1859 13036
rect 4937 13002 4953 13036
rect 4987 13002 5003 13036
rect 8069 12998 8085 13032
rect 8119 12998 8135 13032
rect 11213 12998 11229 13032
rect 11263 12998 11279 13032
rect 14415 13002 14431 13036
rect 14465 13002 14481 13036
rect 17559 13002 17575 13036
rect 17609 13002 17625 13036
rect 20691 12998 20707 13032
rect 20741 12998 20757 13032
rect 23835 12998 23851 13032
rect 23885 12998 23901 13032
rect 30077 12932 30112 13134
rect 30150 13016 30166 13050
rect 30342 13016 30358 13050
rect 31375 13009 31391 13043
rect 31567 13009 31583 13043
rect 30077 12898 30166 12932
rect 30342 12898 30358 12932
rect 1742 12884 1878 12888
rect 1742 12870 1782 12884
rect 1840 12870 1878 12884
rect 1742 12824 1758 12870
rect 1862 12824 1878 12870
rect 1742 12802 1878 12824
rect 4886 12884 5022 12888
rect 14364 12884 14500 12888
rect 4886 12870 4926 12884
rect 4984 12870 5022 12884
rect 4886 12824 4902 12870
rect 5006 12824 5022 12870
rect 4886 12802 5022 12824
rect 8018 12880 8154 12884
rect 8018 12866 8058 12880
rect 8116 12866 8154 12880
rect 8018 12820 8034 12866
rect 8138 12820 8154 12866
rect 8018 12798 8154 12820
rect 11162 12880 11298 12884
rect 11162 12866 11202 12880
rect 11260 12866 11298 12880
rect 11162 12820 11178 12866
rect 11282 12820 11298 12866
rect 11162 12798 11298 12820
rect 14364 12870 14404 12884
rect 14462 12870 14500 12884
rect 14364 12824 14380 12870
rect 14484 12824 14500 12870
rect 14364 12802 14500 12824
rect 17508 12884 17644 12888
rect 17508 12870 17548 12884
rect 17606 12870 17644 12884
rect 17508 12824 17524 12870
rect 17628 12824 17644 12870
rect 17508 12802 17644 12824
rect 20640 12880 20776 12884
rect 20640 12866 20680 12880
rect 20738 12866 20776 12880
rect 20640 12820 20656 12866
rect 20760 12820 20776 12866
rect 20640 12798 20776 12820
rect 23784 12880 23920 12884
rect 23784 12866 23824 12880
rect 23882 12866 23920 12880
rect 23784 12820 23800 12866
rect 23904 12820 23920 12866
rect 31274 12862 31290 12896
rect 31324 12862 31340 12896
rect 31375 12891 31391 12925
rect 31567 12891 31583 12925
rect 23784 12798 23920 12820
rect 30150 12780 30166 12814
rect 30342 12780 30358 12814
rect 30643 12707 30659 12741
rect 31035 12707 31051 12741
rect 31207 12711 31273 12727
rect 29950 12650 29966 12684
rect 30342 12650 30358 12684
rect 31207 12677 31223 12711
rect 31257 12677 31273 12711
rect 31207 12660 31273 12677
rect 30988 12623 31133 12624
rect 30643 12589 30659 12623
rect 31035 12605 31133 12623
rect 31035 12589 31134 12605
rect 31375 12589 31391 12623
rect 30988 12588 31134 12589
rect 31767 12588 31869 12623
rect 29950 12532 29966 12566
rect 30342 12532 30358 12566
rect 31093 12550 31134 12588
rect 31093 12516 31421 12550
rect 30643 12471 30659 12505
rect 31035 12471 31051 12505
rect 1708 12382 1936 12400
rect 1708 12306 1724 12382
rect 1920 12306 1936 12382
rect 1708 12290 1936 12306
rect 4852 12382 5080 12400
rect 4852 12306 4868 12382
rect 5064 12306 5080 12382
rect 4852 12290 5080 12306
rect 7984 12378 8212 12396
rect 7984 12302 8000 12378
rect 8196 12302 8212 12378
rect 7984 12286 8212 12302
rect 11128 12378 11356 12396
rect 11128 12302 11144 12378
rect 11340 12302 11356 12378
rect 11128 12286 11356 12302
rect 14330 12382 14558 12400
rect 14330 12306 14346 12382
rect 14542 12306 14558 12382
rect 14330 12290 14558 12306
rect 17474 12382 17702 12400
rect 17474 12306 17490 12382
rect 17686 12306 17702 12382
rect 17474 12290 17702 12306
rect 20606 12378 20834 12396
rect 20606 12302 20622 12378
rect 20818 12302 20834 12378
rect 20606 12286 20834 12302
rect 23750 12378 23978 12396
rect 23750 12302 23766 12378
rect 23962 12302 23978 12378
rect 23750 12286 23978 12302
rect 29675 12383 29767 12417
rect 29950 12414 29966 12448
rect 30342 12414 30358 12448
rect 31093 12389 31134 12516
rect 31375 12505 31421 12516
rect 31375 12471 31391 12505
rect 31767 12471 31783 12505
rect 31307 12445 31341 12461
rect 31307 12395 31341 12411
rect 30988 12387 31134 12389
rect 29675 12261 29695 12383
rect 29739 12331 29767 12383
rect 30643 12353 30659 12387
rect 31035 12353 31134 12387
rect 31375 12353 31391 12387
rect 31767 12353 31783 12387
rect 29749 12293 29767 12331
rect 29739 12261 29767 12293
rect 29675 12215 29767 12261
rect 29878 12296 29966 12330
rect 30342 12296 30358 12330
rect 983 12164 1253 12203
rect 983 12112 1017 12164
rect 510 11962 780 11999
rect 510 11912 544 11962
rect 510 11720 544 11736
rect 628 11912 662 11928
rect 628 11682 662 11736
rect 746 11912 780 11962
rect 746 11720 780 11736
rect 864 11912 898 11928
rect 864 11682 898 11736
rect 983 11720 1017 11736
rect 1101 12112 1135 12128
rect 628 11643 898 11682
rect 1101 11685 1135 11736
rect 1219 12112 1253 12164
rect 1456 12164 1726 12203
rect 1219 11720 1253 11736
rect 1337 12112 1371 12128
rect 1337 11685 1371 11736
rect 1456 12112 1490 12164
rect 1456 11720 1490 11736
rect 1574 12112 1608 12128
rect 1574 11685 1608 11736
rect 1692 12112 1726 12164
rect 1928 12164 2198 12203
rect 1692 11720 1726 11736
rect 1810 12112 1844 12128
rect 1810 11685 1844 11736
rect 1928 12112 1962 12164
rect 1928 11720 1962 11736
rect 2046 12112 2080 12128
rect 2046 11685 2080 11736
rect 2164 12112 2198 12164
rect 2395 12165 2665 12204
rect 2164 11720 2198 11736
rect 2277 12112 2311 12128
rect 2277 11685 2311 11736
rect 2395 12112 2429 12165
rect 2395 11720 2429 11736
rect 2513 12112 2547 12128
rect 2513 11685 2547 11736
rect 2631 12112 2665 12165
rect 4127 12164 4397 12203
rect 4127 12112 4161 12164
rect 2836 11963 3106 12002
rect 2631 11720 2665 11736
rect 2718 11912 2752 11928
rect 1101 11646 2547 11685
rect 2718 11685 2752 11736
rect 2836 11912 2870 11963
rect 2836 11720 2870 11736
rect 2954 11912 2988 11928
rect 2954 11685 2988 11736
rect 3072 11912 3106 11963
rect 3072 11720 3106 11736
rect 3654 11962 3924 11999
rect 3654 11912 3688 11962
rect 3654 11720 3688 11736
rect 3772 11912 3806 11928
rect 2718 11646 2988 11685
rect 3772 11682 3806 11736
rect 3890 11912 3924 11962
rect 3890 11720 3924 11736
rect 4008 11912 4042 11928
rect 4008 11682 4042 11736
rect 4127 11720 4161 11736
rect 4245 12112 4279 12128
rect 3772 11643 4042 11682
rect 4245 11685 4279 11736
rect 4363 12112 4397 12164
rect 4600 12164 4870 12203
rect 4363 11720 4397 11736
rect 4481 12112 4515 12128
rect 4481 11685 4515 11736
rect 4600 12112 4634 12164
rect 4600 11720 4634 11736
rect 4718 12112 4752 12128
rect 4718 11685 4752 11736
rect 4836 12112 4870 12164
rect 5072 12164 5342 12203
rect 4836 11720 4870 11736
rect 4954 12112 4988 12128
rect 4954 11685 4988 11736
rect 5072 12112 5106 12164
rect 5072 11720 5106 11736
rect 5190 12112 5224 12128
rect 5190 11685 5224 11736
rect 5308 12112 5342 12164
rect 5539 12165 5809 12204
rect 5308 11720 5342 11736
rect 5421 12112 5455 12128
rect 5421 11685 5455 11736
rect 5539 12112 5573 12165
rect 5539 11720 5573 11736
rect 5657 12112 5691 12128
rect 5657 11685 5691 11736
rect 5775 12112 5809 12165
rect 7259 12160 7529 12199
rect 7259 12108 7293 12160
rect 5980 11963 6250 12002
rect 5775 11720 5809 11736
rect 5862 11912 5896 11928
rect 4245 11646 5691 11685
rect 5862 11685 5896 11736
rect 5980 11912 6014 11963
rect 5980 11720 6014 11736
rect 6098 11912 6132 11928
rect 6098 11685 6132 11736
rect 6216 11912 6250 11963
rect 6216 11720 6250 11736
rect 6786 11958 7056 11995
rect 6786 11908 6820 11958
rect 6786 11716 6820 11732
rect 6904 11908 6938 11924
rect 5862 11646 6132 11685
rect 6904 11678 6938 11732
rect 7022 11908 7056 11958
rect 7022 11716 7056 11732
rect 7140 11908 7174 11924
rect 7140 11678 7174 11732
rect 7259 11716 7293 11732
rect 7377 12108 7411 12124
rect 6904 11639 7174 11678
rect 7377 11681 7411 11732
rect 7495 12108 7529 12160
rect 7732 12160 8002 12199
rect 7495 11716 7529 11732
rect 7613 12108 7647 12124
rect 7613 11681 7647 11732
rect 7732 12108 7766 12160
rect 7732 11716 7766 11732
rect 7850 12108 7884 12124
rect 7850 11681 7884 11732
rect 7968 12108 8002 12160
rect 8204 12160 8474 12199
rect 7968 11716 8002 11732
rect 8086 12108 8120 12124
rect 8086 11681 8120 11732
rect 8204 12108 8238 12160
rect 8204 11716 8238 11732
rect 8322 12108 8356 12124
rect 8322 11681 8356 11732
rect 8440 12108 8474 12160
rect 8671 12161 8941 12200
rect 8440 11716 8474 11732
rect 8553 12108 8587 12124
rect 8553 11681 8587 11732
rect 8671 12108 8705 12161
rect 8671 11716 8705 11732
rect 8789 12108 8823 12124
rect 8789 11681 8823 11732
rect 8907 12108 8941 12161
rect 10403 12160 10673 12199
rect 10403 12108 10437 12160
rect 9112 11959 9382 11998
rect 8907 11716 8941 11732
rect 8994 11908 9028 11924
rect 7377 11642 8823 11681
rect 8994 11681 9028 11732
rect 9112 11908 9146 11959
rect 9112 11716 9146 11732
rect 9230 11908 9264 11924
rect 9230 11681 9264 11732
rect 9348 11908 9382 11959
rect 9348 11716 9382 11732
rect 9930 11958 10200 11995
rect 9930 11908 9964 11958
rect 9930 11716 9964 11732
rect 10048 11908 10082 11924
rect 8994 11642 9264 11681
rect 10048 11678 10082 11732
rect 10166 11908 10200 11958
rect 10166 11716 10200 11732
rect 10284 11908 10318 11924
rect 10284 11678 10318 11732
rect 10403 11716 10437 11732
rect 10521 12108 10555 12124
rect 10048 11639 10318 11678
rect 10521 11681 10555 11732
rect 10639 12108 10673 12160
rect 10876 12160 11146 12199
rect 10639 11716 10673 11732
rect 10757 12108 10791 12124
rect 10757 11681 10791 11732
rect 10876 12108 10910 12160
rect 10876 11716 10910 11732
rect 10994 12108 11028 12124
rect 10994 11681 11028 11732
rect 11112 12108 11146 12160
rect 11348 12160 11618 12199
rect 11112 11716 11146 11732
rect 11230 12108 11264 12124
rect 11230 11681 11264 11732
rect 11348 12108 11382 12160
rect 11348 11716 11382 11732
rect 11466 12108 11500 12124
rect 11466 11681 11500 11732
rect 11584 12108 11618 12160
rect 11815 12161 12085 12200
rect 11584 11716 11618 11732
rect 11697 12108 11731 12124
rect 11697 11681 11731 11732
rect 11815 12108 11849 12161
rect 11815 11716 11849 11732
rect 11933 12108 11967 12124
rect 11933 11681 11967 11732
rect 12051 12108 12085 12161
rect 13605 12164 13875 12203
rect 13605 12112 13639 12164
rect 12256 11959 12526 11998
rect 12051 11716 12085 11732
rect 12138 11908 12172 11924
rect 10521 11642 11967 11681
rect 12138 11681 12172 11732
rect 12256 11908 12290 11959
rect 12256 11716 12290 11732
rect 12374 11908 12408 11924
rect 12374 11681 12408 11732
rect 12492 11908 12526 11959
rect 12492 11716 12526 11732
rect 13132 11962 13402 11999
rect 13132 11912 13166 11962
rect 13132 11720 13166 11736
rect 13250 11912 13284 11928
rect 12138 11642 12408 11681
rect 13250 11682 13284 11736
rect 13368 11912 13402 11962
rect 13368 11720 13402 11736
rect 13486 11912 13520 11928
rect 13486 11682 13520 11736
rect 13605 11720 13639 11736
rect 13723 12112 13757 12128
rect 13250 11643 13520 11682
rect 13723 11685 13757 11736
rect 13841 12112 13875 12164
rect 14078 12164 14348 12203
rect 13841 11720 13875 11736
rect 13959 12112 13993 12128
rect 13959 11685 13993 11736
rect 14078 12112 14112 12164
rect 14078 11720 14112 11736
rect 14196 12112 14230 12128
rect 14196 11685 14230 11736
rect 14314 12112 14348 12164
rect 14550 12164 14820 12203
rect 14314 11720 14348 11736
rect 14432 12112 14466 12128
rect 14432 11685 14466 11736
rect 14550 12112 14584 12164
rect 14550 11720 14584 11736
rect 14668 12112 14702 12128
rect 14668 11685 14702 11736
rect 14786 12112 14820 12164
rect 15017 12165 15287 12204
rect 14786 11720 14820 11736
rect 14899 12112 14933 12128
rect 14899 11685 14933 11736
rect 15017 12112 15051 12165
rect 15017 11720 15051 11736
rect 15135 12112 15169 12128
rect 15135 11685 15169 11736
rect 15253 12112 15287 12165
rect 16749 12164 17019 12203
rect 16749 12112 16783 12164
rect 15458 11963 15728 12002
rect 15253 11720 15287 11736
rect 15340 11912 15374 11928
rect 13723 11646 15169 11685
rect 15340 11685 15374 11736
rect 15458 11912 15492 11963
rect 15458 11720 15492 11736
rect 15576 11912 15610 11928
rect 15576 11685 15610 11736
rect 15694 11912 15728 11963
rect 15694 11720 15728 11736
rect 16276 11962 16546 11999
rect 16276 11912 16310 11962
rect 16276 11720 16310 11736
rect 16394 11912 16428 11928
rect 15340 11646 15610 11685
rect 16394 11682 16428 11736
rect 16512 11912 16546 11962
rect 16512 11720 16546 11736
rect 16630 11912 16664 11928
rect 16630 11682 16664 11736
rect 16749 11720 16783 11736
rect 16867 12112 16901 12128
rect 16394 11643 16664 11682
rect 16867 11685 16901 11736
rect 16985 12112 17019 12164
rect 17222 12164 17492 12203
rect 16985 11720 17019 11736
rect 17103 12112 17137 12128
rect 17103 11685 17137 11736
rect 17222 12112 17256 12164
rect 17222 11720 17256 11736
rect 17340 12112 17374 12128
rect 17340 11685 17374 11736
rect 17458 12112 17492 12164
rect 17694 12164 17964 12203
rect 17458 11720 17492 11736
rect 17576 12112 17610 12128
rect 17576 11685 17610 11736
rect 17694 12112 17728 12164
rect 17694 11720 17728 11736
rect 17812 12112 17846 12128
rect 17812 11685 17846 11736
rect 17930 12112 17964 12164
rect 18161 12165 18431 12204
rect 17930 11720 17964 11736
rect 18043 12112 18077 12128
rect 18043 11685 18077 11736
rect 18161 12112 18195 12165
rect 18161 11720 18195 11736
rect 18279 12112 18313 12128
rect 18279 11685 18313 11736
rect 18397 12112 18431 12165
rect 19881 12160 20151 12199
rect 19881 12108 19915 12160
rect 18602 11963 18872 12002
rect 18397 11720 18431 11736
rect 18484 11912 18518 11928
rect 16867 11646 18313 11685
rect 18484 11685 18518 11736
rect 18602 11912 18636 11963
rect 18602 11720 18636 11736
rect 18720 11912 18754 11928
rect 18720 11685 18754 11736
rect 18838 11912 18872 11963
rect 18838 11720 18872 11736
rect 19408 11958 19678 11995
rect 19408 11908 19442 11958
rect 19408 11716 19442 11732
rect 19526 11908 19560 11924
rect 18484 11646 18754 11685
rect 19526 11678 19560 11732
rect 19644 11908 19678 11958
rect 19644 11716 19678 11732
rect 19762 11908 19796 11924
rect 19762 11678 19796 11732
rect 19881 11716 19915 11732
rect 19999 12108 20033 12124
rect 19526 11639 19796 11678
rect 19999 11681 20033 11732
rect 20117 12108 20151 12160
rect 20354 12160 20624 12199
rect 20117 11716 20151 11732
rect 20235 12108 20269 12124
rect 20235 11681 20269 11732
rect 20354 12108 20388 12160
rect 20354 11716 20388 11732
rect 20472 12108 20506 12124
rect 20472 11681 20506 11732
rect 20590 12108 20624 12160
rect 20826 12160 21096 12199
rect 20590 11716 20624 11732
rect 20708 12108 20742 12124
rect 20708 11681 20742 11732
rect 20826 12108 20860 12160
rect 20826 11716 20860 11732
rect 20944 12108 20978 12124
rect 20944 11681 20978 11732
rect 21062 12108 21096 12160
rect 21293 12161 21563 12200
rect 21062 11716 21096 11732
rect 21175 12108 21209 12124
rect 21175 11681 21209 11732
rect 21293 12108 21327 12161
rect 21293 11716 21327 11732
rect 21411 12108 21445 12124
rect 21411 11681 21445 11732
rect 21529 12108 21563 12161
rect 23025 12160 23295 12199
rect 23025 12108 23059 12160
rect 21734 11959 22004 11998
rect 21529 11716 21563 11732
rect 21616 11908 21650 11924
rect 19999 11642 21445 11681
rect 21616 11681 21650 11732
rect 21734 11908 21768 11959
rect 21734 11716 21768 11732
rect 21852 11908 21886 11924
rect 21852 11681 21886 11732
rect 21970 11908 22004 11959
rect 21970 11716 22004 11732
rect 22552 11958 22822 11995
rect 22552 11908 22586 11958
rect 22552 11716 22586 11732
rect 22670 11908 22704 11924
rect 21616 11642 21886 11681
rect 22670 11678 22704 11732
rect 22788 11908 22822 11958
rect 22788 11716 22822 11732
rect 22906 11908 22940 11924
rect 22906 11678 22940 11732
rect 23025 11716 23059 11732
rect 23143 12108 23177 12124
rect 22670 11639 22940 11678
rect 23143 11681 23177 11732
rect 23261 12108 23295 12160
rect 23498 12160 23768 12199
rect 23261 11716 23295 11732
rect 23379 12108 23413 12124
rect 23379 11681 23413 11732
rect 23498 12108 23532 12160
rect 23498 11716 23532 11732
rect 23616 12108 23650 12124
rect 23616 11681 23650 11732
rect 23734 12108 23768 12160
rect 23970 12160 24240 12199
rect 23734 11716 23768 11732
rect 23852 12108 23886 12124
rect 23852 11681 23886 11732
rect 23970 12108 24004 12160
rect 23970 11716 24004 11732
rect 24088 12108 24122 12124
rect 24088 11681 24122 11732
rect 24206 12108 24240 12160
rect 24437 12161 24707 12200
rect 24206 11716 24240 11732
rect 24319 12108 24353 12124
rect 24319 11681 24353 11732
rect 24437 12108 24471 12161
rect 24437 11716 24471 11732
rect 24555 12108 24589 12124
rect 24555 11681 24589 11732
rect 24673 12108 24707 12161
rect 29878 12094 29913 12296
rect 30643 12235 30659 12269
rect 31035 12235 31051 12269
rect 29950 12178 29966 12212
rect 30342 12178 30358 12212
rect 31093 12151 31134 12353
rect 31306 12327 31340 12343
rect 31306 12277 31340 12293
rect 31375 12235 31391 12269
rect 31767 12235 31783 12269
rect 31834 12152 31869 12588
rect 31939 12433 32027 12449
rect 31939 12393 31955 12433
rect 31939 12301 31955 12343
rect 32011 12301 32027 12433
rect 31939 12285 32027 12301
rect 30643 12117 30659 12151
rect 31035 12117 31134 12151
rect 31375 12117 31391 12151
rect 31767 12117 31869 12152
rect 30989 12115 31134 12117
rect 29878 12060 29966 12094
rect 30342 12060 30358 12094
rect 30643 11999 30659 12033
rect 31035 11999 31051 12033
rect 24878 11959 25148 11998
rect 24673 11716 24707 11732
rect 24760 11908 24794 11924
rect 23143 11642 24589 11681
rect 24760 11681 24794 11732
rect 24878 11908 24912 11959
rect 24878 11716 24912 11732
rect 24996 11908 25030 11924
rect 24996 11681 25030 11732
rect 25114 11908 25148 11959
rect 29950 11942 29966 11976
rect 30342 11942 30358 11976
rect 30150 11813 30166 11847
rect 30342 11813 30358 11847
rect 30521 11761 30555 11767
rect 25114 11716 25148 11732
rect 30150 11695 30166 11729
rect 30342 11695 30358 11729
rect 30521 11701 30555 11707
rect 24760 11642 25030 11681
rect 30150 11577 30166 11611
rect 30342 11577 30358 11611
rect 660 11528 676 11562
rect 710 11528 726 11562
rect 1986 11521 2020 11537
rect 3804 11528 3820 11562
rect 3854 11528 3870 11562
rect 1986 11471 2020 11487
rect 5130 11521 5164 11537
rect 6936 11524 6952 11558
rect 6986 11524 7002 11558
rect 5130 11471 5164 11487
rect 8262 11517 8296 11533
rect 10080 11524 10096 11558
rect 10130 11524 10146 11558
rect 8262 11467 8296 11483
rect 11406 11517 11440 11533
rect 13282 11528 13298 11562
rect 13332 11528 13348 11562
rect 11406 11467 11440 11483
rect 14608 11521 14642 11537
rect 16426 11528 16442 11562
rect 16476 11528 16492 11562
rect 14608 11471 14642 11487
rect 17752 11521 17786 11537
rect 19558 11524 19574 11558
rect 19608 11524 19624 11558
rect 17752 11471 17786 11487
rect 20884 11517 20918 11533
rect 22702 11524 22718 11558
rect 22752 11524 22768 11558
rect 20884 11467 20918 11483
rect 24028 11517 24062 11533
rect 31093 11529 31134 12115
rect 31207 12063 31273 12080
rect 31207 12029 31223 12063
rect 31257 12029 31273 12063
rect 31207 12013 31273 12029
rect 31275 11739 31291 11773
rect 31325 11739 31341 11773
rect 31375 11711 31391 11745
rect 31567 11711 31583 11745
rect 31375 11593 31391 11627
rect 31567 11593 31583 11627
rect 24028 11467 24062 11483
rect 30150 11459 30166 11493
rect 30342 11459 30358 11493
rect 1840 11422 1932 11435
rect 1840 11367 1856 11422
rect 1916 11367 1932 11422
rect 1840 11350 1932 11367
rect 2925 11421 3017 11438
rect 2925 11366 2941 11421
rect 3001 11366 3017 11421
rect 2925 11353 3017 11366
rect 4984 11422 5076 11435
rect 4984 11367 5000 11422
rect 5060 11367 5076 11422
rect 4984 11350 5076 11367
rect 6069 11421 6161 11438
rect 6069 11366 6085 11421
rect 6145 11366 6161 11421
rect 6069 11353 6161 11366
rect 8116 11418 8208 11431
rect 8116 11363 8132 11418
rect 8192 11363 8208 11418
rect 8116 11346 8208 11363
rect 9201 11417 9293 11434
rect 9201 11362 9217 11417
rect 9277 11362 9293 11417
rect 9201 11349 9293 11362
rect 9468 11418 9525 11422
rect 9468 11358 9472 11418
rect 9521 11358 9525 11418
rect 9468 11354 9525 11358
rect 11260 11418 11352 11431
rect 11260 11363 11276 11418
rect 11336 11363 11352 11418
rect 11260 11346 11352 11363
rect 12345 11417 12437 11434
rect 12345 11362 12361 11417
rect 12421 11362 12437 11417
rect 12345 11349 12437 11362
rect 14462 11422 14554 11435
rect 14462 11367 14478 11422
rect 14538 11367 14554 11422
rect 14462 11350 14554 11367
rect 15547 11421 15639 11438
rect 15547 11366 15563 11421
rect 15623 11366 15639 11421
rect 15547 11353 15639 11366
rect 17606 11422 17698 11435
rect 17606 11367 17622 11422
rect 17682 11367 17698 11422
rect 17606 11350 17698 11367
rect 18691 11421 18783 11438
rect 18691 11366 18707 11421
rect 18767 11366 18783 11421
rect 18691 11353 18783 11366
rect 20738 11418 20830 11431
rect 20738 11363 20754 11418
rect 20814 11363 20830 11418
rect 20738 11346 20830 11363
rect 21823 11417 21915 11434
rect 21823 11362 21839 11417
rect 21899 11362 21915 11417
rect 21823 11349 21915 11362
rect 23882 11418 23974 11431
rect 23882 11363 23898 11418
rect 23958 11363 23974 11418
rect 23882 11346 23974 11363
rect 24967 11417 25059 11434
rect 24967 11362 24983 11417
rect 25043 11362 25059 11417
rect 24967 11349 25059 11362
rect 1632 11291 1666 11307
rect 1632 11241 1666 11257
rect 3192 11306 3249 11310
rect 3192 11246 3196 11306
rect 3245 11246 3249 11306
rect 3192 11242 3249 11246
rect 4776 11291 4810 11307
rect 4776 11241 4810 11257
rect 6336 11306 6393 11310
rect 6336 11246 6340 11306
rect 6389 11246 6393 11306
rect 6336 11242 6393 11246
rect 7908 11287 7942 11303
rect 7908 11237 7942 11253
rect 9468 11302 9525 11306
rect 9468 11242 9472 11302
rect 9521 11242 9525 11302
rect 9468 11238 9525 11242
rect 11052 11287 11086 11303
rect 11052 11237 11086 11253
rect 12612 11302 12669 11306
rect 12612 11242 12616 11302
rect 12665 11242 12669 11302
rect 12612 11238 12669 11242
rect 14254 11291 14288 11307
rect 14254 11241 14288 11257
rect 15814 11306 15871 11310
rect 15814 11246 15818 11306
rect 15867 11246 15871 11306
rect 15814 11242 15871 11246
rect 17398 11291 17432 11307
rect 17398 11241 17432 11257
rect 18958 11306 19015 11310
rect 18958 11246 18962 11306
rect 19011 11246 19015 11306
rect 18958 11242 19015 11246
rect 20530 11287 20564 11303
rect 20530 11237 20564 11253
rect 22090 11302 22147 11306
rect 22090 11242 22094 11302
rect 22143 11242 22147 11302
rect 22090 11238 22147 11242
rect 23674 11287 23708 11303
rect 23674 11237 23708 11253
rect 25234 11302 25291 11306
rect 25234 11242 25238 11302
rect 25287 11242 25291 11302
rect 25234 11238 25291 11242
rect 1958 11137 2050 11150
rect 1958 11082 1974 11137
rect 2034 11082 2050 11137
rect 1958 11065 2050 11082
rect 3192 11138 3249 11142
rect 3192 11078 3196 11138
rect 3245 11078 3249 11138
rect 3192 11074 3249 11078
rect 5102 11137 5194 11150
rect 5102 11082 5118 11137
rect 5178 11082 5194 11137
rect 5102 11065 5194 11082
rect 6336 11138 6393 11142
rect 6336 11078 6340 11138
rect 6389 11078 6393 11138
rect 6336 11074 6393 11078
rect 8234 11133 8326 11146
rect 8234 11078 8250 11133
rect 8310 11078 8326 11133
rect 8234 11061 8326 11078
rect 9468 11134 9525 11138
rect 9468 11074 9472 11134
rect 9521 11074 9525 11134
rect 9468 11070 9525 11074
rect 11378 11133 11470 11146
rect 11378 11078 11394 11133
rect 11454 11078 11470 11133
rect 11378 11061 11470 11078
rect 12612 11134 12669 11138
rect 12612 11074 12616 11134
rect 12665 11074 12669 11134
rect 12612 11070 12669 11074
rect 14580 11137 14672 11150
rect 14580 11082 14596 11137
rect 14656 11082 14672 11137
rect 14580 11065 14672 11082
rect 15814 11138 15871 11142
rect 15814 11078 15818 11138
rect 15867 11078 15871 11138
rect 15814 11074 15871 11078
rect 17724 11137 17816 11150
rect 17724 11082 17740 11137
rect 17800 11082 17816 11137
rect 17724 11065 17816 11082
rect 18958 11138 19015 11142
rect 18958 11078 18962 11138
rect 19011 11078 19015 11138
rect 18958 11074 19015 11078
rect 20856 11133 20948 11146
rect 20856 11078 20872 11133
rect 20932 11078 20948 11133
rect 20856 11061 20948 11078
rect 22090 11134 22147 11138
rect 22090 11074 22094 11134
rect 22143 11074 22147 11134
rect 22090 11070 22147 11074
rect 24000 11133 24092 11146
rect 24000 11078 24016 11133
rect 24076 11078 24092 11133
rect 24000 11061 24092 11078
rect 25234 11134 25291 11138
rect 25234 11074 25238 11134
rect 25287 11074 25291 11134
rect 25234 11070 25291 11074
rect 30075 11066 30164 11100
rect 30340 11066 30356 11100
rect 1751 10901 1785 10917
rect 1751 10851 1785 10867
rect 4895 10901 4929 10917
rect 4895 10851 4929 10867
rect 8027 10897 8061 10913
rect 8027 10847 8061 10863
rect 11171 10897 11205 10913
rect 11171 10847 11205 10863
rect 14373 10901 14407 10917
rect 14373 10851 14407 10867
rect 17517 10901 17551 10917
rect 17517 10851 17551 10867
rect 20649 10897 20683 10913
rect 20649 10847 20683 10863
rect 23793 10897 23827 10913
rect 23793 10847 23827 10863
rect 30075 10864 30110 11066
rect 30148 10948 30164 10982
rect 30340 10948 30356 10982
rect 31373 10941 31389 10975
rect 31565 10941 31581 10975
rect 30075 10830 30164 10864
rect 30340 10830 30356 10864
rect 1378 10779 1412 10795
rect 1378 10587 1412 10603
rect 1496 10791 1530 10795
rect 1574 10791 1608 10795
rect 1496 10779 1608 10791
rect 1530 10603 1574 10779
rect 1496 10591 1574 10603
rect 1496 10587 1530 10591
rect 1574 10387 1608 10403
rect 1692 10779 1726 10795
rect 1692 10387 1726 10403
rect 1810 10779 1844 10795
rect 1810 10387 1844 10403
rect 1928 10779 1962 10795
rect 1928 10387 1962 10403
rect 2046 10791 2080 10795
rect 2120 10791 2154 10795
rect 2046 10779 2154 10791
rect 2080 10603 2120 10779
rect 2080 10591 2154 10603
rect 2120 10587 2154 10591
rect 2238 10779 2272 10795
rect 2238 10587 2272 10603
rect 4522 10779 4556 10795
rect 4522 10587 4556 10603
rect 4640 10791 4674 10795
rect 4718 10791 4752 10795
rect 4640 10779 4752 10791
rect 4674 10603 4718 10779
rect 4640 10591 4718 10603
rect 4640 10587 4674 10591
rect 2046 10387 2080 10403
rect 4718 10387 4752 10403
rect 4836 10779 4870 10795
rect 4836 10387 4870 10403
rect 4954 10779 4988 10795
rect 4954 10387 4988 10403
rect 5072 10779 5106 10795
rect 5072 10387 5106 10403
rect 5190 10791 5224 10795
rect 5264 10791 5298 10795
rect 5190 10779 5298 10791
rect 5224 10603 5264 10779
rect 5224 10591 5298 10603
rect 5264 10587 5298 10591
rect 5382 10779 5416 10795
rect 5382 10587 5416 10603
rect 7654 10775 7688 10791
rect 7654 10583 7688 10599
rect 7772 10787 7806 10791
rect 7850 10787 7884 10791
rect 7772 10775 7884 10787
rect 7806 10599 7850 10775
rect 7772 10587 7850 10599
rect 7772 10583 7806 10587
rect 5190 10387 5224 10403
rect 7850 10383 7884 10399
rect 7968 10775 8002 10791
rect 7968 10383 8002 10399
rect 8086 10775 8120 10791
rect 8086 10383 8120 10399
rect 8204 10775 8238 10791
rect 8204 10383 8238 10399
rect 8322 10787 8356 10791
rect 8396 10787 8430 10791
rect 8322 10775 8430 10787
rect 8356 10599 8396 10775
rect 8356 10587 8430 10599
rect 8396 10583 8430 10587
rect 8514 10775 8548 10791
rect 8514 10583 8548 10599
rect 10798 10775 10832 10791
rect 10798 10583 10832 10599
rect 10916 10787 10950 10791
rect 10994 10787 11028 10791
rect 10916 10775 11028 10787
rect 10950 10599 10994 10775
rect 10916 10587 10994 10599
rect 10916 10583 10950 10587
rect 8322 10383 8356 10399
rect 10994 10383 11028 10399
rect 11112 10775 11146 10791
rect 11112 10383 11146 10399
rect 11230 10775 11264 10791
rect 11230 10383 11264 10399
rect 11348 10775 11382 10791
rect 11348 10383 11382 10399
rect 11466 10787 11500 10791
rect 11540 10787 11574 10791
rect 11466 10775 11574 10787
rect 11500 10599 11540 10775
rect 11500 10587 11574 10599
rect 11540 10583 11574 10587
rect 11658 10775 11692 10791
rect 11658 10583 11692 10599
rect 14000 10779 14034 10795
rect 14000 10587 14034 10603
rect 14118 10791 14152 10795
rect 14196 10791 14230 10795
rect 14118 10779 14230 10791
rect 14152 10603 14196 10779
rect 14118 10591 14196 10603
rect 14118 10587 14152 10591
rect 11466 10383 11500 10399
rect 14196 10387 14230 10403
rect 14314 10779 14348 10795
rect 14314 10387 14348 10403
rect 14432 10779 14466 10795
rect 14432 10387 14466 10403
rect 14550 10779 14584 10795
rect 14550 10387 14584 10403
rect 14668 10791 14702 10795
rect 14742 10791 14776 10795
rect 14668 10779 14776 10791
rect 14702 10603 14742 10779
rect 14702 10591 14776 10603
rect 14742 10587 14776 10591
rect 14860 10779 14894 10795
rect 14860 10587 14894 10603
rect 17144 10779 17178 10795
rect 17144 10587 17178 10603
rect 17262 10791 17296 10795
rect 17340 10791 17374 10795
rect 17262 10779 17374 10791
rect 17296 10603 17340 10779
rect 17262 10591 17340 10603
rect 17262 10587 17296 10591
rect 14668 10387 14702 10403
rect 17340 10387 17374 10403
rect 17458 10779 17492 10795
rect 17458 10387 17492 10403
rect 17576 10779 17610 10795
rect 17576 10387 17610 10403
rect 17694 10779 17728 10795
rect 17694 10387 17728 10403
rect 17812 10791 17846 10795
rect 17886 10791 17920 10795
rect 17812 10779 17920 10791
rect 17846 10603 17886 10779
rect 17846 10591 17920 10603
rect 17886 10587 17920 10591
rect 18004 10779 18038 10795
rect 31272 10794 31288 10828
rect 31322 10794 31338 10828
rect 31373 10823 31389 10857
rect 31565 10823 31581 10857
rect 18004 10587 18038 10603
rect 20276 10775 20310 10791
rect 20276 10583 20310 10599
rect 20394 10787 20428 10791
rect 20472 10787 20506 10791
rect 20394 10775 20506 10787
rect 20428 10599 20472 10775
rect 20394 10587 20472 10599
rect 20394 10583 20428 10587
rect 17812 10387 17846 10403
rect 20472 10383 20506 10399
rect 20590 10775 20624 10791
rect 20590 10383 20624 10399
rect 20708 10775 20742 10791
rect 20708 10383 20742 10399
rect 20826 10775 20860 10791
rect 20826 10383 20860 10399
rect 20944 10787 20978 10791
rect 21018 10787 21052 10791
rect 20944 10775 21052 10787
rect 20978 10599 21018 10775
rect 20978 10587 21052 10599
rect 21018 10583 21052 10587
rect 21136 10775 21170 10791
rect 21136 10583 21170 10599
rect 23420 10775 23454 10791
rect 23420 10583 23454 10599
rect 23538 10787 23572 10791
rect 23616 10787 23650 10791
rect 23538 10775 23650 10787
rect 23572 10599 23616 10775
rect 23538 10587 23616 10599
rect 23538 10583 23572 10587
rect 20944 10383 20978 10399
rect 23616 10383 23650 10399
rect 23734 10775 23768 10791
rect 23734 10383 23768 10399
rect 23852 10775 23886 10791
rect 23852 10383 23886 10399
rect 23970 10775 24004 10791
rect 23970 10383 24004 10399
rect 24088 10787 24122 10791
rect 24162 10787 24196 10791
rect 24088 10775 24196 10787
rect 24122 10599 24162 10775
rect 24122 10587 24196 10599
rect 24162 10583 24196 10587
rect 24280 10775 24314 10791
rect 30148 10712 30164 10746
rect 30340 10712 30356 10746
rect 30641 10639 30657 10673
rect 31033 10639 31049 10673
rect 31205 10643 31271 10659
rect 24280 10583 24314 10599
rect 29948 10582 29964 10616
rect 30340 10582 30356 10616
rect 31205 10609 31221 10643
rect 31255 10609 31271 10643
rect 31205 10592 31271 10609
rect 30986 10555 31131 10556
rect 30641 10521 30657 10555
rect 31033 10537 31131 10555
rect 31033 10521 31132 10537
rect 31373 10521 31389 10555
rect 30986 10520 31132 10521
rect 31765 10520 31867 10555
rect 29948 10464 29964 10498
rect 30340 10464 30356 10498
rect 31091 10482 31132 10520
rect 31091 10448 31419 10482
rect 30641 10403 30657 10437
rect 31033 10403 31049 10437
rect 24088 10383 24122 10399
rect 29673 10315 29765 10349
rect 29948 10346 29964 10380
rect 30340 10346 30356 10380
rect 31091 10321 31132 10448
rect 31373 10437 31419 10448
rect 31373 10403 31389 10437
rect 31765 10403 31781 10437
rect 31305 10377 31339 10393
rect 31305 10327 31339 10343
rect 30986 10319 31132 10321
rect 1793 10268 1809 10302
rect 1843 10268 1859 10302
rect 4937 10268 4953 10302
rect 4987 10268 5003 10302
rect 8069 10264 8085 10298
rect 8119 10264 8135 10298
rect 11213 10264 11229 10298
rect 11263 10264 11279 10298
rect 14415 10268 14431 10302
rect 14465 10268 14481 10302
rect 17559 10268 17575 10302
rect 17609 10268 17625 10302
rect 20691 10264 20707 10298
rect 20741 10264 20757 10298
rect 23835 10264 23851 10298
rect 23885 10264 23901 10298
rect 29673 10193 29693 10315
rect 29737 10263 29765 10315
rect 30641 10285 30657 10319
rect 31033 10285 31132 10319
rect 31373 10285 31389 10319
rect 31765 10285 31781 10319
rect 29747 10225 29765 10263
rect 29737 10193 29765 10225
rect 1742 10150 1878 10154
rect 1742 10136 1782 10150
rect 1840 10136 1878 10150
rect 1742 10090 1758 10136
rect 1862 10090 1878 10136
rect 1742 10068 1878 10090
rect 4886 10150 5022 10154
rect 14364 10150 14500 10154
rect 4886 10136 4926 10150
rect 4984 10136 5022 10150
rect 4886 10090 4902 10136
rect 5006 10090 5022 10136
rect 4886 10068 5022 10090
rect 8018 10146 8154 10150
rect 8018 10132 8058 10146
rect 8116 10132 8154 10146
rect 8018 10086 8034 10132
rect 8138 10086 8154 10132
rect 8018 10064 8154 10086
rect 11162 10146 11298 10150
rect 11162 10132 11202 10146
rect 11260 10132 11298 10146
rect 11162 10086 11178 10132
rect 11282 10086 11298 10132
rect 11162 10064 11298 10086
rect 14364 10136 14404 10150
rect 14462 10136 14500 10150
rect 14364 10090 14380 10136
rect 14484 10090 14500 10136
rect 14364 10068 14500 10090
rect 17508 10150 17644 10154
rect 17508 10136 17548 10150
rect 17606 10136 17644 10150
rect 17508 10090 17524 10136
rect 17628 10090 17644 10136
rect 17508 10068 17644 10090
rect 20640 10146 20776 10150
rect 20640 10132 20680 10146
rect 20738 10132 20776 10146
rect 20640 10086 20656 10132
rect 20760 10086 20776 10132
rect 20640 10064 20776 10086
rect 23784 10146 23920 10150
rect 29673 10147 29765 10193
rect 29876 10228 29964 10262
rect 30340 10228 30356 10262
rect 23784 10132 23824 10146
rect 23882 10132 23920 10146
rect 23784 10086 23800 10132
rect 23904 10086 23920 10132
rect 23784 10064 23920 10086
rect 29876 10026 29911 10228
rect 30641 10167 30657 10201
rect 31033 10167 31049 10201
rect 29948 10110 29964 10144
rect 30340 10110 30356 10144
rect 31091 10083 31132 10285
rect 31304 10259 31338 10275
rect 31304 10209 31338 10225
rect 31373 10167 31389 10201
rect 31765 10167 31781 10201
rect 31832 10084 31867 10520
rect 31937 10365 32025 10381
rect 31937 10325 31953 10365
rect 31937 10233 31953 10275
rect 32009 10233 32025 10365
rect 31937 10217 32025 10233
rect 30641 10049 30657 10083
rect 31033 10049 31132 10083
rect 31373 10049 31389 10083
rect 31765 10049 31867 10084
rect 30987 10047 31132 10049
rect 29876 9992 29964 10026
rect 30340 9992 30356 10026
rect 30641 9931 30657 9965
rect 31033 9931 31049 9965
rect 29948 9874 29964 9908
rect 30340 9874 30356 9908
rect 30148 9745 30164 9779
rect 30340 9745 30356 9779
rect 30519 9693 30553 9699
rect 1718 9650 1946 9668
rect 1718 9574 1734 9650
rect 1930 9574 1946 9650
rect 1718 9558 1946 9574
rect 4862 9650 5090 9668
rect 4862 9574 4878 9650
rect 5074 9574 5090 9650
rect 4862 9558 5090 9574
rect 7994 9646 8222 9664
rect 7994 9570 8010 9646
rect 8206 9570 8222 9646
rect 7994 9554 8222 9570
rect 11138 9646 11366 9664
rect 11138 9570 11154 9646
rect 11350 9570 11366 9646
rect 11138 9554 11366 9570
rect 14340 9650 14568 9668
rect 14340 9574 14356 9650
rect 14552 9574 14568 9650
rect 14340 9558 14568 9574
rect 17484 9650 17712 9668
rect 17484 9574 17500 9650
rect 17696 9574 17712 9650
rect 17484 9558 17712 9574
rect 20616 9646 20844 9664
rect 20616 9570 20632 9646
rect 20828 9570 20844 9646
rect 20616 9554 20844 9570
rect 23760 9646 23988 9664
rect 23760 9570 23776 9646
rect 23972 9570 23988 9646
rect 30148 9627 30164 9661
rect 30340 9627 30356 9661
rect 30519 9633 30553 9639
rect 23760 9554 23988 9570
rect 30148 9509 30164 9543
rect 30340 9509 30356 9543
rect 993 9432 1263 9471
rect 993 9380 1027 9432
rect 520 9230 790 9267
rect 520 9180 554 9230
rect 520 8988 554 9004
rect 638 9180 672 9196
rect 638 8950 672 9004
rect 756 9180 790 9230
rect 756 8988 790 9004
rect 874 9180 908 9196
rect 874 8950 908 9004
rect 993 8988 1027 9004
rect 1111 9380 1145 9396
rect 638 8911 908 8950
rect 1111 8953 1145 9004
rect 1229 9380 1263 9432
rect 1466 9432 1736 9471
rect 1229 8988 1263 9004
rect 1347 9380 1381 9396
rect 1347 8953 1381 9004
rect 1466 9380 1500 9432
rect 1466 8988 1500 9004
rect 1584 9380 1618 9396
rect 1584 8953 1618 9004
rect 1702 9380 1736 9432
rect 1938 9432 2208 9471
rect 1702 8988 1736 9004
rect 1820 9380 1854 9396
rect 1820 8953 1854 9004
rect 1938 9380 1972 9432
rect 1938 8988 1972 9004
rect 2056 9380 2090 9396
rect 2056 8953 2090 9004
rect 2174 9380 2208 9432
rect 2405 9433 2675 9472
rect 2174 8988 2208 9004
rect 2287 9380 2321 9396
rect 2287 8953 2321 9004
rect 2405 9380 2439 9433
rect 2405 8988 2439 9004
rect 2523 9380 2557 9396
rect 2523 8953 2557 9004
rect 2641 9380 2675 9433
rect 4137 9432 4407 9471
rect 4137 9380 4171 9432
rect 2846 9231 3116 9270
rect 2641 8988 2675 9004
rect 2728 9180 2762 9196
rect 1111 8914 2557 8953
rect 2728 8953 2762 9004
rect 2846 9180 2880 9231
rect 2846 8988 2880 9004
rect 2964 9180 2998 9196
rect 2964 8953 2998 9004
rect 3082 9180 3116 9231
rect 3082 8988 3116 9004
rect 3664 9230 3934 9267
rect 3664 9180 3698 9230
rect 3664 8988 3698 9004
rect 3782 9180 3816 9196
rect 2728 8914 2998 8953
rect 3782 8950 3816 9004
rect 3900 9180 3934 9230
rect 3900 8988 3934 9004
rect 4018 9180 4052 9196
rect 4018 8950 4052 9004
rect 4137 8988 4171 9004
rect 4255 9380 4289 9396
rect 3782 8911 4052 8950
rect 4255 8953 4289 9004
rect 4373 9380 4407 9432
rect 4610 9432 4880 9471
rect 4373 8988 4407 9004
rect 4491 9380 4525 9396
rect 4491 8953 4525 9004
rect 4610 9380 4644 9432
rect 4610 8988 4644 9004
rect 4728 9380 4762 9396
rect 4728 8953 4762 9004
rect 4846 9380 4880 9432
rect 5082 9432 5352 9471
rect 4846 8988 4880 9004
rect 4964 9380 4998 9396
rect 4964 8953 4998 9004
rect 5082 9380 5116 9432
rect 5082 8988 5116 9004
rect 5200 9380 5234 9396
rect 5200 8953 5234 9004
rect 5318 9380 5352 9432
rect 5549 9433 5819 9472
rect 5318 8988 5352 9004
rect 5431 9380 5465 9396
rect 5431 8953 5465 9004
rect 5549 9380 5583 9433
rect 5549 8988 5583 9004
rect 5667 9380 5701 9396
rect 5667 8953 5701 9004
rect 5785 9380 5819 9433
rect 7269 9428 7539 9467
rect 7269 9376 7303 9428
rect 5990 9231 6260 9270
rect 5785 8988 5819 9004
rect 5872 9180 5906 9196
rect 4255 8914 5701 8953
rect 5872 8953 5906 9004
rect 5990 9180 6024 9231
rect 5990 8988 6024 9004
rect 6108 9180 6142 9196
rect 6108 8953 6142 9004
rect 6226 9180 6260 9231
rect 6226 8988 6260 9004
rect 6796 9226 7066 9263
rect 6796 9176 6830 9226
rect 6796 8984 6830 9000
rect 6914 9176 6948 9192
rect 5872 8914 6142 8953
rect 6914 8946 6948 9000
rect 7032 9176 7066 9226
rect 7032 8984 7066 9000
rect 7150 9176 7184 9192
rect 7150 8946 7184 9000
rect 7269 8984 7303 9000
rect 7387 9376 7421 9392
rect 6914 8907 7184 8946
rect 7387 8949 7421 9000
rect 7505 9376 7539 9428
rect 7742 9428 8012 9467
rect 7505 8984 7539 9000
rect 7623 9376 7657 9392
rect 7623 8949 7657 9000
rect 7742 9376 7776 9428
rect 7742 8984 7776 9000
rect 7860 9376 7894 9392
rect 7860 8949 7894 9000
rect 7978 9376 8012 9428
rect 8214 9428 8484 9467
rect 7978 8984 8012 9000
rect 8096 9376 8130 9392
rect 8096 8949 8130 9000
rect 8214 9376 8248 9428
rect 8214 8984 8248 9000
rect 8332 9376 8366 9392
rect 8332 8949 8366 9000
rect 8450 9376 8484 9428
rect 8681 9429 8951 9468
rect 8450 8984 8484 9000
rect 8563 9376 8597 9392
rect 8563 8949 8597 9000
rect 8681 9376 8715 9429
rect 8681 8984 8715 9000
rect 8799 9376 8833 9392
rect 8799 8949 8833 9000
rect 8917 9376 8951 9429
rect 10413 9428 10683 9467
rect 10413 9376 10447 9428
rect 9122 9227 9392 9266
rect 8917 8984 8951 9000
rect 9004 9176 9038 9192
rect 7387 8910 8833 8949
rect 9004 8949 9038 9000
rect 9122 9176 9156 9227
rect 9122 8984 9156 9000
rect 9240 9176 9274 9192
rect 9240 8949 9274 9000
rect 9358 9176 9392 9227
rect 9358 8984 9392 9000
rect 9940 9226 10210 9263
rect 9940 9176 9974 9226
rect 9940 8984 9974 9000
rect 10058 9176 10092 9192
rect 9004 8910 9274 8949
rect 10058 8946 10092 9000
rect 10176 9176 10210 9226
rect 10176 8984 10210 9000
rect 10294 9176 10328 9192
rect 10294 8946 10328 9000
rect 10413 8984 10447 9000
rect 10531 9376 10565 9392
rect 10058 8907 10328 8946
rect 10531 8949 10565 9000
rect 10649 9376 10683 9428
rect 10886 9428 11156 9467
rect 10649 8984 10683 9000
rect 10767 9376 10801 9392
rect 10767 8949 10801 9000
rect 10886 9376 10920 9428
rect 10886 8984 10920 9000
rect 11004 9376 11038 9392
rect 11004 8949 11038 9000
rect 11122 9376 11156 9428
rect 11358 9428 11628 9467
rect 11122 8984 11156 9000
rect 11240 9376 11274 9392
rect 11240 8949 11274 9000
rect 11358 9376 11392 9428
rect 11358 8984 11392 9000
rect 11476 9376 11510 9392
rect 11476 8949 11510 9000
rect 11594 9376 11628 9428
rect 11825 9429 12095 9468
rect 11594 8984 11628 9000
rect 11707 9376 11741 9392
rect 11707 8949 11741 9000
rect 11825 9376 11859 9429
rect 11825 8984 11859 9000
rect 11943 9376 11977 9392
rect 11943 8949 11977 9000
rect 12061 9376 12095 9429
rect 13615 9432 13885 9471
rect 13615 9380 13649 9432
rect 12266 9227 12536 9266
rect 12061 8984 12095 9000
rect 12148 9176 12182 9192
rect 10531 8910 11977 8949
rect 12148 8949 12182 9000
rect 12266 9176 12300 9227
rect 12266 8984 12300 9000
rect 12384 9176 12418 9192
rect 12384 8949 12418 9000
rect 12502 9176 12536 9227
rect 12502 8984 12536 9000
rect 13142 9230 13412 9267
rect 13142 9180 13176 9230
rect 13142 8988 13176 9004
rect 13260 9180 13294 9196
rect 12148 8910 12418 8949
rect 13260 8950 13294 9004
rect 13378 9180 13412 9230
rect 13378 8988 13412 9004
rect 13496 9180 13530 9196
rect 13496 8950 13530 9004
rect 13615 8988 13649 9004
rect 13733 9380 13767 9396
rect 13260 8911 13530 8950
rect 13733 8953 13767 9004
rect 13851 9380 13885 9432
rect 14088 9432 14358 9471
rect 13851 8988 13885 9004
rect 13969 9380 14003 9396
rect 13969 8953 14003 9004
rect 14088 9380 14122 9432
rect 14088 8988 14122 9004
rect 14206 9380 14240 9396
rect 14206 8953 14240 9004
rect 14324 9380 14358 9432
rect 14560 9432 14830 9471
rect 14324 8988 14358 9004
rect 14442 9380 14476 9396
rect 14442 8953 14476 9004
rect 14560 9380 14594 9432
rect 14560 8988 14594 9004
rect 14678 9380 14712 9396
rect 14678 8953 14712 9004
rect 14796 9380 14830 9432
rect 15027 9433 15297 9472
rect 14796 8988 14830 9004
rect 14909 9380 14943 9396
rect 14909 8953 14943 9004
rect 15027 9380 15061 9433
rect 15027 8988 15061 9004
rect 15145 9380 15179 9396
rect 15145 8953 15179 9004
rect 15263 9380 15297 9433
rect 16759 9432 17029 9471
rect 16759 9380 16793 9432
rect 15468 9231 15738 9270
rect 15263 8988 15297 9004
rect 15350 9180 15384 9196
rect 13733 8914 15179 8953
rect 15350 8953 15384 9004
rect 15468 9180 15502 9231
rect 15468 8988 15502 9004
rect 15586 9180 15620 9196
rect 15586 8953 15620 9004
rect 15704 9180 15738 9231
rect 15704 8988 15738 9004
rect 16286 9230 16556 9267
rect 16286 9180 16320 9230
rect 16286 8988 16320 9004
rect 16404 9180 16438 9196
rect 15350 8914 15620 8953
rect 16404 8950 16438 9004
rect 16522 9180 16556 9230
rect 16522 8988 16556 9004
rect 16640 9180 16674 9196
rect 16640 8950 16674 9004
rect 16759 8988 16793 9004
rect 16877 9380 16911 9396
rect 16404 8911 16674 8950
rect 16877 8953 16911 9004
rect 16995 9380 17029 9432
rect 17232 9432 17502 9471
rect 16995 8988 17029 9004
rect 17113 9380 17147 9396
rect 17113 8953 17147 9004
rect 17232 9380 17266 9432
rect 17232 8988 17266 9004
rect 17350 9380 17384 9396
rect 17350 8953 17384 9004
rect 17468 9380 17502 9432
rect 17704 9432 17974 9471
rect 17468 8988 17502 9004
rect 17586 9380 17620 9396
rect 17586 8953 17620 9004
rect 17704 9380 17738 9432
rect 17704 8988 17738 9004
rect 17822 9380 17856 9396
rect 17822 8953 17856 9004
rect 17940 9380 17974 9432
rect 18171 9433 18441 9472
rect 17940 8988 17974 9004
rect 18053 9380 18087 9396
rect 18053 8953 18087 9004
rect 18171 9380 18205 9433
rect 18171 8988 18205 9004
rect 18289 9380 18323 9396
rect 18289 8953 18323 9004
rect 18407 9380 18441 9433
rect 19891 9428 20161 9467
rect 19891 9376 19925 9428
rect 18612 9231 18882 9270
rect 18407 8988 18441 9004
rect 18494 9180 18528 9196
rect 16877 8914 18323 8953
rect 18494 8953 18528 9004
rect 18612 9180 18646 9231
rect 18612 8988 18646 9004
rect 18730 9180 18764 9196
rect 18730 8953 18764 9004
rect 18848 9180 18882 9231
rect 18848 8988 18882 9004
rect 19418 9226 19688 9263
rect 19418 9176 19452 9226
rect 19418 8984 19452 9000
rect 19536 9176 19570 9192
rect 18494 8914 18764 8953
rect 19536 8946 19570 9000
rect 19654 9176 19688 9226
rect 19654 8984 19688 9000
rect 19772 9176 19806 9192
rect 19772 8946 19806 9000
rect 19891 8984 19925 9000
rect 20009 9376 20043 9392
rect 19536 8907 19806 8946
rect 20009 8949 20043 9000
rect 20127 9376 20161 9428
rect 20364 9428 20634 9467
rect 20127 8984 20161 9000
rect 20245 9376 20279 9392
rect 20245 8949 20279 9000
rect 20364 9376 20398 9428
rect 20364 8984 20398 9000
rect 20482 9376 20516 9392
rect 20482 8949 20516 9000
rect 20600 9376 20634 9428
rect 20836 9428 21106 9467
rect 20600 8984 20634 9000
rect 20718 9376 20752 9392
rect 20718 8949 20752 9000
rect 20836 9376 20870 9428
rect 20836 8984 20870 9000
rect 20954 9376 20988 9392
rect 20954 8949 20988 9000
rect 21072 9376 21106 9428
rect 21303 9429 21573 9468
rect 21072 8984 21106 9000
rect 21185 9376 21219 9392
rect 21185 8949 21219 9000
rect 21303 9376 21337 9429
rect 21303 8984 21337 9000
rect 21421 9376 21455 9392
rect 21421 8949 21455 9000
rect 21539 9376 21573 9429
rect 23035 9428 23305 9467
rect 23035 9376 23069 9428
rect 21744 9227 22014 9266
rect 21539 8984 21573 9000
rect 21626 9176 21660 9192
rect 20009 8910 21455 8949
rect 21626 8949 21660 9000
rect 21744 9176 21778 9227
rect 21744 8984 21778 9000
rect 21862 9176 21896 9192
rect 21862 8949 21896 9000
rect 21980 9176 22014 9227
rect 21980 8984 22014 9000
rect 22562 9226 22832 9263
rect 22562 9176 22596 9226
rect 22562 8984 22596 9000
rect 22680 9176 22714 9192
rect 21626 8910 21896 8949
rect 22680 8946 22714 9000
rect 22798 9176 22832 9226
rect 22798 8984 22832 9000
rect 22916 9176 22950 9192
rect 22916 8946 22950 9000
rect 23035 8984 23069 9000
rect 23153 9376 23187 9392
rect 22680 8907 22950 8946
rect 23153 8949 23187 9000
rect 23271 9376 23305 9428
rect 23508 9428 23778 9467
rect 23271 8984 23305 9000
rect 23389 9376 23423 9392
rect 23389 8949 23423 9000
rect 23508 9376 23542 9428
rect 23508 8984 23542 9000
rect 23626 9376 23660 9392
rect 23626 8949 23660 9000
rect 23744 9376 23778 9428
rect 23980 9428 24250 9467
rect 23744 8984 23778 9000
rect 23862 9376 23896 9392
rect 23862 8949 23896 9000
rect 23980 9376 24014 9428
rect 23980 8984 24014 9000
rect 24098 9376 24132 9392
rect 24098 8949 24132 9000
rect 24216 9376 24250 9428
rect 24447 9429 24717 9468
rect 31091 9461 31132 10047
rect 31205 9995 31271 10012
rect 31205 9961 31221 9995
rect 31255 9961 31271 9995
rect 31205 9945 31271 9961
rect 31273 9671 31289 9705
rect 31323 9671 31339 9705
rect 31373 9643 31389 9677
rect 31565 9643 31581 9677
rect 31373 9525 31389 9559
rect 31565 9525 31581 9559
rect 24216 8984 24250 9000
rect 24329 9376 24363 9392
rect 24329 8949 24363 9000
rect 24447 9376 24481 9429
rect 24447 8984 24481 9000
rect 24565 9376 24599 9392
rect 24565 8949 24599 9000
rect 24683 9376 24717 9429
rect 30148 9391 30164 9425
rect 30340 9391 30356 9425
rect 24888 9227 25158 9266
rect 24683 8984 24717 9000
rect 24770 9176 24804 9192
rect 23153 8910 24599 8949
rect 24770 8949 24804 9000
rect 24888 9176 24922 9227
rect 24888 8984 24922 9000
rect 25006 9176 25040 9192
rect 25006 8949 25040 9000
rect 25124 9176 25158 9227
rect 25124 8984 25158 9000
rect 30077 8997 30166 9031
rect 30342 8997 30358 9031
rect 24770 8910 25040 8949
rect 670 8796 686 8830
rect 720 8796 736 8830
rect 1996 8789 2030 8805
rect 3814 8796 3830 8830
rect 3864 8796 3880 8830
rect 1996 8739 2030 8755
rect 5140 8789 5174 8805
rect 6946 8792 6962 8826
rect 6996 8792 7012 8826
rect 5140 8739 5174 8755
rect 8272 8785 8306 8801
rect 10090 8792 10106 8826
rect 10140 8792 10156 8826
rect 8272 8735 8306 8751
rect 11416 8785 11450 8801
rect 13292 8796 13308 8830
rect 13342 8796 13358 8830
rect 11416 8735 11450 8751
rect 14618 8789 14652 8805
rect 16436 8796 16452 8830
rect 16486 8796 16502 8830
rect 14618 8739 14652 8755
rect 17762 8789 17796 8805
rect 19568 8792 19584 8826
rect 19618 8792 19634 8826
rect 17762 8739 17796 8755
rect 20894 8785 20928 8801
rect 22712 8792 22728 8826
rect 22762 8792 22778 8826
rect 20894 8735 20928 8751
rect 24038 8785 24072 8801
rect 30077 8795 30112 8997
rect 30150 8879 30166 8913
rect 30342 8879 30358 8913
rect 31375 8872 31391 8906
rect 31567 8872 31583 8906
rect 30077 8761 30166 8795
rect 30342 8761 30358 8795
rect 24038 8735 24072 8751
rect 31274 8725 31290 8759
rect 31324 8725 31340 8759
rect 31375 8754 31391 8788
rect 31567 8754 31583 8788
rect 1850 8690 1942 8703
rect 1850 8635 1866 8690
rect 1926 8635 1942 8690
rect 1850 8618 1942 8635
rect 2935 8689 3027 8706
rect 2935 8634 2951 8689
rect 3011 8634 3027 8689
rect 2935 8621 3027 8634
rect 3202 8690 3259 8694
rect 3202 8630 3206 8690
rect 3255 8630 3259 8690
rect 3202 8626 3259 8630
rect 4994 8690 5086 8703
rect 4994 8635 5010 8690
rect 5070 8635 5086 8690
rect 4994 8618 5086 8635
rect 6079 8689 6171 8706
rect 6079 8634 6095 8689
rect 6155 8634 6171 8689
rect 6079 8621 6171 8634
rect 6346 8690 6403 8694
rect 6346 8630 6350 8690
rect 6399 8630 6403 8690
rect 6346 8626 6403 8630
rect 8126 8686 8218 8699
rect 8126 8631 8142 8686
rect 8202 8631 8218 8686
rect 8126 8614 8218 8631
rect 9211 8685 9303 8702
rect 9211 8630 9227 8685
rect 9287 8630 9303 8685
rect 9211 8617 9303 8630
rect 9478 8686 9535 8690
rect 9478 8626 9482 8686
rect 9531 8626 9535 8686
rect 9478 8622 9535 8626
rect 11270 8686 11362 8699
rect 11270 8631 11286 8686
rect 11346 8631 11362 8686
rect 11270 8614 11362 8631
rect 12355 8685 12447 8702
rect 14472 8690 14564 8703
rect 12355 8630 12371 8685
rect 12431 8630 12447 8685
rect 12355 8617 12447 8630
rect 12622 8686 12679 8690
rect 12622 8626 12626 8686
rect 12675 8626 12679 8686
rect 12622 8622 12679 8626
rect 14472 8635 14488 8690
rect 14548 8635 14564 8690
rect 14472 8618 14564 8635
rect 15557 8689 15649 8706
rect 15557 8634 15573 8689
rect 15633 8634 15649 8689
rect 15557 8621 15649 8634
rect 15824 8690 15881 8694
rect 15824 8630 15828 8690
rect 15877 8630 15881 8690
rect 15824 8626 15881 8630
rect 17616 8690 17708 8703
rect 17616 8635 17632 8690
rect 17692 8635 17708 8690
rect 17616 8618 17708 8635
rect 18701 8689 18793 8706
rect 18701 8634 18717 8689
rect 18777 8634 18793 8689
rect 18701 8621 18793 8634
rect 18968 8690 19025 8694
rect 18968 8630 18972 8690
rect 19021 8630 19025 8690
rect 18968 8626 19025 8630
rect 20748 8686 20840 8699
rect 20748 8631 20764 8686
rect 20824 8631 20840 8686
rect 20748 8614 20840 8631
rect 21833 8685 21925 8702
rect 21833 8630 21849 8685
rect 21909 8630 21925 8685
rect 21833 8617 21925 8630
rect 22100 8686 22157 8690
rect 22100 8626 22104 8686
rect 22153 8626 22157 8686
rect 22100 8622 22157 8626
rect 23892 8686 23984 8699
rect 23892 8631 23908 8686
rect 23968 8631 23984 8686
rect 23892 8614 23984 8631
rect 24977 8685 25069 8702
rect 24977 8630 24993 8685
rect 25053 8630 25069 8685
rect 24977 8617 25069 8630
rect 25244 8686 25301 8690
rect 25244 8626 25248 8686
rect 25297 8626 25301 8686
rect 30150 8643 30166 8677
rect 30342 8643 30358 8677
rect 25244 8622 25301 8626
rect 1642 8559 1676 8575
rect 1642 8509 1676 8525
rect 3202 8574 3259 8578
rect 6346 8576 6403 8578
rect 3202 8514 3206 8574
rect 3255 8514 3479 8574
rect 3202 8510 3479 8514
rect 1968 8405 2060 8418
rect 1968 8350 1984 8405
rect 2044 8350 2060 8405
rect 1968 8333 2060 8350
rect 3202 8406 3259 8410
rect 3202 8346 3206 8406
rect 3255 8346 3259 8406
rect 3202 8342 3259 8346
rect 1761 8169 1795 8185
rect 1761 8119 1795 8135
rect 1388 8047 1422 8063
rect 1388 7855 1422 7871
rect 1506 8059 1540 8063
rect 1584 8059 1618 8063
rect 1506 8047 1618 8059
rect 1540 7871 1584 8047
rect 1506 7859 1584 7871
rect 1506 7855 1540 7859
rect 1584 7655 1618 7671
rect 1702 8047 1736 8063
rect 1702 7655 1736 7671
rect 1820 8047 1854 8063
rect 1820 7655 1854 7671
rect 1938 8047 1972 8063
rect 1938 7655 1972 7671
rect 2056 8059 2090 8063
rect 2130 8059 2164 8063
rect 2056 8047 2164 8059
rect 2090 7871 2130 8047
rect 2090 7859 2164 7871
rect 2130 7855 2164 7859
rect 2248 8047 2282 8063
rect 2248 7855 2282 7871
rect 2056 7655 2090 7671
rect 1803 7536 1819 7570
rect 1853 7536 1869 7570
rect 1752 7418 1888 7422
rect 1752 7404 1792 7418
rect 1850 7404 1888 7418
rect 1752 7358 1768 7404
rect 1872 7358 1888 7404
rect 1752 7336 1888 7358
rect 3415 6954 3479 8510
rect 4786 8559 4820 8575
rect 4786 8509 4820 8525
rect 6346 8574 6619 8576
rect 15824 8575 15881 8578
rect 18968 8576 19025 8578
rect 6346 8514 6350 8574
rect 6399 8514 6619 8574
rect 9478 8573 9535 8574
rect 6346 8512 6619 8514
rect 6346 8510 6403 8512
rect 5112 8405 5204 8418
rect 5112 8350 5128 8405
rect 5188 8350 5204 8405
rect 5112 8333 5204 8350
rect 6346 8406 6403 8410
rect 6346 8346 6350 8406
rect 6399 8346 6403 8406
rect 6346 8342 6403 8346
rect 4905 8169 4939 8185
rect 4905 8119 4939 8135
rect 4532 8047 4566 8063
rect 4532 7855 4566 7871
rect 4650 8059 4684 8063
rect 4728 8059 4762 8063
rect 4650 8047 4762 8059
rect 4684 7871 4728 8047
rect 4650 7859 4728 7871
rect 4650 7855 4684 7859
rect 4728 7655 4762 7671
rect 4846 8047 4880 8063
rect 4846 7655 4880 7671
rect 4964 8047 4998 8063
rect 4964 7655 4998 7671
rect 5082 8047 5116 8063
rect 5082 7655 5116 7671
rect 5200 8059 5234 8063
rect 5274 8059 5308 8063
rect 5200 8047 5308 8059
rect 5234 7871 5274 8047
rect 5234 7859 5308 7871
rect 5274 7855 5308 7859
rect 5392 8047 5426 8063
rect 5392 7855 5426 7871
rect 5200 7655 5234 7671
rect 4947 7536 4963 7570
rect 4997 7536 5013 7570
rect 4896 7418 5032 7422
rect 4896 7404 4936 7418
rect 4994 7404 5032 7418
rect 4896 7358 4912 7404
rect 5016 7358 5032 7404
rect 4896 7336 5032 7358
rect 6555 7052 6619 8512
rect 7918 8555 7952 8571
rect 7918 8505 7952 8521
rect 9478 8570 9761 8573
rect 12622 8572 12679 8574
rect 9478 8510 9482 8570
rect 9531 8510 9761 8570
rect 9478 8509 9761 8510
rect 9478 8506 9535 8509
rect 8244 8401 8336 8414
rect 8244 8346 8260 8401
rect 8320 8346 8336 8401
rect 8244 8329 8336 8346
rect 9478 8402 9535 8406
rect 9478 8342 9482 8402
rect 9531 8342 9535 8402
rect 9478 8338 9535 8342
rect 8037 8165 8071 8181
rect 8037 8115 8071 8131
rect 7664 8043 7698 8059
rect 7664 7851 7698 7867
rect 7782 8055 7816 8059
rect 7860 8055 7894 8059
rect 7782 8043 7894 8055
rect 7816 7867 7860 8043
rect 7782 7855 7860 7867
rect 7782 7851 7816 7855
rect 7860 7651 7894 7667
rect 7978 8043 8012 8059
rect 7978 7651 8012 7667
rect 8096 8043 8130 8059
rect 8096 7651 8130 7667
rect 8214 8043 8248 8059
rect 8214 7651 8248 7667
rect 8332 8055 8366 8059
rect 8406 8055 8440 8059
rect 8332 8043 8440 8055
rect 8366 7867 8406 8043
rect 8366 7855 8440 7867
rect 8406 7851 8440 7855
rect 8524 8043 8558 8059
rect 8524 7851 8558 7867
rect 8332 7651 8366 7667
rect 8079 7532 8095 7566
rect 8129 7532 8145 7566
rect 8028 7414 8164 7418
rect 8028 7400 8068 7414
rect 8126 7400 8164 7414
rect 8028 7354 8044 7400
rect 8148 7354 8164 7400
rect 8028 7332 8164 7354
rect 9697 7175 9761 8509
rect 11062 8555 11096 8571
rect 11062 8505 11096 8521
rect 12621 8570 12923 8572
rect 12621 8510 12626 8570
rect 12675 8510 12923 8570
rect 12621 8508 12923 8510
rect 14264 8559 14298 8575
rect 14264 8509 14298 8525
rect 15824 8574 16097 8575
rect 15824 8514 15828 8574
rect 15877 8514 16097 8574
rect 15824 8511 16097 8514
rect 15824 8510 15881 8511
rect 12622 8506 12679 8508
rect 11388 8401 11480 8414
rect 11388 8346 11404 8401
rect 11464 8346 11480 8401
rect 11388 8329 11480 8346
rect 12622 8402 12679 8406
rect 12622 8342 12626 8402
rect 12675 8342 12679 8402
rect 12622 8338 12679 8342
rect 11181 8165 11215 8181
rect 11181 8115 11215 8131
rect 10808 8043 10842 8059
rect 10808 7851 10842 7867
rect 10926 8055 10960 8059
rect 11004 8055 11038 8059
rect 10926 8043 11038 8055
rect 10960 7867 11004 8043
rect 10926 7855 11004 7867
rect 10926 7851 10960 7855
rect 11004 7651 11038 7667
rect 11122 8043 11156 8059
rect 11122 7651 11156 7667
rect 11240 8043 11274 8059
rect 11240 7651 11274 7667
rect 11358 8043 11392 8059
rect 11358 7651 11392 7667
rect 11476 8055 11510 8059
rect 11550 8055 11584 8059
rect 11476 8043 11584 8055
rect 11510 7867 11550 8043
rect 11510 7855 11584 7867
rect 11550 7851 11584 7855
rect 11668 8043 11702 8059
rect 11668 7851 11702 7867
rect 11476 7651 11510 7667
rect 11223 7532 11239 7566
rect 11273 7532 11289 7566
rect 11172 7414 11308 7418
rect 11172 7400 11212 7414
rect 11270 7400 11308 7414
rect 11172 7354 11188 7400
rect 11292 7354 11308 7400
rect 11172 7332 11308 7354
rect 12859 7273 12923 8508
rect 14590 8405 14682 8418
rect 14590 8350 14606 8405
rect 14666 8350 14682 8405
rect 14590 8333 14682 8350
rect 15824 8406 15881 8410
rect 15824 8346 15828 8406
rect 15877 8346 15881 8406
rect 15824 8342 15881 8346
rect 14383 8169 14417 8185
rect 14383 8119 14417 8135
rect 14010 8047 14044 8063
rect 14010 7855 14044 7871
rect 14128 8059 14162 8063
rect 14206 8059 14240 8063
rect 14128 8047 14240 8059
rect 14162 7871 14206 8047
rect 14128 7859 14206 7871
rect 14128 7855 14162 7859
rect 14206 7655 14240 7671
rect 14324 8047 14358 8063
rect 14324 7655 14358 7671
rect 14442 8047 14476 8063
rect 14442 7655 14476 7671
rect 14560 8047 14594 8063
rect 14560 7655 14594 7671
rect 14678 8059 14712 8063
rect 14752 8059 14786 8063
rect 14678 8047 14786 8059
rect 14712 7871 14752 8047
rect 14712 7859 14786 7871
rect 14752 7855 14786 7859
rect 14870 8047 14904 8063
rect 14870 7855 14904 7871
rect 14678 7655 14712 7671
rect 14425 7536 14441 7570
rect 14475 7536 14491 7570
rect 14374 7418 14510 7422
rect 14374 7404 14414 7418
rect 14472 7404 14510 7418
rect 14374 7358 14390 7404
rect 14494 7358 14510 7404
rect 14374 7336 14510 7358
rect 12859 7209 15337 7273
rect 9697 7111 13260 7175
rect 6555 6988 11182 7052
rect 3415 6890 9131 6954
rect 3213 6751 3427 6755
rect 3213 6689 3253 6751
rect 3393 6689 3427 6751
rect 3213 6671 3427 6689
rect 3951 6751 4165 6755
rect 3951 6689 3991 6751
rect 4131 6689 4165 6751
rect 3951 6671 4165 6689
rect 4689 6751 4903 6755
rect 4689 6689 4729 6751
rect 4869 6689 4903 6751
rect 4689 6671 4903 6689
rect 5427 6751 5641 6755
rect 5427 6689 5467 6751
rect 5607 6689 5641 6751
rect 5427 6671 5641 6689
rect 6167 6751 6381 6755
rect 6167 6689 6207 6751
rect 6347 6689 6381 6751
rect 6167 6671 6381 6689
rect 6909 6751 7123 6755
rect 6909 6689 6949 6751
rect 7089 6689 7123 6751
rect 6909 6671 7123 6689
rect 7647 6751 7861 6755
rect 7647 6689 7687 6751
rect 7827 6689 7861 6751
rect 7647 6671 7861 6689
rect 8385 6753 8599 6757
rect 8385 6691 8425 6753
rect 8565 6691 8599 6753
rect 8385 6673 8599 6691
rect 3129 6601 3399 6635
rect 3129 6545 3163 6601
rect 3129 6353 3163 6369
rect 3247 6545 3281 6561
rect 3247 6353 3281 6369
rect 3365 6545 3399 6601
rect 3867 6601 4137 6635
rect 3365 6353 3399 6369
rect 3483 6545 3517 6561
rect 3483 6353 3517 6369
rect 3867 6545 3901 6601
rect 3867 6353 3901 6369
rect 3985 6545 4019 6561
rect 3985 6353 4019 6369
rect 4103 6545 4137 6601
rect 4605 6601 4875 6635
rect 4103 6353 4137 6369
rect 4221 6545 4255 6561
rect 4221 6353 4255 6369
rect 4605 6545 4639 6601
rect 4605 6353 4639 6369
rect 4723 6545 4757 6561
rect 4723 6353 4757 6369
rect 4841 6545 4875 6601
rect 5343 6601 5613 6635
rect 4841 6353 4875 6369
rect 4959 6545 4993 6561
rect 4959 6353 4993 6369
rect 5343 6545 5377 6601
rect 5343 6353 5377 6369
rect 5461 6545 5495 6561
rect 5461 6353 5495 6369
rect 5579 6545 5613 6601
rect 6083 6601 6353 6635
rect 5579 6353 5613 6369
rect 5697 6545 5731 6561
rect 5697 6353 5731 6369
rect 6083 6545 6117 6601
rect 6083 6353 6117 6369
rect 6201 6545 6235 6561
rect 6201 6353 6235 6369
rect 6319 6545 6353 6601
rect 6825 6601 7095 6635
rect 6319 6353 6353 6369
rect 6437 6545 6471 6561
rect 6437 6353 6471 6369
rect 6825 6547 6859 6601
rect 6825 6355 6859 6371
rect 6943 6547 6977 6563
rect 6943 6355 6977 6371
rect 7061 6547 7095 6601
rect 7563 6601 7833 6635
rect 7061 6355 7095 6371
rect 7179 6547 7213 6563
rect 7179 6355 7213 6371
rect 7563 6551 7597 6601
rect 7563 6359 7597 6375
rect 7681 6551 7715 6567
rect 7681 6359 7715 6375
rect 7799 6551 7833 6601
rect 8301 6603 8571 6637
rect 7799 6359 7833 6375
rect 7917 6551 7951 6567
rect 7917 6359 7951 6375
rect 8301 6547 8335 6603
rect 8301 6355 8335 6371
rect 8419 6547 8453 6563
rect 8419 6355 8453 6371
rect 8537 6547 8571 6603
rect 8537 6355 8571 6371
rect 8655 6547 8689 6563
rect 8655 6355 8689 6371
rect 3291 6229 3307 6263
rect 3341 6229 3357 6263
rect 3525 6223 3641 6269
rect 4029 6229 4045 6263
rect 4079 6229 4095 6263
rect 4262 6223 4399 6269
rect 4767 6229 4783 6263
rect 4817 6229 5189 6263
rect 5505 6229 5521 6263
rect 5555 6229 5887 6263
rect 6245 6229 6261 6263
rect 6295 6229 6710 6263
rect 6987 6229 7003 6263
rect 7037 6229 7439 6263
rect 7725 6229 7741 6263
rect 7775 6229 8159 6263
rect 8463 6231 8479 6265
rect 8513 6231 8759 6265
rect 4810 6228 5189 6229
rect 3247 6163 3281 6179
rect 3247 5971 3281 5987
rect 3365 6163 3399 6179
rect 3365 5971 3399 5987
rect 3295 5871 3479 5891
rect 3295 5801 3315 5871
rect 3459 5801 3479 5871
rect 3295 5795 3479 5801
rect 3577 4004 3641 6223
rect 3985 6163 4019 6179
rect 3985 5971 4019 5987
rect 4103 6163 4137 6179
rect 4103 5971 4137 5987
rect 4033 5871 4217 5891
rect 4033 5801 4053 5871
rect 4197 5801 4217 5871
rect 4033 5795 4217 5801
rect -2012 3398 235 3421
rect -2012 3361 -1976 3398
rect -1883 3361 151 3398
rect -2012 3354 151 3361
rect 205 3354 235 3398
rect -2012 3334 235 3354
rect 3577 3404 3642 4004
rect 4334 3502 4398 6223
rect 4723 6159 4757 6175
rect 4723 5967 4757 5983
rect 4841 6159 4875 6175
rect 4841 5967 4875 5983
rect 4771 5871 4955 5891
rect 4771 5801 4791 5871
rect 4935 5801 4955 5871
rect 4771 5795 4955 5801
rect 5125 3643 5189 6228
rect 5461 6159 5495 6175
rect 5461 5967 5495 5983
rect 5579 6159 5613 6175
rect 5579 5967 5613 5983
rect 5509 5871 5693 5891
rect 5509 5801 5529 5871
rect 5673 5801 5693 5871
rect 5509 5795 5693 5801
rect 5823 3741 5887 6229
rect 6201 6159 6235 6175
rect 6201 5967 6235 5983
rect 6319 6159 6353 6175
rect 6319 5967 6353 5983
rect 6249 5871 6433 5891
rect 6249 5801 6269 5871
rect 6413 5801 6433 5871
rect 6249 5795 6433 5801
rect 6646 3849 6710 6229
rect 6943 6159 6977 6175
rect 6943 5967 6977 5983
rect 7061 6159 7095 6175
rect 7061 5967 7095 5983
rect 6991 5871 7175 5891
rect 6991 5801 7011 5871
rect 7155 5801 7175 5871
rect 6991 5795 7175 5801
rect 7375 3947 7439 6229
rect 7681 6163 7715 6179
rect 7681 5971 7715 5987
rect 7799 6163 7833 6179
rect 7799 5971 7833 5987
rect 7729 5871 7913 5891
rect 7729 5801 7749 5871
rect 7893 5801 7913 5871
rect 7729 5795 7913 5801
rect 8095 4056 8159 6229
rect 8419 6161 8453 6177
rect 8419 5969 8453 5985
rect 8537 6161 8571 6177
rect 8537 5969 8571 5985
rect 8467 5873 8651 5893
rect 8467 5803 8487 5873
rect 8631 5803 8651 5873
rect 8467 5797 8651 5803
rect 8695 4154 8759 6231
rect 9067 5308 9131 6890
rect 9989 6706 10191 6726
rect 9989 6662 10035 6706
rect 10157 6662 10191 6706
rect 9989 6652 10067 6662
rect 10105 6652 10191 6662
rect 9989 6634 10191 6652
rect 9834 6488 10104 6523
rect 9716 6435 9750 6451
rect 9233 6235 9267 6251
rect 9233 6043 9267 6059
rect 9351 6235 9385 6251
rect 9351 6043 9385 6059
rect 9469 6235 9503 6251
rect 9469 6043 9503 6059
rect 9587 6235 9621 6251
rect 9587 6043 9621 6059
rect 9716 6043 9750 6059
rect 9834 6435 9868 6488
rect 9834 6043 9868 6059
rect 9952 6435 9986 6451
rect 9952 6043 9986 6059
rect 10070 6435 10104 6488
rect 10070 6043 10104 6059
rect 10188 6435 10222 6451
rect 10188 6043 10222 6059
rect 10306 6435 10340 6451
rect 10306 6043 10340 6059
rect 10424 6435 10458 6451
rect 10672 6289 10942 6324
rect 10424 6043 10458 6059
rect 10554 6235 10588 6251
rect 10554 6043 10588 6059
rect 10672 6235 10706 6289
rect 10672 6043 10706 6059
rect 10790 6235 10824 6251
rect 10790 6043 10824 6059
rect 10908 6235 10942 6289
rect 10908 6043 10942 6059
rect 9475 5846 9481 5880
rect 9535 5846 9541 5880
rect 9773 5742 9807 5758
rect 9891 5742 9925 5758
rect 9773 5350 9807 5366
rect 9889 5366 9891 5412
rect 9067 5267 9201 5308
rect 9889 5308 9925 5366
rect 10009 5742 10043 5758
rect 10009 5350 10043 5366
rect 10127 5742 10161 5758
rect 10245 5742 10279 5758
rect 10161 5366 10163 5413
rect 10127 5308 10163 5366
rect 10363 5742 10397 5758
rect 10245 5350 10279 5366
rect 10362 5366 10363 5413
rect 10481 5742 10515 5758
rect 10397 5366 10398 5413
rect 10362 5308 10398 5366
rect 10869 5631 10935 5640
rect 10481 5350 10515 5366
rect 9303 5268 10398 5308
rect 11118 5306 11182 6988
rect 12057 6704 12259 6724
rect 12057 6660 12103 6704
rect 12225 6660 12259 6704
rect 12057 6650 12135 6660
rect 12173 6650 12259 6660
rect 12057 6632 12259 6650
rect 11902 6486 12172 6521
rect 11784 6433 11818 6449
rect 11301 6233 11335 6249
rect 11301 6041 11335 6057
rect 11419 6233 11453 6249
rect 11419 6041 11453 6057
rect 11537 6233 11571 6249
rect 11537 6041 11571 6057
rect 11655 6233 11689 6249
rect 11655 6041 11689 6057
rect 11784 6041 11818 6057
rect 11902 6433 11936 6486
rect 11902 6041 11936 6057
rect 12020 6433 12054 6449
rect 12020 6041 12054 6057
rect 12138 6433 12172 6486
rect 12138 6041 12172 6057
rect 12256 6433 12290 6449
rect 12256 6041 12290 6057
rect 12374 6433 12408 6449
rect 12374 6041 12408 6057
rect 12492 6433 12526 6449
rect 12740 6287 13010 6322
rect 12492 6041 12526 6057
rect 12622 6233 12656 6249
rect 12622 6041 12656 6057
rect 12740 6233 12774 6287
rect 12740 6041 12774 6057
rect 12858 6233 12892 6249
rect 12858 6041 12892 6057
rect 12976 6233 13010 6287
rect 12976 6041 13010 6057
rect 11543 5844 11549 5878
rect 11603 5844 11609 5878
rect 11841 5740 11875 5756
rect 11959 5740 11993 5756
rect 11841 5348 11875 5364
rect 11957 5364 11959 5410
rect 9303 5267 10379 5268
rect 9787 5178 9854 5194
rect 9787 5144 9803 5178
rect 9837 5144 9854 5178
rect 9787 5128 9854 5144
rect 9513 5110 9547 5126
rect 9513 5060 9547 5076
rect 10051 5061 10067 5095
rect 10101 5061 10117 5095
rect 10169 5060 10185 5094
rect 10219 5060 10235 5094
rect 10290 5026 10324 5267
rect 11118 5265 11269 5306
rect 11957 5306 11993 5364
rect 12077 5740 12111 5756
rect 12077 5348 12111 5364
rect 12195 5740 12229 5756
rect 12313 5740 12347 5756
rect 12229 5364 12231 5411
rect 12195 5306 12231 5364
rect 12431 5740 12465 5756
rect 12313 5348 12347 5364
rect 12430 5364 12431 5411
rect 12549 5740 12583 5756
rect 12465 5364 12466 5411
rect 12430 5306 12466 5364
rect 12549 5348 12583 5364
rect 11371 5266 12466 5306
rect 13196 5308 13260 7111
rect 14126 6706 14328 6726
rect 14126 6662 14172 6706
rect 14294 6662 14328 6706
rect 14126 6652 14204 6662
rect 14242 6652 14328 6662
rect 14126 6634 14328 6652
rect 13971 6488 14241 6523
rect 13853 6435 13887 6451
rect 13370 6235 13404 6251
rect 13370 6043 13404 6059
rect 13488 6235 13522 6251
rect 13488 6043 13522 6059
rect 13606 6235 13640 6251
rect 13606 6043 13640 6059
rect 13724 6235 13758 6251
rect 13724 6043 13758 6059
rect 13853 6043 13887 6059
rect 13971 6435 14005 6488
rect 13971 6043 14005 6059
rect 14089 6435 14123 6451
rect 14089 6043 14123 6059
rect 14207 6435 14241 6488
rect 14207 6043 14241 6059
rect 14325 6435 14359 6451
rect 14325 6043 14359 6059
rect 14443 6435 14477 6451
rect 14443 6043 14477 6059
rect 14561 6435 14595 6451
rect 14809 6289 15079 6324
rect 14561 6043 14595 6059
rect 14691 6235 14725 6251
rect 14691 6043 14725 6059
rect 14809 6235 14843 6289
rect 14809 6043 14843 6059
rect 14927 6235 14961 6251
rect 14927 6043 14961 6059
rect 15045 6235 15079 6289
rect 15045 6043 15079 6059
rect 13612 5846 13618 5880
rect 13672 5846 13678 5880
rect 13910 5742 13944 5758
rect 14028 5742 14062 5758
rect 13910 5350 13944 5366
rect 14026 5366 14028 5412
rect 13196 5267 13338 5308
rect 11371 5265 12447 5266
rect 10434 5178 10501 5194
rect 10434 5144 10451 5178
rect 10485 5144 10501 5178
rect 10434 5128 10501 5144
rect 11855 5176 11922 5192
rect 11855 5142 11871 5176
rect 11905 5142 11922 5176
rect 10636 5111 10670 5127
rect 11855 5126 11922 5142
rect 10636 5061 10670 5077
rect 11581 5108 11615 5124
rect 11581 5058 11615 5074
rect 12119 5059 12135 5093
rect 12169 5059 12185 5093
rect 12237 5058 12253 5092
rect 12287 5058 12303 5092
rect 9367 5010 9401 5026
rect 9367 4818 9401 4834
rect 9485 5010 9519 5026
rect 9485 4818 9519 4834
rect 9891 5010 9925 5026
rect 10009 5010 10043 5026
rect 9891 4567 9926 4634
rect 10009 4618 10043 4634
rect 10127 5010 10161 5026
rect 10127 4618 10161 4634
rect 10245 5010 10324 5026
rect 10279 4980 10324 5010
rect 10363 5010 10397 5026
rect 10665 5010 10699 5026
rect 10665 4818 10699 4834
rect 10783 5010 10817 5026
rect 12358 5024 12392 5265
rect 14026 5308 14062 5366
rect 14146 5742 14180 5758
rect 14146 5350 14180 5366
rect 14264 5742 14298 5758
rect 14382 5742 14416 5758
rect 14298 5366 14300 5413
rect 14264 5308 14300 5366
rect 14500 5742 14534 5758
rect 14382 5350 14416 5366
rect 14499 5366 14500 5413
rect 14618 5742 14652 5758
rect 14534 5366 14535 5413
rect 14499 5308 14535 5366
rect 14618 5350 14652 5366
rect 13440 5268 14535 5308
rect 15273 5306 15337 7209
rect 16033 7246 16097 8511
rect 17408 8559 17442 8575
rect 17408 8509 17442 8525
rect 18968 8574 19223 8576
rect 18968 8514 18972 8574
rect 19021 8514 19223 8574
rect 22100 8572 22157 8574
rect 18968 8512 19223 8514
rect 18968 8510 19025 8512
rect 17734 8405 17826 8418
rect 17734 8350 17750 8405
rect 17810 8350 17826 8405
rect 17734 8333 17826 8350
rect 18968 8406 19025 8410
rect 18968 8346 18972 8406
rect 19021 8346 19025 8406
rect 18968 8342 19025 8346
rect 17527 8169 17561 8185
rect 17527 8119 17561 8135
rect 19159 8072 19223 8512
rect 20540 8555 20574 8571
rect 20540 8505 20574 8521
rect 22100 8570 22353 8572
rect 22100 8510 22104 8570
rect 22153 8510 22353 8570
rect 22100 8508 22353 8510
rect 22100 8506 22157 8508
rect 20866 8401 20958 8414
rect 20866 8346 20882 8401
rect 20942 8346 20958 8401
rect 20866 8329 20958 8346
rect 22100 8402 22157 8406
rect 22100 8342 22104 8402
rect 22153 8342 22157 8402
rect 22100 8338 22157 8342
rect 20659 8165 20693 8181
rect 20659 8115 20693 8131
rect 17154 8047 17188 8063
rect 17154 7855 17188 7871
rect 17272 8059 17306 8063
rect 17350 8059 17384 8063
rect 17272 8047 17384 8059
rect 17306 7871 17350 8047
rect 17272 7859 17350 7871
rect 17272 7855 17306 7859
rect 17350 7655 17384 7671
rect 17468 8047 17502 8063
rect 17468 7655 17502 7671
rect 17586 8047 17620 8063
rect 17586 7655 17620 7671
rect 17704 8047 17738 8063
rect 17704 7655 17738 7671
rect 17822 8059 17856 8063
rect 17896 8059 17930 8063
rect 17822 8047 17930 8059
rect 17856 7871 17896 8047
rect 17856 7859 17930 7871
rect 17896 7855 17930 7859
rect 18014 8047 18048 8063
rect 19159 8008 19484 8072
rect 18014 7855 18048 7871
rect 17822 7655 17856 7671
rect 17569 7536 17585 7570
rect 17619 7536 17635 7570
rect 17518 7418 17654 7422
rect 17518 7404 17558 7418
rect 17616 7404 17654 7418
rect 17518 7358 17534 7404
rect 17638 7358 17654 7404
rect 17518 7336 17654 7358
rect 16033 7182 17403 7246
rect 16194 6704 16396 6724
rect 16194 6660 16240 6704
rect 16362 6660 16396 6704
rect 16194 6650 16272 6660
rect 16310 6650 16396 6660
rect 16194 6632 16396 6650
rect 16039 6486 16309 6521
rect 15921 6433 15955 6449
rect 15438 6233 15472 6249
rect 15438 6041 15472 6057
rect 15556 6233 15590 6249
rect 15556 6041 15590 6057
rect 15674 6233 15708 6249
rect 15674 6041 15708 6057
rect 15792 6233 15826 6249
rect 15792 6041 15826 6057
rect 15921 6041 15955 6057
rect 16039 6433 16073 6486
rect 16039 6041 16073 6057
rect 16157 6433 16191 6449
rect 16157 6041 16191 6057
rect 16275 6433 16309 6486
rect 16275 6041 16309 6057
rect 16393 6433 16427 6449
rect 16393 6041 16427 6057
rect 16511 6433 16545 6449
rect 16511 6041 16545 6057
rect 16629 6433 16663 6449
rect 16877 6287 17147 6322
rect 16629 6041 16663 6057
rect 16759 6233 16793 6249
rect 16759 6041 16793 6057
rect 16877 6233 16911 6287
rect 16877 6041 16911 6057
rect 16995 6233 17029 6249
rect 16995 6041 17029 6057
rect 17113 6233 17147 6287
rect 17113 6041 17147 6057
rect 15680 5844 15686 5878
rect 15740 5844 15746 5878
rect 15978 5740 16012 5756
rect 16096 5740 16130 5756
rect 15978 5348 16012 5364
rect 16094 5364 16096 5410
rect 13440 5267 14516 5268
rect 12502 5176 12569 5192
rect 12502 5142 12519 5176
rect 12553 5142 12569 5176
rect 12502 5126 12569 5142
rect 13924 5178 13991 5194
rect 13924 5144 13940 5178
rect 13974 5144 13991 5178
rect 13924 5128 13991 5144
rect 12704 5109 12738 5125
rect 12704 5059 12738 5075
rect 13650 5110 13684 5126
rect 13650 5060 13684 5076
rect 14188 5061 14204 5095
rect 14238 5061 14254 5095
rect 14306 5060 14322 5094
rect 14356 5060 14372 5094
rect 14427 5026 14461 5267
rect 15273 5265 15406 5306
rect 16094 5306 16130 5364
rect 16214 5740 16248 5756
rect 16214 5348 16248 5364
rect 16332 5740 16366 5756
rect 16450 5740 16484 5756
rect 16366 5364 16368 5411
rect 16332 5306 16368 5364
rect 16568 5740 16602 5756
rect 16450 5348 16484 5364
rect 16567 5364 16568 5411
rect 16686 5740 16720 5756
rect 16602 5364 16603 5411
rect 16567 5306 16603 5364
rect 16686 5348 16720 5364
rect 15508 5266 16603 5306
rect 17338 5319 17403 7182
rect 18263 6704 18465 6724
rect 18263 6660 18309 6704
rect 18431 6660 18465 6704
rect 18263 6650 18341 6660
rect 18379 6650 18465 6660
rect 18263 6632 18465 6650
rect 18108 6486 18378 6521
rect 17990 6433 18024 6449
rect 17507 6233 17541 6249
rect 17507 6041 17541 6057
rect 17625 6233 17659 6249
rect 17625 6041 17659 6057
rect 17743 6233 17777 6249
rect 17743 6041 17777 6057
rect 17861 6233 17895 6249
rect 17861 6041 17895 6057
rect 17990 6041 18024 6057
rect 18108 6433 18142 6486
rect 18108 6041 18142 6057
rect 18226 6433 18260 6449
rect 18226 6041 18260 6057
rect 18344 6433 18378 6486
rect 18344 6041 18378 6057
rect 18462 6433 18496 6449
rect 18462 6041 18496 6057
rect 18580 6433 18614 6449
rect 18580 6041 18614 6057
rect 18698 6433 18732 6449
rect 18946 6287 19216 6322
rect 18698 6041 18732 6057
rect 18828 6233 18862 6249
rect 18828 6041 18862 6057
rect 18946 6233 18980 6287
rect 18946 6041 18980 6057
rect 19064 6233 19098 6249
rect 19064 6041 19098 6057
rect 19182 6233 19216 6287
rect 19182 6041 19216 6057
rect 17749 5844 17755 5878
rect 17809 5844 17815 5878
rect 18047 5740 18081 5756
rect 18165 5740 18199 5756
rect 18047 5348 18081 5364
rect 18163 5364 18165 5410
rect 15508 5265 16584 5266
rect 14571 5178 14638 5194
rect 14571 5144 14588 5178
rect 14622 5144 14638 5178
rect 14571 5128 14638 5144
rect 15992 5176 16059 5192
rect 15992 5142 16008 5176
rect 16042 5142 16059 5176
rect 14773 5111 14807 5127
rect 15992 5126 16059 5142
rect 14773 5061 14807 5077
rect 15718 5108 15752 5124
rect 15718 5058 15752 5074
rect 16256 5059 16272 5093
rect 16306 5059 16322 5093
rect 16374 5058 16390 5092
rect 16424 5058 16440 5092
rect 10783 4818 10817 4834
rect 11435 5008 11469 5024
rect 11435 4816 11469 4832
rect 11553 5008 11587 5024
rect 11553 4816 11587 4832
rect 11959 5008 11993 5024
rect 10245 4618 10279 4634
rect 10362 4567 10397 4634
rect 9891 4532 10397 4567
rect 12077 5008 12111 5024
rect 11959 4565 11994 4632
rect 12077 4616 12111 4632
rect 12195 5008 12229 5024
rect 12195 4616 12229 4632
rect 12313 5008 12392 5024
rect 12347 4978 12392 5008
rect 12431 5008 12465 5024
rect 12733 5008 12767 5024
rect 12733 4816 12767 4832
rect 12851 5008 12885 5024
rect 12851 4816 12885 4832
rect 13504 5010 13538 5026
rect 13504 4818 13538 4834
rect 13622 5010 13656 5026
rect 13622 4818 13656 4834
rect 14028 5010 14062 5026
rect 12313 4616 12347 4632
rect 12430 4565 12465 4632
rect 11959 4530 12465 4565
rect 14146 5010 14180 5026
rect 14028 4567 14063 4634
rect 14146 4618 14180 4634
rect 14264 5010 14298 5026
rect 14264 4618 14298 4634
rect 14382 5010 14461 5026
rect 14416 4980 14461 5010
rect 14500 5010 14534 5026
rect 14802 5010 14836 5026
rect 14802 4818 14836 4834
rect 14920 5010 14954 5026
rect 16495 5024 16529 5265
rect 17338 5255 17475 5319
rect 18163 5306 18199 5364
rect 18283 5740 18317 5756
rect 18283 5348 18317 5364
rect 18401 5740 18435 5756
rect 18519 5740 18553 5756
rect 18435 5364 18437 5411
rect 18401 5306 18437 5364
rect 18637 5740 18671 5756
rect 18519 5348 18553 5364
rect 18636 5364 18637 5411
rect 18755 5740 18789 5756
rect 18671 5364 18672 5411
rect 18636 5306 18672 5364
rect 18755 5348 18789 5364
rect 17577 5266 18672 5306
rect 19420 5315 19484 8008
rect 20286 8043 20320 8059
rect 20286 7851 20320 7867
rect 20404 8055 20438 8059
rect 20482 8055 20516 8059
rect 20404 8043 20516 8055
rect 20438 7867 20482 8043
rect 20404 7855 20482 7867
rect 20404 7851 20438 7855
rect 20482 7651 20516 7667
rect 20600 8043 20634 8059
rect 20600 7651 20634 7667
rect 20718 8043 20752 8059
rect 20718 7651 20752 7667
rect 20836 8043 20870 8059
rect 20836 7651 20870 7667
rect 20954 8055 20988 8059
rect 21028 8055 21062 8059
rect 20954 8043 21062 8055
rect 20988 7867 21028 8043
rect 20988 7855 21062 7867
rect 21028 7851 21062 7855
rect 21146 8043 21180 8059
rect 21146 7851 21180 7867
rect 20954 7651 20988 7667
rect 20701 7532 20717 7566
rect 20751 7532 20767 7566
rect 20650 7414 20786 7418
rect 20650 7400 20690 7414
rect 20748 7400 20786 7414
rect 20650 7354 20666 7400
rect 20770 7354 20786 7400
rect 20650 7332 20786 7354
rect 22289 6928 22353 8508
rect 23684 8555 23718 8571
rect 23684 8505 23718 8521
rect 25244 8570 25301 8574
rect 25465 8570 25581 8571
rect 30643 8570 30659 8604
rect 31035 8570 31051 8604
rect 31207 8574 31273 8590
rect 25244 8510 25248 8570
rect 25297 8510 25581 8570
rect 29950 8513 29966 8547
rect 30342 8513 30358 8547
rect 31207 8540 31223 8574
rect 31257 8540 31273 8574
rect 31207 8523 31273 8540
rect 25244 8506 25581 8510
rect 24010 8401 24102 8414
rect 24010 8346 24026 8401
rect 24086 8346 24102 8401
rect 24010 8329 24102 8346
rect 25244 8402 25301 8406
rect 25244 8342 25248 8402
rect 25297 8342 25301 8402
rect 25244 8338 25301 8342
rect 23803 8165 23837 8181
rect 23803 8115 23837 8131
rect 23430 8043 23464 8059
rect 23430 7851 23464 7867
rect 23548 8055 23582 8059
rect 23626 8055 23660 8059
rect 23548 8043 23660 8055
rect 23582 7867 23626 8043
rect 23548 7855 23626 7867
rect 23548 7851 23582 7855
rect 23626 7651 23660 7667
rect 23744 8043 23778 8059
rect 23744 7651 23778 7667
rect 23862 8043 23896 8059
rect 23862 7651 23896 7667
rect 23980 8043 24014 8059
rect 23980 7651 24014 7667
rect 24098 8055 24132 8059
rect 24172 8055 24206 8059
rect 24098 8043 24206 8055
rect 24132 7867 24172 8043
rect 24132 7855 24206 7867
rect 24172 7851 24206 7855
rect 24290 8043 24324 8059
rect 24290 7851 24324 7867
rect 24098 7651 24132 7667
rect 23845 7532 23861 7566
rect 23895 7532 23911 7566
rect 23794 7414 23930 7418
rect 23794 7400 23834 7414
rect 23892 7400 23930 7414
rect 23794 7354 23810 7400
rect 23914 7354 23930 7400
rect 23794 7332 23930 7354
rect 25516 6944 25580 8506
rect 30988 8486 31133 8487
rect 30643 8452 30659 8486
rect 31035 8468 31133 8486
rect 31035 8452 31134 8468
rect 31375 8452 31391 8486
rect 30988 8451 31134 8452
rect 31767 8451 31869 8486
rect 29950 8395 29966 8429
rect 30342 8395 30358 8429
rect 31093 8413 31134 8451
rect 31093 8379 31421 8413
rect 30643 8334 30659 8368
rect 31035 8334 31051 8368
rect 29675 8246 29767 8280
rect 29950 8277 29966 8311
rect 30342 8277 30358 8311
rect 31093 8252 31134 8379
rect 31375 8368 31421 8379
rect 31375 8334 31391 8368
rect 31767 8334 31783 8368
rect 31307 8308 31341 8324
rect 31307 8258 31341 8274
rect 30988 8250 31134 8252
rect 29675 8124 29695 8246
rect 29739 8194 29767 8246
rect 30643 8216 30659 8250
rect 31035 8216 31134 8250
rect 31375 8216 31391 8250
rect 31767 8216 31783 8250
rect 29749 8156 29767 8194
rect 29739 8124 29767 8156
rect 29675 8078 29767 8124
rect 29878 8159 29966 8193
rect 30342 8159 30358 8193
rect 29878 7957 29913 8159
rect 30643 8098 30659 8132
rect 31035 8098 31051 8132
rect 29950 8041 29966 8075
rect 30342 8041 30358 8075
rect 31093 8014 31134 8216
rect 31306 8190 31340 8206
rect 31306 8140 31340 8156
rect 31375 8098 31391 8132
rect 31767 8098 31783 8132
rect 31834 8015 31869 8451
rect 31939 8296 32027 8312
rect 31939 8256 31955 8296
rect 31939 8164 31955 8206
rect 32011 8164 32027 8296
rect 31939 8148 32027 8164
rect 30643 7980 30659 8014
rect 31035 7980 31134 8014
rect 31375 7980 31391 8014
rect 31767 7980 31869 8015
rect 30989 7978 31134 7980
rect 29878 7923 29966 7957
rect 30342 7923 30358 7957
rect 30643 7862 30659 7896
rect 31035 7862 31051 7896
rect 29950 7805 29966 7839
rect 30342 7805 30358 7839
rect 30150 7676 30166 7710
rect 30342 7676 30358 7710
rect 30521 7624 30555 7630
rect 30150 7558 30166 7592
rect 30342 7558 30358 7592
rect 30521 7564 30555 7570
rect 30150 7440 30166 7474
rect 30342 7440 30358 7474
rect 31093 7392 31134 7978
rect 31207 7926 31273 7943
rect 31207 7892 31223 7926
rect 31257 7892 31273 7926
rect 31207 7876 31273 7892
rect 31275 7602 31291 7636
rect 31325 7602 31341 7636
rect 31375 7574 31391 7608
rect 31567 7574 31583 7608
rect 31375 7456 31391 7490
rect 31567 7456 31583 7490
rect 30150 7322 30166 7356
rect 30342 7322 30358 7356
rect 21515 6864 22353 6928
rect 23581 6880 25580 6944
rect 30075 6929 30164 6963
rect 30340 6929 30356 6963
rect 33364 6941 33458 21486
rect 33511 9477 33601 21936
rect 20331 6702 20533 6722
rect 20331 6658 20377 6702
rect 20499 6658 20533 6702
rect 20331 6648 20409 6658
rect 20447 6648 20533 6658
rect 20331 6630 20533 6648
rect 20176 6484 20446 6519
rect 20058 6431 20092 6447
rect 19575 6231 19609 6247
rect 19575 6039 19609 6055
rect 19693 6231 19727 6247
rect 19693 6039 19727 6055
rect 19811 6231 19845 6247
rect 19811 6039 19845 6055
rect 19929 6231 19963 6247
rect 19929 6039 19963 6055
rect 20058 6039 20092 6055
rect 20176 6431 20210 6484
rect 20176 6039 20210 6055
rect 20294 6431 20328 6447
rect 20294 6039 20328 6055
rect 20412 6431 20446 6484
rect 20412 6039 20446 6055
rect 20530 6431 20564 6447
rect 20530 6039 20564 6055
rect 20648 6431 20682 6447
rect 20648 6039 20682 6055
rect 20766 6431 20800 6447
rect 21014 6285 21284 6320
rect 20766 6039 20800 6055
rect 20896 6231 20930 6247
rect 20896 6039 20930 6055
rect 21014 6231 21048 6285
rect 21014 6039 21048 6055
rect 21132 6231 21166 6247
rect 21132 6039 21166 6055
rect 21250 6231 21284 6285
rect 21250 6039 21284 6055
rect 19817 5842 19823 5876
rect 19877 5842 19883 5876
rect 20115 5738 20149 5754
rect 20233 5738 20267 5754
rect 20115 5346 20149 5362
rect 20231 5362 20233 5408
rect 17577 5265 18653 5266
rect 16639 5176 16706 5192
rect 16639 5142 16656 5176
rect 16690 5142 16706 5176
rect 16639 5126 16706 5142
rect 18061 5176 18128 5192
rect 18061 5142 18077 5176
rect 18111 5142 18128 5176
rect 18061 5126 18128 5142
rect 16841 5109 16875 5125
rect 16841 5059 16875 5075
rect 17787 5108 17821 5124
rect 17787 5058 17821 5074
rect 18325 5059 18341 5093
rect 18375 5059 18391 5093
rect 18443 5058 18459 5092
rect 18493 5058 18509 5092
rect 18564 5024 18598 5265
rect 19420 5251 19543 5315
rect 20231 5304 20267 5362
rect 20351 5738 20385 5754
rect 20351 5346 20385 5362
rect 20469 5738 20503 5754
rect 20587 5738 20621 5754
rect 20503 5362 20505 5409
rect 20469 5304 20505 5362
rect 20705 5738 20739 5754
rect 20587 5346 20621 5362
rect 20704 5362 20705 5409
rect 20823 5738 20857 5754
rect 20739 5362 20740 5409
rect 20704 5304 20740 5362
rect 20823 5346 20857 5362
rect 19645 5264 20740 5304
rect 21516 5306 21572 6864
rect 22400 6704 22602 6724
rect 22400 6660 22446 6704
rect 22568 6660 22602 6704
rect 22400 6650 22478 6660
rect 22516 6650 22602 6660
rect 22400 6632 22602 6650
rect 22245 6486 22515 6521
rect 22127 6433 22161 6449
rect 21644 6233 21678 6249
rect 21644 6041 21678 6057
rect 21762 6233 21796 6249
rect 21762 6041 21796 6057
rect 21880 6233 21914 6249
rect 21880 6041 21914 6057
rect 21998 6233 22032 6249
rect 21998 6041 22032 6057
rect 22127 6041 22161 6057
rect 22245 6433 22279 6486
rect 22245 6041 22279 6057
rect 22363 6433 22397 6449
rect 22363 6041 22397 6057
rect 22481 6433 22515 6486
rect 22481 6041 22515 6057
rect 22599 6433 22633 6449
rect 22599 6041 22633 6057
rect 22717 6433 22751 6449
rect 22717 6041 22751 6057
rect 22835 6433 22869 6449
rect 23083 6287 23353 6322
rect 22835 6041 22869 6057
rect 22965 6233 22999 6249
rect 22965 6041 22999 6057
rect 23083 6233 23117 6287
rect 23083 6041 23117 6057
rect 23201 6233 23235 6249
rect 23201 6041 23235 6057
rect 23319 6233 23353 6287
rect 23319 6041 23353 6057
rect 21886 5844 21892 5878
rect 21946 5844 21952 5878
rect 22184 5740 22218 5756
rect 22302 5740 22336 5756
rect 22184 5348 22218 5364
rect 22300 5364 22302 5410
rect 21516 5265 21612 5306
rect 19645 5263 20721 5264
rect 18708 5176 18775 5192
rect 18708 5142 18725 5176
rect 18759 5142 18775 5176
rect 18708 5126 18775 5142
rect 20129 5174 20196 5190
rect 20129 5140 20145 5174
rect 20179 5140 20196 5174
rect 18910 5109 18944 5125
rect 20129 5124 20196 5140
rect 18910 5059 18944 5075
rect 19855 5106 19889 5122
rect 19855 5056 19889 5072
rect 20393 5057 20409 5091
rect 20443 5057 20459 5091
rect 20511 5056 20527 5090
rect 20561 5056 20577 5090
rect 14920 4818 14954 4834
rect 15572 5008 15606 5024
rect 15572 4816 15606 4832
rect 15690 5008 15724 5024
rect 15690 4816 15724 4832
rect 16096 5008 16130 5024
rect 14382 4618 14416 4634
rect 14499 4567 14534 4634
rect 14028 4532 14534 4567
rect 16214 5008 16248 5024
rect 16096 4565 16131 4632
rect 16214 4616 16248 4632
rect 16332 5008 16366 5024
rect 16332 4616 16366 4632
rect 16450 5008 16529 5024
rect 16484 4978 16529 5008
rect 16568 5008 16602 5024
rect 16870 5008 16904 5024
rect 16870 4816 16904 4832
rect 16988 5008 17022 5024
rect 16988 4816 17022 4832
rect 17641 5008 17675 5024
rect 17641 4816 17675 4832
rect 17759 5008 17793 5024
rect 17759 4816 17793 4832
rect 18165 5008 18199 5024
rect 16450 4616 16484 4632
rect 16567 4565 16602 4632
rect 16096 4530 16602 4565
rect 18283 5008 18317 5024
rect 18165 4565 18200 4632
rect 18283 4616 18317 4632
rect 18401 5008 18435 5024
rect 18401 4616 18435 4632
rect 18519 5008 18598 5024
rect 18553 4978 18598 5008
rect 18637 5008 18671 5024
rect 18939 5008 18973 5024
rect 18939 4816 18973 4832
rect 19057 5008 19091 5024
rect 20632 5022 20666 5263
rect 22300 5306 22336 5364
rect 22420 5740 22454 5756
rect 22420 5348 22454 5364
rect 22538 5740 22572 5756
rect 22656 5740 22690 5756
rect 22572 5364 22574 5411
rect 22538 5306 22574 5364
rect 22774 5740 22808 5756
rect 22656 5348 22690 5364
rect 22773 5364 22774 5411
rect 22892 5740 22926 5756
rect 22808 5364 22809 5411
rect 22773 5306 22809 5364
rect 22892 5348 22926 5364
rect 21714 5266 22809 5306
rect 23581 5317 23645 6880
rect 30075 6727 30110 6929
rect 30148 6811 30164 6845
rect 30340 6811 30356 6845
rect 31373 6804 31389 6838
rect 31565 6804 31581 6838
rect 24468 6702 24670 6722
rect 24468 6658 24514 6702
rect 24636 6658 24670 6702
rect 30075 6693 30164 6727
rect 30340 6693 30356 6727
rect 24468 6648 24546 6658
rect 24584 6648 24670 6658
rect 31272 6657 31288 6691
rect 31322 6657 31338 6691
rect 31373 6686 31389 6720
rect 31565 6686 31581 6720
rect 24468 6630 24670 6648
rect 30148 6575 30164 6609
rect 30340 6575 30356 6609
rect 24313 6484 24583 6519
rect 30641 6502 30657 6536
rect 31033 6502 31049 6536
rect 31205 6506 31271 6522
rect 24195 6431 24229 6447
rect 23712 6231 23746 6247
rect 23712 6039 23746 6055
rect 23830 6231 23864 6247
rect 23830 6039 23864 6055
rect 23948 6231 23982 6247
rect 23948 6039 23982 6055
rect 24066 6231 24100 6247
rect 24066 6039 24100 6055
rect 24195 6039 24229 6055
rect 24313 6431 24347 6484
rect 24313 6039 24347 6055
rect 24431 6431 24465 6447
rect 24431 6039 24465 6055
rect 24549 6431 24583 6484
rect 24549 6039 24583 6055
rect 24667 6431 24701 6447
rect 24667 6039 24701 6055
rect 24785 6431 24819 6447
rect 24785 6039 24819 6055
rect 24903 6431 24937 6447
rect 29948 6445 29964 6479
rect 30340 6445 30356 6479
rect 31205 6472 31221 6506
rect 31255 6472 31271 6506
rect 31205 6455 31271 6472
rect 30986 6418 31131 6419
rect 30641 6384 30657 6418
rect 31033 6400 31131 6418
rect 31033 6384 31132 6400
rect 31373 6384 31389 6418
rect 30986 6383 31132 6384
rect 31765 6383 31867 6418
rect 29948 6327 29964 6361
rect 30340 6327 30356 6361
rect 31091 6345 31132 6383
rect 25151 6285 25421 6320
rect 31091 6311 31419 6345
rect 24903 6039 24937 6055
rect 25033 6231 25067 6247
rect 25033 6039 25067 6055
rect 25151 6231 25185 6285
rect 25151 6039 25185 6055
rect 25269 6231 25303 6247
rect 25269 6039 25303 6055
rect 25387 6231 25421 6285
rect 30641 6266 30657 6300
rect 31033 6266 31049 6300
rect 25387 6039 25421 6055
rect 29673 6178 29765 6212
rect 29948 6209 29964 6243
rect 30340 6209 30356 6243
rect 31091 6184 31132 6311
rect 31373 6300 31419 6311
rect 31373 6266 31389 6300
rect 31765 6266 31781 6300
rect 31305 6240 31339 6256
rect 31305 6190 31339 6206
rect 30986 6182 31132 6184
rect 29673 6056 29693 6178
rect 29737 6126 29765 6178
rect 30641 6148 30657 6182
rect 31033 6148 31132 6182
rect 31373 6148 31389 6182
rect 31765 6148 31781 6182
rect 29747 6088 29765 6126
rect 29737 6056 29765 6088
rect 29673 6010 29765 6056
rect 29876 6091 29964 6125
rect 30340 6091 30356 6125
rect 29876 5889 29911 6091
rect 30641 6030 30657 6064
rect 31033 6030 31049 6064
rect 29948 5973 29964 6007
rect 30340 5973 30356 6007
rect 31091 5946 31132 6148
rect 31304 6122 31338 6138
rect 31304 6072 31338 6088
rect 31373 6030 31389 6064
rect 31765 6030 31781 6064
rect 31832 5947 31867 6383
rect 31937 6228 32025 6244
rect 31937 6188 31953 6228
rect 31937 6096 31953 6138
rect 32009 6096 32025 6228
rect 31937 6080 32025 6096
rect 30641 5912 30657 5946
rect 31033 5912 31132 5946
rect 31373 5912 31389 5946
rect 31765 5912 31867 5947
rect 30987 5910 31132 5912
rect 23954 5842 23960 5876
rect 24014 5842 24020 5876
rect 29876 5855 29964 5889
rect 30340 5855 30356 5889
rect 30641 5794 30657 5828
rect 31033 5794 31049 5828
rect 24252 5738 24286 5754
rect 24370 5738 24404 5754
rect 24252 5346 24286 5362
rect 24368 5362 24370 5408
rect 21714 5265 22790 5266
rect 20776 5174 20843 5190
rect 20776 5140 20793 5174
rect 20827 5140 20843 5174
rect 20776 5124 20843 5140
rect 22198 5176 22265 5192
rect 22198 5142 22214 5176
rect 22248 5142 22265 5176
rect 22198 5126 22265 5142
rect 20978 5107 21012 5123
rect 20978 5057 21012 5073
rect 21924 5108 21958 5124
rect 21924 5058 21958 5074
rect 22462 5059 22478 5093
rect 22512 5059 22528 5093
rect 22580 5058 22596 5092
rect 22630 5058 22646 5092
rect 22701 5024 22735 5265
rect 23581 5253 23680 5317
rect 24368 5304 24404 5362
rect 24488 5738 24522 5754
rect 24488 5346 24522 5362
rect 24606 5738 24640 5754
rect 24724 5738 24758 5754
rect 24640 5362 24642 5409
rect 24606 5304 24642 5362
rect 24842 5738 24876 5754
rect 24724 5346 24758 5362
rect 24841 5362 24842 5409
rect 24960 5738 24994 5754
rect 24876 5362 24877 5409
rect 24841 5304 24877 5362
rect 29948 5737 29964 5771
rect 30340 5737 30356 5771
rect 25414 5636 25451 5696
rect 25386 5580 25451 5636
rect 30148 5608 30164 5642
rect 30340 5608 30356 5642
rect 24960 5346 24994 5362
rect 23782 5264 24877 5304
rect 23782 5263 24858 5264
rect 22845 5176 22912 5192
rect 22845 5142 22862 5176
rect 22896 5142 22912 5176
rect 22845 5126 22912 5142
rect 24266 5174 24333 5190
rect 24266 5140 24282 5174
rect 24316 5140 24333 5174
rect 23047 5109 23081 5125
rect 24266 5124 24333 5140
rect 23047 5059 23081 5075
rect 23992 5106 24026 5122
rect 23992 5056 24026 5072
rect 24530 5057 24546 5091
rect 24580 5057 24596 5091
rect 24648 5056 24664 5090
rect 24698 5056 24714 5090
rect 19057 4816 19091 4832
rect 19709 5006 19743 5022
rect 19709 4814 19743 4830
rect 19827 5006 19861 5022
rect 19827 4814 19861 4830
rect 20233 5006 20267 5022
rect 18519 4616 18553 4632
rect 18636 4565 18671 4632
rect 18165 4530 18671 4565
rect 20351 5006 20385 5022
rect 20233 4563 20268 4630
rect 20351 4614 20385 4630
rect 20469 5006 20503 5022
rect 20469 4614 20503 4630
rect 20587 5006 20666 5022
rect 20621 4976 20666 5006
rect 20705 5006 20739 5022
rect 21007 5006 21041 5022
rect 21007 4814 21041 4830
rect 21125 5006 21159 5022
rect 21125 4814 21159 4830
rect 21778 5008 21812 5024
rect 21778 4816 21812 4832
rect 21896 5008 21930 5024
rect 21896 4816 21930 4832
rect 22302 5008 22336 5024
rect 20587 4614 20621 4630
rect 20704 4563 20739 4630
rect 20233 4528 20739 4563
rect 22420 5008 22454 5024
rect 22302 4565 22337 4632
rect 22420 4616 22454 4632
rect 22538 5008 22572 5024
rect 22538 4616 22572 4632
rect 22656 5008 22735 5024
rect 22690 4978 22735 5008
rect 22774 5008 22808 5024
rect 23076 5008 23110 5024
rect 23076 4816 23110 4832
rect 23194 5008 23228 5024
rect 24769 5022 24803 5263
rect 24913 5174 24980 5190
rect 24913 5140 24930 5174
rect 24964 5140 24980 5174
rect 24913 5124 24980 5140
rect 25115 5107 25149 5123
rect 25115 5057 25149 5073
rect 23194 4816 23228 4832
rect 23846 5006 23880 5022
rect 23846 4814 23880 4830
rect 23964 5006 23998 5022
rect 23964 4814 23998 4830
rect 24370 5006 24404 5022
rect 22656 4616 22690 4632
rect 22773 4565 22808 4632
rect 22302 4530 22808 4565
rect 24488 5006 24522 5022
rect 24370 4563 24405 4630
rect 24488 4614 24522 4630
rect 24606 5006 24640 5022
rect 24606 4614 24640 4630
rect 24724 5006 24803 5022
rect 24758 4976 24803 5006
rect 24842 5006 24876 5022
rect 25144 5006 25178 5022
rect 25144 4814 25178 4830
rect 25262 5006 25296 5022
rect 25262 4814 25296 4830
rect 24724 4614 24758 4630
rect 24841 4563 24876 4630
rect 24370 4528 24876 4563
rect 10059 4446 10117 4462
rect 10167 4446 10223 4462
rect 10059 4390 10075 4446
rect 10207 4390 10223 4446
rect 10059 4374 10223 4390
rect 12127 4444 12185 4460
rect 12235 4444 12291 4460
rect 12127 4388 12143 4444
rect 12275 4388 12291 4444
rect 12127 4372 12291 4388
rect 14196 4446 14254 4462
rect 14304 4446 14360 4462
rect 14196 4390 14212 4446
rect 14344 4390 14360 4446
rect 14196 4374 14360 4390
rect 16264 4444 16322 4460
rect 16372 4444 16428 4460
rect 16264 4388 16280 4444
rect 16412 4388 16428 4444
rect 16264 4372 16428 4388
rect 18333 4444 18391 4460
rect 18441 4444 18497 4460
rect 18333 4388 18349 4444
rect 18481 4388 18497 4444
rect 18333 4372 18497 4388
rect 20401 4442 20459 4458
rect 20509 4442 20565 4458
rect 20401 4386 20417 4442
rect 20549 4386 20565 4442
rect 20401 4370 20565 4386
rect 22470 4444 22528 4460
rect 22578 4444 22634 4460
rect 22470 4388 22486 4444
rect 22618 4388 22634 4444
rect 22470 4372 22634 4388
rect 24538 4442 24596 4458
rect 24646 4442 24702 4458
rect 24538 4386 24554 4442
rect 24686 4386 24702 4442
rect 24538 4370 24702 4386
rect 25387 4154 25451 5580
rect 30519 5556 30553 5562
rect 30148 5490 30164 5524
rect 30340 5490 30356 5524
rect 30519 5496 30553 5502
rect 30148 5372 30164 5406
rect 30340 5372 30356 5406
rect 31091 5324 31132 5910
rect 31205 5858 31271 5875
rect 31205 5824 31221 5858
rect 31255 5824 31271 5858
rect 31205 5808 31271 5824
rect 31273 5534 31289 5568
rect 31323 5534 31339 5568
rect 31373 5506 31389 5540
rect 31565 5506 31581 5540
rect 31373 5388 31389 5422
rect 31565 5388 31581 5422
rect 30148 5254 30164 5288
rect 30340 5254 30356 5288
rect 30075 4860 30164 4894
rect 30340 4860 30356 4894
rect 30075 4658 30110 4860
rect 30148 4742 30164 4776
rect 30340 4742 30356 4776
rect 31373 4735 31389 4769
rect 31565 4735 31581 4769
rect 30075 4624 30164 4658
rect 30340 4624 30356 4658
rect 31272 4588 31288 4622
rect 31322 4588 31338 4622
rect 31373 4617 31389 4651
rect 31565 4617 31581 4651
rect 30148 4506 30164 4540
rect 30340 4506 30356 4540
rect 30641 4433 30657 4467
rect 31033 4433 31049 4467
rect 31205 4437 31271 4453
rect 29948 4376 29964 4410
rect 30340 4376 30356 4410
rect 31205 4403 31221 4437
rect 31255 4403 31271 4437
rect 31205 4386 31271 4403
rect 30986 4349 31131 4350
rect 30641 4315 30657 4349
rect 31033 4331 31131 4349
rect 31033 4315 31132 4331
rect 31373 4315 31389 4349
rect 30986 4314 31132 4315
rect 31765 4314 31867 4349
rect 29948 4258 29964 4292
rect 30340 4258 30356 4292
rect 31091 4276 31132 4314
rect 31091 4242 31419 4276
rect 30641 4197 30657 4231
rect 31033 4197 31049 4231
rect 8695 4090 25451 4154
rect 29673 4109 29765 4143
rect 29948 4140 29964 4174
rect 30340 4140 30356 4174
rect 31091 4115 31132 4242
rect 31373 4231 31419 4242
rect 31373 4197 31389 4231
rect 31765 4197 31781 4231
rect 31305 4171 31339 4187
rect 31305 4121 31339 4137
rect 30986 4113 31132 4115
rect 8095 4055 23401 4056
rect 8095 4004 23350 4055
rect 8095 3992 23401 4004
rect 29673 3987 29693 4109
rect 29737 4057 29765 4109
rect 30641 4079 30657 4113
rect 31033 4079 31132 4113
rect 31373 4079 31389 4113
rect 31765 4079 31781 4113
rect 29747 4019 29765 4057
rect 29737 3987 29765 4019
rect 7375 3896 21319 3947
rect 29673 3941 29765 3987
rect 29876 4022 29964 4056
rect 30340 4022 30356 4056
rect 7375 3883 21366 3896
rect 21303 3882 21366 3883
rect 6646 3847 19328 3849
rect 6646 3793 19272 3847
rect 19319 3793 19328 3847
rect 6646 3785 19328 3793
rect 29876 3820 29911 4022
rect 30641 3961 30657 3995
rect 31033 3961 31049 3995
rect 29948 3904 29964 3938
rect 30340 3904 30356 3938
rect 31091 3877 31132 4079
rect 31304 4053 31338 4069
rect 31304 4003 31338 4019
rect 31373 3961 31389 3995
rect 31765 3961 31781 3995
rect 31832 3878 31867 4314
rect 31937 4159 32025 4175
rect 31937 4119 31953 4159
rect 31937 4027 31953 4069
rect 32009 4027 32025 4159
rect 31937 4011 32025 4027
rect 30641 3843 30657 3877
rect 31033 3843 31132 3877
rect 31373 3843 31389 3877
rect 31765 3843 31867 3878
rect 30987 3841 31132 3843
rect 29876 3786 29964 3820
rect 30340 3786 30356 3820
rect 5823 3737 17229 3741
rect 5823 3686 17179 3737
rect 30641 3725 30657 3759
rect 31033 3725 31049 3759
rect 5823 3677 17229 3686
rect 29948 3668 29964 3702
rect 30340 3668 30356 3702
rect 5125 3642 15158 3643
rect 5125 3589 15107 3642
rect 5125 3579 15158 3589
rect 30148 3539 30164 3573
rect 30340 3539 30356 3573
rect 4334 3498 13065 3502
rect 4334 3447 13011 3498
rect 13055 3447 13065 3498
rect 30519 3487 30553 3493
rect 4334 3438 13065 3447
rect 30148 3421 30164 3455
rect 30340 3421 30356 3455
rect 30519 3427 30553 3433
rect 3577 3403 10987 3404
rect 3577 3349 10934 3403
rect 3577 3340 10987 3349
rect 10906 3339 10987 3340
rect 30148 3303 30164 3337
rect 30340 3303 30356 3337
rect 31091 3255 31132 3841
rect 31205 3789 31271 3806
rect 31205 3755 31221 3789
rect 31255 3755 31271 3789
rect 31205 3739 31271 3755
rect 31273 3465 31289 3499
rect 31323 3465 31339 3499
rect 31373 3437 31389 3471
rect 31565 3437 31581 3471
rect 31373 3319 31389 3353
rect 31565 3319 31581 3353
rect 30148 3185 30164 3219
rect 30340 3185 30356 3219
rect -1538 3158 227 3175
rect -1538 3122 -1506 3158
rect -1414 3150 227 3158
rect -1414 3122 150 3150
rect -1538 3106 150 3122
rect 204 3106 227 3150
rect -1538 3101 227 3106
rect -1538 3088 -1357 3101
rect 108 3091 227 3101
rect -1277 3057 -1104 3067
rect -1277 3044 226 3057
rect -1277 3001 -1246 3044
rect -1166 3034 226 3044
rect -1166 3001 149 3034
rect -1277 2990 149 3001
rect 203 2990 226 3034
rect -1277 2986 226 2990
rect 115 2972 226 2986
rect 32680 3000 32760 3005
rect -1063 2934 -887 2950
rect 32680 2938 32681 3000
rect 32747 2938 32760 3000
rect -1063 2933 226 2934
rect -1063 2876 -1030 2933
rect -952 2910 226 2933
rect -952 2876 149 2910
rect -1063 2866 149 2876
rect 203 2866 226 2910
rect -1063 2851 226 2866
rect -2397 2802 -1888 2803
rect -2430 2746 -1888 2802
rect 30073 2792 30162 2826
rect 30338 2792 30354 2826
rect -2430 2662 22140 2746
rect -2429 2623 22140 2662
rect 3 1452 107 2623
rect 1430 2398 1658 2416
rect 1430 2322 1446 2398
rect 1642 2322 1658 2398
rect 1430 2306 1658 2322
rect 701 2181 971 2220
rect 701 2128 735 2181
rect 260 1979 530 2018
rect 260 1928 294 1979
rect 260 1736 294 1752
rect 378 1928 412 1944
rect 378 1701 412 1752
rect 496 1928 530 1979
rect 496 1736 530 1752
rect 614 1928 648 1944
rect 614 1701 648 1752
rect 701 1736 735 1752
rect 819 2128 853 2144
rect 378 1662 648 1701
rect 819 1701 853 1752
rect 937 2128 971 2181
rect 1168 2180 1438 2219
rect 937 1736 971 1752
rect 1055 2128 1089 2144
rect 1055 1701 1089 1752
rect 1168 2128 1202 2180
rect 1168 1736 1202 1752
rect 1286 2128 1320 2144
rect 1286 1701 1320 1752
rect 1404 2128 1438 2180
rect 1640 2180 1910 2219
rect 1404 1736 1438 1752
rect 1522 2128 1556 2144
rect 1522 1701 1556 1752
rect 1640 2128 1674 2180
rect 1640 1736 1674 1752
rect 1758 2128 1792 2144
rect 1758 1701 1792 1752
rect 1876 2128 1910 2180
rect 2113 2180 2383 2219
rect 1876 1736 1910 1752
rect 1995 2128 2029 2144
rect 1995 1701 2029 1752
rect 2113 2128 2147 2180
rect 2113 1736 2147 1752
rect 2231 2128 2265 2144
rect 2231 1701 2265 1752
rect 2349 2128 2383 2180
rect 2586 1978 2856 2015
rect 2349 1736 2383 1752
rect 2468 1928 2502 1944
rect 819 1662 2265 1701
rect 2468 1698 2502 1752
rect 2586 1928 2620 1978
rect 2586 1736 2620 1752
rect 2704 1928 2738 1944
rect 2704 1698 2738 1752
rect 2822 1928 2856 1978
rect 2822 1736 2856 1752
rect 2468 1659 2738 1698
rect 1346 1537 1380 1553
rect 2640 1544 2656 1578
rect 2690 1544 2706 1578
rect 1346 1487 1380 1503
rect 3 1438 192 1452
rect 3 1378 121 1438
rect 170 1378 192 1438
rect 3 1363 192 1378
rect 349 1437 441 1454
rect 3143 1453 3238 2623
rect 4574 2398 4802 2416
rect 4574 2322 4590 2398
rect 4786 2322 4802 2398
rect 4574 2306 4802 2322
rect 3845 2181 4115 2220
rect 3845 2128 3879 2181
rect 3404 1979 3674 2018
rect 3404 1928 3438 1979
rect 3404 1736 3438 1752
rect 3522 1928 3556 1944
rect 3522 1701 3556 1752
rect 3640 1928 3674 1979
rect 3640 1736 3674 1752
rect 3758 1928 3792 1944
rect 3758 1701 3792 1752
rect 3845 1736 3879 1752
rect 3963 2128 3997 2144
rect 3522 1662 3792 1701
rect 3963 1701 3997 1752
rect 4081 2128 4115 2181
rect 4312 2180 4582 2219
rect 4081 1736 4115 1752
rect 4199 2128 4233 2144
rect 4199 1701 4233 1752
rect 4312 2128 4346 2180
rect 4312 1736 4346 1752
rect 4430 2128 4464 2144
rect 4430 1701 4464 1752
rect 4548 2128 4582 2180
rect 4784 2180 5054 2219
rect 4548 1736 4582 1752
rect 4666 2128 4700 2144
rect 4666 1701 4700 1752
rect 4784 2128 4818 2180
rect 4784 1736 4818 1752
rect 4902 2128 4936 2144
rect 4902 1701 4936 1752
rect 5020 2128 5054 2180
rect 5257 2180 5527 2219
rect 5020 1736 5054 1752
rect 5139 2128 5173 2144
rect 5139 1701 5173 1752
rect 5257 2128 5291 2180
rect 5257 1736 5291 1752
rect 5375 2128 5409 2144
rect 5375 1701 5409 1752
rect 5493 2128 5527 2180
rect 5730 1978 6000 2015
rect 5493 1736 5527 1752
rect 5612 1928 5646 1944
rect 3963 1662 5409 1701
rect 5612 1698 5646 1752
rect 5730 1928 5764 1978
rect 5730 1736 5764 1752
rect 5848 1928 5882 1944
rect 5848 1698 5882 1752
rect 5966 1928 6000 1978
rect 5966 1736 6000 1752
rect 5612 1659 5882 1698
rect 4490 1537 4524 1553
rect 5784 1544 5800 1578
rect 5834 1544 5850 1578
rect 4490 1487 4524 1503
rect 6275 1454 6374 2623
rect 7706 2402 7934 2420
rect 7706 2326 7722 2402
rect 7918 2326 7934 2402
rect 7706 2310 7934 2326
rect 6977 2185 7247 2224
rect 6977 2132 7011 2185
rect 6536 1983 6806 2022
rect 6536 1932 6570 1983
rect 6536 1740 6570 1756
rect 6654 1932 6688 1948
rect 6654 1705 6688 1756
rect 6772 1932 6806 1983
rect 6772 1740 6806 1756
rect 6890 1932 6924 1948
rect 6890 1705 6924 1756
rect 6977 1740 7011 1756
rect 7095 2132 7129 2148
rect 6654 1666 6924 1705
rect 7095 1705 7129 1756
rect 7213 2132 7247 2185
rect 7444 2184 7714 2223
rect 7213 1740 7247 1756
rect 7331 2132 7365 2148
rect 7331 1705 7365 1756
rect 7444 2132 7478 2184
rect 7444 1740 7478 1756
rect 7562 2132 7596 2148
rect 7562 1705 7596 1756
rect 7680 2132 7714 2184
rect 7916 2184 8186 2223
rect 7680 1740 7714 1756
rect 7798 2132 7832 2148
rect 7798 1705 7832 1756
rect 7916 2132 7950 2184
rect 7916 1740 7950 1756
rect 8034 2132 8068 2148
rect 8034 1705 8068 1756
rect 8152 2132 8186 2184
rect 8389 2184 8659 2223
rect 8152 1740 8186 1756
rect 8271 2132 8305 2148
rect 8271 1705 8305 1756
rect 8389 2132 8423 2184
rect 8389 1740 8423 1756
rect 8507 2132 8541 2148
rect 8507 1705 8541 1756
rect 8625 2132 8659 2184
rect 8862 1982 9132 2019
rect 8625 1740 8659 1756
rect 8744 1932 8778 1948
rect 7095 1666 8541 1705
rect 8744 1702 8778 1756
rect 8862 1932 8896 1982
rect 8862 1740 8896 1756
rect 8980 1932 9014 1948
rect 8980 1702 9014 1756
rect 9098 1932 9132 1982
rect 9098 1740 9132 1756
rect 8744 1663 9014 1702
rect 7622 1541 7656 1557
rect 8916 1548 8932 1582
rect 8966 1548 8982 1582
rect 7622 1491 7656 1507
rect 349 1382 365 1437
rect 425 1382 441 1437
rect 349 1369 441 1382
rect 1434 1438 1526 1451
rect 1434 1383 1450 1438
rect 1510 1383 1526 1438
rect 1434 1366 1526 1383
rect 3143 1438 3331 1453
rect 3143 1378 3265 1438
rect 3314 1378 3331 1438
rect 3143 1364 3331 1378
rect 3493 1437 3585 1454
rect 3493 1382 3509 1437
rect 3569 1382 3585 1437
rect 3493 1369 3585 1382
rect 4578 1438 4670 1451
rect 4578 1383 4594 1438
rect 4654 1383 4670 1438
rect 4578 1366 4670 1383
rect 6275 1442 6464 1454
rect 6275 1382 6397 1442
rect 6446 1382 6464 1442
rect 6275 1366 6464 1382
rect 6625 1441 6717 1458
rect 9420 1456 9519 2623
rect 10850 2402 11078 2420
rect 10850 2326 10866 2402
rect 11062 2326 11078 2402
rect 10850 2310 11078 2326
rect 10121 2185 10391 2224
rect 10121 2132 10155 2185
rect 9680 1983 9950 2022
rect 9680 1932 9714 1983
rect 9680 1740 9714 1756
rect 9798 1932 9832 1948
rect 9798 1705 9832 1756
rect 9916 1932 9950 1983
rect 9916 1740 9950 1756
rect 10034 1932 10068 1948
rect 10034 1705 10068 1756
rect 10121 1740 10155 1756
rect 10239 2132 10273 2148
rect 9798 1666 10068 1705
rect 10239 1705 10273 1756
rect 10357 2132 10391 2185
rect 10588 2184 10858 2223
rect 10357 1740 10391 1756
rect 10475 2132 10509 2148
rect 10475 1705 10509 1756
rect 10588 2132 10622 2184
rect 10588 1740 10622 1756
rect 10706 2132 10740 2148
rect 10706 1705 10740 1756
rect 10824 2132 10858 2184
rect 11060 2184 11330 2223
rect 10824 1740 10858 1756
rect 10942 2132 10976 2148
rect 10942 1705 10976 1756
rect 11060 2132 11094 2184
rect 11060 1740 11094 1756
rect 11178 2132 11212 2148
rect 11178 1705 11212 1756
rect 11296 2132 11330 2184
rect 11533 2184 11803 2223
rect 11296 1740 11330 1756
rect 11415 2132 11449 2148
rect 11415 1705 11449 1756
rect 11533 2132 11567 2184
rect 11533 1740 11567 1756
rect 11651 2132 11685 2148
rect 11651 1705 11685 1756
rect 11769 2132 11803 2184
rect 12006 1982 12276 2019
rect 11769 1740 11803 1756
rect 11888 1932 11922 1948
rect 10239 1666 11685 1705
rect 11888 1702 11922 1756
rect 12006 1932 12040 1982
rect 12006 1740 12040 1756
rect 12124 1932 12158 1948
rect 12124 1702 12158 1756
rect 12242 1932 12276 1982
rect 12242 1740 12276 1756
rect 11888 1663 12158 1702
rect 10766 1541 10800 1557
rect 12060 1548 12076 1582
rect 12110 1548 12126 1582
rect 10766 1491 10800 1507
rect 6625 1386 6641 1441
rect 6701 1386 6717 1441
rect 6625 1373 6717 1386
rect 7710 1442 7802 1455
rect 7710 1387 7726 1442
rect 7786 1387 7802 1442
rect 7710 1370 7802 1387
rect 9420 1442 9612 1456
rect 9420 1382 9541 1442
rect 9590 1382 9612 1442
rect 9420 1365 9612 1382
rect 9769 1441 9861 1458
rect 9769 1386 9785 1441
rect 9845 1386 9861 1441
rect 9769 1373 9861 1386
rect 10854 1442 10946 1455
rect 10854 1387 10870 1442
rect 10930 1387 10946 1442
rect 12620 1454 12719 2623
rect 14052 2398 14280 2416
rect 14052 2322 14068 2398
rect 14264 2322 14280 2398
rect 14052 2306 14280 2322
rect 13323 2181 13593 2220
rect 13323 2128 13357 2181
rect 12882 1979 13152 2018
rect 12882 1928 12916 1979
rect 12882 1736 12916 1752
rect 13000 1928 13034 1944
rect 13000 1701 13034 1752
rect 13118 1928 13152 1979
rect 13118 1736 13152 1752
rect 13236 1928 13270 1944
rect 13236 1701 13270 1752
rect 13323 1736 13357 1752
rect 13441 2128 13475 2144
rect 13000 1662 13270 1701
rect 13441 1701 13475 1752
rect 13559 2128 13593 2181
rect 13790 2180 14060 2219
rect 13559 1736 13593 1752
rect 13677 2128 13711 2144
rect 13677 1701 13711 1752
rect 13790 2128 13824 2180
rect 13790 1736 13824 1752
rect 13908 2128 13942 2144
rect 13908 1701 13942 1752
rect 14026 2128 14060 2180
rect 14262 2180 14532 2219
rect 14026 1736 14060 1752
rect 14144 2128 14178 2144
rect 14144 1701 14178 1752
rect 14262 2128 14296 2180
rect 14262 1736 14296 1752
rect 14380 2128 14414 2144
rect 14380 1701 14414 1752
rect 14498 2128 14532 2180
rect 14735 2180 15005 2219
rect 14498 1736 14532 1752
rect 14617 2128 14651 2144
rect 14617 1701 14651 1752
rect 14735 2128 14769 2180
rect 14735 1736 14769 1752
rect 14853 2128 14887 2144
rect 14853 1701 14887 1752
rect 14971 2128 15005 2180
rect 15208 1978 15478 2015
rect 14971 1736 15005 1752
rect 15090 1928 15124 1944
rect 13441 1662 14887 1701
rect 15090 1698 15124 1752
rect 15208 1928 15242 1978
rect 15208 1736 15242 1752
rect 15326 1928 15360 1944
rect 15326 1698 15360 1752
rect 15444 1928 15478 1978
rect 15444 1736 15478 1752
rect 15090 1659 15360 1698
rect 13968 1537 14002 1553
rect 15262 1544 15278 1578
rect 15312 1544 15328 1578
rect 13968 1487 14002 1503
rect 12620 1438 12811 1454
rect 12620 1399 12743 1438
rect 10854 1370 10946 1387
rect 12621 1378 12743 1399
rect 12792 1378 12811 1438
rect 9496 1364 9612 1365
rect 12621 1364 12811 1378
rect 12971 1437 13063 1454
rect 15765 1453 15864 2623
rect 17196 2398 17424 2416
rect 17196 2322 17212 2398
rect 17408 2322 17424 2398
rect 17196 2306 17424 2322
rect 16467 2181 16737 2220
rect 16467 2128 16501 2181
rect 16026 1979 16296 2018
rect 16026 1928 16060 1979
rect 16026 1736 16060 1752
rect 16144 1928 16178 1944
rect 16144 1701 16178 1752
rect 16262 1928 16296 1979
rect 16262 1736 16296 1752
rect 16380 1928 16414 1944
rect 16380 1701 16414 1752
rect 16467 1736 16501 1752
rect 16585 2128 16619 2144
rect 16144 1662 16414 1701
rect 16585 1701 16619 1752
rect 16703 2128 16737 2181
rect 16934 2180 17204 2219
rect 16703 1736 16737 1752
rect 16821 2128 16855 2144
rect 16821 1701 16855 1752
rect 16934 2128 16968 2180
rect 16934 1736 16968 1752
rect 17052 2128 17086 2144
rect 17052 1701 17086 1752
rect 17170 2128 17204 2180
rect 17406 2180 17676 2219
rect 17170 1736 17204 1752
rect 17288 2128 17322 2144
rect 17288 1701 17322 1752
rect 17406 2128 17440 2180
rect 17406 1736 17440 1752
rect 17524 2128 17558 2144
rect 17524 1701 17558 1752
rect 17642 2128 17676 2180
rect 17879 2180 18149 2219
rect 17642 1736 17676 1752
rect 17761 2128 17795 2144
rect 17761 1701 17795 1752
rect 17879 2128 17913 2180
rect 17879 1736 17913 1752
rect 17997 2128 18031 2144
rect 17997 1701 18031 1752
rect 18115 2128 18149 2180
rect 18352 1978 18622 2015
rect 18115 1736 18149 1752
rect 18234 1928 18268 1944
rect 16585 1662 18031 1701
rect 18234 1698 18268 1752
rect 18352 1928 18386 1978
rect 18352 1736 18386 1752
rect 18470 1928 18504 1944
rect 18470 1698 18504 1752
rect 18588 1928 18622 1978
rect 18588 1736 18622 1752
rect 18234 1659 18504 1698
rect 17112 1537 17146 1553
rect 18406 1544 18422 1578
rect 18456 1544 18472 1578
rect 17112 1487 17146 1503
rect 18897 1464 18996 2623
rect 20328 2402 20556 2420
rect 20328 2326 20344 2402
rect 20540 2326 20556 2402
rect 20328 2310 20556 2326
rect 19599 2185 19869 2224
rect 19599 2132 19633 2185
rect 19158 1983 19428 2022
rect 19158 1932 19192 1983
rect 19158 1740 19192 1756
rect 19276 1932 19310 1948
rect 19276 1705 19310 1756
rect 19394 1932 19428 1983
rect 19394 1740 19428 1756
rect 19512 1932 19546 1948
rect 19512 1705 19546 1756
rect 19599 1740 19633 1756
rect 19717 2132 19751 2148
rect 19276 1666 19546 1705
rect 19717 1705 19751 1756
rect 19835 2132 19869 2185
rect 20066 2184 20336 2223
rect 19835 1740 19869 1756
rect 19953 2132 19987 2148
rect 19953 1705 19987 1756
rect 20066 2132 20100 2184
rect 20066 1740 20100 1756
rect 20184 2132 20218 2148
rect 20184 1705 20218 1756
rect 20302 2132 20336 2184
rect 20538 2184 20808 2223
rect 20302 1740 20336 1756
rect 20420 2132 20454 2148
rect 20420 1705 20454 1756
rect 20538 2132 20572 2184
rect 20538 1740 20572 1756
rect 20656 2132 20690 2148
rect 20656 1705 20690 1756
rect 20774 2132 20808 2184
rect 21011 2184 21281 2223
rect 20774 1740 20808 1756
rect 20893 2132 20927 2148
rect 20893 1705 20927 1756
rect 21011 2132 21045 2184
rect 21011 1740 21045 1756
rect 21129 2132 21163 2148
rect 21129 1705 21163 1756
rect 21247 2132 21281 2184
rect 21484 1982 21754 2019
rect 21247 1740 21281 1756
rect 21366 1932 21400 1948
rect 19717 1666 21163 1705
rect 21366 1702 21400 1756
rect 21484 1932 21518 1982
rect 21484 1740 21518 1756
rect 21602 1932 21636 1948
rect 21602 1702 21636 1756
rect 21720 1932 21754 1982
rect 21720 1740 21754 1756
rect 21366 1663 21636 1702
rect 20244 1541 20278 1557
rect 21538 1548 21554 1582
rect 21588 1548 21604 1582
rect 20244 1491 20278 1507
rect 12971 1382 12987 1437
rect 13047 1382 13063 1437
rect 12971 1369 13063 1382
rect 14056 1438 14148 1451
rect 14056 1383 14072 1438
rect 14132 1383 14148 1438
rect 14056 1366 14148 1383
rect 15765 1438 15954 1453
rect 15765 1378 15887 1438
rect 15936 1378 15954 1438
rect 15765 1363 15954 1378
rect 16115 1437 16207 1454
rect 16115 1382 16131 1437
rect 16191 1382 16207 1437
rect 16115 1369 16207 1382
rect 17200 1438 17292 1451
rect 17200 1383 17216 1438
rect 17276 1383 17292 1438
rect 17200 1366 17292 1383
rect 18897 1442 19085 1464
rect 18897 1382 19019 1442
rect 19068 1382 19085 1442
rect 18897 1364 19085 1382
rect 19247 1441 19339 1458
rect 22040 1457 22139 2623
rect 30073 2590 30108 2792
rect 30146 2674 30162 2708
rect 30338 2674 30354 2708
rect 31371 2667 31387 2701
rect 31563 2667 31579 2701
rect 30073 2556 30162 2590
rect 30338 2556 30354 2590
rect 31270 2520 31286 2554
rect 31320 2520 31336 2554
rect 31371 2549 31387 2583
rect 31563 2549 31579 2583
rect 30146 2438 30162 2472
rect 30338 2438 30354 2472
rect 23472 2402 23700 2420
rect 23472 2326 23488 2402
rect 23684 2326 23700 2402
rect 30639 2365 30655 2399
rect 31031 2365 31047 2399
rect 31203 2369 31269 2385
rect 23472 2310 23700 2326
rect 29946 2308 29962 2342
rect 30338 2308 30354 2342
rect 31203 2335 31219 2369
rect 31253 2335 31269 2369
rect 31203 2318 31269 2335
rect 30984 2281 31129 2282
rect 30639 2247 30655 2281
rect 31031 2263 31129 2281
rect 31031 2247 31130 2263
rect 31371 2247 31387 2281
rect 30984 2246 31130 2247
rect 31763 2246 31865 2281
rect 22743 2185 23013 2224
rect 22743 2132 22777 2185
rect 22302 1983 22572 2022
rect 22302 1932 22336 1983
rect 22302 1740 22336 1756
rect 22420 1932 22454 1948
rect 22420 1705 22454 1756
rect 22538 1932 22572 1983
rect 22538 1740 22572 1756
rect 22656 1932 22690 1948
rect 22656 1705 22690 1756
rect 22743 1740 22777 1756
rect 22861 2132 22895 2148
rect 22420 1666 22690 1705
rect 22861 1705 22895 1756
rect 22979 2132 23013 2185
rect 23210 2184 23480 2223
rect 22979 1740 23013 1756
rect 23097 2132 23131 2148
rect 23097 1705 23131 1756
rect 23210 2132 23244 2184
rect 23210 1740 23244 1756
rect 23328 2132 23362 2148
rect 23328 1705 23362 1756
rect 23446 2132 23480 2184
rect 23682 2184 23952 2223
rect 23446 1740 23480 1756
rect 23564 2132 23598 2148
rect 23564 1705 23598 1756
rect 23682 2132 23716 2184
rect 23682 1740 23716 1756
rect 23800 2132 23834 2148
rect 23800 1705 23834 1756
rect 23918 2132 23952 2184
rect 24155 2184 24425 2223
rect 29946 2190 29962 2224
rect 30338 2190 30354 2224
rect 31089 2208 31130 2246
rect 23918 1740 23952 1756
rect 24037 2132 24071 2148
rect 24037 1705 24071 1756
rect 24155 2132 24189 2184
rect 24155 1740 24189 1756
rect 24273 2132 24307 2148
rect 24273 1705 24307 1756
rect 24391 2132 24425 2184
rect 31089 2174 31417 2208
rect 30639 2129 30655 2163
rect 31031 2129 31047 2163
rect 29671 2041 29763 2075
rect 29946 2072 29962 2106
rect 30338 2072 30354 2106
rect 31089 2047 31130 2174
rect 31371 2163 31417 2174
rect 31371 2129 31387 2163
rect 31763 2129 31779 2163
rect 31303 2103 31337 2119
rect 31303 2053 31337 2069
rect 30984 2045 31130 2047
rect 24628 1982 24898 2019
rect 24391 1740 24425 1756
rect 24510 1932 24544 1948
rect 22861 1666 24307 1705
rect 24510 1702 24544 1756
rect 24628 1932 24662 1982
rect 24628 1740 24662 1756
rect 24746 1932 24780 1948
rect 24746 1702 24780 1756
rect 24864 1932 24898 1982
rect 29671 1919 29691 2041
rect 29735 1989 29763 2041
rect 30639 2011 30655 2045
rect 31031 2011 31130 2045
rect 31371 2011 31387 2045
rect 31763 2011 31779 2045
rect 29745 1951 29763 1989
rect 29735 1919 29763 1951
rect 29671 1873 29763 1919
rect 29874 1954 29962 1988
rect 30338 1954 30354 1988
rect 24864 1740 24898 1756
rect 29874 1752 29909 1954
rect 30639 1893 30655 1927
rect 31031 1893 31047 1927
rect 29946 1836 29962 1870
rect 30338 1836 30354 1870
rect 31089 1809 31130 2011
rect 31302 1985 31336 2001
rect 31302 1935 31336 1951
rect 31371 1893 31387 1927
rect 31763 1893 31779 1927
rect 31830 1810 31865 2246
rect 31935 2091 32023 2107
rect 31935 2051 31951 2091
rect 31935 1959 31951 2001
rect 32007 1959 32023 2091
rect 31935 1943 32023 1959
rect 30639 1775 30655 1809
rect 31031 1775 31130 1809
rect 31371 1775 31387 1809
rect 31763 1775 31865 1810
rect 30985 1773 31130 1775
rect 29874 1718 29962 1752
rect 30338 1718 30354 1752
rect 24510 1663 24780 1702
rect 30639 1657 30655 1691
rect 31031 1657 31047 1691
rect 29946 1600 29962 1634
rect 30338 1600 30354 1634
rect 23388 1541 23422 1557
rect 24682 1548 24698 1582
rect 24732 1548 24748 1582
rect 23388 1491 23422 1507
rect 30146 1471 30162 1505
rect 30338 1471 30354 1505
rect 19247 1386 19263 1441
rect 19323 1386 19339 1441
rect 19247 1373 19339 1386
rect 20332 1442 20424 1455
rect 20332 1387 20348 1442
rect 20408 1387 20424 1442
rect 20332 1370 20424 1387
rect 22040 1442 22233 1457
rect 22040 1382 22163 1442
rect 22212 1382 22233 1442
rect 22040 1371 22233 1382
rect 22391 1441 22483 1458
rect 22391 1386 22407 1441
rect 22467 1386 22483 1441
rect 22391 1373 22483 1386
rect 23476 1442 23568 1455
rect 23476 1387 23492 1442
rect 23552 1387 23568 1442
rect 30517 1419 30551 1425
rect 22107 1368 22233 1371
rect 23476 1370 23568 1387
rect 30146 1353 30162 1387
rect 30338 1353 30354 1387
rect 30517 1359 30551 1365
rect 6393 1326 6450 1330
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 1700 1307 1734 1323
rect 1700 1257 1734 1273
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 4844 1307 4878 1323
rect 4844 1257 4878 1273
rect 6393 1266 6397 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 7976 1311 8010 1327
rect 7976 1261 8010 1277
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 11120 1311 11154 1327
rect 19015 1326 19072 1330
rect 11120 1261 11154 1277
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 14322 1307 14356 1323
rect 14322 1257 14356 1273
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 17466 1307 17500 1323
rect 17466 1257 17500 1273
rect 19015 1266 19019 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 20598 1311 20632 1327
rect 20598 1261 20632 1277
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 23742 1311 23776 1327
rect 23742 1261 23776 1277
rect 30146 1235 30162 1269
rect 30338 1235 30354 1269
rect 31089 1187 31130 1773
rect 31203 1721 31269 1738
rect 31203 1687 31219 1721
rect 31253 1687 31269 1721
rect 31203 1671 31269 1687
rect 31271 1397 31287 1431
rect 31321 1397 31337 1431
rect 31371 1369 31387 1403
rect 31563 1369 31579 1403
rect 31371 1251 31387 1285
rect 31563 1251 31579 1285
rect 1316 1153 1408 1166
rect 1316 1098 1332 1153
rect 1392 1098 1408 1153
rect 1316 1081 1408 1098
rect 4460 1153 4552 1166
rect 4460 1098 4476 1153
rect 4536 1098 4552 1153
rect 4460 1081 4552 1098
rect 7592 1157 7684 1170
rect 7592 1102 7608 1157
rect 7668 1102 7684 1157
rect 7592 1085 7684 1102
rect 10736 1157 10828 1170
rect 10736 1102 10752 1157
rect 10812 1102 10828 1157
rect 10736 1085 10828 1102
rect 13938 1153 14030 1166
rect 13938 1098 13954 1153
rect 14014 1098 14030 1153
rect 13938 1081 14030 1098
rect 17082 1153 17174 1166
rect 17082 1098 17098 1153
rect 17158 1098 17174 1153
rect 17082 1081 17174 1098
rect 20214 1157 20306 1170
rect 20214 1102 20230 1157
rect 20290 1102 20306 1157
rect 20214 1085 20306 1102
rect 23358 1157 23450 1170
rect 23358 1102 23374 1157
rect 23434 1102 23450 1157
rect 30146 1117 30162 1151
rect 30338 1117 30354 1151
rect 23358 1085 23450 1102
rect 1581 917 1615 933
rect 1581 867 1615 883
rect 4725 917 4759 933
rect 4725 867 4759 883
rect 7857 921 7891 937
rect 7857 871 7891 887
rect 11001 921 11035 937
rect 11001 871 11035 887
rect 14203 917 14237 933
rect 14203 867 14237 883
rect 17347 917 17381 933
rect 17347 867 17381 883
rect 20479 921 20513 937
rect 20479 871 20513 887
rect 23623 921 23657 937
rect 23623 871 23657 887
rect 32528 921 32614 933
rect 32528 866 32534 921
rect 32604 866 32614 921
rect 1094 795 1128 811
rect 1094 603 1128 619
rect 1212 807 1246 811
rect 1286 807 1320 811
rect 1212 795 1320 807
rect 1246 619 1286 795
rect 1212 607 1286 619
rect 1212 603 1246 607
rect 1286 403 1320 419
rect 1404 795 1438 811
rect 1404 403 1438 419
rect 1522 795 1556 811
rect 1522 403 1556 419
rect 1640 795 1674 811
rect 1640 403 1674 419
rect 1758 807 1792 811
rect 1836 807 1870 811
rect 1758 795 1870 807
rect 1792 619 1836 795
rect 1792 607 1870 619
rect 1836 603 1870 607
rect 1954 795 1988 811
rect 1954 603 1988 619
rect 4238 795 4272 811
rect 4238 603 4272 619
rect 4356 807 4390 811
rect 4430 807 4464 811
rect 4356 795 4464 807
rect 4390 619 4430 795
rect 4356 607 4430 619
rect 4356 603 4390 607
rect 1758 403 1792 419
rect 4430 403 4464 419
rect 4548 795 4582 811
rect 4548 403 4582 419
rect 4666 795 4700 811
rect 4666 403 4700 419
rect 4784 795 4818 811
rect 4784 403 4818 419
rect 4902 807 4936 811
rect 4980 807 5014 811
rect 4902 795 5014 807
rect 4936 619 4980 795
rect 4936 607 5014 619
rect 4980 603 5014 607
rect 5098 795 5132 811
rect 5098 603 5132 619
rect 7370 799 7404 815
rect 7370 607 7404 623
rect 7488 811 7522 815
rect 7562 811 7596 815
rect 7488 799 7596 811
rect 7522 623 7562 799
rect 7488 611 7562 623
rect 7488 607 7522 611
rect 4902 403 4936 419
rect 7562 407 7596 423
rect 7680 799 7714 815
rect 7680 407 7714 423
rect 7798 799 7832 815
rect 7798 407 7832 423
rect 7916 799 7950 815
rect 7916 407 7950 423
rect 8034 811 8068 815
rect 8112 811 8146 815
rect 8034 799 8146 811
rect 8068 623 8112 799
rect 8068 611 8146 623
rect 8112 607 8146 611
rect 8230 799 8264 815
rect 8230 607 8264 623
rect 10514 799 10548 815
rect 10514 607 10548 623
rect 10632 811 10666 815
rect 10706 811 10740 815
rect 10632 799 10740 811
rect 10666 623 10706 799
rect 10632 611 10706 623
rect 10632 607 10666 611
rect 8034 407 8068 423
rect 10706 407 10740 423
rect 10824 799 10858 815
rect 10824 407 10858 423
rect 10942 799 10976 815
rect 10942 407 10976 423
rect 11060 799 11094 815
rect 11060 407 11094 423
rect 11178 811 11212 815
rect 11256 811 11290 815
rect 11178 799 11290 811
rect 11212 623 11256 799
rect 11212 611 11290 623
rect 11256 607 11290 611
rect 11374 799 11408 815
rect 11374 607 11408 623
rect 13716 795 13750 811
rect 13716 603 13750 619
rect 13834 807 13868 811
rect 13908 807 13942 811
rect 13834 795 13942 807
rect 13868 619 13908 795
rect 13834 607 13908 619
rect 13834 603 13868 607
rect 11178 407 11212 423
rect 13908 403 13942 419
rect 14026 795 14060 811
rect 14026 403 14060 419
rect 14144 795 14178 811
rect 14144 403 14178 419
rect 14262 795 14296 811
rect 14262 403 14296 419
rect 14380 807 14414 811
rect 14458 807 14492 811
rect 14380 795 14492 807
rect 14414 619 14458 795
rect 14414 607 14492 619
rect 14458 603 14492 607
rect 14576 795 14610 811
rect 14576 603 14610 619
rect 16860 795 16894 811
rect 16860 603 16894 619
rect 16978 807 17012 811
rect 17052 807 17086 811
rect 16978 795 17086 807
rect 17012 619 17052 795
rect 16978 607 17052 619
rect 16978 603 17012 607
rect 14380 403 14414 419
rect 17052 403 17086 419
rect 17170 795 17204 811
rect 17170 403 17204 419
rect 17288 795 17322 811
rect 17288 403 17322 419
rect 17406 795 17440 811
rect 17406 403 17440 419
rect 17524 807 17558 811
rect 17602 807 17636 811
rect 17524 795 17636 807
rect 17558 619 17602 795
rect 17558 607 17636 619
rect 17602 603 17636 607
rect 17720 795 17754 811
rect 17720 603 17754 619
rect 19992 799 20026 815
rect 19992 607 20026 623
rect 20110 811 20144 815
rect 20184 811 20218 815
rect 20110 799 20218 811
rect 20144 623 20184 799
rect 20110 611 20184 623
rect 20110 607 20144 611
rect 17524 403 17558 419
rect 20184 407 20218 423
rect 20302 799 20336 815
rect 20302 407 20336 423
rect 20420 799 20454 815
rect 20420 407 20454 423
rect 20538 799 20572 815
rect 20538 407 20572 423
rect 20656 811 20690 815
rect 20734 811 20768 815
rect 20656 799 20768 811
rect 20690 623 20734 799
rect 20690 611 20768 623
rect 20734 607 20768 611
rect 20852 799 20886 815
rect 20852 607 20886 623
rect 23136 799 23170 815
rect 23136 607 23170 623
rect 23254 811 23288 815
rect 23328 811 23362 815
rect 23254 799 23362 811
rect 23288 623 23328 799
rect 23254 611 23328 623
rect 23254 607 23288 611
rect 20656 407 20690 423
rect 23328 407 23362 423
rect 23446 799 23480 815
rect 23446 407 23480 423
rect 23564 799 23598 815
rect 23564 407 23598 423
rect 23682 799 23716 815
rect 23682 407 23716 423
rect 23800 811 23834 815
rect 23878 811 23912 815
rect 23800 799 23912 811
rect 23834 623 23878 799
rect 23834 611 23912 623
rect 23878 607 23912 611
rect 23996 799 24030 815
rect 23996 607 24030 623
rect 30075 723 30164 757
rect 30340 723 30356 757
rect 30075 521 30110 723
rect 30148 605 30164 639
rect 30340 605 30356 639
rect 31373 598 31389 632
rect 31565 598 31581 632
rect 30075 487 30164 521
rect 30340 487 30356 521
rect 31272 451 31288 485
rect 31322 451 31338 485
rect 31373 480 31389 514
rect 31565 480 31581 514
rect 23800 407 23834 423
rect 30148 369 30164 403
rect 30340 369 30356 403
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 30641 296 30657 330
rect 31033 296 31049 330
rect 31205 300 31271 316
rect 29948 239 29964 273
rect 30340 239 30356 273
rect 31205 266 31221 300
rect 31255 266 31271 300
rect 31205 249 31271 266
rect 30986 212 31131 213
rect 30641 178 30657 212
rect 31033 194 31131 212
rect 31033 178 31132 194
rect 31373 178 31389 212
rect 30986 177 31132 178
rect 31765 177 31867 212
rect 7764 170 7900 174
rect 1488 166 1624 170
rect 1488 152 1526 166
rect 1584 152 1624 166
rect 1488 106 1504 152
rect 1608 106 1624 152
rect 1488 84 1624 106
rect 4632 166 4768 170
rect 4632 152 4670 166
rect 4728 152 4768 166
rect 4632 106 4648 152
rect 4752 106 4768 152
rect 4632 84 4768 106
rect 7764 156 7802 170
rect 7860 156 7900 170
rect 7764 110 7780 156
rect 7884 110 7900 156
rect 7764 88 7900 110
rect 10908 170 11044 174
rect 20386 170 20522 174
rect 10908 156 10946 170
rect 11004 156 11044 170
rect 10908 110 10924 156
rect 11028 110 11044 156
rect 10908 88 11044 110
rect 14110 166 14246 170
rect 14110 152 14148 166
rect 14206 152 14246 166
rect 14110 106 14126 152
rect 14230 106 14246 152
rect 14110 84 14246 106
rect 17254 166 17390 170
rect 17254 152 17292 166
rect 17350 152 17390 166
rect 17254 106 17270 152
rect 17374 106 17390 152
rect 17254 84 17390 106
rect 20386 156 20424 170
rect 20482 156 20522 170
rect 20386 110 20402 156
rect 20506 110 20522 156
rect 20386 88 20522 110
rect 23530 170 23666 174
rect 23530 156 23568 170
rect 23626 156 23666 170
rect 23530 110 23546 156
rect 23650 110 23666 156
rect 29948 121 29964 155
rect 30340 121 30356 155
rect 31091 139 31132 177
rect 23530 88 23666 110
rect 31091 105 31419 139
rect 30641 60 30657 94
rect 31033 60 31049 94
rect 29673 -28 29765 6
rect 29948 3 29964 37
rect 30340 3 30356 37
rect 31091 -22 31132 105
rect 31373 94 31419 105
rect 31373 60 31389 94
rect 31765 60 31781 94
rect 31305 34 31339 50
rect 31305 -16 31339 0
rect 30986 -24 31132 -22
rect 29673 -150 29693 -28
rect 29737 -80 29765 -28
rect 30641 -58 30657 -24
rect 31033 -58 31132 -24
rect 31373 -58 31389 -24
rect 31765 -58 31781 -24
rect 29747 -118 29765 -80
rect 29737 -150 29765 -118
rect 29673 -196 29765 -150
rect 29876 -115 29964 -81
rect 30340 -115 30356 -81
rect 29876 -317 29911 -115
rect 30641 -176 30657 -142
rect 31033 -176 31049 -142
rect 29948 -233 29964 -199
rect 30340 -233 30356 -199
rect 31091 -260 31132 -58
rect 31304 -84 31338 -68
rect 31304 -134 31338 -118
rect 31373 -176 31389 -142
rect 31765 -176 31781 -142
rect 31832 -259 31867 177
rect 31937 22 32025 38
rect 31937 -18 31953 22
rect 31937 -110 31953 -68
rect 32009 -110 32025 22
rect 31937 -126 32025 -110
rect 30641 -294 30657 -260
rect 31033 -294 31132 -260
rect 31373 -294 31389 -260
rect 31765 -294 31867 -259
rect 30987 -296 31132 -294
rect 29876 -351 29964 -317
rect 30340 -351 30356 -317
rect 30641 -412 30657 -378
rect 31033 -412 31049 -378
rect 29948 -469 29964 -435
rect 30340 -469 30356 -435
rect 30148 -598 30164 -564
rect 30340 -598 30356 -564
rect 30519 -650 30553 -644
rect 30148 -716 30164 -682
rect 30340 -716 30356 -682
rect 30519 -710 30553 -704
rect 30148 -834 30164 -800
rect 30340 -834 30356 -800
rect 31091 -882 31132 -296
rect 31205 -348 31271 -331
rect 31205 -382 31221 -348
rect 31255 -382 31271 -348
rect 31205 -398 31271 -382
rect 31273 -672 31289 -638
rect 31323 -672 31339 -638
rect 31373 -700 31389 -666
rect 31565 -700 31581 -666
rect 31373 -818 31389 -784
rect 31565 -818 31581 -784
rect 30148 -952 30164 -918
rect 30340 -952 30356 -918
rect -2374 -995 -1865 -991
rect -2442 -1067 -1865 -995
rect -2442 -1190 22177 -1067
rect 30 -2440 135 -1190
rect 1462 -1494 1690 -1476
rect 1462 -1570 1478 -1494
rect 1674 -1570 1690 -1494
rect 1462 -1586 1690 -1570
rect 733 -1711 1003 -1672
rect 733 -1764 767 -1711
rect 292 -1913 562 -1874
rect 292 -1964 326 -1913
rect 292 -2156 326 -2140
rect 410 -1964 444 -1948
rect 410 -2191 444 -2140
rect 528 -1964 562 -1913
rect 528 -2156 562 -2140
rect 646 -1964 680 -1948
rect 646 -2191 680 -2140
rect 733 -2156 767 -2140
rect 851 -1764 885 -1748
rect 410 -2230 680 -2191
rect 851 -2191 885 -2140
rect 969 -1764 1003 -1711
rect 1200 -1712 1470 -1673
rect 969 -2156 1003 -2140
rect 1087 -1764 1121 -1748
rect 1087 -2191 1121 -2140
rect 1200 -1764 1234 -1712
rect 1200 -2156 1234 -2140
rect 1318 -1764 1352 -1748
rect 1318 -2191 1352 -2140
rect 1436 -1764 1470 -1712
rect 1672 -1712 1942 -1673
rect 1436 -2156 1470 -2140
rect 1554 -1764 1588 -1748
rect 1554 -2191 1588 -2140
rect 1672 -1764 1706 -1712
rect 1672 -2156 1706 -2140
rect 1790 -1764 1824 -1748
rect 1790 -2191 1824 -2140
rect 1908 -1764 1942 -1712
rect 2145 -1712 2415 -1673
rect 1908 -2156 1942 -2140
rect 2027 -1764 2061 -1748
rect 2027 -2191 2061 -2140
rect 2145 -1764 2179 -1712
rect 2145 -2156 2179 -2140
rect 2263 -1764 2297 -1748
rect 2263 -2191 2297 -2140
rect 2381 -1764 2415 -1712
rect 2618 -1914 2888 -1877
rect 2381 -2156 2415 -2140
rect 2500 -1964 2534 -1948
rect 851 -2230 2297 -2191
rect 2500 -2194 2534 -2140
rect 2618 -1964 2652 -1914
rect 2618 -2156 2652 -2140
rect 2736 -1964 2770 -1948
rect 2736 -2194 2770 -2140
rect 2854 -1964 2888 -1914
rect 2854 -2156 2888 -2140
rect 2500 -2233 2770 -2194
rect 1378 -2355 1412 -2339
rect 2672 -2348 2688 -2314
rect 2722 -2348 2738 -2314
rect 1378 -2405 1412 -2389
rect 3174 -2437 3279 -1190
rect 4606 -1494 4834 -1476
rect 4606 -1570 4622 -1494
rect 4818 -1570 4834 -1494
rect 4606 -1586 4834 -1570
rect 3877 -1711 4147 -1672
rect 3877 -1764 3911 -1711
rect 3436 -1913 3706 -1874
rect 3436 -1964 3470 -1913
rect 3436 -2156 3470 -2140
rect 3554 -1964 3588 -1948
rect 3554 -2191 3588 -2140
rect 3672 -1964 3706 -1913
rect 3672 -2156 3706 -2140
rect 3790 -1964 3824 -1948
rect 3790 -2191 3824 -2140
rect 3877 -2156 3911 -2140
rect 3995 -1764 4029 -1748
rect 3554 -2230 3824 -2191
rect 3995 -2191 4029 -2140
rect 4113 -1764 4147 -1711
rect 4344 -1712 4614 -1673
rect 4113 -2156 4147 -2140
rect 4231 -1764 4265 -1748
rect 4231 -2191 4265 -2140
rect 4344 -1764 4378 -1712
rect 4344 -2156 4378 -2140
rect 4462 -1764 4496 -1748
rect 4462 -2191 4496 -2140
rect 4580 -1764 4614 -1712
rect 4816 -1712 5086 -1673
rect 4580 -2156 4614 -2140
rect 4698 -1764 4732 -1748
rect 4698 -2191 4732 -2140
rect 4816 -1764 4850 -1712
rect 4816 -2156 4850 -2140
rect 4934 -1764 4968 -1748
rect 4934 -2191 4968 -2140
rect 5052 -1764 5086 -1712
rect 5289 -1712 5559 -1673
rect 5052 -2156 5086 -2140
rect 5171 -1764 5205 -1748
rect 5171 -2191 5205 -2140
rect 5289 -1764 5323 -1712
rect 5289 -2156 5323 -2140
rect 5407 -1764 5441 -1748
rect 5407 -2191 5441 -2140
rect 5525 -1764 5559 -1712
rect 5762 -1914 6032 -1877
rect 5525 -2156 5559 -2140
rect 5644 -1964 5678 -1948
rect 3995 -2230 5441 -2191
rect 5644 -2194 5678 -2140
rect 5762 -1964 5796 -1914
rect 5762 -2156 5796 -2140
rect 5880 -1964 5914 -1948
rect 5880 -2194 5914 -2140
rect 5998 -1964 6032 -1914
rect 5998 -2156 6032 -2140
rect 5644 -2233 5914 -2194
rect 4522 -2355 4556 -2339
rect 5816 -2348 5832 -2314
rect 5866 -2348 5882 -2314
rect 4522 -2405 4556 -2389
rect 6308 -2429 6413 -1190
rect 7738 -1490 7966 -1472
rect 7738 -1566 7754 -1490
rect 7950 -1566 7966 -1490
rect 7738 -1582 7966 -1566
rect 7009 -1707 7279 -1668
rect 7009 -1760 7043 -1707
rect 6568 -1909 6838 -1870
rect 6568 -1960 6602 -1909
rect 6568 -2152 6602 -2136
rect 6686 -1960 6720 -1944
rect 6686 -2187 6720 -2136
rect 6804 -1960 6838 -1909
rect 6804 -2152 6838 -2136
rect 6922 -1960 6956 -1944
rect 6922 -2187 6956 -2136
rect 7009 -2152 7043 -2136
rect 7127 -1760 7161 -1744
rect 6686 -2226 6956 -2187
rect 7127 -2187 7161 -2136
rect 7245 -1760 7279 -1707
rect 7476 -1708 7746 -1669
rect 7245 -2152 7279 -2136
rect 7363 -1760 7397 -1744
rect 7363 -2187 7397 -2136
rect 7476 -1760 7510 -1708
rect 7476 -2152 7510 -2136
rect 7594 -1760 7628 -1744
rect 7594 -2187 7628 -2136
rect 7712 -1760 7746 -1708
rect 7948 -1708 8218 -1669
rect 7712 -2152 7746 -2136
rect 7830 -1760 7864 -1744
rect 7830 -2187 7864 -2136
rect 7948 -1760 7982 -1708
rect 7948 -2152 7982 -2136
rect 8066 -1760 8100 -1744
rect 8066 -2187 8100 -2136
rect 8184 -1760 8218 -1708
rect 8421 -1708 8691 -1669
rect 8184 -2152 8218 -2136
rect 8303 -1760 8337 -1744
rect 8303 -2187 8337 -2136
rect 8421 -1760 8455 -1708
rect 8421 -2152 8455 -2136
rect 8539 -1760 8573 -1744
rect 8539 -2187 8573 -2136
rect 8657 -1760 8691 -1708
rect 8894 -1910 9164 -1873
rect 8657 -2152 8691 -2136
rect 8776 -1960 8810 -1944
rect 7127 -2226 8573 -2187
rect 8776 -2190 8810 -2136
rect 8894 -1960 8928 -1910
rect 8894 -2152 8928 -2136
rect 9012 -1960 9046 -1944
rect 9012 -2190 9046 -2136
rect 9130 -1960 9164 -1910
rect 9130 -2152 9164 -2136
rect 8776 -2229 9046 -2190
rect 7654 -2351 7688 -2335
rect 8948 -2344 8964 -2310
rect 8998 -2344 9014 -2310
rect 7654 -2401 7688 -2385
rect 30 -2454 220 -2440
rect 30 -2514 153 -2454
rect 202 -2514 220 -2454
rect 30 -2532 220 -2514
rect 381 -2455 473 -2438
rect 381 -2510 397 -2455
rect 457 -2510 473 -2455
rect 381 -2523 473 -2510
rect 1466 -2454 1558 -2441
rect 1466 -2509 1482 -2454
rect 1542 -2509 1558 -2454
rect 1466 -2526 1558 -2509
rect 3174 -2454 3379 -2437
rect 3174 -2514 3297 -2454
rect 3346 -2514 3379 -2454
rect 3174 -2532 3379 -2514
rect 3525 -2455 3617 -2438
rect 3525 -2510 3541 -2455
rect 3601 -2510 3617 -2455
rect 3525 -2523 3617 -2510
rect 4610 -2454 4702 -2441
rect 4610 -2509 4626 -2454
rect 4686 -2509 4702 -2454
rect 4610 -2526 4702 -2509
rect 6308 -2450 6503 -2429
rect 9451 -2432 9556 -1190
rect 10882 -1490 11110 -1472
rect 10882 -1566 10898 -1490
rect 11094 -1566 11110 -1490
rect 10882 -1582 11110 -1566
rect 10153 -1707 10423 -1668
rect 10153 -1760 10187 -1707
rect 9712 -1909 9982 -1870
rect 9712 -1960 9746 -1909
rect 9712 -2152 9746 -2136
rect 9830 -1960 9864 -1944
rect 9830 -2187 9864 -2136
rect 9948 -1960 9982 -1909
rect 9948 -2152 9982 -2136
rect 10066 -1960 10100 -1944
rect 10066 -2187 10100 -2136
rect 10153 -2152 10187 -2136
rect 10271 -1760 10305 -1744
rect 9830 -2226 10100 -2187
rect 10271 -2187 10305 -2136
rect 10389 -1760 10423 -1707
rect 10620 -1708 10890 -1669
rect 10389 -2152 10423 -2136
rect 10507 -1760 10541 -1744
rect 10507 -2187 10541 -2136
rect 10620 -1760 10654 -1708
rect 10620 -2152 10654 -2136
rect 10738 -1760 10772 -1744
rect 10738 -2187 10772 -2136
rect 10856 -1760 10890 -1708
rect 11092 -1708 11362 -1669
rect 10856 -2152 10890 -2136
rect 10974 -1760 11008 -1744
rect 10974 -2187 11008 -2136
rect 11092 -1760 11126 -1708
rect 11092 -2152 11126 -2136
rect 11210 -1760 11244 -1744
rect 11210 -2187 11244 -2136
rect 11328 -1760 11362 -1708
rect 11565 -1708 11835 -1669
rect 11328 -2152 11362 -2136
rect 11447 -1760 11481 -1744
rect 11447 -2187 11481 -2136
rect 11565 -1760 11599 -1708
rect 11565 -2152 11599 -2136
rect 11683 -1760 11717 -1744
rect 11683 -2187 11717 -2136
rect 11801 -1760 11835 -1708
rect 12038 -1910 12308 -1873
rect 11801 -2152 11835 -2136
rect 11920 -1960 11954 -1944
rect 10271 -2226 11717 -2187
rect 11920 -2190 11954 -2136
rect 12038 -1960 12072 -1910
rect 12038 -2152 12072 -2136
rect 12156 -1960 12190 -1944
rect 12156 -2190 12190 -2136
rect 12274 -1960 12308 -1910
rect 12274 -2152 12308 -2136
rect 11920 -2229 12190 -2190
rect 10798 -2351 10832 -2335
rect 12092 -2344 12108 -2310
rect 12142 -2344 12158 -2310
rect 10798 -2401 10832 -2385
rect 12652 -2432 12757 -1190
rect 14084 -1494 14312 -1476
rect 14084 -1570 14100 -1494
rect 14296 -1570 14312 -1494
rect 14084 -1586 14312 -1570
rect 13355 -1711 13625 -1672
rect 13355 -1764 13389 -1711
rect 12914 -1913 13184 -1874
rect 12914 -1964 12948 -1913
rect 12914 -2156 12948 -2140
rect 13032 -1964 13066 -1948
rect 13032 -2191 13066 -2140
rect 13150 -1964 13184 -1913
rect 13150 -2156 13184 -2140
rect 13268 -1964 13302 -1948
rect 13268 -2191 13302 -2140
rect 13355 -2156 13389 -2140
rect 13473 -1764 13507 -1748
rect 13032 -2230 13302 -2191
rect 13473 -2191 13507 -2140
rect 13591 -1764 13625 -1711
rect 13822 -1712 14092 -1673
rect 13591 -2156 13625 -2140
rect 13709 -1764 13743 -1748
rect 13709 -2191 13743 -2140
rect 13822 -1764 13856 -1712
rect 13822 -2156 13856 -2140
rect 13940 -1764 13974 -1748
rect 13940 -2191 13974 -2140
rect 14058 -1764 14092 -1712
rect 14294 -1712 14564 -1673
rect 14058 -2156 14092 -2140
rect 14176 -1764 14210 -1748
rect 14176 -2191 14210 -2140
rect 14294 -1764 14328 -1712
rect 14294 -2156 14328 -2140
rect 14412 -1764 14446 -1748
rect 14412 -2191 14446 -2140
rect 14530 -1764 14564 -1712
rect 14767 -1712 15037 -1673
rect 14530 -2156 14564 -2140
rect 14649 -1764 14683 -1748
rect 14649 -2191 14683 -2140
rect 14767 -1764 14801 -1712
rect 14767 -2156 14801 -2140
rect 14885 -1764 14919 -1748
rect 14885 -2191 14919 -2140
rect 15003 -1764 15037 -1712
rect 15240 -1914 15510 -1877
rect 15003 -2156 15037 -2140
rect 15122 -1964 15156 -1948
rect 13473 -2230 14919 -2191
rect 15122 -2194 15156 -2140
rect 15240 -1964 15274 -1914
rect 15240 -2156 15274 -2140
rect 15358 -1964 15392 -1948
rect 15358 -2194 15392 -2140
rect 15476 -1964 15510 -1914
rect 15476 -2156 15510 -2140
rect 15122 -2233 15392 -2194
rect 14000 -2355 14034 -2339
rect 15294 -2348 15310 -2314
rect 15344 -2348 15360 -2314
rect 14000 -2405 14034 -2389
rect 15798 -2431 15903 -1190
rect 17228 -1494 17456 -1476
rect 17228 -1570 17244 -1494
rect 17440 -1570 17456 -1494
rect 17228 -1586 17456 -1570
rect 16499 -1711 16769 -1672
rect 16499 -1764 16533 -1711
rect 16058 -1913 16328 -1874
rect 16058 -1964 16092 -1913
rect 16058 -2156 16092 -2140
rect 16176 -1964 16210 -1948
rect 16176 -2191 16210 -2140
rect 16294 -1964 16328 -1913
rect 16294 -2156 16328 -2140
rect 16412 -1964 16446 -1948
rect 16412 -2191 16446 -2140
rect 16499 -2156 16533 -2140
rect 16617 -1764 16651 -1748
rect 16176 -2230 16446 -2191
rect 16617 -2191 16651 -2140
rect 16735 -1764 16769 -1711
rect 16966 -1712 17236 -1673
rect 16735 -2156 16769 -2140
rect 16853 -1764 16887 -1748
rect 16853 -2191 16887 -2140
rect 16966 -1764 17000 -1712
rect 16966 -2156 17000 -2140
rect 17084 -1764 17118 -1748
rect 17084 -2191 17118 -2140
rect 17202 -1764 17236 -1712
rect 17438 -1712 17708 -1673
rect 17202 -2156 17236 -2140
rect 17320 -1764 17354 -1748
rect 17320 -2191 17354 -2140
rect 17438 -1764 17472 -1712
rect 17438 -2156 17472 -2140
rect 17556 -1764 17590 -1748
rect 17556 -2191 17590 -2140
rect 17674 -1764 17708 -1712
rect 17911 -1712 18181 -1673
rect 17674 -2156 17708 -2140
rect 17793 -1764 17827 -1748
rect 17793 -2191 17827 -2140
rect 17911 -1764 17945 -1712
rect 17911 -2156 17945 -2140
rect 18029 -1764 18063 -1748
rect 18029 -2191 18063 -2140
rect 18147 -1764 18181 -1712
rect 18384 -1914 18654 -1877
rect 18147 -2156 18181 -2140
rect 18266 -1964 18300 -1948
rect 16617 -2230 18063 -2191
rect 18266 -2194 18300 -2140
rect 18384 -1964 18418 -1914
rect 18384 -2156 18418 -2140
rect 18502 -1964 18536 -1948
rect 18502 -2194 18536 -2140
rect 18620 -1964 18654 -1914
rect 18620 -2156 18654 -2140
rect 18266 -2233 18536 -2194
rect 17144 -2355 17178 -2339
rect 18438 -2348 18454 -2314
rect 18488 -2348 18504 -2314
rect 17144 -2405 17178 -2389
rect 18930 -2428 19035 -1190
rect 20360 -1490 20588 -1472
rect 20360 -1566 20376 -1490
rect 20572 -1566 20588 -1490
rect 20360 -1582 20588 -1566
rect 19631 -1707 19901 -1668
rect 19631 -1760 19665 -1707
rect 19190 -1909 19460 -1870
rect 19190 -1960 19224 -1909
rect 19190 -2152 19224 -2136
rect 19308 -1960 19342 -1944
rect 19308 -2187 19342 -2136
rect 19426 -1960 19460 -1909
rect 19426 -2152 19460 -2136
rect 19544 -1960 19578 -1944
rect 19544 -2187 19578 -2136
rect 19631 -2152 19665 -2136
rect 19749 -1760 19783 -1744
rect 19308 -2226 19578 -2187
rect 19749 -2187 19783 -2136
rect 19867 -1760 19901 -1707
rect 20098 -1708 20368 -1669
rect 19867 -2152 19901 -2136
rect 19985 -1760 20019 -1744
rect 19985 -2187 20019 -2136
rect 20098 -1760 20132 -1708
rect 20098 -2152 20132 -2136
rect 20216 -1760 20250 -1744
rect 20216 -2187 20250 -2136
rect 20334 -1760 20368 -1708
rect 20570 -1708 20840 -1669
rect 20334 -2152 20368 -2136
rect 20452 -1760 20486 -1744
rect 20452 -2187 20486 -2136
rect 20570 -1760 20604 -1708
rect 20570 -2152 20604 -2136
rect 20688 -1760 20722 -1744
rect 20688 -2187 20722 -2136
rect 20806 -1760 20840 -1708
rect 21043 -1708 21313 -1669
rect 20806 -2152 20840 -2136
rect 20925 -1760 20959 -1744
rect 20925 -2187 20959 -2136
rect 21043 -1760 21077 -1708
rect 21043 -2152 21077 -2136
rect 21161 -1760 21195 -1744
rect 21161 -2187 21195 -2136
rect 21279 -1760 21313 -1708
rect 21516 -1910 21786 -1873
rect 21279 -2152 21313 -2136
rect 21398 -1960 21432 -1944
rect 19749 -2226 21195 -2187
rect 21398 -2190 21432 -2136
rect 21516 -1960 21550 -1910
rect 21516 -2152 21550 -2136
rect 21634 -1960 21668 -1944
rect 21634 -2190 21668 -2136
rect 21752 -1960 21786 -1910
rect 21752 -2152 21786 -2136
rect 21398 -2229 21668 -2190
rect 20276 -2351 20310 -2335
rect 21570 -2344 21586 -2310
rect 21620 -2344 21636 -2310
rect 20276 -2401 20310 -2385
rect 6308 -2510 6429 -2450
rect 6478 -2510 6503 -2450
rect 6308 -2525 6503 -2510
rect 6657 -2451 6749 -2434
rect 6657 -2506 6673 -2451
rect 6733 -2506 6749 -2451
rect 6657 -2519 6749 -2506
rect 7742 -2450 7834 -2437
rect 7742 -2505 7758 -2450
rect 7818 -2505 7834 -2450
rect 7742 -2522 7834 -2505
rect 9451 -2450 9644 -2432
rect 9451 -2510 9573 -2450
rect 9622 -2510 9644 -2450
rect 9451 -2528 9644 -2510
rect 9801 -2451 9893 -2434
rect 9801 -2506 9817 -2451
rect 9877 -2506 9893 -2451
rect 9801 -2519 9893 -2506
rect 10886 -2450 10978 -2437
rect 10886 -2505 10902 -2450
rect 10962 -2505 10978 -2450
rect 10886 -2522 10978 -2505
rect 12652 -2454 12850 -2432
rect 12652 -2514 12775 -2454
rect 12824 -2514 12850 -2454
rect 12652 -2531 12850 -2514
rect 13003 -2455 13095 -2438
rect 13003 -2510 13019 -2455
rect 13079 -2510 13095 -2455
rect 13003 -2523 13095 -2510
rect 14088 -2454 14180 -2441
rect 14088 -2509 14104 -2454
rect 14164 -2509 14180 -2454
rect 14088 -2526 14180 -2509
rect 15798 -2454 16000 -2431
rect 15798 -2514 15919 -2454
rect 15968 -2514 16000 -2454
rect 12699 -2532 12850 -2531
rect 15798 -2531 16000 -2514
rect 16147 -2455 16239 -2438
rect 16147 -2510 16163 -2455
rect 16223 -2510 16239 -2455
rect 16147 -2523 16239 -2510
rect 17232 -2454 17324 -2441
rect 17232 -2509 17248 -2454
rect 17308 -2509 17324 -2454
rect 17232 -2526 17324 -2509
rect 18930 -2450 19119 -2428
rect 22072 -2433 22177 -1190
rect 30073 -1345 30162 -1311
rect 30338 -1345 30354 -1311
rect 23504 -1490 23732 -1472
rect 23504 -1566 23520 -1490
rect 23716 -1566 23732 -1490
rect 23504 -1582 23732 -1566
rect 30073 -1547 30108 -1345
rect 30146 -1463 30162 -1429
rect 30338 -1463 30354 -1429
rect 31371 -1470 31387 -1436
rect 31563 -1470 31579 -1436
rect 30073 -1581 30162 -1547
rect 30338 -1581 30354 -1547
rect 31270 -1617 31286 -1583
rect 31320 -1617 31336 -1583
rect 31371 -1588 31387 -1554
rect 31563 -1588 31579 -1554
rect 22775 -1707 23045 -1668
rect 22775 -1760 22809 -1707
rect 22334 -1909 22604 -1870
rect 22334 -1960 22368 -1909
rect 22334 -2152 22368 -2136
rect 22452 -1960 22486 -1944
rect 22452 -2187 22486 -2136
rect 22570 -1960 22604 -1909
rect 22570 -2152 22604 -2136
rect 22688 -1960 22722 -1944
rect 22688 -2187 22722 -2136
rect 22775 -2152 22809 -2136
rect 22893 -1760 22927 -1744
rect 22452 -2226 22722 -2187
rect 22893 -2187 22927 -2136
rect 23011 -1760 23045 -1707
rect 23242 -1708 23512 -1669
rect 23011 -2152 23045 -2136
rect 23129 -1760 23163 -1744
rect 23129 -2187 23163 -2136
rect 23242 -1760 23276 -1708
rect 23242 -2152 23276 -2136
rect 23360 -1760 23394 -1744
rect 23360 -2187 23394 -2136
rect 23478 -1760 23512 -1708
rect 23714 -1708 23984 -1669
rect 23478 -2152 23512 -2136
rect 23596 -1760 23630 -1744
rect 23596 -2187 23630 -2136
rect 23714 -1760 23748 -1708
rect 23714 -2152 23748 -2136
rect 23832 -1760 23866 -1744
rect 23832 -2187 23866 -2136
rect 23950 -1760 23984 -1708
rect 24187 -1708 24457 -1669
rect 30146 -1699 30162 -1665
rect 30338 -1699 30354 -1665
rect 23950 -2152 23984 -2136
rect 24069 -1760 24103 -1744
rect 24069 -2187 24103 -2136
rect 24187 -1760 24221 -1708
rect 24187 -2152 24221 -2136
rect 24305 -1760 24339 -1744
rect 24305 -2187 24339 -2136
rect 24423 -1760 24457 -1708
rect 30639 -1772 30655 -1738
rect 31031 -1772 31047 -1738
rect 31203 -1768 31269 -1752
rect 29946 -1829 29962 -1795
rect 30338 -1829 30354 -1795
rect 31203 -1802 31219 -1768
rect 31253 -1802 31269 -1768
rect 31203 -1819 31269 -1802
rect 30984 -1856 31129 -1855
rect 24660 -1910 24930 -1873
rect 30639 -1890 30655 -1856
rect 31031 -1874 31129 -1856
rect 31031 -1890 31130 -1874
rect 31371 -1890 31387 -1856
rect 30984 -1891 31130 -1890
rect 31763 -1891 31865 -1856
rect 24423 -2152 24457 -2136
rect 24542 -1960 24576 -1944
rect 22893 -2226 24339 -2187
rect 24542 -2190 24576 -2136
rect 24660 -1960 24694 -1910
rect 24660 -2152 24694 -2136
rect 24778 -1960 24812 -1944
rect 24778 -2190 24812 -2136
rect 24896 -1960 24930 -1910
rect 29946 -1947 29962 -1913
rect 30338 -1947 30354 -1913
rect 31089 -1929 31130 -1891
rect 31089 -1963 31417 -1929
rect 30639 -2008 30655 -1974
rect 31031 -2008 31047 -1974
rect 24896 -2152 24930 -2136
rect 29671 -2096 29763 -2062
rect 29946 -2065 29962 -2031
rect 30338 -2065 30354 -2031
rect 31089 -2090 31130 -1963
rect 31371 -1974 31417 -1963
rect 31371 -2008 31387 -1974
rect 31763 -2008 31779 -1974
rect 31303 -2034 31337 -2018
rect 31303 -2084 31337 -2068
rect 30984 -2092 31130 -2090
rect 24542 -2229 24812 -2190
rect 29671 -2218 29691 -2096
rect 29735 -2148 29763 -2096
rect 30639 -2126 30655 -2092
rect 31031 -2126 31130 -2092
rect 31371 -2126 31387 -2092
rect 31763 -2126 31779 -2092
rect 29745 -2186 29763 -2148
rect 29735 -2218 29763 -2186
rect 29671 -2264 29763 -2218
rect 29874 -2183 29962 -2149
rect 30338 -2183 30354 -2149
rect 23420 -2351 23454 -2335
rect 24714 -2344 24730 -2310
rect 24764 -2344 24780 -2310
rect 23420 -2401 23454 -2385
rect 29874 -2385 29909 -2183
rect 30639 -2244 30655 -2210
rect 31031 -2244 31047 -2210
rect 29946 -2301 29962 -2267
rect 30338 -2301 30354 -2267
rect 31089 -2328 31130 -2126
rect 31302 -2152 31336 -2136
rect 31302 -2202 31336 -2186
rect 31371 -2244 31387 -2210
rect 31763 -2244 31779 -2210
rect 31830 -2327 31865 -1891
rect 31935 -2046 32023 -2030
rect 31935 -2086 31951 -2046
rect 31935 -2178 31951 -2136
rect 32007 -2178 32023 -2046
rect 31935 -2194 32023 -2178
rect 30639 -2362 30655 -2328
rect 31031 -2362 31130 -2328
rect 31371 -2362 31387 -2328
rect 31763 -2362 31865 -2327
rect 30985 -2364 31130 -2362
rect 29874 -2419 29962 -2385
rect 30338 -2419 30354 -2385
rect 18930 -2510 19051 -2450
rect 19100 -2510 19119 -2450
rect 18930 -2527 19119 -2510
rect 19279 -2451 19371 -2434
rect 19279 -2506 19295 -2451
rect 19355 -2506 19371 -2451
rect 19279 -2519 19371 -2506
rect 20364 -2450 20456 -2437
rect 20364 -2505 20380 -2450
rect 20440 -2505 20456 -2450
rect 20364 -2522 20456 -2505
rect 22072 -2450 22259 -2433
rect 22072 -2510 22195 -2450
rect 22244 -2510 22259 -2450
rect 18968 -2528 19119 -2527
rect 22072 -2528 22259 -2510
rect 22423 -2451 22515 -2434
rect 22423 -2506 22439 -2451
rect 22499 -2506 22515 -2451
rect 22423 -2519 22515 -2506
rect 23508 -2450 23600 -2437
rect 23508 -2505 23524 -2450
rect 23584 -2505 23600 -2450
rect 30639 -2480 30655 -2446
rect 31031 -2480 31047 -2446
rect 23508 -2522 23600 -2505
rect 15798 -2532 15903 -2531
rect 29946 -2537 29962 -2503
rect 30338 -2537 30354 -2503
rect 1732 -2585 1766 -2569
rect 1732 -2635 1766 -2619
rect 4876 -2585 4910 -2569
rect 4876 -2635 4910 -2619
rect 8008 -2581 8042 -2565
rect 8008 -2631 8042 -2615
rect 11152 -2581 11186 -2565
rect 11152 -2631 11186 -2615
rect 14354 -2585 14388 -2569
rect 14354 -2635 14388 -2619
rect 17498 -2585 17532 -2569
rect 17498 -2635 17532 -2619
rect 20630 -2581 20664 -2565
rect 20630 -2631 20664 -2615
rect 23774 -2581 23808 -2565
rect 23774 -2631 23808 -2615
rect 30146 -2666 30162 -2632
rect 30338 -2666 30354 -2632
rect 30517 -2718 30551 -2712
rect 1348 -2739 1440 -2726
rect 1348 -2794 1364 -2739
rect 1424 -2794 1440 -2739
rect 1348 -2811 1440 -2794
rect 4492 -2739 4584 -2726
rect 4492 -2794 4508 -2739
rect 4568 -2794 4584 -2739
rect 4492 -2811 4584 -2794
rect 7624 -2735 7716 -2722
rect 7624 -2790 7640 -2735
rect 7700 -2790 7716 -2735
rect 7624 -2807 7716 -2790
rect 10768 -2735 10860 -2722
rect 10768 -2790 10784 -2735
rect 10844 -2790 10860 -2735
rect 10768 -2807 10860 -2790
rect 13970 -2739 14062 -2726
rect 13970 -2794 13986 -2739
rect 14046 -2794 14062 -2739
rect 13970 -2811 14062 -2794
rect 17114 -2739 17206 -2726
rect 17114 -2794 17130 -2739
rect 17190 -2794 17206 -2739
rect 17114 -2811 17206 -2794
rect 20246 -2735 20338 -2722
rect 20246 -2790 20262 -2735
rect 20322 -2790 20338 -2735
rect 20246 -2807 20338 -2790
rect 23390 -2735 23482 -2722
rect 23390 -2790 23406 -2735
rect 23466 -2790 23482 -2735
rect 30146 -2784 30162 -2750
rect 30338 -2784 30354 -2750
rect 30517 -2778 30551 -2772
rect 23390 -2807 23482 -2790
rect 30146 -2902 30162 -2868
rect 30338 -2902 30354 -2868
rect 31089 -2950 31130 -2364
rect 31203 -2416 31269 -2399
rect 31203 -2450 31219 -2416
rect 31253 -2450 31269 -2416
rect 31203 -2466 31269 -2450
rect 31271 -2740 31287 -2706
rect 31321 -2740 31337 -2706
rect 32528 -2716 32614 866
rect 32680 -2178 32760 2938
rect 33365 922 33458 6941
rect 33510 6708 33601 9477
rect 33658 9510 33743 22360
rect 33812 10840 33883 22803
rect 39614 22679 39648 22695
rect 39732 22871 39766 22887
rect 39732 22679 39766 22695
rect 39850 22871 39884 22887
rect 39850 22679 39884 22695
rect 39968 22871 40002 22887
rect 39968 22679 40002 22695
rect 40086 22871 40120 22887
rect 40086 22679 40120 22695
rect 40204 22871 40238 22887
rect 40204 22679 40238 22695
rect 40322 22871 40356 22887
rect 40322 22679 40356 22695
rect 40440 22871 40474 22921
rect 40440 22679 40474 22695
rect 40558 22871 40592 22887
rect 40558 22679 40592 22695
rect 40676 22871 40710 22921
rect 40676 22679 40710 22695
rect 43720 22942 43945 23018
rect 43720 22793 43799 22942
rect 43866 22793 43945 22942
rect 46953 22918 47223 22952
rect 43720 22687 43945 22793
rect 46127 22868 46161 22884
rect 46127 22676 46161 22692
rect 46245 22868 46279 22884
rect 46245 22676 46279 22692
rect 46363 22868 46397 22884
rect 46363 22676 46397 22692
rect 46481 22868 46515 22884
rect 46481 22676 46515 22692
rect 46599 22868 46633 22884
rect 46599 22676 46633 22692
rect 46717 22868 46751 22884
rect 46717 22676 46751 22692
rect 46835 22868 46869 22884
rect 46835 22676 46869 22692
rect 46953 22868 46987 22918
rect 46953 22676 46987 22692
rect 47071 22868 47105 22884
rect 47071 22676 47105 22692
rect 47189 22868 47223 22918
rect 47189 22676 47223 22692
rect 50233 22939 50458 23015
rect 50233 22790 50312 22939
rect 50379 22790 50458 22939
rect 53487 22913 53757 22947
rect 50233 22684 50458 22790
rect 52661 22863 52695 22879
rect 52661 22671 52695 22687
rect 52779 22863 52813 22879
rect 52779 22671 52813 22687
rect 52897 22863 52931 22879
rect 52897 22671 52931 22687
rect 53015 22863 53049 22879
rect 53015 22671 53049 22687
rect 53133 22863 53167 22879
rect 53133 22671 53167 22687
rect 53251 22863 53285 22879
rect 53251 22671 53285 22687
rect 53369 22863 53403 22879
rect 53369 22671 53403 22687
rect 53487 22863 53521 22913
rect 53487 22671 53521 22687
rect 53605 22863 53639 22879
rect 53605 22671 53639 22687
rect 53723 22863 53757 22913
rect 53723 22671 53757 22687
rect 56767 22934 56992 23010
rect 56767 22785 56846 22934
rect 56913 22785 56992 22934
rect 60045 22917 60315 22951
rect 56767 22679 56992 22785
rect 59219 22867 59253 22883
rect 59219 22675 59253 22691
rect 59337 22867 59371 22883
rect 59337 22675 59371 22691
rect 59455 22867 59489 22883
rect 59455 22675 59489 22691
rect 59573 22867 59607 22883
rect 59573 22675 59607 22691
rect 59691 22867 59725 22883
rect 59691 22675 59725 22691
rect 59809 22867 59843 22883
rect 59809 22675 59843 22691
rect 59927 22867 59961 22883
rect 59927 22675 59961 22691
rect 60045 22867 60079 22917
rect 60045 22675 60079 22691
rect 60163 22867 60197 22883
rect 60163 22675 60197 22691
rect 60281 22867 60315 22917
rect 60281 22675 60315 22691
rect 63325 22938 63550 23014
rect 63325 22789 63404 22938
rect 63471 22789 63550 22938
rect 63325 22683 63550 22789
rect 40365 22601 40381 22635
rect 40415 22601 40431 22635
rect 46878 22598 46894 22632
rect 46928 22598 46944 22632
rect 53412 22593 53428 22627
rect 53462 22593 53478 22627
rect 59970 22597 59986 22631
rect 60020 22597 60036 22631
rect 40247 22484 40263 22518
rect 40297 22484 40313 22518
rect 41916 22507 42186 22542
rect 41562 22454 41596 22470
rect 39851 22434 39885 22450
rect 39851 22042 39885 22058
rect 39969 22434 40003 22450
rect 39969 22042 40003 22058
rect 40087 22434 40121 22450
rect 40204 22434 40238 22450
rect 40204 22242 40238 22258
rect 40322 22434 40356 22450
rect 40322 22242 40356 22258
rect 41078 22308 41348 22343
rect 41078 22254 41112 22308
rect 40087 22042 40121 22058
rect 40374 22108 40623 22151
rect 40374 22018 40421 22108
rect 40584 22018 40623 22108
rect 41078 22062 41112 22078
rect 41196 22254 41230 22270
rect 41196 22062 41230 22078
rect 41314 22254 41348 22308
rect 41314 22062 41348 22078
rect 41432 22254 41466 22270
rect 41432 22062 41466 22078
rect 41562 22062 41596 22078
rect 41680 22454 41714 22470
rect 41680 22062 41714 22078
rect 41798 22454 41832 22470
rect 41798 22062 41832 22078
rect 41916 22454 41950 22507
rect 41916 22062 41950 22078
rect 42034 22454 42068 22470
rect 42034 22062 42068 22078
rect 42152 22454 42186 22507
rect 43814 22507 44084 22542
rect 42152 22062 42186 22078
rect 42270 22454 42304 22470
rect 43460 22454 43494 22470
rect 42976 22308 43246 22343
rect 42270 22062 42304 22078
rect 42399 22254 42433 22270
rect 42399 22062 42433 22078
rect 42517 22254 42551 22270
rect 42517 22062 42551 22078
rect 42635 22254 42669 22270
rect 42635 22062 42669 22078
rect 42753 22254 42787 22270
rect 42753 22062 42787 22078
rect 42976 22254 43010 22308
rect 42976 22062 43010 22078
rect 43094 22254 43128 22270
rect 43094 22062 43128 22078
rect 43212 22254 43246 22308
rect 43212 22062 43246 22078
rect 43330 22254 43364 22270
rect 43330 22062 43364 22078
rect 43460 22062 43494 22078
rect 43578 22454 43612 22470
rect 43578 22062 43612 22078
rect 43696 22454 43730 22470
rect 43696 22062 43730 22078
rect 43814 22454 43848 22507
rect 43814 22062 43848 22078
rect 43932 22454 43966 22470
rect 43932 22062 43966 22078
rect 44050 22454 44084 22507
rect 46760 22481 46776 22515
rect 46810 22481 46826 22515
rect 48429 22504 48699 22539
rect 44050 22062 44084 22078
rect 44168 22454 44202 22470
rect 48075 22451 48109 22467
rect 46364 22431 46398 22447
rect 44168 22062 44202 22078
rect 44297 22254 44331 22270
rect 44297 22062 44331 22078
rect 44415 22254 44449 22270
rect 44415 22062 44449 22078
rect 44533 22254 44567 22270
rect 44533 22062 44567 22078
rect 44651 22254 44685 22270
rect 44651 22062 44685 22078
rect 46364 22039 46398 22055
rect 46482 22431 46516 22447
rect 46482 22039 46516 22055
rect 46600 22431 46634 22447
rect 46717 22431 46751 22447
rect 46717 22239 46751 22255
rect 46835 22431 46869 22447
rect 46835 22239 46869 22255
rect 47591 22305 47861 22340
rect 47591 22251 47625 22305
rect 46600 22039 46634 22055
rect 46887 22105 47136 22148
rect 39894 21974 39910 22008
rect 39944 21974 39960 22008
rect 40012 21974 40028 22008
rect 40062 21974 40078 22008
rect 40374 21979 40623 22018
rect 46887 22015 46934 22105
rect 47097 22015 47136 22105
rect 47591 22059 47625 22075
rect 47709 22251 47743 22267
rect 47709 22059 47743 22075
rect 47827 22251 47861 22305
rect 47827 22059 47861 22075
rect 47945 22251 47979 22267
rect 47945 22059 47979 22075
rect 48075 22059 48109 22075
rect 48193 22451 48227 22467
rect 48193 22059 48227 22075
rect 48311 22451 48345 22467
rect 48311 22059 48345 22075
rect 48429 22451 48463 22504
rect 48429 22059 48463 22075
rect 48547 22451 48581 22467
rect 48547 22059 48581 22075
rect 48665 22451 48699 22504
rect 50327 22504 50597 22539
rect 48665 22059 48699 22075
rect 48783 22451 48817 22467
rect 49973 22451 50007 22467
rect 49489 22305 49759 22340
rect 48783 22059 48817 22075
rect 48912 22251 48946 22267
rect 48912 22059 48946 22075
rect 49030 22251 49064 22267
rect 49030 22059 49064 22075
rect 49148 22251 49182 22267
rect 49148 22059 49182 22075
rect 49266 22251 49300 22267
rect 49266 22059 49300 22075
rect 49489 22251 49523 22305
rect 49489 22059 49523 22075
rect 49607 22251 49641 22267
rect 49607 22059 49641 22075
rect 49725 22251 49759 22305
rect 49725 22059 49759 22075
rect 49843 22251 49877 22267
rect 49843 22059 49877 22075
rect 49973 22059 50007 22075
rect 50091 22451 50125 22467
rect 50091 22059 50125 22075
rect 50209 22451 50243 22467
rect 50209 22059 50243 22075
rect 50327 22451 50361 22504
rect 50327 22059 50361 22075
rect 50445 22451 50479 22467
rect 50445 22059 50479 22075
rect 50563 22451 50597 22504
rect 53294 22476 53310 22510
rect 53344 22476 53360 22510
rect 54963 22499 55233 22534
rect 50563 22059 50597 22075
rect 50681 22451 50715 22467
rect 54609 22446 54643 22462
rect 52898 22426 52932 22442
rect 50681 22059 50715 22075
rect 50810 22251 50844 22267
rect 50810 22059 50844 22075
rect 50928 22251 50962 22267
rect 50928 22059 50962 22075
rect 51046 22251 51080 22267
rect 51046 22059 51080 22075
rect 51164 22251 51198 22267
rect 51164 22059 51198 22075
rect 52898 22034 52932 22050
rect 53016 22426 53050 22442
rect 53016 22034 53050 22050
rect 53134 22426 53168 22442
rect 53251 22426 53285 22442
rect 53251 22234 53285 22250
rect 53369 22426 53403 22442
rect 53369 22234 53403 22250
rect 54125 22300 54395 22335
rect 54125 22246 54159 22300
rect 53134 22034 53168 22050
rect 53421 22100 53670 22143
rect 46407 21971 46423 22005
rect 46457 21971 46473 22005
rect 46525 21971 46541 22005
rect 46575 21971 46591 22005
rect 46887 21976 47136 22015
rect 53421 22010 53468 22100
rect 53631 22010 53670 22100
rect 54125 22054 54159 22070
rect 54243 22246 54277 22262
rect 54243 22054 54277 22070
rect 54361 22246 54395 22300
rect 54361 22054 54395 22070
rect 54479 22246 54513 22262
rect 54479 22054 54513 22070
rect 54609 22054 54643 22070
rect 54727 22446 54761 22462
rect 54727 22054 54761 22070
rect 54845 22446 54879 22462
rect 54845 22054 54879 22070
rect 54963 22446 54997 22499
rect 54963 22054 54997 22070
rect 55081 22446 55115 22462
rect 55081 22054 55115 22070
rect 55199 22446 55233 22499
rect 56861 22499 57131 22534
rect 55199 22054 55233 22070
rect 55317 22446 55351 22462
rect 56507 22446 56541 22462
rect 56023 22300 56293 22335
rect 55317 22054 55351 22070
rect 55446 22246 55480 22262
rect 55446 22054 55480 22070
rect 55564 22246 55598 22262
rect 55564 22054 55598 22070
rect 55682 22246 55716 22262
rect 55682 22054 55716 22070
rect 55800 22246 55834 22262
rect 55800 22054 55834 22070
rect 56023 22246 56057 22300
rect 56023 22054 56057 22070
rect 56141 22246 56175 22262
rect 56141 22054 56175 22070
rect 56259 22246 56293 22300
rect 56259 22054 56293 22070
rect 56377 22246 56411 22262
rect 56377 22054 56411 22070
rect 56507 22054 56541 22070
rect 56625 22446 56659 22462
rect 56625 22054 56659 22070
rect 56743 22446 56777 22462
rect 56743 22054 56777 22070
rect 56861 22446 56895 22499
rect 56861 22054 56895 22070
rect 56979 22446 57013 22462
rect 56979 22054 57013 22070
rect 57097 22446 57131 22499
rect 59852 22480 59868 22514
rect 59902 22480 59918 22514
rect 61521 22503 61791 22538
rect 57097 22054 57131 22070
rect 57215 22446 57249 22462
rect 61167 22450 61201 22466
rect 59456 22430 59490 22446
rect 57215 22054 57249 22070
rect 57344 22246 57378 22262
rect 57344 22054 57378 22070
rect 57462 22246 57496 22262
rect 57462 22054 57496 22070
rect 57580 22246 57614 22262
rect 57580 22054 57614 22070
rect 57698 22246 57732 22262
rect 57698 22054 57732 22070
rect 59456 22038 59490 22054
rect 59574 22430 59608 22446
rect 59574 22038 59608 22054
rect 59692 22430 59726 22446
rect 59809 22430 59843 22446
rect 59809 22238 59843 22254
rect 59927 22430 59961 22446
rect 59927 22238 59961 22254
rect 60683 22304 60953 22339
rect 60683 22250 60717 22304
rect 59692 22038 59726 22054
rect 59979 22104 60228 22147
rect 52941 21966 52957 22000
rect 52991 21966 53007 22000
rect 53059 21966 53075 22000
rect 53109 21966 53125 22000
rect 53421 21971 53670 22010
rect 59979 22014 60026 22104
rect 60189 22014 60228 22104
rect 60683 22058 60717 22074
rect 60801 22250 60835 22266
rect 60801 22058 60835 22074
rect 60919 22250 60953 22304
rect 60919 22058 60953 22074
rect 61037 22250 61071 22266
rect 61037 22058 61071 22074
rect 61167 22058 61201 22074
rect 61285 22450 61319 22466
rect 61285 22058 61319 22074
rect 61403 22450 61437 22466
rect 61403 22058 61437 22074
rect 61521 22450 61555 22503
rect 61521 22058 61555 22074
rect 61639 22450 61673 22466
rect 61639 22058 61673 22074
rect 61757 22450 61791 22503
rect 63419 22503 63689 22538
rect 61757 22058 61791 22074
rect 61875 22450 61909 22466
rect 63065 22450 63099 22466
rect 62581 22304 62851 22339
rect 61875 22058 61909 22074
rect 62004 22250 62038 22266
rect 62004 22058 62038 22074
rect 62122 22250 62156 22266
rect 62122 22058 62156 22074
rect 62240 22250 62274 22266
rect 62240 22058 62274 22074
rect 62358 22250 62392 22266
rect 62358 22058 62392 22074
rect 62581 22250 62615 22304
rect 62581 22058 62615 22074
rect 62699 22250 62733 22266
rect 62699 22058 62733 22074
rect 62817 22250 62851 22304
rect 62817 22058 62851 22074
rect 62935 22250 62969 22266
rect 62935 22058 62969 22074
rect 63065 22058 63099 22074
rect 63183 22450 63217 22466
rect 63183 22058 63217 22074
rect 63301 22450 63335 22466
rect 63301 22058 63335 22074
rect 63419 22450 63453 22503
rect 63419 22058 63453 22074
rect 63537 22450 63571 22466
rect 63537 22058 63571 22074
rect 63655 22450 63689 22503
rect 63655 22058 63689 22074
rect 63773 22450 63807 22466
rect 68599 22300 68722 22316
rect 63773 22058 63807 22074
rect 63902 22250 63936 22266
rect 63902 22058 63936 22074
rect 64020 22250 64054 22266
rect 64020 22058 64054 22074
rect 64138 22250 64172 22266
rect 64138 22058 64172 22074
rect 64256 22250 64290 22266
rect 64256 22058 64290 22074
rect 68599 22235 68618 22300
rect 68701 22235 68722 22300
rect 59499 21970 59515 22004
rect 59549 21970 59565 22004
rect 59617 21970 59633 22004
rect 59667 21970 59683 22004
rect 59979 21975 60228 22014
rect 42542 21840 42576 21856
rect 49055 21837 49089 21853
rect 42542 21790 42576 21806
rect 44632 21819 44699 21835
rect 44632 21785 44649 21819
rect 44683 21785 44699 21819
rect 55589 21832 55623 21848
rect 49055 21787 49089 21803
rect 51145 21816 51212 21832
rect 41505 21761 41539 21777
rect 40004 21681 40227 21757
rect 40004 21532 40083 21681
rect 40150 21532 40227 21681
rect 40004 21426 40227 21532
rect 41623 21761 41657 21777
rect 41505 21369 41539 21385
rect 41622 21385 41623 21432
rect 41741 21761 41775 21777
rect 41657 21385 41658 21432
rect 40435 21317 40705 21351
rect 39609 21267 39643 21283
rect 39609 21075 39643 21091
rect 39727 21267 39761 21283
rect 39727 21075 39761 21091
rect 39845 21267 39879 21283
rect 39845 21075 39879 21091
rect 39963 21267 39997 21283
rect 39963 21075 39997 21091
rect 40081 21267 40115 21283
rect 40081 21075 40115 21091
rect 40199 21267 40233 21283
rect 40199 21075 40233 21091
rect 40317 21267 40351 21283
rect 40317 21075 40351 21091
rect 40435 21267 40469 21317
rect 40435 21075 40469 21091
rect 40553 21267 40587 21283
rect 40553 21075 40587 21091
rect 40671 21267 40705 21317
rect 41622 21327 41658 21385
rect 41859 21761 41893 21777
rect 41741 21369 41775 21385
rect 41857 21385 41859 21432
rect 41857 21327 41893 21385
rect 41977 21761 42011 21777
rect 41977 21369 42011 21385
rect 42095 21761 42129 21777
rect 42213 21761 42247 21777
rect 42129 21385 42131 21431
rect 42095 21327 42131 21385
rect 42213 21369 42247 21385
rect 43403 21761 43437 21777
rect 43521 21761 43555 21777
rect 43403 21369 43437 21385
rect 43520 21385 43521 21432
rect 43639 21761 43673 21777
rect 43555 21385 43556 21432
rect 42718 21327 43215 21345
rect 41622 21324 43215 21327
rect 41622 21290 43163 21324
rect 43197 21290 43215 21324
rect 41622 21287 43215 21290
rect 43520 21327 43556 21385
rect 43757 21761 43791 21777
rect 43639 21369 43673 21385
rect 43755 21385 43757 21432
rect 43755 21327 43791 21385
rect 43875 21761 43909 21777
rect 43875 21369 43909 21385
rect 43993 21761 44027 21777
rect 44111 21761 44145 21777
rect 44632 21769 44699 21785
rect 51145 21782 51162 21816
rect 51196 21782 51212 21816
rect 62147 21836 62181 21852
rect 55589 21782 55623 21798
rect 57679 21811 57746 21827
rect 44027 21385 44029 21431
rect 43993 21327 44029 21385
rect 48018 21758 48052 21774
rect 46517 21678 46740 21754
rect 46517 21529 46596 21678
rect 46663 21529 46740 21678
rect 46517 21423 46740 21529
rect 44111 21369 44145 21385
rect 48136 21758 48170 21774
rect 48018 21366 48052 21382
rect 48135 21382 48136 21429
rect 48254 21758 48288 21774
rect 48170 21382 48171 21429
rect 44616 21356 44716 21357
rect 44616 21327 44904 21356
rect 43520 21287 44904 21327
rect 41641 21286 43215 21287
rect 43539 21286 44904 21287
rect 41519 21197 41586 21213
rect 41519 21163 41535 21197
rect 41569 21163 41586 21197
rect 41519 21147 41586 21163
rect 40671 21075 40705 21091
rect 41350 21130 41384 21146
rect 41350 21080 41384 21096
rect 41696 21045 41730 21286
rect 42718 21269 43215 21286
rect 42166 21197 42233 21213
rect 42166 21163 42183 21197
rect 42217 21163 42233 21197
rect 42166 21147 42233 21163
rect 43417 21197 43484 21213
rect 43417 21163 43433 21197
rect 43467 21163 43484 21197
rect 43417 21147 43484 21163
rect 42473 21129 42507 21145
rect 41785 21079 41801 21113
rect 41835 21079 41851 21113
rect 41903 21080 41919 21114
rect 41953 21080 41969 21114
rect 42473 21079 42507 21095
rect 43248 21130 43282 21146
rect 43248 21080 43282 21096
rect 43594 21045 43628 21286
rect 44616 21281 44904 21286
rect 46948 21314 47218 21348
rect 44616 21258 44906 21281
rect 44616 21257 44716 21258
rect 44062 21198 44129 21214
rect 44062 21164 44079 21198
rect 44113 21164 44129 21198
rect 44062 21148 44129 21164
rect 44371 21129 44405 21145
rect 43683 21079 43699 21113
rect 43733 21079 43749 21113
rect 43801 21080 43817 21114
rect 43851 21080 43867 21114
rect 44371 21079 44405 21095
rect 40360 20997 40376 21031
rect 40410 20997 40426 21031
rect 41203 21029 41237 21045
rect 40242 20880 40258 20914
rect 40292 20880 40308 20914
rect 39846 20830 39880 20846
rect 39846 20438 39880 20454
rect 39964 20830 39998 20846
rect 39964 20438 39998 20454
rect 40082 20830 40116 20846
rect 40199 20830 40233 20846
rect 40199 20638 40233 20654
rect 40317 20830 40351 20846
rect 41203 20837 41237 20853
rect 41321 21029 41355 21045
rect 41321 20837 41355 20853
rect 41623 21029 41657 21045
rect 40317 20638 40351 20654
rect 41696 21029 41775 21045
rect 41696 20999 41741 21029
rect 41623 20586 41658 20653
rect 41741 20637 41775 20653
rect 41859 21029 41893 21045
rect 41859 20637 41893 20653
rect 41977 21029 42011 21045
rect 42095 21029 42129 21045
rect 42501 21029 42535 21045
rect 42501 20837 42535 20853
rect 42619 21029 42653 21045
rect 42619 20837 42653 20853
rect 43101 21029 43135 21045
rect 43101 20837 43135 20853
rect 43219 21029 43253 21045
rect 43219 20837 43253 20853
rect 43521 21029 43555 21045
rect 41977 20637 42011 20653
rect 42094 20586 42129 20653
rect 41623 20551 42129 20586
rect 43594 21029 43673 21045
rect 43594 20999 43639 21029
rect 43521 20586 43556 20653
rect 43639 20637 43673 20653
rect 43757 21029 43791 21045
rect 43757 20637 43791 20653
rect 43875 21029 43909 21045
rect 43993 21029 44027 21045
rect 44399 21029 44433 21045
rect 44399 20837 44433 20853
rect 44517 21029 44551 21045
rect 44517 20837 44551 20853
rect 43875 20637 43909 20653
rect 43992 20586 44027 20653
rect 43521 20551 44027 20586
rect 40082 20438 40116 20454
rect 40369 20504 40618 20547
rect 40369 20414 40416 20504
rect 40579 20414 40618 20504
rect 39889 20370 39905 20404
rect 39939 20370 39955 20404
rect 40007 20370 40023 20404
rect 40057 20370 40073 20404
rect 40369 20375 40618 20414
rect 41794 20344 41966 20391
rect 41794 20181 41833 20344
rect 41923 20181 41966 20344
rect 41794 20141 41966 20181
rect 44765 19641 44906 21258
rect 46122 21264 46156 21280
rect 46122 21072 46156 21088
rect 46240 21264 46274 21280
rect 46240 21072 46274 21088
rect 46358 21264 46392 21280
rect 46358 21072 46392 21088
rect 46476 21264 46510 21280
rect 46476 21072 46510 21088
rect 46594 21264 46628 21280
rect 46594 21072 46628 21088
rect 46712 21264 46746 21280
rect 46712 21072 46746 21088
rect 46830 21264 46864 21280
rect 46830 21072 46864 21088
rect 46948 21264 46982 21314
rect 46948 21072 46982 21088
rect 47066 21264 47100 21280
rect 47066 21072 47100 21088
rect 47184 21264 47218 21314
rect 48135 21324 48171 21382
rect 48372 21758 48406 21774
rect 48254 21366 48288 21382
rect 48370 21382 48372 21429
rect 48370 21324 48406 21382
rect 48490 21758 48524 21774
rect 48490 21366 48524 21382
rect 48608 21758 48642 21774
rect 48726 21758 48760 21774
rect 48642 21382 48644 21428
rect 48608 21324 48644 21382
rect 48726 21366 48760 21382
rect 49916 21758 49950 21774
rect 50034 21758 50068 21774
rect 49916 21366 49950 21382
rect 50033 21382 50034 21429
rect 50152 21758 50186 21774
rect 50068 21382 50069 21429
rect 49231 21324 49728 21342
rect 48135 21321 49728 21324
rect 48135 21287 49676 21321
rect 49710 21287 49728 21321
rect 48135 21284 49728 21287
rect 50033 21324 50069 21382
rect 50270 21758 50304 21774
rect 50152 21366 50186 21382
rect 50268 21382 50270 21429
rect 50268 21324 50304 21382
rect 50388 21758 50422 21774
rect 50388 21366 50422 21382
rect 50506 21758 50540 21774
rect 50624 21758 50658 21774
rect 51145 21766 51212 21782
rect 57679 21777 57696 21811
rect 57730 21777 57746 21811
rect 62147 21786 62181 21802
rect 64237 21815 64304 21831
rect 50540 21382 50542 21428
rect 50506 21324 50542 21382
rect 54552 21753 54586 21769
rect 53051 21673 53274 21749
rect 53051 21524 53130 21673
rect 53197 21524 53274 21673
rect 53051 21418 53274 21524
rect 50624 21366 50658 21382
rect 54670 21753 54704 21769
rect 54552 21361 54586 21377
rect 54669 21377 54670 21424
rect 54788 21753 54822 21769
rect 54704 21377 54705 21424
rect 51129 21353 51229 21354
rect 51129 21324 51417 21353
rect 50033 21312 51417 21324
rect 50033 21284 51418 21312
rect 48154 21283 49728 21284
rect 50052 21283 51418 21284
rect 48032 21194 48099 21210
rect 48032 21160 48048 21194
rect 48082 21160 48099 21194
rect 48032 21144 48099 21160
rect 47184 21072 47218 21088
rect 47863 21127 47897 21143
rect 47863 21077 47897 21093
rect 48209 21042 48243 21283
rect 49231 21266 49728 21283
rect 48679 21194 48746 21210
rect 48679 21160 48696 21194
rect 48730 21160 48746 21194
rect 48679 21144 48746 21160
rect 49930 21194 49997 21210
rect 49930 21160 49946 21194
rect 49980 21160 49997 21194
rect 49930 21144 49997 21160
rect 48986 21126 49020 21142
rect 48298 21076 48314 21110
rect 48348 21076 48364 21110
rect 48416 21077 48432 21111
rect 48466 21077 48482 21111
rect 48986 21076 49020 21092
rect 49761 21127 49795 21143
rect 49761 21077 49795 21093
rect 50107 21042 50141 21283
rect 51129 21255 51418 21283
rect 53482 21309 53752 21343
rect 51129 21254 51229 21255
rect 50575 21195 50642 21211
rect 50575 21161 50592 21195
rect 50626 21161 50642 21195
rect 50575 21145 50642 21161
rect 50884 21126 50918 21142
rect 50196 21076 50212 21110
rect 50246 21076 50262 21110
rect 50314 21077 50330 21111
rect 50364 21077 50380 21111
rect 50884 21076 50918 21092
rect 46873 20994 46889 21028
rect 46923 20994 46939 21028
rect 47716 21026 47750 21042
rect 46755 20877 46771 20911
rect 46805 20877 46821 20911
rect 46359 20827 46393 20843
rect 46359 20435 46393 20451
rect 46477 20827 46511 20843
rect 46477 20435 46511 20451
rect 46595 20827 46629 20843
rect 46712 20827 46746 20843
rect 46712 20635 46746 20651
rect 46830 20827 46864 20843
rect 47716 20834 47750 20850
rect 47834 21026 47868 21042
rect 47834 20834 47868 20850
rect 48136 21026 48170 21042
rect 46830 20635 46864 20651
rect 48209 21026 48288 21042
rect 48209 20996 48254 21026
rect 48136 20583 48171 20650
rect 48254 20634 48288 20650
rect 48372 21026 48406 21042
rect 48372 20634 48406 20650
rect 48490 21026 48524 21042
rect 48608 21026 48642 21042
rect 49014 21026 49048 21042
rect 49014 20834 49048 20850
rect 49132 21026 49166 21042
rect 49132 20834 49166 20850
rect 49614 21026 49648 21042
rect 49614 20834 49648 20850
rect 49732 21026 49766 21042
rect 49732 20834 49766 20850
rect 50034 21026 50068 21042
rect 48490 20634 48524 20650
rect 48607 20583 48642 20650
rect 48136 20548 48642 20583
rect 50107 21026 50186 21042
rect 50107 20996 50152 21026
rect 50034 20583 50069 20650
rect 50152 20634 50186 20650
rect 50270 21026 50304 21042
rect 50270 20634 50304 20650
rect 50388 21026 50422 21042
rect 50506 21026 50540 21042
rect 50912 21026 50946 21042
rect 50912 20834 50946 20850
rect 51030 21026 51064 21042
rect 51030 20834 51064 20850
rect 50388 20634 50422 20650
rect 50505 20583 50540 20650
rect 50034 20548 50540 20583
rect 46595 20435 46629 20451
rect 46882 20501 47131 20544
rect 46882 20411 46929 20501
rect 47092 20411 47131 20501
rect 46402 20367 46418 20401
rect 46452 20367 46468 20401
rect 46520 20367 46536 20401
rect 46570 20367 46586 20401
rect 46882 20372 47131 20411
rect 48307 20341 48479 20388
rect 48307 20178 48346 20341
rect 48436 20178 48479 20341
rect 48307 20138 48479 20178
rect 51290 19828 51418 21255
rect 52656 21259 52690 21275
rect 52656 21067 52690 21083
rect 52774 21259 52808 21275
rect 52774 21067 52808 21083
rect 52892 21259 52926 21275
rect 52892 21067 52926 21083
rect 53010 21259 53044 21275
rect 53010 21067 53044 21083
rect 53128 21259 53162 21275
rect 53128 21067 53162 21083
rect 53246 21259 53280 21275
rect 53246 21067 53280 21083
rect 53364 21259 53398 21275
rect 53364 21067 53398 21083
rect 53482 21259 53516 21309
rect 53482 21067 53516 21083
rect 53600 21259 53634 21275
rect 53600 21067 53634 21083
rect 53718 21259 53752 21309
rect 54669 21319 54705 21377
rect 54906 21753 54940 21769
rect 54788 21361 54822 21377
rect 54904 21377 54906 21424
rect 54904 21319 54940 21377
rect 55024 21753 55058 21769
rect 55024 21361 55058 21377
rect 55142 21753 55176 21769
rect 55260 21753 55294 21769
rect 55176 21377 55178 21423
rect 55142 21319 55178 21377
rect 55260 21361 55294 21377
rect 56450 21753 56484 21769
rect 56568 21753 56602 21769
rect 56450 21361 56484 21377
rect 56567 21377 56568 21424
rect 56686 21753 56720 21769
rect 56602 21377 56603 21424
rect 55765 21319 56262 21337
rect 54669 21316 56262 21319
rect 54669 21282 56210 21316
rect 56244 21282 56262 21316
rect 54669 21279 56262 21282
rect 56567 21319 56603 21377
rect 56804 21753 56838 21769
rect 56686 21361 56720 21377
rect 56802 21377 56804 21424
rect 56802 21319 56838 21377
rect 56922 21753 56956 21769
rect 56922 21361 56956 21377
rect 57040 21753 57074 21769
rect 57158 21753 57192 21769
rect 57679 21761 57746 21777
rect 64237 21781 64254 21815
rect 64288 21781 64304 21815
rect 61110 21757 61144 21773
rect 57074 21377 57076 21423
rect 57040 21319 57076 21377
rect 59609 21677 59832 21753
rect 59609 21528 59688 21677
rect 59755 21528 59832 21677
rect 59609 21422 59832 21528
rect 57158 21361 57192 21377
rect 61228 21757 61262 21773
rect 61110 21365 61144 21381
rect 61227 21381 61228 21428
rect 61346 21757 61380 21773
rect 61262 21381 61263 21428
rect 57663 21348 57763 21349
rect 57663 21319 57951 21348
rect 56567 21295 57951 21319
rect 60040 21313 60310 21347
rect 56567 21279 57952 21295
rect 54688 21278 56262 21279
rect 56586 21278 57952 21279
rect 54566 21189 54633 21205
rect 54566 21155 54582 21189
rect 54616 21155 54633 21189
rect 54566 21139 54633 21155
rect 53718 21067 53752 21083
rect 54397 21122 54431 21138
rect 54397 21072 54431 21088
rect 54743 21037 54777 21278
rect 55765 21261 56262 21278
rect 55213 21189 55280 21205
rect 55213 21155 55230 21189
rect 55264 21155 55280 21189
rect 55213 21139 55280 21155
rect 56464 21189 56531 21205
rect 56464 21155 56480 21189
rect 56514 21155 56531 21189
rect 56464 21139 56531 21155
rect 55520 21121 55554 21137
rect 54832 21071 54848 21105
rect 54882 21071 54898 21105
rect 54950 21072 54966 21106
rect 55000 21072 55016 21106
rect 55520 21071 55554 21087
rect 56295 21122 56329 21138
rect 56295 21072 56329 21088
rect 56641 21037 56675 21278
rect 57663 21250 57952 21278
rect 57663 21249 57763 21250
rect 57109 21190 57176 21206
rect 57109 21156 57126 21190
rect 57160 21156 57176 21190
rect 57109 21140 57176 21156
rect 57418 21121 57452 21137
rect 56730 21071 56746 21105
rect 56780 21071 56796 21105
rect 56848 21072 56864 21106
rect 56898 21072 56914 21106
rect 57418 21071 57452 21087
rect 53407 20989 53423 21023
rect 53457 20989 53473 21023
rect 54250 21021 54284 21037
rect 53289 20872 53305 20906
rect 53339 20872 53355 20906
rect 52893 20822 52927 20838
rect 52893 20430 52927 20446
rect 53011 20822 53045 20838
rect 53011 20430 53045 20446
rect 53129 20822 53163 20838
rect 53246 20822 53280 20838
rect 53246 20630 53280 20646
rect 53364 20822 53398 20838
rect 54250 20829 54284 20845
rect 54368 21021 54402 21037
rect 54368 20829 54402 20845
rect 54670 21021 54704 21037
rect 53364 20630 53398 20646
rect 54743 21021 54822 21037
rect 54743 20991 54788 21021
rect 54670 20578 54705 20645
rect 54788 20629 54822 20645
rect 54906 21021 54940 21037
rect 54906 20629 54940 20645
rect 55024 21021 55058 21037
rect 55142 21021 55176 21037
rect 55548 21021 55582 21037
rect 55548 20829 55582 20845
rect 55666 21021 55700 21037
rect 55666 20829 55700 20845
rect 56148 21021 56182 21037
rect 56148 20829 56182 20845
rect 56266 21021 56300 21037
rect 56266 20829 56300 20845
rect 56568 21021 56602 21037
rect 55024 20629 55058 20645
rect 55141 20578 55176 20645
rect 54670 20543 55176 20578
rect 56641 21021 56720 21037
rect 56641 20991 56686 21021
rect 56568 20578 56603 20645
rect 56686 20629 56720 20645
rect 56804 21021 56838 21037
rect 56804 20629 56838 20645
rect 56922 21021 56956 21037
rect 57040 21021 57074 21037
rect 57446 21021 57480 21037
rect 57446 20829 57480 20845
rect 57564 21021 57598 21037
rect 57564 20829 57598 20845
rect 56922 20629 56956 20645
rect 57039 20578 57074 20645
rect 56568 20543 57074 20578
rect 53129 20430 53163 20446
rect 53416 20496 53665 20539
rect 53416 20406 53463 20496
rect 53626 20406 53665 20496
rect 52936 20362 52952 20396
rect 52986 20362 53002 20396
rect 53054 20362 53070 20396
rect 53104 20362 53120 20396
rect 53416 20367 53665 20406
rect 54841 20336 55013 20383
rect 54841 20173 54880 20336
rect 54970 20173 55013 20336
rect 54841 20133 55013 20173
rect 57818 19977 57952 21250
rect 59214 21263 59248 21279
rect 59214 21071 59248 21087
rect 59332 21263 59366 21279
rect 59332 21071 59366 21087
rect 59450 21263 59484 21279
rect 59450 21071 59484 21087
rect 59568 21263 59602 21279
rect 59568 21071 59602 21087
rect 59686 21263 59720 21279
rect 59686 21071 59720 21087
rect 59804 21263 59838 21279
rect 59804 21071 59838 21087
rect 59922 21263 59956 21279
rect 59922 21071 59956 21087
rect 60040 21263 60074 21313
rect 60040 21071 60074 21087
rect 60158 21263 60192 21279
rect 60158 21071 60192 21087
rect 60276 21263 60310 21313
rect 61227 21323 61263 21381
rect 61464 21757 61498 21773
rect 61346 21365 61380 21381
rect 61462 21381 61464 21428
rect 61462 21323 61498 21381
rect 61582 21757 61616 21773
rect 61582 21365 61616 21381
rect 61700 21757 61734 21773
rect 61818 21757 61852 21773
rect 61734 21381 61736 21427
rect 61700 21323 61736 21381
rect 61818 21365 61852 21381
rect 63008 21757 63042 21773
rect 63126 21757 63160 21773
rect 63008 21365 63042 21381
rect 63125 21381 63126 21428
rect 63244 21757 63278 21773
rect 63160 21381 63161 21428
rect 62323 21323 62820 21341
rect 61227 21320 62820 21323
rect 61227 21286 62768 21320
rect 62802 21286 62820 21320
rect 61227 21283 62820 21286
rect 63125 21323 63161 21381
rect 63362 21757 63396 21773
rect 63244 21365 63278 21381
rect 63360 21381 63362 21428
rect 63360 21323 63396 21381
rect 63480 21757 63514 21773
rect 63480 21365 63514 21381
rect 63598 21757 63632 21773
rect 63716 21757 63750 21773
rect 64237 21765 64304 21781
rect 63632 21381 63634 21427
rect 63598 21323 63634 21381
rect 63716 21365 63750 21381
rect 64221 21352 64321 21353
rect 64400 21352 66075 21353
rect 64221 21342 66075 21352
rect 64221 21323 65917 21342
rect 63125 21283 65917 21323
rect 61246 21282 62820 21283
rect 63144 21282 65917 21283
rect 61124 21193 61191 21209
rect 61124 21159 61140 21193
rect 61174 21159 61191 21193
rect 61124 21143 61191 21159
rect 60276 21071 60310 21087
rect 60955 21126 60989 21142
rect 60955 21076 60989 21092
rect 61301 21041 61335 21282
rect 62323 21265 62820 21282
rect 61771 21193 61838 21209
rect 61771 21159 61788 21193
rect 61822 21159 61838 21193
rect 61771 21143 61838 21159
rect 63022 21193 63089 21209
rect 63022 21159 63038 21193
rect 63072 21159 63089 21193
rect 63022 21143 63089 21159
rect 62078 21125 62112 21141
rect 61390 21075 61406 21109
rect 61440 21075 61456 21109
rect 61508 21076 61524 21110
rect 61558 21076 61574 21110
rect 62078 21075 62112 21091
rect 62853 21126 62887 21142
rect 62853 21076 62887 21092
rect 63199 21041 63233 21282
rect 64221 21264 65917 21282
rect 66062 21264 66075 21342
rect 64221 21256 66075 21264
rect 64221 21254 64509 21256
rect 64221 21253 64321 21254
rect 63667 21194 63734 21210
rect 63667 21160 63684 21194
rect 63718 21160 63734 21194
rect 63667 21144 63734 21160
rect 63976 21125 64010 21141
rect 63288 21075 63304 21109
rect 63338 21075 63354 21109
rect 63406 21076 63422 21110
rect 63456 21076 63472 21110
rect 63976 21075 64010 21091
rect 59965 20993 59981 21027
rect 60015 20993 60031 21027
rect 60808 21025 60842 21041
rect 59847 20876 59863 20910
rect 59897 20876 59913 20910
rect 59451 20826 59485 20842
rect 59451 20434 59485 20450
rect 59569 20826 59603 20842
rect 59569 20434 59603 20450
rect 59687 20826 59721 20842
rect 59804 20826 59838 20842
rect 59804 20634 59838 20650
rect 59922 20826 59956 20842
rect 60808 20833 60842 20849
rect 60926 21025 60960 21041
rect 60926 20833 60960 20849
rect 61228 21025 61262 21041
rect 59922 20634 59956 20650
rect 61301 21025 61380 21041
rect 61301 20995 61346 21025
rect 61228 20582 61263 20649
rect 61346 20633 61380 20649
rect 61464 21025 61498 21041
rect 61464 20633 61498 20649
rect 61582 21025 61616 21041
rect 61700 21025 61734 21041
rect 62106 21025 62140 21041
rect 62106 20833 62140 20849
rect 62224 21025 62258 21041
rect 62224 20833 62258 20849
rect 62706 21025 62740 21041
rect 62706 20833 62740 20849
rect 62824 21025 62858 21041
rect 62824 20833 62858 20849
rect 63126 21025 63160 21041
rect 61582 20633 61616 20649
rect 61699 20582 61734 20649
rect 61228 20547 61734 20582
rect 63199 21025 63278 21041
rect 63199 20995 63244 21025
rect 63126 20582 63161 20649
rect 63244 20633 63278 20649
rect 63362 21025 63396 21041
rect 63362 20633 63396 20649
rect 63480 21025 63514 21041
rect 63598 21025 63632 21041
rect 64004 21025 64038 21041
rect 64004 20833 64038 20849
rect 64122 21025 64156 21041
rect 64122 20833 64156 20849
rect 63480 20633 63514 20649
rect 63597 20582 63632 20649
rect 63126 20547 63632 20582
rect 59687 20434 59721 20450
rect 59974 20500 60223 20543
rect 59974 20410 60021 20500
rect 60184 20410 60223 20500
rect 59494 20366 59510 20400
rect 59544 20366 59560 20400
rect 59612 20366 59628 20400
rect 59662 20366 59678 20400
rect 59974 20371 60223 20410
rect 61399 20340 61571 20387
rect 61399 20177 61438 20340
rect 61528 20177 61571 20340
rect 61399 20137 61571 20177
rect 57818 19976 66583 19977
rect 57818 19962 66589 19976
rect 57818 19890 66434 19962
rect 66569 19890 66589 19962
rect 57818 19882 66589 19890
rect 57818 19878 66583 19882
rect 57818 19874 57952 19878
rect 51287 19812 67151 19828
rect 51287 19722 67002 19812
rect 67132 19722 67151 19812
rect 51287 19705 67151 19722
rect 68599 19641 68722 22235
rect 68936 22235 71573 22317
rect 68936 22091 69053 22235
rect 71485 22200 71573 22235
rect 71485 22151 71499 22200
rect 71559 22151 71573 22200
rect 71485 22135 71573 22151
rect 68936 20363 69055 22091
rect 70635 22027 70725 22061
rect 70901 22027 70917 22061
rect 70635 21825 70674 22027
rect 71199 21956 71284 21972
rect 70709 21909 70725 21943
rect 70901 21909 70991 21943
rect 70635 21791 70725 21825
rect 70901 21791 70917 21825
rect 70952 21707 70991 21909
rect 71199 21896 71216 21956
rect 71271 21896 71284 21956
rect 71199 21880 71284 21896
rect 70709 21673 70725 21707
rect 70901 21673 70991 21707
rect 70433 21586 70525 21620
rect 70901 21586 70917 21620
rect 70433 21384 70472 21586
rect 70509 21468 70525 21502
rect 70901 21468 70991 21502
rect 70433 21350 70525 21384
rect 70901 21350 70917 21384
rect 70952 21266 70991 21468
rect 70509 21232 70525 21266
rect 70901 21232 70991 21266
rect 70434 21119 70525 21153
rect 70901 21119 70917 21153
rect 70434 20917 70473 21119
rect 70952 21035 70991 21232
rect 71842 21193 71858 21227
rect 72034 21193 72050 21227
rect 71842 21075 71858 21109
rect 72034 21075 72050 21109
rect 71846 21035 72046 21075
rect 70509 21001 70525 21035
rect 70901 21001 70991 21035
rect 70237 20875 70347 20891
rect 70434 20883 70525 20917
rect 70901 20883 70917 20917
rect 70237 20679 70255 20875
rect 70331 20679 70347 20875
rect 70952 20799 70991 21001
rect 71487 20989 71572 21005
rect 71842 21001 71858 21035
rect 72234 21001 72250 21035
rect 71100 20941 71116 20975
rect 71150 20941 71166 20975
rect 71487 20929 71500 20989
rect 71555 20929 71572 20989
rect 71487 20913 71572 20929
rect 70509 20765 70525 20799
rect 70901 20765 70991 20799
rect 71202 20871 71287 20887
rect 71842 20883 71858 20917
rect 72234 20883 72250 20917
rect 71202 20811 71215 20871
rect 71270 20811 71287 20871
rect 72483 20817 72569 20833
rect 71202 20795 71287 20811
rect 71842 20765 71858 20799
rect 72234 20765 72250 20799
rect 72335 20798 72369 20814
rect 70237 20663 70347 20679
rect 70434 20647 70525 20681
rect 70901 20647 70917 20681
rect 70434 20445 70473 20647
rect 70952 20563 70991 20765
rect 72335 20748 72369 20764
rect 72483 20795 72501 20817
rect 71720 20706 71736 20740
rect 71770 20706 71786 20740
rect 72483 20737 72487 20795
rect 72483 20713 72501 20737
rect 72547 20713 72569 20817
rect 72483 20697 72569 20713
rect 71842 20647 71858 20681
rect 72234 20647 72250 20681
rect 71330 20587 71346 20621
rect 71380 20587 71396 20621
rect 70509 20529 70525 20563
rect 70901 20529 70991 20563
rect 71842 20529 71858 20563
rect 72234 20529 72250 20563
rect 70434 20411 70525 20445
rect 70901 20411 70917 20445
rect 68936 19847 69054 20363
rect 70952 20326 70991 20529
rect 71846 20485 72046 20529
rect 71842 20451 71858 20485
rect 72034 20451 72050 20485
rect 71842 20333 71858 20367
rect 72034 20333 72050 20367
rect 70509 20292 70525 20326
rect 70901 20292 70991 20326
rect 70434 20174 70525 20208
rect 70901 20174 70917 20208
rect 70434 19972 70473 20174
rect 70952 20090 70991 20292
rect 70509 20056 70525 20090
rect 70901 20056 70991 20090
rect 70434 19938 70525 19972
rect 70901 19938 70917 19972
rect 44765 19520 68722 19641
rect 44765 19519 68718 19520
rect 44765 19517 44904 19519
rect 68932 19483 69056 19847
rect 70709 19819 70725 19853
rect 70901 19819 70994 19853
rect 39573 19381 39796 19457
rect 39573 19232 39650 19381
rect 39717 19232 39796 19381
rect 39573 19126 39796 19232
rect 40720 19381 40943 19457
rect 40720 19232 40797 19381
rect 40864 19232 40943 19381
rect 40446 19167 40480 19183
rect 40446 19117 40480 19133
rect 40720 19126 40943 19232
rect 43202 19327 43425 19403
rect 43202 19178 43279 19327
rect 43346 19178 43425 19327
rect 41576 19161 41610 19177
rect 41576 19111 41610 19127
rect 43202 19072 43425 19178
rect 46131 19377 46354 19453
rect 46131 19228 46208 19377
rect 46275 19228 46354 19377
rect 46131 19122 46354 19228
rect 47278 19377 47501 19453
rect 47278 19228 47355 19377
rect 47422 19228 47501 19377
rect 47004 19163 47038 19179
rect 47004 19113 47038 19129
rect 47278 19122 47501 19228
rect 49760 19323 49983 19399
rect 49760 19174 49837 19323
rect 49904 19174 49983 19323
rect 48134 19157 48168 19173
rect 48134 19107 48168 19123
rect 49760 19068 49983 19174
rect 52665 19382 52888 19458
rect 52665 19233 52742 19382
rect 52809 19233 52888 19382
rect 52665 19127 52888 19233
rect 53812 19382 54035 19458
rect 53812 19233 53889 19382
rect 53956 19233 54035 19382
rect 53538 19168 53572 19184
rect 53538 19118 53572 19134
rect 53812 19127 54035 19233
rect 56294 19328 56517 19404
rect 56294 19179 56371 19328
rect 56438 19179 56517 19328
rect 54668 19162 54702 19178
rect 54668 19112 54702 19128
rect 56294 19073 56517 19179
rect 59178 19385 59401 19461
rect 59178 19236 59255 19385
rect 59322 19236 59401 19385
rect 59178 19130 59401 19236
rect 60325 19385 60548 19461
rect 64602 19441 69056 19483
rect 70638 19701 70725 19735
rect 70901 19701 70917 19735
rect 70638 19499 70675 19701
rect 70955 19617 70994 19819
rect 70709 19583 70725 19617
rect 70901 19583 70994 19617
rect 71075 19665 71109 19681
rect 71075 19615 71109 19631
rect 70638 19465 70725 19499
rect 70901 19465 70917 19499
rect 60325 19236 60402 19385
rect 60469 19236 60548 19385
rect 60051 19171 60085 19187
rect 60051 19121 60085 19137
rect 60325 19130 60548 19236
rect 62807 19331 63030 19407
rect 62807 19182 62884 19331
rect 62951 19182 63030 19331
rect 61181 19165 61215 19181
rect 61181 19115 61215 19131
rect 62807 19076 63030 19182
rect 64602 19358 69058 19441
rect 40446 19047 40480 19063
rect 39611 18989 39645 19005
rect 39611 18597 39645 18613
rect 39729 18989 39763 19005
rect 39729 18597 39763 18613
rect 39847 18989 39881 19005
rect 39847 18597 39881 18613
rect 39965 18989 39999 19005
rect 39965 18597 39999 18613
rect 40083 18989 40117 19005
rect 40083 18597 40117 18613
rect 40201 18989 40235 19005
rect 40201 18597 40235 18613
rect 40319 18989 40353 19005
rect 40446 18997 40480 19013
rect 41576 19043 41610 19059
rect 40319 18597 40353 18613
rect 40753 18985 40787 19001
rect 40753 18593 40787 18609
rect 40871 18985 40905 19001
rect 40871 18593 40905 18609
rect 40989 18985 41023 19001
rect 40989 18593 41023 18609
rect 41107 18985 41141 19001
rect 41107 18593 41141 18609
rect 41225 18985 41259 19001
rect 41225 18593 41259 18609
rect 41343 18985 41377 19001
rect 41343 18593 41377 18609
rect 41461 18985 41495 19001
rect 41576 18993 41610 19009
rect 47004 19043 47038 19059
rect 42724 18963 42994 18997
rect 42724 18913 42758 18963
rect 42724 18721 42758 18737
rect 42842 18913 42876 18929
rect 42842 18721 42876 18737
rect 42960 18913 42994 18963
rect 46169 18985 46203 19001
rect 42960 18721 42994 18737
rect 43078 18913 43112 18929
rect 43078 18721 43112 18737
rect 43196 18913 43230 18929
rect 43196 18721 43230 18737
rect 43314 18913 43348 18929
rect 43314 18721 43348 18737
rect 43432 18913 43466 18929
rect 43432 18721 43466 18737
rect 43550 18913 43584 18929
rect 43550 18721 43584 18737
rect 43668 18913 43702 18929
rect 43668 18721 43702 18737
rect 43786 18913 43820 18929
rect 43786 18721 43820 18737
rect 43003 18643 43019 18677
rect 43053 18643 43069 18677
rect 41461 18593 41495 18609
rect 46169 18593 46203 18609
rect 46287 18985 46321 19001
rect 46287 18593 46321 18609
rect 46405 18985 46439 19001
rect 46405 18593 46439 18609
rect 46523 18985 46557 19001
rect 46523 18593 46557 18609
rect 46641 18985 46675 19001
rect 46641 18593 46675 18609
rect 46759 18985 46793 19001
rect 46759 18593 46793 18609
rect 46877 18985 46911 19001
rect 47004 18993 47038 19009
rect 48134 19039 48168 19055
rect 53538 19048 53572 19064
rect 46877 18593 46911 18609
rect 47311 18981 47345 18997
rect 47311 18589 47345 18605
rect 47429 18981 47463 18997
rect 47429 18589 47463 18605
rect 47547 18981 47581 18997
rect 47547 18589 47581 18605
rect 47665 18981 47699 18997
rect 47665 18589 47699 18605
rect 47783 18981 47817 18997
rect 47783 18589 47817 18605
rect 47901 18981 47935 18997
rect 47901 18589 47935 18605
rect 48019 18981 48053 18997
rect 48134 18989 48168 19005
rect 49282 18959 49552 18993
rect 49282 18909 49316 18959
rect 49282 18717 49316 18733
rect 49400 18909 49434 18925
rect 49400 18717 49434 18733
rect 49518 18909 49552 18959
rect 52703 18990 52737 19006
rect 49518 18717 49552 18733
rect 49636 18909 49670 18925
rect 49636 18717 49670 18733
rect 49754 18909 49788 18925
rect 49754 18717 49788 18733
rect 49872 18909 49906 18925
rect 49872 18717 49906 18733
rect 49990 18909 50024 18925
rect 49990 18717 50024 18733
rect 50108 18909 50142 18925
rect 50108 18717 50142 18733
rect 50226 18909 50260 18925
rect 50226 18717 50260 18733
rect 50344 18909 50378 18925
rect 50344 18717 50378 18733
rect 49561 18639 49577 18673
rect 49611 18639 49627 18673
rect 48019 18589 48053 18605
rect 52703 18598 52737 18614
rect 52821 18990 52855 19006
rect 52821 18598 52855 18614
rect 52939 18990 52973 19006
rect 52939 18598 52973 18614
rect 53057 18990 53091 19006
rect 53057 18598 53091 18614
rect 53175 18990 53209 19006
rect 53175 18598 53209 18614
rect 53293 18990 53327 19006
rect 53293 18598 53327 18614
rect 53411 18990 53445 19006
rect 53538 18998 53572 19014
rect 54668 19044 54702 19060
rect 53411 18598 53445 18614
rect 53845 18986 53879 19002
rect 53845 18594 53879 18610
rect 53963 18986 53997 19002
rect 53963 18594 53997 18610
rect 54081 18986 54115 19002
rect 54081 18594 54115 18610
rect 54199 18986 54233 19002
rect 54199 18594 54233 18610
rect 54317 18986 54351 19002
rect 54317 18594 54351 18610
rect 54435 18986 54469 19002
rect 54435 18594 54469 18610
rect 54553 18986 54587 19002
rect 54668 18994 54702 19010
rect 60051 19051 60085 19067
rect 55816 18964 56086 18998
rect 55816 18914 55850 18964
rect 55816 18722 55850 18738
rect 55934 18914 55968 18930
rect 55934 18722 55968 18738
rect 56052 18914 56086 18964
rect 59216 18993 59250 19009
rect 56052 18722 56086 18738
rect 56170 18914 56204 18930
rect 56170 18722 56204 18738
rect 56288 18914 56322 18930
rect 56288 18722 56322 18738
rect 56406 18914 56440 18930
rect 56406 18722 56440 18738
rect 56524 18914 56558 18930
rect 56524 18722 56558 18738
rect 56642 18914 56676 18930
rect 56642 18722 56676 18738
rect 56760 18914 56794 18930
rect 56760 18722 56794 18738
rect 56878 18914 56912 18930
rect 56878 18722 56912 18738
rect 56095 18644 56111 18678
rect 56145 18644 56161 18678
rect 54553 18594 54587 18610
rect 59216 18601 59250 18617
rect 59334 18993 59368 19009
rect 59334 18601 59368 18617
rect 59452 18993 59486 19009
rect 59452 18601 59486 18617
rect 59570 18993 59604 19009
rect 59570 18601 59604 18617
rect 59688 18993 59722 19009
rect 59688 18601 59722 18617
rect 59806 18993 59840 19009
rect 59806 18601 59840 18617
rect 59924 18993 59958 19009
rect 60051 19001 60085 19017
rect 61181 19047 61215 19063
rect 59924 18601 59958 18617
rect 60358 18989 60392 19005
rect 60358 18597 60392 18613
rect 60476 18989 60510 19005
rect 60476 18597 60510 18613
rect 60594 18989 60628 19005
rect 60594 18597 60628 18613
rect 60712 18989 60746 19005
rect 60712 18597 60746 18613
rect 60830 18989 60864 19005
rect 60830 18597 60864 18613
rect 60948 18989 60982 19005
rect 60948 18597 60982 18613
rect 61066 18989 61100 19005
rect 61181 18997 61215 19013
rect 62329 18967 62599 19001
rect 62329 18917 62363 18967
rect 62329 18725 62363 18741
rect 62447 18917 62481 18933
rect 62447 18725 62481 18741
rect 62565 18917 62599 18967
rect 62565 18725 62599 18741
rect 62683 18917 62717 18933
rect 62683 18725 62717 18741
rect 62801 18917 62835 18933
rect 62801 18725 62835 18741
rect 62919 18917 62953 18933
rect 62919 18725 62953 18741
rect 63037 18917 63071 18933
rect 63037 18725 63071 18741
rect 63155 18917 63189 18933
rect 63155 18725 63189 18741
rect 63273 18917 63307 18933
rect 63273 18725 63307 18741
rect 63391 18917 63425 18933
rect 63391 18725 63425 18741
rect 62608 18647 62624 18681
rect 62658 18647 62674 18681
rect 61066 18597 61100 18613
rect 43121 18526 43137 18560
rect 43171 18526 43187 18560
rect 49679 18522 49695 18556
rect 49729 18522 49745 18556
rect 56213 18527 56229 18561
rect 56263 18527 56279 18561
rect 62726 18530 62742 18564
rect 62776 18530 62792 18564
rect 43078 18476 43112 18492
rect 40098 18257 40114 18291
rect 40148 18257 40164 18291
rect 41240 18253 41256 18287
rect 41290 18253 41306 18287
rect 43078 18284 43112 18300
rect 43196 18476 43230 18492
rect 43196 18284 43230 18300
rect 43313 18476 43347 18492
rect 39536 18206 39570 18222
rect 39536 18014 39570 18030
rect 39654 18206 39688 18222
rect 39654 18014 39688 18030
rect 39772 18206 39806 18222
rect 39772 18014 39806 18030
rect 39890 18206 39924 18222
rect 39890 18014 39924 18030
rect 40055 18206 40089 18222
rect 40055 18014 40089 18030
rect 40173 18206 40207 18222
rect 40173 18014 40207 18030
rect 40291 18206 40325 18222
rect 40291 18014 40325 18030
rect 40409 18206 40443 18222
rect 40409 18014 40443 18030
rect 40678 18202 40712 18218
rect 40678 18010 40712 18026
rect 40796 18202 40830 18218
rect 40796 18010 40830 18026
rect 40914 18202 40948 18218
rect 40914 18010 40948 18026
rect 41032 18202 41066 18218
rect 41032 18010 41066 18026
rect 41197 18202 41231 18218
rect 41197 18010 41231 18026
rect 41315 18202 41349 18218
rect 41315 18010 41349 18026
rect 41433 18202 41467 18218
rect 41433 18010 41467 18026
rect 41551 18202 41585 18218
rect 41551 18010 41585 18026
rect 42811 18150 43060 18193
rect 42811 18060 42850 18150
rect 43013 18060 43060 18150
rect 43313 18084 43347 18100
rect 43431 18476 43465 18492
rect 43431 18084 43465 18100
rect 43549 18476 43583 18492
rect 49636 18472 49670 18488
rect 46656 18253 46672 18287
rect 46706 18253 46722 18287
rect 47798 18249 47814 18283
rect 47848 18249 47864 18283
rect 49636 18280 49670 18296
rect 49754 18472 49788 18488
rect 49754 18280 49788 18296
rect 49871 18472 49905 18488
rect 43549 18084 43583 18100
rect 46094 18202 46128 18218
rect 42811 18021 43060 18060
rect 43356 18016 43372 18050
rect 43406 18016 43422 18050
rect 43474 18016 43490 18050
rect 43524 18016 43540 18050
rect 46094 18010 46128 18026
rect 46212 18202 46246 18218
rect 46212 18010 46246 18026
rect 46330 18202 46364 18218
rect 46330 18010 46364 18026
rect 46448 18202 46482 18218
rect 46448 18010 46482 18026
rect 46613 18202 46647 18218
rect 46613 18010 46647 18026
rect 46731 18202 46765 18218
rect 46731 18010 46765 18026
rect 46849 18202 46883 18218
rect 46849 18010 46883 18026
rect 46967 18202 47001 18218
rect 46967 18010 47001 18026
rect 47236 18198 47270 18214
rect 47236 18006 47270 18022
rect 47354 18198 47388 18214
rect 47354 18006 47388 18022
rect 47472 18198 47506 18214
rect 47472 18006 47506 18022
rect 47590 18198 47624 18214
rect 47590 18006 47624 18022
rect 47755 18198 47789 18214
rect 47755 18006 47789 18022
rect 47873 18198 47907 18214
rect 47873 18006 47907 18022
rect 47991 18198 48025 18214
rect 47991 18006 48025 18022
rect 48109 18198 48143 18214
rect 48109 18006 48143 18022
rect 49369 18146 49618 18189
rect 49369 18056 49408 18146
rect 49571 18056 49618 18146
rect 49871 18080 49905 18096
rect 49989 18472 50023 18488
rect 49989 18080 50023 18096
rect 50107 18472 50141 18488
rect 56170 18477 56204 18493
rect 53190 18258 53206 18292
rect 53240 18258 53256 18292
rect 54332 18254 54348 18288
rect 54382 18254 54398 18288
rect 56170 18285 56204 18301
rect 56288 18477 56322 18493
rect 56288 18285 56322 18301
rect 56405 18477 56439 18493
rect 50107 18080 50141 18096
rect 52628 18207 52662 18223
rect 49369 18017 49618 18056
rect 49914 18012 49930 18046
rect 49964 18012 49980 18046
rect 50032 18012 50048 18046
rect 50082 18012 50098 18046
rect 52628 18015 52662 18031
rect 52746 18207 52780 18223
rect 52746 18015 52780 18031
rect 52864 18207 52898 18223
rect 52864 18015 52898 18031
rect 52982 18207 53016 18223
rect 52982 18015 53016 18031
rect 53147 18207 53181 18223
rect 53147 18015 53181 18031
rect 53265 18207 53299 18223
rect 53265 18015 53299 18031
rect 53383 18207 53417 18223
rect 53383 18015 53417 18031
rect 53501 18207 53535 18223
rect 53501 18015 53535 18031
rect 53770 18203 53804 18219
rect 53770 18011 53804 18027
rect 53888 18203 53922 18219
rect 53888 18011 53922 18027
rect 54006 18203 54040 18219
rect 54006 18011 54040 18027
rect 54124 18203 54158 18219
rect 54124 18011 54158 18027
rect 54289 18203 54323 18219
rect 54289 18011 54323 18027
rect 54407 18203 54441 18219
rect 54407 18011 54441 18027
rect 54525 18203 54559 18219
rect 54525 18011 54559 18027
rect 54643 18203 54677 18219
rect 54643 18011 54677 18027
rect 55903 18151 56152 18194
rect 55903 18061 55942 18151
rect 56105 18061 56152 18151
rect 56405 18085 56439 18101
rect 56523 18477 56557 18493
rect 56523 18085 56557 18101
rect 56641 18477 56675 18493
rect 62683 18480 62717 18496
rect 59703 18261 59719 18295
rect 59753 18261 59769 18295
rect 60845 18257 60861 18291
rect 60895 18257 60911 18291
rect 62683 18288 62717 18304
rect 62801 18480 62835 18496
rect 62801 18288 62835 18304
rect 62918 18480 62952 18496
rect 56641 18085 56675 18101
rect 59141 18210 59175 18226
rect 55903 18022 56152 18061
rect 56448 18017 56464 18051
rect 56498 18017 56514 18051
rect 56566 18017 56582 18051
rect 56616 18017 56632 18051
rect 59141 18018 59175 18034
rect 59259 18210 59293 18226
rect 59259 18018 59293 18034
rect 59377 18210 59411 18226
rect 59377 18018 59411 18034
rect 59495 18210 59529 18226
rect 59495 18018 59529 18034
rect 59660 18210 59694 18226
rect 59660 18018 59694 18034
rect 59778 18210 59812 18226
rect 59778 18018 59812 18034
rect 59896 18210 59930 18226
rect 59896 18018 59930 18034
rect 60014 18210 60048 18226
rect 60014 18018 60048 18034
rect 60283 18206 60317 18222
rect 60283 18014 60317 18030
rect 60401 18206 60435 18222
rect 60401 18014 60435 18030
rect 60519 18206 60553 18222
rect 60519 18014 60553 18030
rect 60637 18206 60671 18222
rect 60637 18014 60671 18030
rect 60802 18206 60836 18222
rect 60802 18014 60836 18030
rect 60920 18206 60954 18222
rect 60920 18014 60954 18030
rect 61038 18206 61072 18222
rect 61038 18014 61072 18030
rect 61156 18206 61190 18222
rect 61156 18014 61190 18030
rect 62416 18154 62665 18197
rect 62416 18064 62455 18154
rect 62618 18064 62665 18154
rect 62918 18088 62952 18104
rect 63036 18480 63070 18496
rect 63036 18088 63070 18104
rect 63154 18480 63188 18496
rect 63154 18088 63188 18104
rect 62416 18025 62665 18064
rect 62961 18020 62977 18054
rect 63011 18020 63027 18054
rect 63079 18020 63095 18054
rect 63129 18020 63145 18054
rect 40256 17777 40428 17824
rect 40256 17614 40299 17777
rect 40389 17614 40428 17777
rect 40256 17575 40428 17614
rect 41398 17779 41570 17826
rect 41398 17616 41441 17779
rect 41531 17616 41570 17779
rect 46814 17773 46986 17820
rect 41398 17577 41570 17616
rect 43188 17677 43411 17753
rect 43188 17528 43265 17677
rect 43332 17528 43411 17677
rect 43188 17422 43411 17528
rect 44457 17571 44746 17618
rect 46814 17610 46857 17773
rect 46947 17610 46986 17773
rect 46814 17571 46986 17610
rect 47956 17775 48128 17822
rect 47956 17612 47999 17775
rect 48089 17612 48128 17775
rect 53348 17778 53520 17825
rect 47956 17573 48128 17612
rect 49746 17673 49969 17749
rect 44457 17462 44496 17571
rect 44607 17462 44746 17571
rect 44457 17450 44746 17462
rect 39475 17334 39700 17410
rect 39475 17185 39554 17334
rect 39621 17185 39700 17334
rect 39475 17079 39700 17185
rect 42710 17313 42980 17347
rect 42710 17263 42744 17313
rect 42710 17071 42744 17087
rect 42828 17263 42862 17279
rect 42828 17071 42862 17087
rect 42946 17263 42980 17313
rect 42946 17071 42980 17087
rect 43064 17263 43098 17279
rect 43064 17071 43098 17087
rect 43182 17263 43216 17279
rect 43182 17071 43216 17087
rect 43300 17263 43334 17279
rect 43300 17071 43334 17087
rect 43418 17263 43452 17279
rect 43418 17071 43452 17087
rect 43536 17263 43570 17279
rect 43536 17071 43570 17087
rect 43654 17263 43688 17279
rect 43654 17071 43688 17087
rect 43772 17263 43806 17279
rect 43772 17071 43806 17087
rect 42989 16993 43005 17027
rect 43039 16993 43055 17027
rect 39336 16899 39606 16934
rect 39218 16846 39252 16862
rect 38735 16646 38769 16662
rect 38735 16454 38769 16470
rect 38853 16646 38887 16662
rect 38853 16454 38887 16470
rect 38971 16646 39005 16662
rect 38971 16454 39005 16470
rect 39089 16646 39123 16662
rect 39089 16454 39123 16470
rect 39218 16454 39252 16470
rect 39336 16846 39370 16899
rect 39336 16454 39370 16470
rect 39454 16846 39488 16862
rect 39454 16454 39488 16470
rect 39572 16846 39606 16899
rect 41234 16899 41504 16934
rect 39572 16454 39606 16470
rect 39690 16846 39724 16862
rect 39690 16454 39724 16470
rect 39808 16846 39842 16862
rect 39808 16454 39842 16470
rect 39926 16846 39960 16862
rect 41116 16846 41150 16862
rect 40174 16700 40444 16735
rect 39926 16454 39960 16470
rect 40056 16646 40090 16662
rect 40056 16454 40090 16470
rect 40174 16646 40208 16700
rect 40174 16454 40208 16470
rect 40292 16646 40326 16662
rect 40292 16454 40326 16470
rect 40410 16646 40444 16700
rect 40410 16454 40444 16470
rect 40633 16646 40667 16662
rect 40633 16454 40667 16470
rect 40751 16646 40785 16662
rect 40751 16454 40785 16470
rect 40869 16646 40903 16662
rect 40869 16454 40903 16470
rect 40987 16646 41021 16662
rect 40987 16454 41021 16470
rect 41116 16454 41150 16470
rect 41234 16846 41268 16899
rect 41234 16454 41268 16470
rect 41352 16846 41386 16862
rect 41352 16454 41386 16470
rect 41470 16846 41504 16899
rect 43107 16876 43123 16910
rect 43157 16876 43173 16910
rect 41470 16454 41504 16470
rect 41588 16846 41622 16862
rect 41588 16454 41622 16470
rect 41706 16846 41740 16862
rect 41706 16454 41740 16470
rect 41824 16846 41858 16862
rect 43064 16826 43098 16842
rect 42072 16700 42342 16735
rect 41824 16454 41858 16470
rect 41954 16646 41988 16662
rect 41954 16454 41988 16470
rect 42072 16646 42106 16700
rect 42072 16454 42106 16470
rect 42190 16646 42224 16662
rect 42190 16454 42224 16470
rect 42308 16646 42342 16700
rect 43064 16634 43098 16650
rect 43182 16826 43216 16842
rect 43182 16634 43216 16650
rect 43299 16826 43333 16842
rect 42308 16454 42342 16470
rect 42797 16500 43046 16543
rect 42797 16410 42836 16500
rect 42999 16410 43046 16500
rect 43299 16434 43333 16450
rect 43417 16826 43451 16842
rect 43417 16434 43451 16450
rect 43535 16826 43569 16842
rect 43535 16434 43569 16450
rect 42797 16371 43046 16410
rect 43342 16366 43358 16400
rect 43392 16366 43408 16400
rect 43460 16366 43476 16400
rect 43510 16366 43526 16400
rect 40844 16232 40878 16248
rect 38721 16211 38788 16227
rect 38721 16177 38737 16211
rect 38771 16177 38788 16211
rect 40844 16182 40878 16198
rect 38721 16161 38788 16177
rect 39275 16153 39309 16169
rect 39393 16153 39427 16169
rect 39275 15761 39309 15777
rect 39391 15777 39393 15823
rect 38704 15748 38804 15749
rect 38648 15719 38804 15748
rect 39391 15719 39427 15777
rect 39511 16153 39545 16169
rect 39511 15761 39545 15777
rect 39629 16153 39663 16169
rect 39747 16153 39781 16169
rect 39663 15777 39665 15824
rect 39629 15719 39665 15777
rect 39865 16153 39899 16169
rect 39747 15761 39781 15777
rect 39864 15777 39865 15824
rect 39983 16153 40017 16169
rect 39899 15777 39900 15824
rect 39864 15719 39900 15777
rect 39983 15761 40017 15777
rect 41173 16153 41207 16169
rect 41291 16153 41325 16169
rect 41173 15761 41207 15777
rect 41289 15777 41291 15823
rect 38648 15679 39900 15719
rect 40205 15719 40702 15737
rect 41289 15719 41325 15777
rect 41409 16153 41443 16169
rect 41409 15761 41443 15777
rect 41527 16153 41561 16169
rect 41645 16153 41679 16169
rect 41561 15777 41563 15824
rect 41527 15719 41563 15777
rect 41763 16153 41797 16169
rect 41645 15761 41679 15777
rect 41762 15777 41763 15824
rect 41881 16153 41915 16169
rect 41797 15777 41798 15824
rect 41762 15719 41798 15777
rect 43193 16073 43416 16149
rect 43193 15924 43270 16073
rect 43337 15924 43416 16073
rect 43193 15818 43416 15924
rect 41881 15761 41915 15777
rect 40205 15716 41798 15719
rect 40205 15682 40223 15716
rect 40257 15682 41798 15716
rect 40205 15679 41798 15682
rect 42715 15709 42985 15743
rect 38648 15678 39881 15679
rect 40205 15678 41779 15679
rect 38648 15650 38804 15678
rect 38704 15649 38804 15650
rect 39291 15590 39358 15606
rect 39291 15556 39307 15590
rect 39341 15556 39358 15590
rect 39291 15540 39358 15556
rect 39015 15521 39049 15537
rect 39015 15471 39049 15487
rect 39553 15472 39569 15506
rect 39603 15472 39619 15506
rect 39671 15471 39687 15505
rect 39721 15471 39737 15505
rect 39792 15437 39826 15678
rect 40205 15661 40702 15678
rect 39936 15589 40003 15605
rect 39936 15555 39953 15589
rect 39987 15555 40003 15589
rect 39936 15539 40003 15555
rect 41187 15589 41254 15605
rect 41187 15555 41203 15589
rect 41237 15555 41254 15589
rect 41187 15539 41254 15555
rect 40138 15522 40172 15538
rect 40138 15472 40172 15488
rect 40913 15521 40947 15537
rect 40913 15471 40947 15487
rect 41451 15472 41467 15506
rect 41501 15472 41517 15506
rect 41569 15471 41585 15505
rect 41619 15471 41635 15505
rect 41690 15437 41724 15678
rect 42715 15659 42749 15709
rect 41834 15589 41901 15605
rect 41834 15555 41851 15589
rect 41885 15555 41901 15589
rect 41834 15539 41901 15555
rect 42036 15522 42070 15538
rect 42036 15472 42070 15488
rect 42715 15467 42749 15483
rect 42833 15659 42867 15675
rect 42833 15467 42867 15483
rect 42951 15659 42985 15709
rect 42951 15467 42985 15483
rect 43069 15659 43103 15675
rect 43069 15467 43103 15483
rect 43187 15659 43221 15675
rect 43187 15467 43221 15483
rect 43305 15659 43339 15675
rect 43305 15467 43339 15483
rect 43423 15659 43457 15675
rect 43423 15467 43457 15483
rect 43541 15659 43575 15675
rect 43541 15467 43575 15483
rect 43659 15659 43693 15675
rect 43659 15467 43693 15483
rect 43777 15659 43811 15675
rect 43777 15467 43811 15483
rect 38869 15421 38903 15437
rect 38869 15229 38903 15245
rect 38987 15421 39021 15437
rect 38987 15229 39021 15245
rect 39393 15421 39427 15437
rect 39511 15421 39545 15437
rect 39393 14978 39428 15045
rect 39511 15029 39545 15045
rect 39629 15421 39663 15437
rect 39629 15029 39663 15045
rect 39747 15421 39826 15437
rect 39781 15391 39826 15421
rect 39865 15421 39899 15437
rect 40167 15421 40201 15437
rect 40167 15229 40201 15245
rect 40285 15421 40319 15437
rect 40285 15229 40319 15245
rect 40767 15421 40801 15437
rect 40767 15229 40801 15245
rect 40885 15421 40919 15437
rect 40885 15229 40919 15245
rect 41291 15421 41325 15437
rect 39747 15029 39781 15045
rect 39864 14978 39899 15045
rect 39393 14943 39899 14978
rect 41409 15421 41443 15437
rect 41291 14978 41326 15045
rect 41409 15029 41443 15045
rect 41527 15421 41561 15437
rect 41527 15029 41561 15045
rect 41645 15421 41724 15437
rect 41679 15391 41724 15421
rect 41763 15421 41797 15437
rect 42065 15421 42099 15437
rect 42065 15229 42099 15245
rect 42183 15421 42217 15437
rect 42994 15389 43010 15423
rect 43044 15389 43060 15423
rect 43112 15272 43128 15306
rect 43162 15272 43178 15306
rect 42183 15229 42217 15245
rect 41645 15029 41679 15045
rect 41762 14978 41797 15045
rect 43069 15222 43103 15238
rect 43069 15030 43103 15046
rect 43187 15222 43221 15238
rect 43187 15030 43221 15046
rect 43304 15222 43338 15238
rect 41291 14943 41797 14978
rect 42802 14896 43051 14939
rect 42802 14806 42841 14896
rect 43004 14806 43051 14896
rect 43304 14830 43338 14846
rect 43422 15222 43456 15238
rect 43422 14830 43456 14846
rect 43540 15222 43574 15238
rect 43540 14830 43574 14846
rect 41454 14736 41626 14783
rect 42802 14767 43051 14806
rect 43347 14762 43363 14796
rect 43397 14762 43413 14796
rect 43465 14762 43481 14796
rect 43515 14762 43531 14796
rect 41454 14573 41497 14736
rect 41587 14573 41626 14736
rect 41454 14533 41626 14573
rect 44609 12703 44746 17450
rect 49746 17524 49823 17673
rect 49890 17524 49969 17673
rect 49746 17418 49969 17524
rect 51013 17559 51310 17617
rect 53348 17615 53391 17778
rect 53481 17615 53520 17778
rect 53348 17576 53520 17615
rect 54490 17780 54662 17827
rect 54490 17617 54533 17780
rect 54623 17617 54662 17780
rect 59861 17781 60033 17828
rect 54490 17578 54662 17617
rect 56280 17678 56503 17754
rect 51013 17462 51059 17559
rect 51162 17462 51310 17559
rect 51013 17446 51310 17462
rect 46033 17330 46258 17406
rect 46033 17181 46112 17330
rect 46179 17181 46258 17330
rect 46033 17075 46258 17181
rect 49268 17309 49538 17343
rect 49268 17259 49302 17309
rect 49268 17067 49302 17083
rect 49386 17259 49420 17275
rect 49386 17067 49420 17083
rect 49504 17259 49538 17309
rect 49504 17067 49538 17083
rect 49622 17259 49656 17275
rect 49622 17067 49656 17083
rect 49740 17259 49774 17275
rect 49740 17067 49774 17083
rect 49858 17259 49892 17275
rect 49858 17067 49892 17083
rect 49976 17259 50010 17275
rect 49976 17067 50010 17083
rect 50094 17259 50128 17275
rect 50094 17067 50128 17083
rect 50212 17259 50246 17275
rect 50212 17067 50246 17083
rect 50330 17259 50364 17275
rect 50330 17067 50364 17083
rect 49547 16989 49563 17023
rect 49597 16989 49613 17023
rect 45894 16895 46164 16930
rect 45776 16842 45810 16858
rect 45293 16642 45327 16658
rect 45293 16450 45327 16466
rect 45411 16642 45445 16658
rect 45411 16450 45445 16466
rect 45529 16642 45563 16658
rect 45529 16450 45563 16466
rect 45647 16642 45681 16658
rect 45647 16450 45681 16466
rect 45776 16450 45810 16466
rect 45894 16842 45928 16895
rect 45894 16450 45928 16466
rect 46012 16842 46046 16858
rect 46012 16450 46046 16466
rect 46130 16842 46164 16895
rect 47792 16895 48062 16930
rect 46130 16450 46164 16466
rect 46248 16842 46282 16858
rect 46248 16450 46282 16466
rect 46366 16842 46400 16858
rect 46366 16450 46400 16466
rect 46484 16842 46518 16858
rect 47674 16842 47708 16858
rect 46732 16696 47002 16731
rect 46484 16450 46518 16466
rect 46614 16642 46648 16658
rect 46614 16450 46648 16466
rect 46732 16642 46766 16696
rect 46732 16450 46766 16466
rect 46850 16642 46884 16658
rect 46850 16450 46884 16466
rect 46968 16642 47002 16696
rect 46968 16450 47002 16466
rect 47191 16642 47225 16658
rect 47191 16450 47225 16466
rect 47309 16642 47343 16658
rect 47309 16450 47343 16466
rect 47427 16642 47461 16658
rect 47427 16450 47461 16466
rect 47545 16642 47579 16658
rect 47545 16450 47579 16466
rect 47674 16450 47708 16466
rect 47792 16842 47826 16895
rect 47792 16450 47826 16466
rect 47910 16842 47944 16858
rect 47910 16450 47944 16466
rect 48028 16842 48062 16895
rect 49665 16872 49681 16906
rect 49715 16872 49731 16906
rect 48028 16450 48062 16466
rect 48146 16842 48180 16858
rect 48146 16450 48180 16466
rect 48264 16842 48298 16858
rect 48264 16450 48298 16466
rect 48382 16842 48416 16858
rect 49622 16822 49656 16838
rect 48630 16696 48900 16731
rect 48382 16450 48416 16466
rect 48512 16642 48546 16658
rect 48512 16450 48546 16466
rect 48630 16642 48664 16696
rect 48630 16450 48664 16466
rect 48748 16642 48782 16658
rect 48748 16450 48782 16466
rect 48866 16642 48900 16696
rect 49622 16630 49656 16646
rect 49740 16822 49774 16838
rect 49740 16630 49774 16646
rect 49857 16822 49891 16838
rect 48866 16450 48900 16466
rect 49355 16496 49604 16539
rect 49355 16406 49394 16496
rect 49557 16406 49604 16496
rect 49857 16430 49891 16446
rect 49975 16822 50009 16838
rect 49975 16430 50009 16446
rect 50093 16822 50127 16838
rect 50093 16430 50127 16446
rect 49355 16367 49604 16406
rect 49900 16362 49916 16396
rect 49950 16362 49966 16396
rect 50018 16362 50034 16396
rect 50068 16362 50084 16396
rect 47402 16228 47436 16244
rect 45279 16207 45346 16223
rect 45279 16173 45295 16207
rect 45329 16173 45346 16207
rect 47402 16178 47436 16194
rect 45279 16157 45346 16173
rect 45833 16149 45867 16165
rect 45951 16149 45985 16165
rect 45833 15757 45867 15773
rect 45949 15773 45951 15819
rect 45262 15744 45362 15745
rect 45206 15715 45362 15744
rect 45949 15715 45985 15773
rect 46069 16149 46103 16165
rect 46069 15757 46103 15773
rect 46187 16149 46221 16165
rect 46305 16149 46339 16165
rect 46221 15773 46223 15820
rect 46187 15715 46223 15773
rect 46423 16149 46457 16165
rect 46305 15757 46339 15773
rect 46422 15773 46423 15820
rect 46541 16149 46575 16165
rect 46457 15773 46458 15820
rect 46422 15715 46458 15773
rect 46541 15757 46575 15773
rect 47731 16149 47765 16165
rect 47849 16149 47883 16165
rect 47731 15757 47765 15773
rect 47847 15773 47849 15819
rect 45206 15675 46458 15715
rect 46763 15715 47260 15733
rect 47847 15715 47883 15773
rect 47967 16149 48001 16165
rect 47967 15757 48001 15773
rect 48085 16149 48119 16165
rect 48203 16149 48237 16165
rect 48119 15773 48121 15820
rect 48085 15715 48121 15773
rect 48321 16149 48355 16165
rect 48203 15757 48237 15773
rect 48320 15773 48321 15820
rect 48439 16149 48473 16165
rect 48355 15773 48356 15820
rect 48320 15715 48356 15773
rect 49751 16069 49974 16145
rect 49751 15920 49828 16069
rect 49895 15920 49974 16069
rect 49751 15814 49974 15920
rect 48439 15757 48473 15773
rect 46763 15712 48356 15715
rect 46763 15678 46781 15712
rect 46815 15678 48356 15712
rect 46763 15675 48356 15678
rect 49273 15705 49543 15739
rect 45206 15674 46439 15675
rect 46763 15674 48337 15675
rect 45206 15646 45362 15674
rect 45262 15645 45362 15646
rect 45849 15586 45916 15602
rect 45849 15552 45865 15586
rect 45899 15552 45916 15586
rect 45849 15536 45916 15552
rect 45573 15517 45607 15533
rect 45573 15467 45607 15483
rect 46111 15468 46127 15502
rect 46161 15468 46177 15502
rect 46229 15467 46245 15501
rect 46279 15467 46295 15501
rect 46350 15433 46384 15674
rect 46763 15657 47260 15674
rect 46494 15585 46561 15601
rect 46494 15551 46511 15585
rect 46545 15551 46561 15585
rect 46494 15535 46561 15551
rect 47745 15585 47812 15601
rect 47745 15551 47761 15585
rect 47795 15551 47812 15585
rect 47745 15535 47812 15551
rect 46696 15518 46730 15534
rect 46696 15468 46730 15484
rect 47471 15517 47505 15533
rect 47471 15467 47505 15483
rect 48009 15468 48025 15502
rect 48059 15468 48075 15502
rect 48127 15467 48143 15501
rect 48177 15467 48193 15501
rect 48248 15433 48282 15674
rect 49273 15655 49307 15705
rect 48392 15585 48459 15601
rect 48392 15551 48409 15585
rect 48443 15551 48459 15585
rect 48392 15535 48459 15551
rect 48594 15518 48628 15534
rect 48594 15468 48628 15484
rect 49273 15463 49307 15479
rect 49391 15655 49425 15671
rect 49391 15463 49425 15479
rect 49509 15655 49543 15705
rect 49509 15463 49543 15479
rect 49627 15655 49661 15671
rect 49627 15463 49661 15479
rect 49745 15655 49779 15671
rect 49745 15463 49779 15479
rect 49863 15655 49897 15671
rect 49863 15463 49897 15479
rect 49981 15655 50015 15671
rect 49981 15463 50015 15479
rect 50099 15655 50133 15671
rect 50099 15463 50133 15479
rect 50217 15655 50251 15671
rect 50217 15463 50251 15479
rect 50335 15655 50369 15671
rect 50335 15463 50369 15479
rect 45427 15417 45461 15433
rect 45427 15225 45461 15241
rect 45545 15417 45579 15433
rect 45545 15225 45579 15241
rect 45951 15417 45985 15433
rect 46069 15417 46103 15433
rect 45951 14974 45986 15041
rect 46069 15025 46103 15041
rect 46187 15417 46221 15433
rect 46187 15025 46221 15041
rect 46305 15417 46384 15433
rect 46339 15387 46384 15417
rect 46423 15417 46457 15433
rect 46725 15417 46759 15433
rect 46725 15225 46759 15241
rect 46843 15417 46877 15433
rect 46843 15225 46877 15241
rect 47325 15417 47359 15433
rect 47325 15225 47359 15241
rect 47443 15417 47477 15433
rect 47443 15225 47477 15241
rect 47849 15417 47883 15433
rect 46305 15025 46339 15041
rect 46422 14974 46457 15041
rect 45951 14939 46457 14974
rect 47967 15417 48001 15433
rect 47849 14974 47884 15041
rect 47967 15025 48001 15041
rect 48085 15417 48119 15433
rect 48085 15025 48119 15041
rect 48203 15417 48282 15433
rect 48237 15387 48282 15417
rect 48321 15417 48355 15433
rect 48623 15417 48657 15433
rect 48623 15225 48657 15241
rect 48741 15417 48775 15433
rect 49552 15385 49568 15419
rect 49602 15385 49618 15419
rect 49670 15268 49686 15302
rect 49720 15268 49736 15302
rect 48741 15225 48775 15241
rect 48203 15025 48237 15041
rect 48320 14974 48355 15041
rect 49627 15218 49661 15234
rect 49627 15026 49661 15042
rect 49745 15218 49779 15234
rect 49745 15026 49779 15042
rect 49862 15218 49896 15234
rect 47849 14939 48355 14974
rect 49360 14892 49609 14935
rect 49360 14802 49399 14892
rect 49562 14802 49609 14892
rect 49862 14826 49896 14842
rect 49980 15218 50014 15234
rect 49980 14826 50014 14842
rect 50098 15218 50132 15234
rect 50098 14826 50132 14842
rect 48012 14732 48184 14779
rect 49360 14763 49609 14802
rect 49905 14758 49921 14792
rect 49955 14758 49971 14792
rect 50023 14758 50039 14792
rect 50073 14758 50089 14792
rect 48012 14569 48055 14732
rect 48145 14569 48184 14732
rect 48012 14529 48184 14569
rect 51189 13036 51310 17446
rect 56280 17529 56357 17678
rect 56424 17529 56503 17678
rect 59861 17618 59904 17781
rect 59994 17618 60033 17781
rect 56280 17423 56503 17529
rect 57547 17563 57833 17617
rect 59861 17579 60033 17618
rect 61003 17783 61175 17830
rect 61003 17620 61046 17783
rect 61136 17620 61175 17783
rect 61003 17581 61175 17620
rect 62793 17681 63016 17757
rect 57547 17471 57595 17563
rect 57693 17471 57833 17563
rect 57547 17452 57833 17471
rect 52567 17335 52792 17411
rect 52567 17186 52646 17335
rect 52713 17186 52792 17335
rect 52567 17080 52792 17186
rect 55802 17314 56072 17348
rect 55802 17264 55836 17314
rect 55802 17072 55836 17088
rect 55920 17264 55954 17280
rect 55920 17072 55954 17088
rect 56038 17264 56072 17314
rect 56038 17072 56072 17088
rect 56156 17264 56190 17280
rect 56156 17072 56190 17088
rect 56274 17264 56308 17280
rect 56274 17072 56308 17088
rect 56392 17264 56426 17280
rect 56392 17072 56426 17088
rect 56510 17264 56544 17280
rect 56510 17072 56544 17088
rect 56628 17264 56662 17280
rect 56628 17072 56662 17088
rect 56746 17264 56780 17280
rect 56746 17072 56780 17088
rect 56864 17264 56898 17280
rect 56864 17072 56898 17088
rect 56081 16994 56097 17028
rect 56131 16994 56147 17028
rect 52428 16900 52698 16935
rect 52310 16847 52344 16863
rect 51827 16647 51861 16663
rect 51827 16455 51861 16471
rect 51945 16647 51979 16663
rect 51945 16455 51979 16471
rect 52063 16647 52097 16663
rect 52063 16455 52097 16471
rect 52181 16647 52215 16663
rect 52181 16455 52215 16471
rect 52310 16455 52344 16471
rect 52428 16847 52462 16900
rect 52428 16455 52462 16471
rect 52546 16847 52580 16863
rect 52546 16455 52580 16471
rect 52664 16847 52698 16900
rect 54326 16900 54596 16935
rect 52664 16455 52698 16471
rect 52782 16847 52816 16863
rect 52782 16455 52816 16471
rect 52900 16847 52934 16863
rect 52900 16455 52934 16471
rect 53018 16847 53052 16863
rect 54208 16847 54242 16863
rect 53266 16701 53536 16736
rect 53018 16455 53052 16471
rect 53148 16647 53182 16663
rect 53148 16455 53182 16471
rect 53266 16647 53300 16701
rect 53266 16455 53300 16471
rect 53384 16647 53418 16663
rect 53384 16455 53418 16471
rect 53502 16647 53536 16701
rect 53502 16455 53536 16471
rect 53725 16647 53759 16663
rect 53725 16455 53759 16471
rect 53843 16647 53877 16663
rect 53843 16455 53877 16471
rect 53961 16647 53995 16663
rect 53961 16455 53995 16471
rect 54079 16647 54113 16663
rect 54079 16455 54113 16471
rect 54208 16455 54242 16471
rect 54326 16847 54360 16900
rect 54326 16455 54360 16471
rect 54444 16847 54478 16863
rect 54444 16455 54478 16471
rect 54562 16847 54596 16900
rect 56199 16877 56215 16911
rect 56249 16877 56265 16911
rect 54562 16455 54596 16471
rect 54680 16847 54714 16863
rect 54680 16455 54714 16471
rect 54798 16847 54832 16863
rect 54798 16455 54832 16471
rect 54916 16847 54950 16863
rect 56156 16827 56190 16843
rect 55164 16701 55434 16736
rect 54916 16455 54950 16471
rect 55046 16647 55080 16663
rect 55046 16455 55080 16471
rect 55164 16647 55198 16701
rect 55164 16455 55198 16471
rect 55282 16647 55316 16663
rect 55282 16455 55316 16471
rect 55400 16647 55434 16701
rect 56156 16635 56190 16651
rect 56274 16827 56308 16843
rect 56274 16635 56308 16651
rect 56391 16827 56425 16843
rect 55400 16455 55434 16471
rect 55889 16501 56138 16544
rect 55889 16411 55928 16501
rect 56091 16411 56138 16501
rect 56391 16435 56425 16451
rect 56509 16827 56543 16843
rect 56509 16435 56543 16451
rect 56627 16827 56661 16843
rect 56627 16435 56661 16451
rect 55889 16372 56138 16411
rect 56434 16367 56450 16401
rect 56484 16367 56500 16401
rect 56552 16367 56568 16401
rect 56602 16367 56618 16401
rect 53936 16233 53970 16249
rect 51813 16212 51880 16228
rect 51813 16178 51829 16212
rect 51863 16178 51880 16212
rect 53936 16183 53970 16199
rect 51813 16162 51880 16178
rect 52367 16154 52401 16170
rect 52485 16154 52519 16170
rect 52367 15762 52401 15778
rect 52483 15778 52485 15824
rect 51796 15749 51896 15750
rect 51740 15720 51896 15749
rect 52483 15720 52519 15778
rect 52603 16154 52637 16170
rect 52603 15762 52637 15778
rect 52721 16154 52755 16170
rect 52839 16154 52873 16170
rect 52755 15778 52757 15825
rect 52721 15720 52757 15778
rect 52957 16154 52991 16170
rect 52839 15762 52873 15778
rect 52956 15778 52957 15825
rect 53075 16154 53109 16170
rect 52991 15778 52992 15825
rect 52956 15720 52992 15778
rect 53075 15762 53109 15778
rect 54265 16154 54299 16170
rect 54383 16154 54417 16170
rect 54265 15762 54299 15778
rect 54381 15778 54383 15824
rect 51740 15680 52992 15720
rect 53297 15720 53794 15738
rect 54381 15720 54417 15778
rect 54501 16154 54535 16170
rect 54501 15762 54535 15778
rect 54619 16154 54653 16170
rect 54737 16154 54771 16170
rect 54653 15778 54655 15825
rect 54619 15720 54655 15778
rect 54855 16154 54889 16170
rect 54737 15762 54771 15778
rect 54854 15778 54855 15825
rect 54973 16154 55007 16170
rect 54889 15778 54890 15825
rect 54854 15720 54890 15778
rect 56285 16074 56508 16150
rect 56285 15925 56362 16074
rect 56429 15925 56508 16074
rect 56285 15819 56508 15925
rect 54973 15762 55007 15778
rect 53297 15717 54890 15720
rect 53297 15683 53315 15717
rect 53349 15683 54890 15717
rect 53297 15680 54890 15683
rect 55807 15710 56077 15744
rect 51740 15679 52973 15680
rect 53297 15679 54871 15680
rect 51740 15651 51896 15679
rect 51796 15650 51896 15651
rect 52383 15591 52450 15607
rect 52383 15557 52399 15591
rect 52433 15557 52450 15591
rect 52383 15541 52450 15557
rect 52107 15522 52141 15538
rect 52107 15472 52141 15488
rect 52645 15473 52661 15507
rect 52695 15473 52711 15507
rect 52763 15472 52779 15506
rect 52813 15472 52829 15506
rect 52884 15438 52918 15679
rect 53297 15662 53794 15679
rect 53028 15590 53095 15606
rect 53028 15556 53045 15590
rect 53079 15556 53095 15590
rect 53028 15540 53095 15556
rect 54279 15590 54346 15606
rect 54279 15556 54295 15590
rect 54329 15556 54346 15590
rect 54279 15540 54346 15556
rect 53230 15523 53264 15539
rect 53230 15473 53264 15489
rect 54005 15522 54039 15538
rect 54005 15472 54039 15488
rect 54543 15473 54559 15507
rect 54593 15473 54609 15507
rect 54661 15472 54677 15506
rect 54711 15472 54727 15506
rect 54782 15438 54816 15679
rect 55807 15660 55841 15710
rect 54926 15590 54993 15606
rect 54926 15556 54943 15590
rect 54977 15556 54993 15590
rect 54926 15540 54993 15556
rect 55128 15523 55162 15539
rect 55128 15473 55162 15489
rect 55807 15468 55841 15484
rect 55925 15660 55959 15676
rect 55925 15468 55959 15484
rect 56043 15660 56077 15710
rect 56043 15468 56077 15484
rect 56161 15660 56195 15676
rect 56161 15468 56195 15484
rect 56279 15660 56313 15676
rect 56279 15468 56313 15484
rect 56397 15660 56431 15676
rect 56397 15468 56431 15484
rect 56515 15660 56549 15676
rect 56515 15468 56549 15484
rect 56633 15660 56667 15676
rect 56633 15468 56667 15484
rect 56751 15660 56785 15676
rect 56751 15468 56785 15484
rect 56869 15660 56903 15676
rect 56869 15468 56903 15484
rect 51961 15422 51995 15438
rect 51961 15230 51995 15246
rect 52079 15422 52113 15438
rect 52079 15230 52113 15246
rect 52485 15422 52519 15438
rect 52603 15422 52637 15438
rect 52485 14979 52520 15046
rect 52603 15030 52637 15046
rect 52721 15422 52755 15438
rect 52721 15030 52755 15046
rect 52839 15422 52918 15438
rect 52873 15392 52918 15422
rect 52957 15422 52991 15438
rect 53259 15422 53293 15438
rect 53259 15230 53293 15246
rect 53377 15422 53411 15438
rect 53377 15230 53411 15246
rect 53859 15422 53893 15438
rect 53859 15230 53893 15246
rect 53977 15422 54011 15438
rect 53977 15230 54011 15246
rect 54383 15422 54417 15438
rect 52839 15030 52873 15046
rect 52956 14979 52991 15046
rect 52485 14944 52991 14979
rect 54501 15422 54535 15438
rect 54383 14979 54418 15046
rect 54501 15030 54535 15046
rect 54619 15422 54653 15438
rect 54619 15030 54653 15046
rect 54737 15422 54816 15438
rect 54771 15392 54816 15422
rect 54855 15422 54889 15438
rect 55157 15422 55191 15438
rect 55157 15230 55191 15246
rect 55275 15422 55309 15438
rect 56086 15390 56102 15424
rect 56136 15390 56152 15424
rect 56204 15273 56220 15307
rect 56254 15273 56270 15307
rect 55275 15230 55309 15246
rect 54737 15030 54771 15046
rect 54854 14979 54889 15046
rect 56161 15223 56195 15239
rect 56161 15031 56195 15047
rect 56279 15223 56313 15239
rect 56279 15031 56313 15047
rect 56396 15223 56430 15239
rect 54383 14944 54889 14979
rect 55894 14897 56143 14940
rect 55894 14807 55933 14897
rect 56096 14807 56143 14897
rect 56396 14831 56430 14847
rect 56514 15223 56548 15239
rect 56514 14831 56548 14847
rect 56632 15223 56666 15239
rect 56632 14831 56666 14847
rect 54546 14737 54718 14784
rect 55894 14768 56143 14807
rect 56439 14763 56455 14797
rect 56489 14763 56505 14797
rect 56557 14763 56573 14797
rect 56607 14763 56623 14797
rect 54546 14574 54589 14737
rect 54679 14574 54718 14737
rect 54546 14534 54718 14574
rect 57709 13561 57833 17452
rect 62793 17532 62870 17681
rect 62937 17532 63016 17681
rect 62793 17426 63016 17532
rect 59080 17338 59305 17414
rect 59080 17189 59159 17338
rect 59226 17189 59305 17338
rect 59080 17083 59305 17189
rect 62315 17317 62585 17351
rect 62315 17267 62349 17317
rect 62315 17075 62349 17091
rect 62433 17267 62467 17283
rect 62433 17075 62467 17091
rect 62551 17267 62585 17317
rect 62551 17075 62585 17091
rect 62669 17267 62703 17283
rect 62669 17075 62703 17091
rect 62787 17267 62821 17283
rect 62787 17075 62821 17091
rect 62905 17267 62939 17283
rect 62905 17075 62939 17091
rect 63023 17267 63057 17283
rect 63023 17075 63057 17091
rect 63141 17267 63175 17283
rect 63141 17075 63175 17091
rect 63259 17267 63293 17283
rect 63259 17075 63293 17091
rect 63377 17267 63411 17283
rect 63377 17075 63411 17091
rect 62594 16997 62610 17031
rect 62644 16997 62660 17031
rect 58941 16903 59211 16938
rect 58823 16850 58857 16866
rect 58340 16650 58374 16666
rect 58340 16458 58374 16474
rect 58458 16650 58492 16666
rect 58458 16458 58492 16474
rect 58576 16650 58610 16666
rect 58576 16458 58610 16474
rect 58694 16650 58728 16666
rect 58694 16458 58728 16474
rect 58823 16458 58857 16474
rect 58941 16850 58975 16903
rect 58941 16458 58975 16474
rect 59059 16850 59093 16866
rect 59059 16458 59093 16474
rect 59177 16850 59211 16903
rect 60839 16903 61109 16938
rect 59177 16458 59211 16474
rect 59295 16850 59329 16866
rect 59295 16458 59329 16474
rect 59413 16850 59447 16866
rect 59413 16458 59447 16474
rect 59531 16850 59565 16866
rect 60721 16850 60755 16866
rect 59779 16704 60049 16739
rect 59531 16458 59565 16474
rect 59661 16650 59695 16666
rect 59661 16458 59695 16474
rect 59779 16650 59813 16704
rect 59779 16458 59813 16474
rect 59897 16650 59931 16666
rect 59897 16458 59931 16474
rect 60015 16650 60049 16704
rect 60015 16458 60049 16474
rect 60238 16650 60272 16666
rect 60238 16458 60272 16474
rect 60356 16650 60390 16666
rect 60356 16458 60390 16474
rect 60474 16650 60508 16666
rect 60474 16458 60508 16474
rect 60592 16650 60626 16666
rect 60592 16458 60626 16474
rect 60721 16458 60755 16474
rect 60839 16850 60873 16903
rect 60839 16458 60873 16474
rect 60957 16850 60991 16866
rect 60957 16458 60991 16474
rect 61075 16850 61109 16903
rect 62712 16880 62728 16914
rect 62762 16880 62778 16914
rect 61075 16458 61109 16474
rect 61193 16850 61227 16866
rect 61193 16458 61227 16474
rect 61311 16850 61345 16866
rect 61311 16458 61345 16474
rect 61429 16850 61463 16866
rect 62669 16830 62703 16846
rect 61677 16704 61947 16739
rect 61429 16458 61463 16474
rect 61559 16650 61593 16666
rect 61559 16458 61593 16474
rect 61677 16650 61711 16704
rect 61677 16458 61711 16474
rect 61795 16650 61829 16666
rect 61795 16458 61829 16474
rect 61913 16650 61947 16704
rect 62669 16638 62703 16654
rect 62787 16830 62821 16846
rect 62787 16638 62821 16654
rect 62904 16830 62938 16846
rect 61913 16458 61947 16474
rect 62402 16504 62651 16547
rect 62402 16414 62441 16504
rect 62604 16414 62651 16504
rect 62904 16438 62938 16454
rect 63022 16830 63056 16846
rect 63022 16438 63056 16454
rect 63140 16830 63174 16846
rect 63140 16438 63174 16454
rect 62402 16375 62651 16414
rect 62947 16370 62963 16404
rect 62997 16370 63013 16404
rect 63065 16370 63081 16404
rect 63115 16370 63131 16404
rect 60449 16236 60483 16252
rect 58326 16215 58393 16231
rect 58326 16181 58342 16215
rect 58376 16181 58393 16215
rect 60449 16186 60483 16202
rect 58326 16165 58393 16181
rect 58880 16157 58914 16173
rect 58998 16157 59032 16173
rect 58880 15765 58914 15781
rect 58996 15781 58998 15827
rect 58309 15752 58409 15753
rect 58253 15723 58409 15752
rect 58996 15723 59032 15781
rect 59116 16157 59150 16173
rect 59116 15765 59150 15781
rect 59234 16157 59268 16173
rect 59352 16157 59386 16173
rect 59268 15781 59270 15828
rect 59234 15723 59270 15781
rect 59470 16157 59504 16173
rect 59352 15765 59386 15781
rect 59469 15781 59470 15828
rect 59588 16157 59622 16173
rect 59504 15781 59505 15828
rect 59469 15723 59505 15781
rect 59588 15765 59622 15781
rect 60778 16157 60812 16173
rect 60896 16157 60930 16173
rect 60778 15765 60812 15781
rect 60894 15781 60896 15827
rect 58253 15683 59505 15723
rect 59810 15723 60307 15741
rect 60894 15723 60930 15781
rect 61014 16157 61048 16173
rect 61014 15765 61048 15781
rect 61132 16157 61166 16173
rect 61250 16157 61284 16173
rect 61166 15781 61168 15828
rect 61132 15723 61168 15781
rect 61368 16157 61402 16173
rect 61250 15765 61284 15781
rect 61367 15781 61368 15828
rect 61486 16157 61520 16173
rect 61402 15781 61403 15828
rect 61367 15723 61403 15781
rect 62798 16077 63021 16153
rect 62798 15928 62875 16077
rect 62942 15928 63021 16077
rect 62798 15822 63021 15928
rect 61486 15765 61520 15781
rect 59810 15720 61403 15723
rect 59810 15686 59828 15720
rect 59862 15686 61403 15720
rect 59810 15683 61403 15686
rect 62320 15713 62590 15747
rect 58253 15682 59486 15683
rect 59810 15682 61384 15683
rect 58253 15654 58409 15682
rect 58309 15653 58409 15654
rect 58896 15594 58963 15610
rect 58896 15560 58912 15594
rect 58946 15560 58963 15594
rect 58896 15544 58963 15560
rect 58620 15525 58654 15541
rect 58620 15475 58654 15491
rect 59158 15476 59174 15510
rect 59208 15476 59224 15510
rect 59276 15475 59292 15509
rect 59326 15475 59342 15509
rect 59397 15441 59431 15682
rect 59810 15665 60307 15682
rect 59541 15593 59608 15609
rect 59541 15559 59558 15593
rect 59592 15559 59608 15593
rect 59541 15543 59608 15559
rect 60792 15593 60859 15609
rect 60792 15559 60808 15593
rect 60842 15559 60859 15593
rect 60792 15543 60859 15559
rect 59743 15526 59777 15542
rect 59743 15476 59777 15492
rect 60518 15525 60552 15541
rect 60518 15475 60552 15491
rect 61056 15476 61072 15510
rect 61106 15476 61122 15510
rect 61174 15475 61190 15509
rect 61224 15475 61240 15509
rect 61295 15441 61329 15682
rect 62320 15663 62354 15713
rect 61439 15593 61506 15609
rect 61439 15559 61456 15593
rect 61490 15559 61506 15593
rect 61439 15543 61506 15559
rect 61641 15526 61675 15542
rect 61641 15476 61675 15492
rect 62320 15471 62354 15487
rect 62438 15663 62472 15679
rect 62438 15471 62472 15487
rect 62556 15663 62590 15713
rect 62556 15471 62590 15487
rect 62674 15663 62708 15679
rect 62674 15471 62708 15487
rect 62792 15663 62826 15679
rect 62792 15471 62826 15487
rect 62910 15663 62944 15679
rect 62910 15471 62944 15487
rect 63028 15663 63062 15679
rect 63028 15471 63062 15487
rect 63146 15663 63180 15679
rect 63146 15471 63180 15487
rect 63264 15663 63298 15679
rect 63264 15471 63298 15487
rect 63382 15663 63416 15679
rect 63382 15471 63416 15487
rect 58474 15425 58508 15441
rect 58474 15233 58508 15249
rect 58592 15425 58626 15441
rect 58592 15233 58626 15249
rect 58998 15425 59032 15441
rect 59116 15425 59150 15441
rect 58998 14982 59033 15049
rect 59116 15033 59150 15049
rect 59234 15425 59268 15441
rect 59234 15033 59268 15049
rect 59352 15425 59431 15441
rect 59386 15395 59431 15425
rect 59470 15425 59504 15441
rect 59772 15425 59806 15441
rect 59772 15233 59806 15249
rect 59890 15425 59924 15441
rect 59890 15233 59924 15249
rect 60372 15425 60406 15441
rect 60372 15233 60406 15249
rect 60490 15425 60524 15441
rect 60490 15233 60524 15249
rect 60896 15425 60930 15441
rect 59352 15033 59386 15049
rect 59469 14982 59504 15049
rect 58998 14947 59504 14982
rect 61014 15425 61048 15441
rect 60896 14982 60931 15049
rect 61014 15033 61048 15049
rect 61132 15425 61166 15441
rect 61132 15033 61166 15049
rect 61250 15425 61329 15441
rect 61284 15395 61329 15425
rect 61368 15425 61402 15441
rect 61670 15425 61704 15441
rect 61670 15233 61704 15249
rect 61788 15425 61822 15441
rect 62599 15393 62615 15427
rect 62649 15393 62665 15427
rect 62717 15276 62733 15310
rect 62767 15276 62783 15310
rect 61788 15233 61822 15249
rect 61250 15033 61284 15049
rect 61367 14982 61402 15049
rect 62674 15226 62708 15242
rect 62674 15034 62708 15050
rect 62792 15226 62826 15242
rect 62792 15034 62826 15050
rect 62909 15226 62943 15242
rect 60896 14947 61402 14982
rect 62407 14900 62656 14943
rect 62407 14810 62446 14900
rect 62609 14810 62656 14900
rect 62909 14834 62943 14850
rect 63027 15226 63061 15242
rect 63027 14834 63061 14850
rect 63145 15226 63179 15242
rect 63145 14834 63179 14850
rect 61059 14740 61231 14787
rect 62407 14771 62656 14810
rect 62952 14766 62968 14800
rect 63002 14766 63018 14800
rect 63070 14766 63086 14800
rect 63120 14766 63136 14800
rect 61059 14577 61102 14740
rect 61192 14577 61231 14740
rect 61059 14537 61231 14577
rect 57708 13155 57834 13561
rect 57708 13097 57742 13155
rect 57810 13097 57834 13155
rect 57708 13066 57834 13097
rect 51189 12980 51217 13036
rect 51288 12980 51310 13036
rect 51189 12954 51310 12980
rect 64602 12925 64700 19358
rect 68233 19149 71573 19170
rect 68233 19086 68260 19149
rect 68309 19086 71573 19149
rect 68233 19084 71573 19086
rect 71486 19056 71573 19084
rect 71486 19007 71499 19056
rect 71559 19007 71573 19056
rect 71486 18985 71573 19007
rect 70635 18883 70725 18917
rect 70901 18883 70917 18917
rect 70635 18681 70674 18883
rect 71199 18812 71284 18828
rect 70709 18765 70725 18799
rect 70901 18765 70991 18799
rect 70635 18647 70725 18681
rect 70901 18647 70917 18681
rect 70952 18563 70991 18765
rect 71199 18752 71216 18812
rect 71271 18752 71284 18812
rect 71199 18736 71284 18752
rect 70709 18529 70725 18563
rect 70901 18529 70991 18563
rect 70433 18442 70525 18476
rect 70901 18442 70917 18476
rect 70433 18240 70472 18442
rect 70509 18324 70525 18358
rect 70901 18324 70991 18358
rect 70433 18206 70525 18240
rect 70901 18206 70917 18240
rect 70952 18122 70991 18324
rect 70509 18088 70525 18122
rect 70901 18088 70991 18122
rect 70434 17975 70525 18009
rect 70901 17975 70917 18009
rect 70434 17773 70473 17975
rect 70952 17891 70991 18088
rect 71842 18049 71858 18083
rect 72034 18049 72050 18083
rect 71842 17931 71858 17965
rect 72034 17931 72050 17965
rect 71846 17891 72046 17931
rect 70509 17857 70525 17891
rect 70901 17857 70991 17891
rect 70237 17731 70347 17747
rect 70434 17739 70525 17773
rect 70901 17739 70917 17773
rect 70237 17535 70255 17731
rect 70331 17535 70347 17731
rect 70952 17655 70991 17857
rect 71487 17845 71572 17861
rect 71842 17857 71858 17891
rect 72234 17857 72250 17891
rect 71100 17797 71116 17831
rect 71150 17797 71166 17831
rect 71487 17785 71500 17845
rect 71555 17785 71572 17845
rect 71487 17769 71572 17785
rect 70509 17621 70525 17655
rect 70901 17621 70991 17655
rect 71202 17727 71287 17743
rect 71842 17739 71858 17773
rect 72234 17739 72250 17773
rect 71202 17667 71215 17727
rect 71270 17667 71287 17727
rect 72483 17673 72569 17689
rect 71202 17651 71287 17667
rect 71842 17621 71858 17655
rect 72234 17621 72250 17655
rect 72335 17654 72369 17670
rect 70237 17519 70347 17535
rect 70434 17503 70525 17537
rect 70901 17503 70917 17537
rect 70434 17301 70473 17503
rect 70952 17419 70991 17621
rect 72335 17604 72369 17620
rect 72483 17651 72501 17673
rect 71720 17562 71736 17596
rect 71770 17562 71786 17596
rect 72483 17593 72487 17651
rect 72483 17569 72501 17593
rect 72547 17569 72569 17673
rect 72483 17553 72569 17569
rect 71842 17503 71858 17537
rect 72234 17503 72250 17537
rect 71330 17443 71346 17477
rect 71380 17443 71396 17477
rect 70509 17385 70525 17419
rect 70901 17385 70991 17419
rect 71842 17385 71858 17419
rect 72234 17385 72250 17419
rect 70434 17267 70525 17301
rect 70901 17267 70917 17301
rect 70952 17182 70991 17385
rect 71846 17341 72046 17385
rect 71842 17307 71858 17341
rect 72034 17307 72050 17341
rect 71842 17189 71858 17223
rect 72034 17189 72050 17223
rect 70509 17148 70525 17182
rect 70901 17148 70991 17182
rect 70434 17030 70525 17064
rect 70901 17030 70917 17064
rect 70434 16828 70473 17030
rect 70952 16946 70991 17148
rect 70509 16912 70525 16946
rect 70901 16912 70991 16946
rect 70434 16794 70525 16828
rect 70901 16794 70917 16828
rect 70709 16675 70725 16709
rect 70901 16675 70994 16709
rect 70638 16557 70725 16591
rect 70901 16557 70917 16591
rect 70638 16355 70675 16557
rect 70955 16473 70994 16675
rect 70709 16439 70725 16473
rect 70901 16439 70994 16473
rect 71075 16521 71109 16537
rect 71075 16471 71109 16487
rect 70638 16321 70725 16355
rect 70901 16321 70917 16355
rect 68537 15948 71570 16029
rect 44609 12658 44641 12703
rect 44720 12658 44746 12703
rect 44609 12635 44746 12658
rect 55062 12397 55230 12413
rect 41859 12377 42027 12393
rect 41859 12307 41875 12377
rect 42011 12307 42027 12377
rect 41859 12291 42027 12307
rect 48408 12376 48576 12392
rect 48408 12306 48424 12376
rect 48560 12306 48576 12376
rect 55062 12327 55078 12397
rect 55214 12327 55230 12397
rect 55062 12311 55230 12327
rect 64604 12365 64698 12925
rect 48408 12290 48576 12306
rect 64604 12293 64610 12365
rect 64688 12293 64698 12365
rect 64604 12288 64698 12293
rect 65857 12323 66301 12329
rect 42396 12187 42666 12221
rect 41570 12137 41604 12153
rect 41570 11945 41604 11961
rect 41688 12137 41722 12153
rect 41688 11945 41722 11961
rect 41806 12137 41840 12153
rect 41806 11945 41840 11961
rect 41924 12137 41958 12153
rect 41924 11945 41958 11961
rect 42042 12137 42076 12153
rect 42042 11945 42076 11961
rect 42160 12137 42194 12153
rect 42160 11945 42194 11961
rect 42278 12137 42312 12153
rect 42278 11945 42312 11961
rect 42396 12137 42430 12187
rect 42396 11945 42430 11961
rect 42514 12137 42548 12153
rect 42514 11945 42548 11961
rect 42632 12137 42666 12187
rect 48945 12186 49215 12220
rect 42632 11945 42666 11961
rect 48119 12136 48153 12152
rect 48119 11944 48153 11960
rect 48237 12136 48271 12152
rect 48237 11944 48271 11960
rect 48355 12136 48389 12152
rect 48355 11944 48389 11960
rect 48473 12136 48507 12152
rect 48473 11944 48507 11960
rect 48591 12136 48625 12152
rect 48591 11944 48625 11960
rect 48709 12136 48743 12152
rect 48709 11944 48743 11960
rect 48827 12136 48861 12152
rect 48827 11944 48861 11960
rect 48945 12136 48979 12186
rect 48945 11944 48979 11960
rect 49063 12136 49097 12152
rect 49063 11944 49097 11960
rect 49181 12136 49215 12186
rect 55599 12207 55869 12241
rect 54773 12157 54807 12173
rect 54773 11965 54807 11981
rect 54891 12157 54925 12173
rect 54891 11965 54925 11981
rect 55009 12157 55043 12173
rect 55009 11965 55043 11981
rect 55127 12157 55161 12173
rect 55127 11965 55161 11981
rect 55245 12157 55279 12173
rect 55245 11965 55279 11981
rect 55363 12157 55397 12173
rect 55363 11965 55397 11981
rect 55481 12157 55515 12173
rect 55481 11965 55515 11981
rect 55599 12157 55633 12207
rect 55599 11965 55633 11981
rect 55717 12157 55751 12173
rect 55717 11965 55751 11981
rect 55835 12157 55869 12207
rect 63715 12230 63883 12246
rect 63715 12160 63731 12230
rect 63867 12160 63883 12230
rect 63715 12144 63883 12160
rect 65857 12123 65868 12323
rect 66289 12123 66301 12323
rect 65857 12117 66301 12123
rect 64252 12040 64522 12074
rect 55835 11965 55869 11981
rect 63426 11990 63460 12006
rect 49181 11944 49215 11960
rect 42321 11867 42337 11901
rect 42371 11867 42387 11901
rect 48870 11866 48886 11900
rect 48920 11866 48936 11900
rect 55524 11887 55540 11921
rect 55574 11887 55590 11921
rect 42203 11750 42219 11784
rect 42253 11750 42269 11784
rect 48752 11749 48768 11783
rect 48802 11749 48818 11783
rect 55406 11770 55422 11804
rect 55456 11770 55472 11804
rect 63426 11798 63460 11814
rect 63544 11990 63578 12006
rect 63544 11798 63578 11814
rect 63662 11990 63696 12006
rect 63662 11798 63696 11814
rect 63780 11990 63814 12006
rect 63780 11798 63814 11814
rect 63898 11990 63932 12006
rect 63898 11798 63932 11814
rect 64016 11990 64050 12006
rect 64016 11798 64050 11814
rect 64134 11990 64168 12006
rect 64134 11798 64168 11814
rect 64252 11990 64286 12040
rect 64252 11798 64286 11814
rect 64370 11990 64404 12006
rect 64370 11798 64404 11814
rect 64488 11990 64522 12040
rect 64488 11798 64522 11814
rect 66072 11838 66342 11873
rect 65718 11785 65752 11801
rect 55010 11720 55044 11736
rect 41807 11700 41841 11716
rect 41807 11308 41841 11324
rect 41925 11700 41959 11716
rect 41925 11308 41959 11324
rect 42043 11700 42077 11716
rect 42160 11700 42194 11716
rect 42160 11508 42194 11524
rect 42278 11700 42312 11716
rect 42278 11508 42312 11524
rect 48356 11699 48390 11715
rect 42043 11308 42077 11324
rect 48356 11307 48390 11323
rect 48474 11699 48508 11715
rect 48474 11307 48508 11323
rect 48592 11699 48626 11715
rect 48709 11699 48743 11715
rect 48709 11507 48743 11523
rect 48827 11699 48861 11715
rect 48827 11507 48861 11523
rect 55010 11328 55044 11344
rect 55128 11720 55162 11736
rect 55128 11328 55162 11344
rect 55246 11720 55280 11736
rect 55363 11720 55397 11736
rect 55363 11528 55397 11544
rect 55481 11720 55515 11736
rect 64177 11720 64193 11754
rect 64227 11720 64243 11754
rect 65234 11639 65504 11674
rect 64059 11603 64075 11637
rect 64109 11603 64125 11637
rect 65234 11585 65268 11639
rect 55481 11528 55515 11544
rect 63663 11553 63697 11569
rect 55246 11328 55280 11344
rect 48592 11307 48626 11323
rect 54872 11296 54943 11298
rect 48041 11274 48321 11279
rect 41850 11240 41866 11274
rect 41900 11240 41916 11274
rect 41968 11240 41984 11274
rect 42018 11240 42034 11274
rect 48041 11228 48269 11274
rect 48318 11228 48321 11274
rect 48399 11239 48415 11273
rect 48449 11239 48465 11273
rect 48517 11239 48533 11273
rect 48567 11239 48583 11273
rect 54872 11248 54876 11296
rect 54937 11248 54943 11296
rect 55053 11260 55069 11294
rect 55103 11260 55119 11294
rect 55171 11260 55187 11294
rect 55221 11260 55237 11294
rect 48041 11223 48321 11228
rect 54872 11235 54943 11248
rect 42083 11169 42251 11187
rect 42083 11113 42099 11169
rect 42233 11113 42251 11169
rect 42083 11097 42251 11113
rect 33812 10784 33824 10840
rect 33812 10777 33883 10784
rect 33961 11022 34069 11025
rect 33961 10972 33985 11022
rect 34046 10972 34069 11022
rect 33658 9495 33885 9510
rect 33658 9425 33781 9495
rect 33855 9425 33885 9495
rect 33658 9410 33885 9425
rect 33661 9409 33885 9410
rect 33961 9330 34069 10972
rect 48041 10941 48094 11223
rect 48632 11168 48800 11186
rect 48632 11112 48648 11168
rect 48782 11112 48800 11168
rect 48632 11096 48800 11112
rect 34120 10888 48094 10941
rect 34120 10449 34211 10888
rect 54872 10853 54935 11235
rect 34250 10849 54935 10853
rect 34250 10795 41688 10849
rect 41737 10795 54935 10849
rect 34250 10787 54935 10795
rect 54969 11206 55030 11211
rect 54969 11168 54978 11206
rect 55023 11168 55030 11206
rect 34250 10623 34360 10787
rect 54969 10742 55030 11168
rect 55286 11189 55454 11207
rect 55286 11133 55302 11189
rect 55436 11133 55454 11189
rect 63663 11161 63697 11177
rect 63781 11553 63815 11569
rect 63781 11161 63815 11177
rect 63899 11553 63933 11569
rect 64016 11553 64050 11569
rect 64016 11361 64050 11377
rect 64134 11553 64168 11569
rect 65234 11393 65268 11409
rect 65352 11585 65386 11601
rect 65352 11393 65386 11409
rect 65470 11585 65504 11639
rect 65470 11393 65504 11409
rect 65588 11585 65622 11601
rect 65588 11393 65622 11409
rect 65718 11393 65752 11409
rect 65836 11785 65870 11801
rect 65836 11393 65870 11409
rect 65954 11785 65988 11801
rect 65954 11393 65988 11409
rect 66072 11785 66106 11838
rect 66072 11393 66106 11409
rect 66190 11785 66224 11801
rect 66190 11393 66224 11409
rect 66308 11785 66342 11838
rect 67316 11822 67484 11838
rect 66308 11393 66342 11409
rect 66426 11785 66460 11801
rect 67316 11752 67332 11822
rect 67468 11752 67484 11822
rect 67316 11736 67484 11752
rect 67853 11632 68123 11666
rect 66426 11393 66460 11409
rect 66555 11585 66589 11601
rect 66555 11393 66589 11409
rect 66673 11585 66707 11601
rect 66673 11393 66707 11409
rect 66791 11585 66825 11601
rect 66791 11393 66825 11409
rect 66909 11585 66943 11601
rect 66909 11393 66943 11409
rect 67027 11582 67061 11598
rect 67027 11390 67061 11406
rect 67145 11582 67179 11598
rect 67145 11390 67179 11406
rect 67263 11582 67297 11598
rect 67263 11390 67297 11406
rect 67381 11582 67415 11598
rect 67381 11390 67415 11406
rect 67499 11582 67533 11598
rect 67499 11390 67533 11406
rect 67617 11582 67651 11598
rect 67617 11390 67651 11406
rect 67735 11582 67769 11598
rect 67735 11390 67769 11406
rect 67853 11582 67887 11632
rect 67853 11390 67887 11406
rect 67971 11582 68005 11598
rect 67971 11390 68005 11406
rect 68089 11582 68123 11632
rect 68089 11390 68123 11406
rect 64134 11361 64168 11377
rect 67778 11312 67794 11346
rect 67828 11312 67844 11346
rect 66886 11227 66920 11243
rect 67660 11195 67676 11229
rect 67710 11195 67726 11229
rect 66886 11177 66920 11193
rect 63899 11161 63933 11177
rect 55286 11117 55454 11133
rect 67264 11145 67298 11161
rect 63706 11093 63722 11127
rect 63756 11093 63772 11127
rect 63824 11093 63840 11127
rect 63874 11093 63890 11127
rect 64963 11121 65305 11127
rect 64963 11053 65213 11121
rect 65293 11053 65305 11121
rect 65480 11108 65536 11125
rect 65480 11074 65486 11108
rect 65520 11074 65536 11108
rect 65480 11057 65536 11074
rect 65661 11092 65695 11108
rect 64963 11047 65305 11053
rect 63939 11022 64107 11040
rect 63939 10966 63955 11022
rect 64089 10966 64107 11022
rect 63939 10950 64107 10966
rect 34120 10404 34138 10449
rect 34195 10404 34211 10449
rect 34120 10397 34211 10404
rect 33961 9329 34089 9330
rect 33950 9315 34089 9329
rect 33950 9248 33965 9315
rect 33951 9231 33965 9248
rect 34078 9231 34089 9315
rect 33510 6688 33883 6708
rect 33510 6607 33778 6688
rect 33872 6607 33883 6688
rect 33510 6591 33883 6607
rect 33365 914 33876 922
rect 33365 832 33779 914
rect 33861 832 33876 914
rect 33365 821 33876 832
rect 32680 -2190 33880 -2178
rect 32680 -2266 33773 -2190
rect 33867 -2266 33880 -2190
rect 32680 -2274 33880 -2266
rect 33951 -2594 34089 9231
rect 34249 913 34360 10623
rect 36506 10676 55030 10742
rect 35195 10477 35363 10493
rect 35195 10407 35211 10477
rect 35347 10407 35363 10477
rect 35195 10391 35363 10407
rect 35732 10287 36002 10321
rect 34906 10237 34940 10253
rect 34906 10045 34940 10061
rect 35024 10237 35058 10253
rect 35024 10045 35058 10061
rect 35142 10237 35176 10253
rect 35142 10045 35176 10061
rect 35260 10237 35294 10253
rect 35260 10045 35294 10061
rect 35378 10237 35412 10253
rect 35378 10045 35412 10061
rect 35496 10237 35530 10253
rect 35496 10045 35530 10061
rect 35614 10237 35648 10253
rect 35614 10045 35648 10061
rect 35732 10237 35766 10287
rect 35732 10045 35766 10061
rect 35850 10237 35884 10253
rect 35850 10045 35884 10061
rect 35968 10237 36002 10287
rect 35968 10045 36002 10061
rect 35657 9967 35673 10001
rect 35707 9967 35723 10001
rect 35539 9850 35555 9884
rect 35589 9850 35605 9884
rect 35143 9800 35177 9816
rect 34249 832 34257 913
rect 34359 832 34360 913
rect 34249 821 34360 832
rect 34395 9493 34498 9501
rect 34395 9417 34403 9493
rect 34492 9417 34498 9493
rect 34395 -2445 34498 9417
rect 35143 9408 35177 9424
rect 35261 9800 35295 9816
rect 35261 9408 35295 9424
rect 35379 9800 35413 9816
rect 35496 9800 35530 9816
rect 35496 9608 35530 9624
rect 35614 9800 35648 9816
rect 35614 9608 35648 9624
rect 35379 9408 35413 9424
rect 35186 9340 35202 9374
rect 35236 9340 35252 9374
rect 35304 9340 35320 9374
rect 35354 9340 35370 9374
rect 34641 9299 34956 9304
rect 34641 9255 34897 9299
rect 34953 9255 34956 9299
rect 34641 9251 34956 9255
rect 35419 9269 35587 9287
rect 34641 3445 34723 9251
rect 35419 9213 35435 9269
rect 35569 9213 35587 9269
rect 35419 9197 35587 9213
rect 35187 7892 35355 7908
rect 35187 7822 35203 7892
rect 35339 7822 35355 7892
rect 35187 7806 35355 7822
rect 35724 7702 35994 7736
rect 34898 7652 34932 7668
rect 34898 7460 34932 7476
rect 35016 7652 35050 7668
rect 35016 7460 35050 7476
rect 35134 7652 35168 7668
rect 35134 7460 35168 7476
rect 35252 7652 35286 7668
rect 35252 7460 35286 7476
rect 35370 7652 35404 7668
rect 35370 7460 35404 7476
rect 35488 7652 35522 7668
rect 35488 7460 35522 7476
rect 35606 7652 35640 7668
rect 35606 7460 35640 7476
rect 35724 7652 35758 7702
rect 35724 7460 35758 7476
rect 35842 7652 35876 7668
rect 35842 7460 35876 7476
rect 35960 7652 35994 7702
rect 35960 7460 35994 7476
rect 35649 7382 35665 7416
rect 35699 7382 35715 7416
rect 35531 7265 35547 7299
rect 35581 7265 35597 7299
rect 35135 7215 35169 7231
rect 35135 6823 35169 6839
rect 35253 7215 35287 7231
rect 35253 6823 35287 6839
rect 35371 7215 35405 7231
rect 35488 7215 35522 7231
rect 35488 7023 35522 7039
rect 35606 7215 35640 7231
rect 35606 7023 35640 7039
rect 35371 6823 35405 6839
rect 35178 6755 35194 6789
rect 35228 6755 35244 6789
rect 35296 6755 35312 6789
rect 35346 6755 35362 6789
rect 35411 6684 35579 6702
rect 35411 6628 35427 6684
rect 35561 6628 35579 6684
rect 35411 6612 35579 6628
rect 35168 4614 35336 4630
rect 35168 4544 35184 4614
rect 35320 4544 35336 4614
rect 35168 4528 35336 4544
rect 35705 4424 35975 4458
rect 34879 4374 34913 4390
rect 34879 4182 34913 4198
rect 34997 4374 35031 4390
rect 34997 4182 35031 4198
rect 35115 4374 35149 4390
rect 35115 4182 35149 4198
rect 35233 4374 35267 4390
rect 35233 4182 35267 4198
rect 35351 4374 35385 4390
rect 35351 4182 35385 4198
rect 35469 4374 35503 4390
rect 35469 4182 35503 4198
rect 35587 4374 35621 4390
rect 35587 4182 35621 4198
rect 35705 4374 35739 4424
rect 35705 4182 35739 4198
rect 35823 4374 35857 4390
rect 35823 4182 35857 4198
rect 35941 4374 35975 4424
rect 35941 4182 35975 4198
rect 35630 4104 35646 4138
rect 35680 4104 35696 4138
rect 35512 3987 35528 4021
rect 35562 3987 35578 4021
rect 35116 3937 35150 3953
rect 35116 3545 35150 3561
rect 35234 3937 35268 3953
rect 35234 3545 35268 3561
rect 35352 3937 35386 3953
rect 35469 3937 35503 3953
rect 35469 3745 35503 3761
rect 35587 3937 35621 3953
rect 35587 3745 35621 3761
rect 35352 3545 35386 3561
rect 35159 3477 35175 3511
rect 35209 3477 35225 3511
rect 35277 3477 35293 3511
rect 35327 3477 35343 3511
rect 34641 3440 34906 3445
rect 34641 3387 34841 3440
rect 34901 3387 34906 3440
rect 34641 3383 34906 3387
rect 35392 3406 35560 3424
rect 35392 3350 35408 3406
rect 35542 3350 35560 3406
rect 35392 3334 35560 3350
rect 35184 1854 35352 1870
rect 35184 1784 35200 1854
rect 35336 1784 35352 1854
rect 35184 1768 35352 1784
rect 35721 1664 35991 1698
rect 34895 1614 34929 1630
rect 34895 1422 34929 1438
rect 35013 1614 35047 1630
rect 35013 1422 35047 1438
rect 35131 1614 35165 1630
rect 35131 1422 35165 1438
rect 35249 1614 35283 1630
rect 35249 1422 35283 1438
rect 35367 1614 35401 1630
rect 35367 1422 35401 1438
rect 35485 1614 35519 1630
rect 35485 1422 35519 1438
rect 35603 1614 35637 1630
rect 35603 1422 35637 1438
rect 35721 1614 35755 1664
rect 35721 1422 35755 1438
rect 35839 1614 35873 1630
rect 35839 1422 35873 1438
rect 35957 1614 35991 1664
rect 35957 1422 35991 1438
rect 35646 1344 35662 1378
rect 35696 1344 35712 1378
rect 35528 1227 35544 1261
rect 35578 1227 35594 1261
rect 35132 1177 35166 1193
rect 35132 785 35166 801
rect 35250 1177 35284 1193
rect 35250 785 35284 801
rect 35368 1177 35402 1193
rect 35485 1177 35519 1193
rect 35485 985 35519 1001
rect 35603 1177 35637 1193
rect 35603 985 35637 1001
rect 35368 785 35402 801
rect 35175 717 35191 751
rect 35225 717 35241 751
rect 35293 717 35309 751
rect 35343 717 35359 751
rect 35408 646 35576 664
rect 35408 590 35424 646
rect 35558 590 35576 646
rect 35408 574 35576 590
rect 34352 -2454 34543 -2445
rect 34352 -2520 34377 -2454
rect 34521 -2520 34543 -2454
rect 34352 -2528 34543 -2520
rect 33951 -2665 33962 -2594
rect 34076 -2665 34089 -2594
rect 33951 -2682 34089 -2665
rect 32528 -2726 33894 -2716
rect 36506 -2717 36633 10676
rect 38191 10385 38414 10460
rect 38191 10384 38271 10385
rect 38191 10235 38270 10384
rect 38338 10236 38414 10385
rect 38337 10235 38414 10236
rect 38191 10129 38414 10235
rect 40673 10438 40896 10514
rect 40673 10289 40752 10438
rect 40819 10435 40896 10438
rect 40673 10286 40753 10289
rect 40820 10286 40896 10435
rect 40006 10218 40040 10234
rect 40006 10168 40040 10184
rect 40673 10183 40896 10286
rect 41820 10438 42043 10514
rect 41820 10437 41899 10438
rect 41820 10288 41895 10437
rect 41966 10289 42043 10438
rect 41962 10288 42043 10289
rect 41136 10224 41170 10240
rect 41136 10174 41170 10190
rect 41820 10183 42043 10288
rect 44740 10473 44963 10548
rect 44740 10472 44820 10473
rect 44740 10323 44819 10472
rect 44887 10324 44963 10473
rect 44886 10323 44963 10324
rect 44740 10217 44963 10323
rect 47222 10526 47445 10602
rect 47222 10377 47301 10526
rect 47368 10524 47445 10526
rect 47222 10375 47303 10377
rect 47370 10375 47445 10524
rect 46555 10306 46589 10322
rect 46555 10256 46589 10272
rect 47222 10271 47445 10375
rect 48369 10526 48592 10602
rect 48369 10377 48447 10526
rect 48515 10377 48592 10526
rect 47685 10312 47719 10328
rect 47685 10262 47719 10278
rect 48369 10271 48592 10377
rect 51394 10404 51617 10480
rect 51394 10254 51473 10404
rect 51540 10254 51617 10404
rect 53876 10459 54099 10534
rect 53876 10310 53954 10459
rect 54021 10458 54099 10459
rect 53876 10309 53955 10310
rect 54022 10309 54099 10458
rect 46555 10188 46589 10204
rect 40006 10100 40040 10116
rect 38622 10020 38892 10054
rect 40006 10050 40040 10066
rect 41136 10104 41170 10120
rect 45171 10108 45441 10142
rect 46555 10138 46589 10154
rect 47685 10192 47719 10208
rect 37796 9970 37830 9986
rect 37796 9778 37830 9794
rect 37914 9970 37948 9986
rect 37914 9778 37948 9794
rect 38032 9970 38066 9986
rect 38032 9778 38066 9794
rect 38150 9970 38184 9986
rect 38150 9778 38184 9794
rect 38268 9970 38302 9986
rect 38268 9778 38302 9794
rect 38386 9970 38420 9986
rect 38386 9778 38420 9794
rect 38504 9970 38538 9986
rect 38504 9778 38538 9794
rect 38622 9970 38656 10020
rect 38622 9778 38656 9794
rect 38740 9970 38774 9986
rect 38740 9778 38774 9794
rect 38858 9970 38892 10020
rect 38858 9778 38892 9794
rect 40121 10042 40155 10058
rect 38547 9700 38563 9734
rect 38597 9700 38613 9734
rect 40121 9650 40155 9666
rect 40239 10042 40273 10058
rect 40239 9650 40273 9666
rect 40357 10042 40391 10058
rect 40357 9650 40391 9666
rect 40475 10042 40509 10058
rect 40475 9650 40509 9666
rect 40593 10042 40627 10058
rect 40593 9650 40627 9666
rect 40711 10042 40745 10058
rect 40711 9650 40745 9666
rect 40829 10042 40863 10058
rect 41136 10054 41170 10070
rect 40829 9650 40863 9666
rect 41263 10046 41297 10062
rect 41263 9654 41297 9670
rect 41381 10046 41415 10062
rect 41381 9654 41415 9670
rect 41499 10046 41533 10062
rect 41499 9654 41533 9670
rect 41617 10046 41651 10062
rect 41617 9654 41651 9670
rect 41735 10046 41769 10062
rect 41735 9654 41769 9670
rect 41853 10046 41887 10062
rect 41853 9654 41887 9670
rect 41971 10046 42005 10062
rect 44345 10058 44379 10074
rect 44345 9866 44379 9882
rect 44463 10058 44497 10074
rect 44463 9866 44497 9882
rect 44581 10058 44615 10074
rect 44581 9866 44615 9882
rect 44699 10058 44733 10074
rect 44699 9866 44733 9882
rect 44817 10058 44851 10074
rect 44817 9866 44851 9882
rect 44935 10058 44969 10074
rect 44935 9866 44969 9882
rect 45053 10058 45087 10074
rect 45053 9866 45087 9882
rect 45171 10058 45205 10108
rect 45171 9866 45205 9882
rect 45289 10058 45323 10074
rect 45289 9866 45323 9882
rect 45407 10058 45441 10108
rect 45407 9866 45441 9882
rect 46670 10130 46704 10146
rect 45096 9788 45112 9822
rect 45146 9788 45162 9822
rect 46670 9738 46704 9754
rect 46788 10130 46822 10146
rect 46788 9738 46822 9754
rect 46906 10130 46940 10146
rect 46906 9738 46940 9754
rect 47024 10130 47058 10146
rect 47024 9738 47058 9754
rect 47142 10130 47176 10146
rect 47142 9738 47176 9754
rect 47260 10130 47294 10146
rect 47260 9738 47294 9754
rect 47378 10130 47412 10146
rect 47685 10142 47719 10158
rect 47378 9738 47412 9754
rect 47812 10134 47846 10150
rect 47812 9742 47846 9758
rect 47930 10134 47964 10150
rect 47930 9742 47964 9758
rect 48048 10134 48082 10150
rect 48048 9742 48082 9758
rect 48166 10134 48200 10150
rect 48166 9742 48200 9758
rect 48284 10134 48318 10150
rect 48284 9742 48318 9758
rect 48402 10134 48436 10150
rect 48402 9742 48436 9758
rect 48520 10134 48554 10150
rect 51394 10149 51617 10254
rect 53209 10238 53243 10254
rect 53209 10188 53243 10204
rect 53876 10203 54099 10309
rect 55023 10458 55246 10534
rect 55023 10309 55101 10458
rect 55169 10309 55246 10458
rect 54339 10244 54373 10260
rect 54339 10194 54373 10210
rect 55023 10203 55246 10309
rect 58019 10472 58242 10548
rect 58019 10323 58093 10472
rect 58165 10323 58242 10472
rect 58019 10217 58242 10323
rect 60501 10526 60724 10602
rect 60501 10524 60580 10526
rect 60501 10375 60577 10524
rect 60647 10377 60724 10526
rect 60644 10375 60724 10377
rect 59834 10306 59868 10322
rect 59834 10256 59868 10272
rect 60501 10271 60724 10375
rect 61648 10530 61871 10602
rect 61648 10381 61726 10530
rect 61793 10526 61871 10530
rect 61648 10377 61727 10381
rect 61794 10377 61871 10526
rect 60964 10312 60998 10328
rect 60964 10262 60998 10278
rect 61648 10271 61871 10377
rect 59834 10188 59868 10204
rect 53209 10120 53243 10136
rect 51825 10040 52095 10074
rect 53209 10070 53243 10086
rect 54339 10124 54373 10140
rect 50999 9990 51033 10006
rect 50999 9798 51033 9814
rect 51117 9990 51151 10006
rect 51117 9798 51151 9814
rect 51235 9990 51269 10006
rect 51235 9798 51269 9814
rect 51353 9990 51387 10006
rect 51353 9798 51387 9814
rect 51471 9990 51505 10006
rect 51471 9798 51505 9814
rect 51589 9990 51623 10006
rect 51589 9798 51623 9814
rect 51707 9990 51741 10006
rect 51707 9798 51741 9814
rect 51825 9990 51859 10040
rect 51825 9798 51859 9814
rect 51943 9990 51977 10006
rect 51943 9798 51977 9814
rect 52061 9990 52095 10040
rect 52061 9798 52095 9814
rect 53324 10062 53358 10078
rect 48520 9742 48554 9758
rect 51750 9720 51766 9754
rect 51800 9720 51816 9754
rect 44978 9671 44994 9705
rect 45028 9671 45044 9705
rect 53324 9670 53358 9686
rect 53442 10062 53476 10078
rect 53442 9670 53476 9686
rect 53560 10062 53594 10078
rect 53560 9670 53594 9686
rect 53678 10062 53712 10078
rect 53678 9670 53712 9686
rect 53796 10062 53830 10078
rect 53796 9670 53830 9686
rect 53914 10062 53948 10078
rect 53914 9670 53948 9686
rect 54032 10062 54066 10078
rect 54339 10074 54373 10090
rect 58450 10108 58720 10142
rect 59834 10138 59868 10154
rect 60964 10192 60998 10208
rect 54032 9670 54066 9686
rect 54466 10066 54500 10082
rect 54466 9674 54500 9690
rect 54584 10066 54618 10082
rect 54584 9674 54618 9690
rect 54702 10066 54736 10082
rect 54702 9674 54736 9690
rect 54820 10066 54854 10082
rect 54820 9674 54854 9690
rect 54938 10066 54972 10082
rect 54938 9674 54972 9690
rect 55056 10066 55090 10082
rect 55056 9674 55090 9690
rect 55174 10066 55208 10082
rect 57624 10058 57658 10074
rect 57624 9866 57658 9882
rect 57742 10058 57776 10074
rect 57742 9866 57776 9882
rect 57860 10058 57894 10074
rect 57860 9866 57894 9882
rect 57978 10058 58012 10074
rect 57978 9866 58012 9882
rect 58096 10058 58130 10074
rect 58096 9866 58130 9882
rect 58214 10058 58248 10074
rect 58214 9866 58248 9882
rect 58332 10058 58366 10074
rect 58332 9866 58366 9882
rect 58450 10058 58484 10108
rect 58450 9866 58484 9882
rect 58568 10058 58602 10074
rect 58568 9866 58602 9882
rect 58686 10058 58720 10108
rect 58686 9866 58720 9882
rect 59949 10130 59983 10146
rect 58375 9788 58391 9822
rect 58425 9788 58441 9822
rect 59949 9738 59983 9754
rect 60067 10130 60101 10146
rect 60067 9738 60101 9754
rect 60185 10130 60219 10146
rect 60185 9738 60219 9754
rect 60303 10130 60337 10146
rect 60303 9738 60337 9754
rect 60421 10130 60455 10146
rect 60421 9738 60455 9754
rect 60539 10130 60573 10146
rect 60539 9738 60573 9754
rect 60657 10130 60691 10146
rect 60964 10142 60998 10158
rect 60657 9738 60691 9754
rect 61091 10134 61125 10150
rect 61091 9742 61125 9758
rect 61209 10134 61243 10150
rect 61209 9742 61243 9758
rect 61327 10134 61361 10150
rect 61327 9742 61361 9758
rect 61445 10134 61479 10150
rect 61445 9742 61479 9758
rect 61563 10134 61597 10150
rect 61563 9742 61597 9758
rect 61681 10134 61715 10150
rect 61681 9742 61715 9758
rect 61799 10134 61833 10150
rect 61799 9742 61833 9758
rect 55174 9674 55208 9690
rect 58257 9671 58273 9705
rect 58307 9671 58323 9705
rect 41971 9654 42005 9670
rect 63710 9659 63878 9675
rect 44582 9621 44616 9637
rect 38429 9583 38445 9617
rect 38479 9583 38495 9617
rect 38033 9533 38067 9549
rect 38033 9141 38067 9157
rect 38151 9533 38185 9549
rect 38151 9141 38185 9157
rect 38269 9533 38303 9549
rect 38386 9533 38420 9549
rect 38386 9341 38420 9357
rect 38504 9533 38538 9549
rect 38504 9341 38538 9357
rect 40310 9310 40326 9344
rect 40360 9310 40376 9344
rect 41452 9314 41468 9348
rect 41502 9314 41518 9348
rect 40031 9259 40065 9275
rect 38269 9141 38303 9157
rect 38556 9207 38805 9250
rect 38556 9117 38603 9207
rect 38766 9117 38805 9207
rect 38076 9073 38092 9107
rect 38126 9073 38142 9107
rect 38194 9073 38210 9107
rect 38244 9073 38260 9107
rect 38556 9078 38805 9117
rect 40031 9067 40065 9083
rect 40149 9259 40183 9275
rect 40149 9067 40183 9083
rect 40267 9259 40301 9275
rect 40267 9067 40301 9083
rect 40385 9259 40419 9275
rect 40385 9067 40419 9083
rect 40550 9259 40584 9275
rect 40550 9067 40584 9083
rect 40668 9259 40702 9275
rect 40668 9067 40702 9083
rect 40786 9259 40820 9275
rect 40786 9067 40820 9083
rect 40904 9259 40938 9275
rect 40904 9067 40938 9083
rect 41173 9263 41207 9279
rect 41173 9071 41207 9087
rect 41291 9263 41325 9279
rect 41291 9071 41325 9087
rect 41409 9263 41443 9279
rect 41409 9071 41443 9087
rect 41527 9263 41561 9279
rect 41527 9071 41561 9087
rect 41692 9263 41726 9279
rect 41692 9071 41726 9087
rect 41810 9263 41844 9279
rect 41810 9071 41844 9087
rect 41928 9263 41962 9279
rect 41928 9071 41962 9087
rect 42046 9263 42080 9279
rect 44582 9229 44616 9245
rect 44700 9621 44734 9637
rect 44700 9229 44734 9245
rect 44818 9621 44852 9637
rect 44935 9621 44969 9637
rect 44935 9429 44969 9445
rect 45053 9621 45087 9637
rect 51632 9603 51648 9637
rect 51682 9603 51698 9637
rect 57861 9621 57895 9637
rect 45053 9429 45087 9445
rect 51236 9553 51270 9569
rect 46859 9398 46875 9432
rect 46909 9398 46925 9432
rect 48001 9402 48017 9436
rect 48051 9402 48067 9436
rect 46580 9347 46614 9363
rect 44818 9229 44852 9245
rect 45105 9295 45354 9338
rect 45105 9205 45152 9295
rect 45315 9205 45354 9295
rect 44625 9161 44641 9195
rect 44675 9161 44691 9195
rect 44743 9161 44759 9195
rect 44793 9161 44809 9195
rect 45105 9166 45354 9205
rect 46580 9155 46614 9171
rect 46698 9347 46732 9363
rect 46698 9155 46732 9171
rect 46816 9347 46850 9363
rect 46816 9155 46850 9171
rect 46934 9347 46968 9363
rect 46934 9155 46968 9171
rect 47099 9347 47133 9363
rect 47099 9155 47133 9171
rect 47217 9347 47251 9363
rect 47217 9155 47251 9171
rect 47335 9347 47369 9363
rect 47335 9155 47369 9171
rect 47453 9347 47487 9363
rect 47453 9155 47487 9171
rect 47722 9351 47756 9367
rect 47722 9159 47756 9175
rect 47840 9351 47874 9367
rect 47840 9159 47874 9175
rect 47958 9351 47992 9367
rect 47958 9159 47992 9175
rect 48076 9351 48110 9367
rect 48076 9159 48110 9175
rect 48241 9351 48275 9367
rect 48241 9159 48275 9175
rect 48359 9351 48393 9367
rect 48359 9159 48393 9175
rect 48477 9351 48511 9367
rect 48477 9159 48511 9175
rect 48595 9351 48629 9367
rect 48595 9159 48629 9175
rect 51236 9161 51270 9177
rect 51354 9553 51388 9569
rect 51354 9161 51388 9177
rect 51472 9553 51506 9569
rect 51589 9553 51623 9569
rect 51589 9361 51623 9377
rect 51707 9553 51741 9569
rect 51707 9361 51741 9377
rect 53513 9330 53529 9364
rect 53563 9330 53579 9364
rect 54655 9334 54671 9368
rect 54705 9334 54721 9368
rect 53234 9279 53268 9295
rect 51472 9161 51506 9177
rect 51759 9227 52008 9270
rect 51759 9137 51806 9227
rect 51969 9137 52008 9227
rect 51279 9093 51295 9127
rect 51329 9093 51345 9127
rect 51397 9093 51413 9127
rect 51447 9093 51463 9127
rect 51759 9098 52008 9137
rect 53234 9087 53268 9103
rect 53352 9279 53386 9295
rect 53352 9087 53386 9103
rect 53470 9279 53504 9295
rect 53470 9087 53504 9103
rect 53588 9279 53622 9295
rect 53588 9087 53622 9103
rect 53753 9279 53787 9295
rect 53753 9087 53787 9103
rect 53871 9279 53905 9295
rect 53871 9087 53905 9103
rect 53989 9279 54023 9295
rect 53989 9087 54023 9103
rect 54107 9279 54141 9295
rect 54107 9087 54141 9103
rect 54376 9283 54410 9299
rect 54376 9091 54410 9107
rect 54494 9283 54528 9299
rect 54494 9091 54528 9107
rect 54612 9283 54646 9299
rect 54612 9091 54646 9107
rect 54730 9283 54764 9299
rect 54730 9091 54764 9107
rect 54895 9283 54929 9299
rect 54895 9091 54929 9107
rect 55013 9283 55047 9299
rect 55013 9091 55047 9107
rect 55131 9283 55165 9299
rect 55131 9091 55165 9107
rect 55249 9283 55283 9299
rect 57861 9229 57895 9245
rect 57979 9621 58013 9637
rect 57979 9229 58013 9245
rect 58097 9621 58131 9637
rect 58214 9621 58248 9637
rect 58214 9429 58248 9445
rect 58332 9621 58366 9637
rect 63710 9589 63726 9659
rect 63862 9589 63878 9659
rect 63710 9573 63878 9589
rect 58332 9429 58366 9445
rect 64247 9469 64517 9503
rect 60138 9398 60154 9432
rect 60188 9398 60204 9432
rect 61280 9402 61296 9436
rect 61330 9402 61346 9436
rect 63421 9419 63455 9435
rect 59859 9347 59893 9363
rect 58097 9229 58131 9245
rect 58384 9295 58633 9338
rect 58384 9205 58431 9295
rect 58594 9205 58633 9295
rect 57904 9161 57920 9195
rect 57954 9161 57970 9195
rect 58022 9161 58038 9195
rect 58072 9161 58088 9195
rect 58384 9166 58633 9205
rect 59859 9155 59893 9171
rect 59977 9347 60011 9363
rect 59977 9155 60011 9171
rect 60095 9347 60129 9363
rect 60095 9155 60129 9171
rect 60213 9347 60247 9363
rect 60213 9155 60247 9171
rect 60378 9347 60412 9363
rect 60378 9155 60412 9171
rect 60496 9347 60530 9363
rect 60496 9155 60530 9171
rect 60614 9347 60648 9363
rect 60614 9155 60648 9171
rect 60732 9347 60766 9363
rect 60732 9155 60766 9171
rect 61001 9351 61035 9367
rect 61001 9159 61035 9175
rect 61119 9351 61153 9367
rect 61119 9159 61153 9175
rect 61237 9351 61271 9367
rect 61237 9159 61271 9175
rect 61355 9351 61389 9367
rect 61355 9159 61389 9175
rect 61520 9351 61554 9367
rect 61520 9159 61554 9175
rect 61638 9351 61672 9367
rect 61638 9159 61672 9175
rect 61756 9351 61790 9367
rect 61756 9159 61790 9175
rect 61874 9351 61908 9367
rect 63421 9227 63455 9243
rect 63539 9419 63573 9435
rect 63539 9227 63573 9243
rect 63657 9419 63691 9435
rect 63657 9227 63691 9243
rect 63775 9419 63809 9435
rect 63775 9227 63809 9243
rect 63893 9419 63927 9435
rect 63893 9227 63927 9243
rect 64011 9419 64045 9435
rect 64011 9227 64045 9243
rect 64129 9419 64163 9435
rect 64129 9227 64163 9243
rect 64247 9419 64281 9469
rect 64247 9227 64281 9243
rect 64365 9419 64399 9435
rect 64365 9227 64399 9243
rect 64483 9419 64517 9469
rect 64483 9227 64517 9243
rect 61874 9159 61908 9175
rect 64172 9149 64188 9183
rect 64222 9149 64238 9183
rect 55249 9091 55283 9107
rect 42046 9071 42080 9087
rect 64054 9032 64070 9066
rect 64104 9032 64120 9066
rect 63658 8982 63692 8998
rect 46595 8924 46767 8971
rect 40046 8836 40218 8883
rect 38205 8734 38428 8810
rect 38205 8585 38283 8734
rect 38351 8585 38428 8734
rect 40046 8673 40085 8836
rect 40175 8673 40218 8836
rect 40046 8634 40218 8673
rect 41188 8834 41360 8881
rect 41188 8671 41227 8834
rect 41317 8671 41360 8834
rect 41188 8632 41360 8671
rect 44754 8822 44977 8898
rect 44754 8673 44833 8822
rect 44900 8821 44977 8822
rect 44754 8672 44834 8673
rect 44901 8672 44977 8821
rect 46595 8761 46634 8924
rect 46724 8761 46767 8924
rect 46595 8722 46767 8761
rect 47737 8922 47909 8969
rect 47737 8759 47776 8922
rect 47866 8759 47909 8922
rect 59874 8924 60046 8971
rect 53249 8856 53421 8903
rect 47737 8720 47909 8759
rect 51408 8755 51631 8830
rect 51408 8754 51488 8755
rect 38205 8479 38428 8585
rect 44754 8567 44977 8672
rect 51408 8605 51487 8754
rect 51555 8606 51631 8755
rect 53249 8693 53288 8856
rect 53378 8693 53421 8856
rect 53249 8654 53421 8693
rect 54391 8854 54563 8901
rect 54391 8691 54430 8854
rect 54520 8691 54563 8854
rect 54391 8652 54563 8691
rect 58033 8822 58256 8898
rect 58033 8673 58112 8822
rect 58179 8821 58256 8822
rect 58033 8672 58116 8673
rect 58183 8672 58256 8821
rect 59874 8761 59913 8924
rect 60003 8761 60046 8924
rect 59874 8759 59917 8761
rect 59984 8759 60046 8761
rect 59874 8722 60046 8759
rect 61016 8922 61188 8969
rect 61016 8759 61055 8922
rect 61145 8759 61188 8922
rect 61016 8720 61188 8759
rect 51554 8605 51631 8606
rect 38636 8370 38906 8404
rect 37810 8320 37844 8336
rect 37810 8128 37844 8144
rect 37928 8320 37962 8336
rect 37928 8128 37962 8144
rect 38046 8320 38080 8336
rect 38046 8128 38080 8144
rect 38164 8320 38198 8336
rect 38164 8128 38198 8144
rect 38282 8320 38316 8336
rect 38282 8128 38316 8144
rect 38400 8320 38434 8336
rect 38400 8128 38434 8144
rect 38518 8320 38552 8336
rect 38518 8128 38552 8144
rect 38636 8320 38670 8370
rect 38636 8128 38670 8144
rect 38754 8320 38788 8336
rect 38754 8128 38788 8144
rect 38872 8320 38906 8370
rect 38872 8128 38906 8144
rect 41916 8392 42141 8467
rect 45185 8458 45455 8492
rect 41916 8242 41995 8392
rect 42062 8242 42141 8392
rect 41916 8136 42141 8242
rect 44359 8408 44393 8424
rect 44359 8216 44393 8232
rect 44477 8408 44511 8424
rect 44477 8216 44511 8232
rect 44595 8408 44629 8424
rect 44595 8216 44629 8232
rect 44713 8408 44747 8424
rect 44713 8216 44747 8232
rect 44831 8408 44865 8424
rect 44831 8216 44865 8232
rect 44949 8408 44983 8424
rect 44949 8216 44983 8232
rect 45067 8408 45101 8424
rect 45067 8216 45101 8232
rect 45185 8408 45219 8458
rect 45185 8216 45219 8232
rect 45303 8408 45337 8424
rect 45303 8216 45337 8232
rect 45421 8408 45455 8458
rect 45421 8216 45455 8232
rect 48465 8479 48690 8555
rect 51408 8499 51631 8605
rect 58033 8567 58256 8672
rect 63658 8590 63692 8606
rect 63776 8982 63810 8998
rect 63776 8590 63810 8606
rect 63894 8982 63928 8998
rect 64011 8982 64045 8998
rect 64011 8790 64045 8806
rect 64129 8982 64163 8998
rect 64129 8790 64163 8806
rect 63894 8590 63928 8606
rect 48465 8330 48544 8479
rect 48616 8330 48690 8479
rect 51839 8390 52109 8424
rect 48465 8224 48690 8330
rect 51013 8340 51047 8356
rect 45110 8138 45126 8172
rect 45160 8138 45176 8172
rect 51013 8148 51047 8164
rect 51131 8340 51165 8356
rect 51131 8148 51165 8164
rect 51249 8340 51283 8356
rect 51249 8148 51283 8164
rect 51367 8340 51401 8356
rect 51367 8148 51401 8164
rect 51485 8340 51519 8356
rect 51485 8148 51519 8164
rect 51603 8340 51637 8356
rect 51603 8148 51637 8164
rect 51721 8340 51755 8356
rect 51721 8148 51755 8164
rect 51839 8340 51873 8390
rect 51839 8148 51873 8164
rect 51957 8340 51991 8356
rect 51957 8148 51991 8164
rect 52075 8340 52109 8390
rect 52075 8148 52109 8164
rect 55119 8411 55344 8487
rect 58464 8458 58734 8492
rect 55119 8407 55198 8411
rect 55119 8258 55195 8407
rect 55265 8262 55344 8411
rect 55262 8258 55344 8262
rect 55119 8156 55344 8258
rect 57638 8408 57672 8424
rect 57638 8216 57672 8232
rect 57756 8408 57790 8424
rect 57756 8216 57790 8232
rect 57874 8408 57908 8424
rect 57874 8216 57908 8232
rect 57992 8408 58026 8424
rect 57992 8216 58026 8232
rect 58110 8408 58144 8424
rect 58110 8216 58144 8232
rect 58228 8408 58262 8424
rect 58228 8216 58262 8232
rect 58346 8408 58380 8424
rect 58346 8216 58380 8232
rect 58464 8408 58498 8458
rect 58464 8216 58498 8232
rect 58582 8408 58616 8424
rect 58582 8216 58616 8232
rect 58700 8408 58734 8458
rect 58700 8216 58734 8232
rect 61744 8479 61969 8555
rect 63701 8522 63717 8556
rect 63751 8522 63767 8556
rect 63819 8522 63835 8556
rect 63869 8522 63885 8556
rect 61744 8327 61823 8479
rect 61890 8327 61969 8479
rect 63934 8451 64102 8469
rect 63934 8395 63950 8451
rect 64084 8395 64102 8451
rect 63934 8379 64102 8395
rect 61744 8224 61969 8327
rect 58389 8138 58405 8172
rect 58439 8138 58455 8172
rect 38561 8050 38577 8084
rect 38611 8050 38627 8084
rect 44992 8021 45008 8055
rect 45042 8021 45058 8055
rect 46661 8044 46931 8079
rect 46307 7991 46341 8007
rect 38443 7933 38459 7967
rect 38493 7933 38509 7967
rect 40112 7956 40382 7991
rect 39758 7903 39792 7919
rect 38047 7883 38081 7899
rect 36901 7543 37161 7545
rect 36899 7514 37161 7543
rect 36899 7404 37008 7514
rect 37126 7404 37161 7514
rect 38047 7491 38081 7507
rect 38165 7883 38199 7899
rect 38165 7491 38199 7507
rect 38283 7883 38317 7899
rect 38400 7883 38434 7899
rect 38400 7691 38434 7707
rect 38518 7883 38552 7899
rect 38518 7691 38552 7707
rect 39274 7757 39544 7792
rect 39274 7703 39308 7757
rect 38283 7491 38317 7507
rect 38570 7557 38819 7600
rect 38570 7467 38617 7557
rect 38780 7467 38819 7557
rect 39274 7511 39308 7527
rect 39392 7703 39426 7719
rect 39392 7511 39426 7527
rect 39510 7703 39544 7757
rect 39510 7511 39544 7527
rect 39628 7703 39662 7719
rect 39628 7511 39662 7527
rect 39758 7511 39792 7527
rect 39876 7903 39910 7919
rect 39876 7511 39910 7527
rect 39994 7903 40028 7919
rect 39994 7511 40028 7527
rect 40112 7903 40146 7956
rect 40112 7511 40146 7527
rect 40230 7903 40264 7919
rect 40230 7511 40264 7527
rect 40348 7903 40382 7956
rect 42010 7956 42280 7991
rect 40348 7511 40382 7527
rect 40466 7903 40500 7919
rect 41656 7903 41690 7919
rect 41172 7757 41442 7792
rect 40466 7511 40500 7527
rect 40595 7703 40629 7719
rect 40595 7511 40629 7527
rect 40713 7703 40747 7719
rect 40713 7511 40747 7527
rect 40831 7703 40865 7719
rect 40831 7511 40865 7527
rect 40949 7703 40983 7719
rect 40949 7511 40983 7527
rect 41172 7703 41206 7757
rect 41172 7511 41206 7527
rect 41290 7703 41324 7719
rect 41290 7511 41324 7527
rect 41408 7703 41442 7757
rect 41408 7511 41442 7527
rect 41526 7703 41560 7719
rect 41526 7511 41560 7527
rect 41656 7511 41690 7527
rect 41774 7903 41808 7919
rect 41774 7511 41808 7527
rect 41892 7903 41926 7919
rect 41892 7511 41926 7527
rect 42010 7903 42044 7956
rect 42010 7511 42044 7527
rect 42128 7903 42162 7919
rect 42128 7511 42162 7527
rect 42246 7903 42280 7956
rect 44596 7971 44630 7987
rect 42246 7511 42280 7527
rect 42364 7903 42398 7919
rect 42364 7511 42398 7527
rect 42493 7703 42527 7719
rect 42493 7511 42527 7527
rect 42611 7703 42645 7719
rect 42611 7511 42645 7527
rect 42729 7703 42763 7719
rect 42729 7511 42763 7527
rect 42847 7703 42881 7719
rect 44596 7579 44630 7595
rect 44714 7971 44748 7987
rect 44714 7579 44748 7595
rect 44832 7971 44866 7987
rect 44949 7971 44983 7987
rect 44949 7779 44983 7795
rect 45067 7971 45101 7987
rect 45067 7779 45101 7795
rect 45823 7845 46093 7880
rect 45823 7791 45857 7845
rect 44832 7579 44866 7595
rect 45119 7645 45368 7688
rect 45119 7555 45166 7645
rect 45329 7555 45368 7645
rect 45823 7599 45857 7615
rect 45941 7791 45975 7807
rect 45941 7599 45975 7615
rect 46059 7791 46093 7845
rect 46059 7599 46093 7615
rect 46177 7791 46211 7807
rect 46177 7599 46211 7615
rect 46307 7599 46341 7615
rect 46425 7991 46459 8007
rect 46425 7599 46459 7615
rect 46543 7991 46577 8007
rect 46543 7599 46577 7615
rect 46661 7991 46695 8044
rect 46661 7599 46695 7615
rect 46779 7991 46813 8007
rect 46779 7599 46813 7615
rect 46897 7991 46931 8044
rect 48559 8044 48829 8079
rect 51764 8070 51780 8104
rect 51814 8070 51830 8104
rect 46897 7599 46931 7615
rect 47015 7991 47049 8007
rect 48205 7991 48239 8007
rect 47721 7845 47991 7880
rect 47015 7599 47049 7615
rect 47144 7791 47178 7807
rect 47144 7599 47178 7615
rect 47262 7791 47296 7807
rect 47262 7599 47296 7615
rect 47380 7791 47414 7807
rect 47380 7599 47414 7615
rect 47498 7791 47532 7807
rect 47498 7599 47532 7615
rect 47721 7791 47755 7845
rect 47721 7599 47755 7615
rect 47839 7791 47873 7807
rect 47839 7599 47873 7615
rect 47957 7791 47991 7845
rect 47957 7599 47991 7615
rect 48075 7791 48109 7807
rect 48075 7599 48109 7615
rect 48205 7599 48239 7615
rect 48323 7991 48357 8007
rect 48323 7599 48357 7615
rect 48441 7991 48475 8007
rect 48441 7599 48475 7615
rect 48559 7991 48593 8044
rect 48559 7599 48593 7615
rect 48677 7991 48711 8007
rect 48677 7599 48711 7615
rect 48795 7991 48829 8044
rect 58271 8021 58287 8055
rect 58321 8021 58337 8055
rect 59940 8044 60210 8079
rect 48795 7599 48829 7615
rect 48913 7991 48947 8007
rect 51646 7953 51662 7987
rect 51696 7953 51712 7987
rect 53315 7976 53585 8011
rect 52961 7923 52995 7939
rect 51250 7903 51284 7919
rect 48913 7599 48947 7615
rect 49042 7791 49076 7807
rect 49042 7599 49076 7615
rect 49160 7791 49194 7807
rect 49160 7599 49194 7615
rect 49278 7791 49312 7807
rect 49278 7599 49312 7615
rect 49396 7791 49430 7807
rect 49396 7599 49430 7615
rect 42847 7511 42881 7527
rect 44639 7511 44655 7545
rect 44689 7511 44705 7545
rect 44757 7511 44773 7545
rect 44807 7511 44823 7545
rect 45119 7516 45368 7555
rect 50144 7543 50370 7565
rect 38090 7423 38106 7457
rect 38140 7423 38156 7457
rect 38208 7423 38224 7457
rect 38258 7423 38274 7457
rect 38570 7428 38819 7467
rect 50144 7426 50210 7543
rect 50349 7426 50370 7543
rect 51250 7511 51284 7527
rect 51368 7903 51402 7919
rect 51368 7511 51402 7527
rect 51486 7903 51520 7919
rect 51603 7903 51637 7919
rect 51603 7711 51637 7727
rect 51721 7903 51755 7919
rect 51721 7711 51755 7727
rect 52477 7777 52747 7812
rect 52477 7723 52511 7777
rect 51486 7511 51520 7527
rect 51773 7577 52022 7620
rect 51773 7487 51820 7577
rect 51983 7487 52022 7577
rect 52477 7531 52511 7547
rect 52595 7723 52629 7739
rect 52595 7531 52629 7547
rect 52713 7723 52747 7777
rect 52713 7531 52747 7547
rect 52831 7723 52865 7739
rect 52831 7531 52865 7547
rect 52961 7531 52995 7547
rect 53079 7923 53113 7939
rect 53079 7531 53113 7547
rect 53197 7923 53231 7939
rect 53197 7531 53231 7547
rect 53315 7923 53349 7976
rect 53315 7531 53349 7547
rect 53433 7923 53467 7939
rect 53433 7531 53467 7547
rect 53551 7923 53585 7976
rect 55213 7976 55483 8011
rect 59586 7991 59620 8007
rect 53551 7531 53585 7547
rect 53669 7923 53703 7939
rect 54859 7923 54893 7939
rect 54375 7777 54645 7812
rect 53669 7531 53703 7547
rect 53798 7723 53832 7739
rect 53798 7531 53832 7547
rect 53916 7723 53950 7739
rect 53916 7531 53950 7547
rect 54034 7723 54068 7739
rect 54034 7531 54068 7547
rect 54152 7723 54186 7739
rect 54152 7531 54186 7547
rect 54375 7723 54409 7777
rect 54375 7531 54409 7547
rect 54493 7723 54527 7739
rect 54493 7531 54527 7547
rect 54611 7723 54645 7777
rect 54611 7531 54645 7547
rect 54729 7723 54763 7739
rect 54729 7531 54763 7547
rect 54859 7531 54893 7547
rect 54977 7923 55011 7939
rect 54977 7531 55011 7547
rect 55095 7923 55129 7939
rect 55095 7531 55129 7547
rect 55213 7923 55247 7976
rect 55213 7531 55247 7547
rect 55331 7923 55365 7939
rect 55331 7531 55365 7547
rect 55449 7923 55483 7976
rect 57875 7971 57909 7987
rect 55449 7531 55483 7547
rect 55567 7923 55601 7939
rect 55567 7531 55601 7547
rect 55696 7723 55730 7739
rect 55696 7531 55730 7547
rect 55814 7723 55848 7739
rect 55814 7531 55848 7547
rect 55932 7723 55966 7739
rect 55932 7531 55966 7547
rect 56050 7723 56084 7739
rect 57875 7579 57909 7595
rect 57993 7971 58027 7987
rect 57993 7579 58027 7595
rect 58111 7971 58145 7987
rect 58228 7971 58262 7987
rect 58228 7779 58262 7795
rect 58346 7971 58380 7987
rect 58346 7779 58380 7795
rect 59102 7845 59372 7880
rect 59102 7791 59136 7845
rect 58111 7579 58145 7595
rect 58398 7645 58647 7688
rect 56050 7531 56084 7547
rect 58398 7555 58445 7645
rect 58608 7555 58647 7645
rect 59102 7599 59136 7615
rect 59220 7791 59254 7807
rect 59220 7599 59254 7615
rect 59338 7791 59372 7845
rect 59338 7599 59372 7615
rect 59456 7791 59490 7807
rect 59456 7599 59490 7615
rect 59586 7599 59620 7615
rect 59704 7991 59738 8007
rect 59704 7599 59738 7615
rect 59822 7991 59856 8007
rect 59822 7599 59856 7615
rect 59940 7991 59974 8044
rect 59940 7599 59974 7615
rect 60058 7991 60092 8007
rect 60058 7599 60092 7615
rect 60176 7991 60210 8044
rect 61838 8044 62108 8079
rect 60176 7599 60210 7615
rect 60294 7991 60328 8007
rect 61484 7991 61518 8007
rect 61000 7845 61270 7880
rect 60294 7599 60328 7615
rect 60423 7791 60457 7807
rect 60423 7599 60457 7615
rect 60541 7791 60575 7807
rect 60541 7599 60575 7615
rect 60659 7791 60693 7807
rect 60659 7599 60693 7615
rect 60777 7791 60811 7807
rect 60777 7599 60811 7615
rect 61000 7791 61034 7845
rect 61000 7599 61034 7615
rect 61118 7791 61152 7807
rect 61118 7599 61152 7615
rect 61236 7791 61270 7845
rect 61236 7599 61270 7615
rect 61354 7791 61388 7807
rect 61354 7599 61388 7615
rect 61484 7599 61518 7615
rect 61602 7991 61636 8007
rect 61602 7599 61636 7615
rect 61720 7991 61754 8007
rect 61720 7599 61754 7615
rect 61838 7991 61872 8044
rect 61838 7599 61872 7615
rect 61956 7991 61990 8007
rect 61956 7599 61990 7615
rect 62074 7991 62108 8044
rect 62074 7599 62108 7615
rect 62192 7991 62226 8007
rect 62192 7599 62226 7615
rect 62321 7791 62355 7807
rect 62321 7599 62355 7615
rect 62439 7791 62473 7807
rect 62439 7599 62473 7615
rect 62557 7791 62591 7807
rect 62557 7599 62591 7615
rect 62675 7791 62709 7807
rect 62675 7599 62709 7615
rect 57918 7511 57934 7545
rect 57968 7511 57984 7545
rect 58036 7511 58052 7545
rect 58086 7511 58102 7545
rect 58398 7516 58647 7555
rect 51293 7443 51309 7477
rect 51343 7443 51359 7477
rect 51411 7443 51427 7477
rect 51461 7443 51477 7477
rect 51773 7448 52022 7487
rect 50144 7414 50370 7426
rect 36899 7394 37161 7404
rect 36899 4996 37063 7394
rect 47287 7377 47321 7393
rect 47287 7327 47321 7343
rect 49377 7356 49444 7372
rect 49377 7322 49394 7356
rect 49428 7322 49444 7356
rect 40738 7289 40772 7305
rect 46250 7298 46284 7314
rect 40738 7239 40772 7255
rect 42828 7268 42895 7284
rect 42828 7234 42845 7268
rect 42879 7234 42895 7268
rect 39701 7210 39735 7226
rect 38200 7130 38423 7206
rect 38200 6981 38279 7130
rect 38346 7128 38423 7130
rect 38200 6979 38281 6981
rect 38348 6979 38423 7128
rect 38200 6875 38423 6979
rect 39819 7210 39853 7226
rect 39701 6818 39735 6834
rect 39818 6834 39819 6881
rect 39937 7210 39971 7226
rect 39853 6834 39854 6881
rect 38631 6766 38901 6800
rect 37805 6716 37839 6732
rect 37805 6524 37839 6540
rect 37923 6716 37957 6732
rect 37923 6524 37957 6540
rect 38041 6716 38075 6732
rect 38041 6524 38075 6540
rect 38159 6716 38193 6732
rect 38159 6524 38193 6540
rect 38277 6716 38311 6732
rect 38277 6524 38311 6540
rect 38395 6716 38429 6732
rect 38395 6524 38429 6540
rect 38513 6716 38547 6732
rect 38513 6524 38547 6540
rect 38631 6716 38665 6766
rect 38631 6524 38665 6540
rect 38749 6716 38783 6732
rect 38749 6524 38783 6540
rect 38867 6716 38901 6766
rect 39818 6776 39854 6834
rect 40055 7210 40089 7226
rect 39937 6818 39971 6834
rect 40053 6834 40055 6881
rect 40053 6776 40089 6834
rect 40173 7210 40207 7226
rect 40173 6818 40207 6834
rect 40291 7210 40325 7226
rect 40409 7210 40443 7226
rect 40325 6834 40327 6880
rect 40291 6776 40327 6834
rect 40409 6818 40443 6834
rect 41599 7210 41633 7226
rect 41717 7210 41751 7226
rect 41599 6818 41633 6834
rect 41716 6834 41717 6881
rect 41835 7210 41869 7226
rect 41751 6834 41752 6881
rect 40914 6776 41411 6794
rect 39818 6773 41411 6776
rect 39818 6739 41359 6773
rect 41393 6739 41411 6773
rect 39818 6736 41411 6739
rect 41716 6776 41752 6834
rect 41953 7210 41987 7226
rect 41835 6818 41869 6834
rect 41951 6834 41953 6881
rect 41951 6776 41987 6834
rect 42071 7210 42105 7226
rect 42071 6818 42105 6834
rect 42189 7210 42223 7226
rect 42307 7210 42341 7226
rect 42828 7218 42895 7234
rect 44749 7221 44972 7294
rect 42223 6834 42225 6880
rect 42189 6776 42225 6834
rect 44749 7072 44826 7221
rect 44893 7218 44972 7221
rect 44749 7069 44828 7072
rect 44895 7069 44972 7218
rect 44749 6963 44972 7069
rect 46368 7298 46402 7314
rect 46250 6906 46284 6922
rect 46367 6922 46368 6969
rect 46486 7298 46520 7314
rect 46402 6922 46403 6969
rect 42307 6818 42341 6834
rect 45180 6854 45450 6888
rect 42812 6776 43075 6806
rect 41716 6736 43075 6776
rect 39837 6735 41411 6736
rect 41735 6735 43075 6736
rect 39715 6646 39782 6662
rect 39715 6612 39731 6646
rect 39765 6612 39782 6646
rect 39715 6596 39782 6612
rect 38867 6524 38901 6540
rect 39546 6579 39580 6595
rect 39546 6529 39580 6545
rect 39892 6494 39926 6735
rect 40914 6718 41411 6735
rect 40362 6646 40429 6662
rect 40362 6612 40379 6646
rect 40413 6612 40429 6646
rect 40362 6596 40429 6612
rect 41613 6646 41680 6662
rect 41613 6612 41629 6646
rect 41663 6612 41680 6646
rect 41613 6596 41680 6612
rect 40669 6578 40703 6594
rect 39981 6528 39997 6562
rect 40031 6528 40047 6562
rect 40099 6529 40115 6563
rect 40149 6529 40165 6563
rect 40669 6528 40703 6544
rect 41444 6579 41478 6595
rect 41444 6529 41478 6545
rect 41790 6494 41824 6735
rect 42812 6706 43075 6735
rect 42258 6647 42325 6663
rect 42258 6613 42275 6647
rect 42309 6613 42325 6647
rect 42258 6597 42325 6613
rect 42567 6578 42601 6594
rect 41879 6528 41895 6562
rect 41929 6528 41945 6562
rect 41997 6529 42013 6563
rect 42047 6529 42063 6563
rect 42567 6528 42601 6544
rect 38556 6446 38572 6480
rect 38606 6446 38622 6480
rect 39399 6478 39433 6494
rect 38438 6329 38454 6363
rect 38488 6329 38504 6363
rect 38042 6279 38076 6295
rect 38042 5887 38076 5903
rect 38160 6279 38194 6295
rect 38160 5887 38194 5903
rect 38278 6279 38312 6295
rect 38395 6279 38429 6295
rect 38395 6087 38429 6103
rect 38513 6279 38547 6295
rect 39399 6286 39433 6302
rect 39517 6478 39551 6494
rect 39517 6286 39551 6302
rect 39819 6478 39853 6494
rect 38513 6087 38547 6103
rect 39892 6478 39971 6494
rect 39892 6448 39937 6478
rect 39819 6035 39854 6102
rect 39937 6086 39971 6102
rect 40055 6478 40089 6494
rect 40055 6086 40089 6102
rect 40173 6478 40207 6494
rect 40291 6478 40325 6494
rect 40697 6478 40731 6494
rect 40697 6286 40731 6302
rect 40815 6478 40849 6494
rect 40815 6286 40849 6302
rect 41297 6478 41331 6494
rect 41297 6286 41331 6302
rect 41415 6478 41449 6494
rect 41415 6286 41449 6302
rect 41717 6478 41751 6494
rect 40173 6086 40207 6102
rect 40290 6035 40325 6102
rect 39819 6000 40325 6035
rect 41790 6478 41869 6494
rect 41790 6448 41835 6478
rect 41717 6035 41752 6102
rect 41835 6086 41869 6102
rect 41953 6478 41987 6494
rect 41953 6086 41987 6102
rect 42071 6478 42105 6494
rect 42189 6478 42223 6494
rect 42595 6478 42629 6494
rect 42595 6286 42629 6302
rect 42713 6478 42747 6494
rect 42713 6286 42747 6302
rect 42071 6086 42105 6102
rect 42188 6035 42223 6102
rect 41717 6000 42223 6035
rect 38278 5887 38312 5903
rect 38565 5953 38814 5996
rect 38565 5863 38612 5953
rect 38775 5863 38814 5953
rect 38085 5819 38101 5853
rect 38135 5819 38151 5853
rect 38203 5819 38219 5853
rect 38253 5819 38269 5853
rect 38565 5824 38814 5863
rect 39990 5793 40162 5840
rect 39990 5630 40029 5793
rect 40119 5630 40162 5793
rect 39990 5590 40162 5630
rect 42943 5248 43075 6706
rect 44354 6804 44388 6820
rect 44354 6612 44388 6628
rect 44472 6804 44506 6820
rect 44472 6612 44506 6628
rect 44590 6804 44624 6820
rect 44590 6612 44624 6628
rect 44708 6804 44742 6820
rect 44708 6612 44742 6628
rect 44826 6804 44860 6820
rect 44826 6612 44860 6628
rect 44944 6804 44978 6820
rect 44944 6612 44978 6628
rect 45062 6804 45096 6820
rect 45062 6612 45096 6628
rect 45180 6804 45214 6854
rect 45180 6612 45214 6628
rect 45298 6804 45332 6820
rect 45298 6612 45332 6628
rect 45416 6804 45450 6854
rect 46367 6864 46403 6922
rect 46604 7298 46638 7314
rect 46486 6906 46520 6922
rect 46602 6922 46604 6969
rect 46602 6864 46638 6922
rect 46722 7298 46756 7314
rect 46722 6906 46756 6922
rect 46840 7298 46874 7314
rect 46958 7298 46992 7314
rect 46874 6922 46876 6968
rect 46840 6864 46876 6922
rect 46958 6906 46992 6922
rect 48148 7298 48182 7314
rect 48266 7298 48300 7314
rect 48148 6906 48182 6922
rect 48265 6922 48266 6969
rect 48384 7298 48418 7314
rect 48300 6922 48301 6969
rect 47463 6864 47960 6882
rect 46367 6861 47960 6864
rect 46367 6827 47908 6861
rect 47942 6827 47960 6861
rect 46367 6824 47960 6827
rect 48265 6864 48301 6922
rect 48502 7298 48536 7314
rect 48384 6906 48418 6922
rect 48500 6922 48502 6969
rect 48500 6864 48536 6922
rect 48620 7298 48654 7314
rect 48620 6906 48654 6922
rect 48738 7298 48772 7314
rect 48856 7298 48890 7314
rect 49377 7306 49444 7322
rect 48772 6922 48774 6968
rect 48738 6864 48774 6922
rect 48856 6906 48890 6922
rect 49361 6893 49461 6894
rect 49361 6864 49517 6893
rect 48265 6824 49517 6864
rect 46386 6823 47960 6824
rect 48284 6823 49517 6824
rect 46264 6734 46331 6750
rect 46264 6700 46280 6734
rect 46314 6700 46331 6734
rect 46264 6684 46331 6700
rect 45416 6612 45450 6628
rect 46095 6667 46129 6683
rect 46095 6617 46129 6633
rect 46441 6582 46475 6823
rect 47463 6806 47960 6823
rect 46911 6734 46978 6750
rect 46911 6700 46928 6734
rect 46962 6700 46978 6734
rect 46911 6684 46978 6700
rect 48162 6734 48229 6750
rect 48162 6700 48178 6734
rect 48212 6700 48229 6734
rect 48162 6684 48229 6700
rect 47218 6666 47252 6682
rect 46530 6616 46546 6650
rect 46580 6616 46596 6650
rect 46648 6617 46664 6651
rect 46698 6617 46714 6651
rect 47218 6616 47252 6632
rect 47993 6667 48027 6683
rect 47993 6617 48027 6633
rect 48339 6582 48373 6823
rect 49361 6795 49517 6823
rect 49361 6794 49461 6795
rect 48807 6735 48874 6751
rect 48807 6701 48824 6735
rect 48858 6701 48874 6735
rect 48807 6685 48874 6701
rect 49116 6666 49150 6682
rect 48428 6616 48444 6650
rect 48478 6616 48494 6650
rect 48546 6617 48562 6651
rect 48596 6617 48612 6651
rect 49116 6616 49150 6632
rect 45105 6534 45121 6568
rect 45155 6534 45171 6568
rect 45948 6566 45982 6582
rect 44987 6417 45003 6451
rect 45037 6417 45053 6451
rect 44591 6367 44625 6383
rect 44591 5975 44625 5991
rect 44709 6367 44743 6383
rect 44709 5975 44743 5991
rect 44827 6367 44861 6383
rect 44944 6367 44978 6383
rect 44944 6175 44978 6191
rect 45062 6367 45096 6383
rect 45948 6374 45982 6390
rect 46066 6566 46100 6582
rect 46066 6374 46100 6390
rect 46368 6566 46402 6582
rect 45062 6175 45096 6191
rect 46441 6566 46520 6582
rect 46441 6536 46486 6566
rect 46368 6123 46403 6190
rect 46486 6174 46520 6190
rect 46604 6566 46638 6582
rect 46604 6174 46638 6190
rect 46722 6566 46756 6582
rect 46840 6566 46874 6582
rect 47246 6566 47280 6582
rect 47246 6374 47280 6390
rect 47364 6566 47398 6582
rect 47364 6374 47398 6390
rect 47846 6566 47880 6582
rect 47846 6374 47880 6390
rect 47964 6566 47998 6582
rect 47964 6374 47998 6390
rect 48266 6566 48300 6582
rect 46722 6174 46756 6190
rect 46839 6123 46874 6190
rect 46368 6088 46874 6123
rect 48339 6566 48418 6582
rect 48339 6536 48384 6566
rect 48266 6123 48301 6190
rect 48384 6174 48418 6190
rect 48502 6566 48536 6582
rect 48502 6174 48536 6190
rect 48620 6566 48654 6582
rect 48738 6566 48772 6582
rect 49144 6566 49178 6582
rect 49144 6374 49178 6390
rect 49262 6566 49296 6582
rect 49262 6374 49296 6390
rect 48620 6174 48654 6190
rect 48737 6123 48772 6190
rect 48266 6088 48772 6123
rect 44827 5975 44861 5991
rect 45114 6041 45363 6084
rect 45114 5951 45161 6041
rect 45324 5951 45363 6041
rect 44634 5907 44650 5941
rect 44684 5907 44700 5941
rect 44752 5907 44768 5941
rect 44802 5907 44818 5941
rect 45114 5912 45363 5951
rect 46539 5881 46711 5928
rect 46539 5718 46578 5881
rect 46668 5718 46711 5881
rect 46539 5678 46711 5718
rect 50145 5478 50308 7414
rect 60566 7377 60600 7393
rect 60566 7327 60600 7343
rect 62656 7356 62723 7372
rect 53941 7309 53975 7325
rect 62656 7322 62673 7356
rect 62707 7322 62723 7356
rect 53941 7259 53975 7275
rect 56031 7288 56098 7304
rect 59529 7298 59563 7314
rect 56031 7254 56048 7288
rect 56082 7254 56098 7288
rect 52904 7230 52938 7246
rect 51403 7152 51626 7226
rect 51403 7150 51483 7152
rect 51403 7001 51482 7150
rect 51550 7003 51626 7152
rect 51549 7001 51626 7003
rect 51403 6895 51626 7001
rect 53022 7230 53056 7246
rect 52904 6838 52938 6854
rect 53021 6854 53022 6901
rect 53140 7230 53174 7246
rect 53056 6854 53057 6901
rect 51834 6786 52104 6820
rect 51008 6736 51042 6752
rect 51008 6544 51042 6560
rect 51126 6736 51160 6752
rect 51126 6544 51160 6560
rect 51244 6736 51278 6752
rect 51244 6544 51278 6560
rect 51362 6736 51396 6752
rect 51362 6544 51396 6560
rect 51480 6736 51514 6752
rect 51480 6544 51514 6560
rect 51598 6736 51632 6752
rect 51598 6544 51632 6560
rect 51716 6736 51750 6752
rect 51716 6544 51750 6560
rect 51834 6736 51868 6786
rect 51834 6544 51868 6560
rect 51952 6736 51986 6752
rect 51952 6544 51986 6560
rect 52070 6736 52104 6786
rect 53021 6796 53057 6854
rect 53258 7230 53292 7246
rect 53140 6838 53174 6854
rect 53256 6854 53258 6901
rect 53256 6796 53292 6854
rect 53376 7230 53410 7246
rect 53376 6838 53410 6854
rect 53494 7230 53528 7246
rect 53612 7230 53646 7246
rect 53528 6854 53530 6900
rect 53494 6796 53530 6854
rect 53612 6838 53646 6854
rect 54802 7230 54836 7246
rect 54920 7230 54954 7246
rect 54802 6838 54836 6854
rect 54919 6854 54920 6901
rect 55038 7230 55072 7246
rect 54954 6854 54955 6901
rect 54117 6796 54614 6814
rect 53021 6793 54614 6796
rect 53021 6759 54562 6793
rect 54596 6759 54614 6793
rect 53021 6756 54614 6759
rect 54919 6796 54955 6854
rect 55156 7230 55190 7246
rect 55038 6838 55072 6854
rect 55154 6854 55156 6901
rect 55154 6796 55190 6854
rect 55274 7230 55308 7246
rect 55274 6838 55308 6854
rect 55392 7230 55426 7246
rect 55510 7230 55544 7246
rect 56031 7238 56098 7254
rect 55426 6854 55428 6900
rect 55392 6796 55428 6854
rect 58028 7218 58251 7294
rect 58028 7069 58107 7218
rect 58174 7213 58251 7218
rect 58028 7064 58108 7069
rect 58175 7064 58251 7213
rect 58028 6963 58251 7064
rect 59647 7298 59681 7314
rect 59529 6906 59563 6922
rect 59646 6922 59647 6969
rect 59765 7298 59799 7314
rect 59681 6922 59682 6969
rect 55510 6838 55544 6854
rect 58459 6854 58729 6888
rect 56625 6827 56734 6833
rect 56101 6826 56734 6827
rect 56015 6824 56734 6826
rect 56015 6796 56632 6824
rect 54919 6756 56632 6796
rect 53040 6755 54614 6756
rect 54938 6755 56632 6756
rect 52918 6666 52985 6682
rect 52918 6632 52934 6666
rect 52968 6632 52985 6666
rect 52918 6616 52985 6632
rect 52070 6544 52104 6560
rect 52749 6599 52783 6615
rect 52749 6549 52783 6565
rect 53095 6514 53129 6755
rect 54117 6738 54614 6755
rect 53565 6666 53632 6682
rect 53565 6632 53582 6666
rect 53616 6632 53632 6666
rect 53565 6616 53632 6632
rect 54816 6666 54883 6682
rect 54816 6632 54832 6666
rect 54866 6632 54883 6666
rect 54816 6616 54883 6632
rect 53872 6598 53906 6614
rect 53184 6548 53200 6582
rect 53234 6548 53250 6582
rect 53302 6549 53318 6583
rect 53352 6549 53368 6583
rect 53872 6548 53906 6564
rect 54647 6599 54681 6615
rect 54647 6549 54681 6565
rect 54993 6514 55027 6755
rect 56015 6726 56632 6755
rect 56101 6725 56632 6726
rect 56625 6724 56632 6725
rect 56728 6724 56734 6824
rect 56625 6718 56734 6724
rect 57633 6804 57667 6820
rect 55461 6667 55528 6683
rect 55461 6633 55478 6667
rect 55512 6633 55528 6667
rect 55461 6617 55528 6633
rect 55770 6598 55804 6614
rect 57633 6612 57667 6628
rect 57751 6804 57785 6820
rect 57751 6612 57785 6628
rect 57869 6804 57903 6820
rect 57869 6612 57903 6628
rect 57987 6804 58021 6820
rect 57987 6612 58021 6628
rect 58105 6804 58139 6820
rect 58105 6612 58139 6628
rect 58223 6804 58257 6820
rect 58223 6612 58257 6628
rect 58341 6804 58375 6820
rect 58341 6612 58375 6628
rect 58459 6804 58493 6854
rect 58459 6612 58493 6628
rect 58577 6804 58611 6820
rect 58577 6612 58611 6628
rect 58695 6804 58729 6854
rect 59646 6864 59682 6922
rect 59883 7298 59917 7314
rect 59765 6906 59799 6922
rect 59881 6922 59883 6969
rect 59881 6864 59917 6922
rect 60001 7298 60035 7314
rect 60001 6906 60035 6922
rect 60119 7298 60153 7314
rect 60237 7298 60271 7314
rect 60153 6922 60155 6968
rect 60119 6864 60155 6922
rect 60237 6906 60271 6922
rect 61427 7298 61461 7314
rect 61545 7298 61579 7314
rect 61427 6906 61461 6922
rect 61544 6922 61545 6969
rect 61663 7298 61697 7314
rect 61579 6922 61580 6969
rect 60742 6864 61239 6882
rect 59646 6861 61239 6864
rect 59646 6827 61187 6861
rect 61221 6827 61239 6861
rect 59646 6824 61239 6827
rect 61544 6864 61580 6922
rect 61781 7298 61815 7314
rect 61663 6906 61697 6922
rect 61779 6922 61781 6969
rect 61779 6864 61815 6922
rect 61899 7298 61933 7314
rect 61899 6906 61933 6922
rect 62017 7298 62051 7314
rect 62135 7298 62169 7314
rect 62656 7306 62723 7322
rect 62051 6922 62053 6968
rect 62017 6864 62053 6922
rect 62135 6906 62169 6922
rect 62640 6893 62740 6894
rect 62640 6864 62796 6893
rect 61544 6824 62796 6864
rect 59665 6823 61239 6824
rect 61563 6823 62796 6824
rect 59543 6734 59610 6750
rect 59543 6700 59559 6734
rect 59593 6700 59610 6734
rect 59543 6684 59610 6700
rect 58695 6612 58729 6628
rect 59374 6667 59408 6683
rect 59374 6617 59408 6633
rect 55082 6548 55098 6582
rect 55132 6548 55148 6582
rect 55200 6549 55216 6583
rect 55250 6549 55266 6583
rect 59720 6582 59754 6823
rect 60742 6806 61239 6823
rect 60190 6734 60257 6750
rect 60190 6700 60207 6734
rect 60241 6700 60257 6734
rect 60190 6684 60257 6700
rect 61441 6734 61508 6750
rect 61441 6700 61457 6734
rect 61491 6700 61508 6734
rect 61441 6684 61508 6700
rect 60497 6666 60531 6682
rect 59809 6616 59825 6650
rect 59859 6616 59875 6650
rect 59927 6617 59943 6651
rect 59977 6617 59993 6651
rect 60497 6616 60531 6632
rect 61272 6667 61306 6683
rect 61272 6617 61306 6633
rect 61618 6582 61652 6823
rect 62640 6795 62796 6823
rect 62640 6794 62740 6795
rect 62086 6735 62153 6751
rect 62086 6701 62103 6735
rect 62137 6701 62153 6735
rect 62086 6685 62153 6701
rect 62395 6666 62429 6682
rect 61707 6616 61723 6650
rect 61757 6616 61773 6650
rect 61825 6617 61841 6651
rect 61875 6617 61891 6651
rect 62395 6616 62429 6632
rect 63710 6626 63878 6642
rect 55770 6548 55804 6564
rect 58384 6534 58400 6568
rect 58434 6534 58450 6568
rect 59227 6566 59261 6582
rect 51759 6466 51775 6500
rect 51809 6466 51825 6500
rect 52602 6498 52636 6514
rect 51641 6349 51657 6383
rect 51691 6349 51707 6383
rect 51245 6299 51279 6315
rect 51245 5907 51279 5923
rect 51363 6299 51397 6315
rect 51363 5907 51397 5923
rect 51481 6299 51515 6315
rect 51598 6299 51632 6315
rect 51598 6107 51632 6123
rect 51716 6299 51750 6315
rect 52602 6306 52636 6322
rect 52720 6498 52754 6514
rect 52720 6306 52754 6322
rect 53022 6498 53056 6514
rect 51716 6107 51750 6123
rect 53095 6498 53174 6514
rect 53095 6468 53140 6498
rect 53022 6055 53057 6122
rect 53140 6106 53174 6122
rect 53258 6498 53292 6514
rect 53258 6106 53292 6122
rect 53376 6498 53410 6514
rect 53494 6498 53528 6514
rect 53900 6498 53934 6514
rect 53900 6306 53934 6322
rect 54018 6498 54052 6514
rect 54018 6306 54052 6322
rect 54500 6498 54534 6514
rect 54500 6306 54534 6322
rect 54618 6498 54652 6514
rect 54618 6306 54652 6322
rect 54920 6498 54954 6514
rect 53376 6106 53410 6122
rect 53493 6055 53528 6122
rect 53022 6020 53528 6055
rect 54993 6498 55072 6514
rect 54993 6468 55038 6498
rect 54920 6055 54955 6122
rect 55038 6106 55072 6122
rect 55156 6498 55190 6514
rect 55156 6106 55190 6122
rect 55274 6498 55308 6514
rect 55392 6498 55426 6514
rect 55798 6498 55832 6514
rect 55798 6306 55832 6322
rect 55916 6498 55950 6514
rect 58266 6417 58282 6451
rect 58316 6417 58332 6451
rect 55916 6306 55950 6322
rect 57870 6367 57904 6383
rect 55274 6106 55308 6122
rect 55391 6055 55426 6122
rect 54920 6020 55426 6055
rect 51481 5907 51515 5923
rect 51768 5973 52017 6016
rect 57870 5975 57904 5991
rect 57988 6367 58022 6383
rect 57988 5975 58022 5991
rect 58106 6367 58140 6383
rect 58223 6367 58257 6383
rect 58223 6175 58257 6191
rect 58341 6367 58375 6383
rect 59227 6374 59261 6390
rect 59345 6566 59379 6582
rect 59345 6374 59379 6390
rect 59647 6566 59681 6582
rect 58341 6175 58375 6191
rect 59720 6566 59799 6582
rect 59720 6536 59765 6566
rect 59647 6123 59682 6190
rect 59765 6174 59799 6190
rect 59883 6566 59917 6582
rect 59883 6174 59917 6190
rect 60001 6566 60035 6582
rect 60119 6566 60153 6582
rect 60525 6566 60559 6582
rect 60525 6374 60559 6390
rect 60643 6566 60677 6582
rect 60643 6374 60677 6390
rect 61125 6566 61159 6582
rect 61125 6374 61159 6390
rect 61243 6566 61277 6582
rect 61243 6374 61277 6390
rect 61545 6566 61579 6582
rect 60001 6174 60035 6190
rect 60118 6123 60153 6190
rect 59647 6088 60153 6123
rect 61618 6566 61697 6582
rect 61618 6536 61663 6566
rect 61545 6123 61580 6190
rect 61663 6174 61697 6190
rect 61781 6566 61815 6582
rect 61781 6174 61815 6190
rect 61899 6566 61933 6582
rect 62017 6566 62051 6582
rect 62423 6566 62457 6582
rect 62423 6374 62457 6390
rect 62541 6566 62575 6582
rect 63710 6556 63726 6626
rect 63862 6556 63878 6626
rect 63710 6540 63878 6556
rect 64247 6436 64517 6470
rect 62541 6374 62575 6390
rect 63421 6386 63455 6402
rect 63421 6194 63455 6210
rect 63539 6386 63573 6402
rect 63539 6194 63573 6210
rect 63657 6386 63691 6402
rect 63657 6194 63691 6210
rect 63775 6386 63809 6402
rect 63775 6194 63809 6210
rect 63893 6386 63927 6402
rect 63893 6194 63927 6210
rect 64011 6386 64045 6402
rect 64011 6194 64045 6210
rect 64129 6386 64163 6402
rect 64129 6194 64163 6210
rect 64247 6386 64281 6436
rect 64247 6194 64281 6210
rect 64365 6386 64399 6402
rect 64365 6194 64399 6210
rect 64483 6386 64517 6436
rect 64483 6194 64517 6210
rect 61899 6174 61933 6190
rect 62016 6123 62051 6190
rect 61545 6088 62051 6123
rect 64172 6116 64188 6150
rect 64222 6116 64238 6150
rect 58106 5975 58140 5991
rect 58393 6041 58642 6084
rect 51768 5883 51815 5973
rect 51978 5883 52017 5973
rect 58393 5951 58440 6041
rect 58603 5951 58642 6041
rect 64054 5999 64070 6033
rect 64104 5999 64120 6033
rect 57913 5907 57929 5941
rect 57963 5907 57979 5941
rect 58031 5907 58047 5941
rect 58081 5907 58097 5941
rect 58393 5912 58642 5951
rect 63658 5949 63692 5965
rect 51288 5839 51304 5873
rect 51338 5839 51354 5873
rect 51406 5839 51422 5873
rect 51456 5839 51472 5873
rect 51768 5844 52017 5883
rect 59818 5881 59990 5928
rect 53193 5813 53365 5860
rect 53193 5650 53232 5813
rect 53322 5650 53365 5813
rect 59818 5718 59857 5881
rect 59947 5718 59990 5881
rect 59818 5678 59990 5718
rect 53193 5610 53365 5650
rect 63658 5557 63692 5573
rect 63776 5949 63810 5965
rect 63776 5557 63810 5573
rect 63894 5949 63928 5965
rect 64011 5949 64045 5965
rect 64011 5757 64045 5773
rect 64129 5949 64163 5965
rect 64129 5757 64163 5773
rect 63894 5557 63928 5573
rect 50145 5410 50189 5478
rect 50259 5410 50308 5478
rect 50145 5394 50308 5410
rect 56141 5503 57413 5530
rect 56141 5404 56172 5503
rect 56278 5404 57281 5503
rect 57387 5404 57413 5503
rect 63701 5489 63717 5523
rect 63751 5489 63767 5523
rect 63819 5489 63835 5523
rect 63869 5489 63885 5523
rect 56141 5377 57413 5404
rect 63934 5418 64102 5436
rect 63934 5362 63950 5418
rect 64084 5362 64102 5418
rect 63934 5346 64102 5362
rect 50163 5250 62435 5251
rect 64963 5250 65082 11047
rect 65779 11092 65813 11108
rect 65661 10700 65695 10716
rect 65778 10716 65779 10763
rect 65897 11092 65931 11108
rect 65813 10716 65814 10763
rect 65778 10658 65814 10716
rect 66015 11092 66049 11108
rect 65897 10700 65931 10716
rect 66013 10716 66015 10763
rect 66013 10658 66049 10716
rect 66133 11092 66167 11108
rect 66133 10700 66167 10716
rect 66251 11092 66285 11108
rect 66369 11092 66403 11108
rect 66285 10716 66287 10762
rect 66251 10658 66287 10716
rect 66531 10887 66601 10891
rect 66531 10796 66535 10887
rect 66597 10796 66601 10887
rect 66531 10791 66601 10796
rect 66369 10700 66403 10716
rect 66546 10658 66587 10791
rect 67264 10753 67298 10769
rect 67382 11145 67416 11161
rect 67382 10753 67416 10769
rect 67500 11145 67534 11161
rect 67617 11145 67651 11161
rect 67617 10953 67651 10969
rect 67735 11145 67769 11161
rect 67735 10953 67769 10969
rect 68537 10898 68655 15948
rect 71481 15924 71570 15948
rect 71481 15875 71495 15924
rect 71555 15875 71570 15924
rect 71481 15859 71570 15875
rect 70631 15751 70721 15785
rect 70897 15751 70913 15785
rect 70631 15549 70670 15751
rect 71195 15680 71280 15696
rect 70705 15633 70721 15667
rect 70897 15633 70987 15667
rect 70631 15515 70721 15549
rect 70897 15515 70913 15549
rect 70948 15431 70987 15633
rect 71195 15620 71212 15680
rect 71267 15620 71280 15680
rect 71195 15604 71280 15620
rect 70705 15397 70721 15431
rect 70897 15397 70987 15431
rect 70429 15310 70521 15344
rect 70897 15310 70913 15344
rect 70429 15108 70468 15310
rect 70505 15192 70521 15226
rect 70897 15192 70987 15226
rect 70429 15074 70521 15108
rect 70897 15074 70913 15108
rect 70948 14990 70987 15192
rect 70505 14956 70521 14990
rect 70897 14956 70987 14990
rect 70430 14843 70521 14877
rect 70897 14843 70913 14877
rect 70430 14641 70469 14843
rect 70948 14759 70987 14956
rect 71838 14917 71854 14951
rect 72030 14917 72046 14951
rect 71838 14799 71854 14833
rect 72030 14799 72046 14833
rect 71842 14759 72042 14799
rect 70505 14725 70521 14759
rect 70897 14725 70987 14759
rect 70233 14599 70343 14615
rect 70430 14607 70521 14641
rect 70897 14607 70913 14641
rect 70233 14403 70251 14599
rect 70327 14403 70343 14599
rect 70948 14523 70987 14725
rect 71483 14713 71568 14729
rect 71838 14725 71854 14759
rect 72230 14725 72246 14759
rect 71096 14665 71112 14699
rect 71146 14665 71162 14699
rect 71483 14653 71496 14713
rect 71551 14653 71568 14713
rect 71483 14637 71568 14653
rect 70505 14489 70521 14523
rect 70897 14489 70987 14523
rect 71198 14595 71283 14611
rect 71838 14607 71854 14641
rect 72230 14607 72246 14641
rect 71198 14535 71211 14595
rect 71266 14535 71283 14595
rect 72479 14541 72565 14557
rect 71198 14519 71283 14535
rect 71838 14489 71854 14523
rect 72230 14489 72246 14523
rect 72331 14522 72365 14538
rect 70233 14387 70343 14403
rect 70430 14371 70521 14405
rect 70897 14371 70913 14405
rect 70430 14169 70469 14371
rect 70948 14287 70987 14489
rect 72331 14472 72365 14488
rect 72479 14519 72497 14541
rect 71716 14430 71732 14464
rect 71766 14430 71782 14464
rect 72479 14461 72483 14519
rect 72479 14437 72497 14461
rect 72543 14437 72565 14541
rect 72479 14421 72565 14437
rect 71838 14371 71854 14405
rect 72230 14371 72246 14405
rect 71326 14311 71342 14345
rect 71376 14311 71392 14345
rect 70505 14253 70521 14287
rect 70897 14253 70987 14287
rect 71838 14253 71854 14287
rect 72230 14253 72246 14287
rect 70430 14135 70521 14169
rect 70897 14135 70913 14169
rect 70948 14050 70987 14253
rect 71842 14209 72042 14253
rect 71838 14175 71854 14209
rect 72030 14175 72046 14209
rect 71838 14057 71854 14091
rect 72030 14057 72046 14091
rect 70505 14016 70521 14050
rect 70897 14016 70987 14050
rect 70430 13898 70521 13932
rect 70897 13898 70913 13932
rect 70430 13696 70469 13898
rect 70948 13814 70987 14016
rect 70505 13780 70521 13814
rect 70897 13780 70987 13814
rect 70430 13662 70521 13696
rect 70897 13662 70913 13696
rect 70705 13543 70721 13577
rect 70897 13543 70990 13577
rect 70634 13425 70721 13459
rect 70897 13425 70913 13459
rect 70634 13223 70671 13425
rect 70951 13341 70990 13543
rect 70705 13307 70721 13341
rect 70897 13307 70990 13341
rect 71071 13389 71105 13405
rect 71071 13339 71105 13355
rect 70634 13189 70721 13223
rect 70897 13189 70913 13223
rect 70631 12607 70721 12641
rect 70897 12607 70913 12641
rect 70631 12405 70670 12607
rect 71195 12536 71280 12552
rect 70705 12489 70721 12523
rect 70897 12489 70987 12523
rect 70631 12371 70721 12405
rect 70897 12371 70913 12405
rect 70948 12287 70987 12489
rect 71195 12476 71212 12536
rect 71267 12476 71280 12536
rect 71195 12460 71280 12476
rect 70705 12253 70721 12287
rect 70897 12253 70987 12287
rect 70429 12166 70521 12200
rect 70897 12166 70913 12200
rect 70429 11964 70468 12166
rect 70505 12048 70521 12082
rect 70897 12048 70987 12082
rect 70429 11930 70521 11964
rect 70897 11930 70913 11964
rect 70948 11846 70987 12048
rect 70505 11812 70521 11846
rect 70897 11812 70987 11846
rect 70430 11699 70521 11733
rect 70897 11699 70913 11733
rect 70430 11497 70469 11699
rect 70948 11615 70987 11812
rect 71838 11773 71854 11807
rect 72030 11773 72046 11807
rect 71838 11655 71854 11689
rect 72030 11655 72046 11689
rect 71842 11615 72042 11655
rect 70505 11581 70521 11615
rect 70897 11581 70987 11615
rect 70233 11455 70343 11471
rect 70430 11463 70521 11497
rect 70897 11463 70913 11497
rect 70233 11259 70251 11455
rect 70327 11259 70343 11455
rect 70948 11379 70987 11581
rect 71483 11569 71568 11585
rect 71838 11581 71854 11615
rect 72230 11581 72246 11615
rect 71096 11521 71112 11555
rect 71146 11521 71162 11555
rect 71483 11509 71496 11569
rect 71551 11509 71568 11569
rect 71483 11493 71568 11509
rect 70505 11345 70521 11379
rect 70897 11345 70987 11379
rect 71198 11451 71283 11467
rect 71838 11463 71854 11497
rect 72230 11463 72246 11497
rect 71198 11391 71211 11451
rect 71266 11391 71283 11451
rect 72479 11397 72565 11413
rect 71198 11375 71283 11391
rect 71838 11345 71854 11379
rect 72230 11345 72246 11379
rect 72331 11378 72365 11394
rect 70233 11243 70343 11259
rect 70430 11227 70521 11261
rect 70897 11227 70913 11261
rect 70430 11025 70469 11227
rect 70948 11143 70987 11345
rect 72331 11328 72365 11344
rect 72479 11375 72497 11397
rect 71716 11286 71732 11320
rect 71766 11286 71782 11320
rect 72479 11317 72483 11375
rect 72479 11293 72497 11317
rect 72543 11293 72565 11397
rect 72479 11277 72565 11293
rect 71838 11227 71854 11261
rect 72230 11227 72246 11261
rect 71326 11167 71342 11201
rect 71376 11167 71392 11201
rect 70505 11109 70521 11143
rect 70897 11109 70987 11143
rect 71838 11109 71854 11143
rect 72230 11109 72246 11143
rect 70430 10991 70521 11025
rect 70897 10991 70913 11025
rect 70948 10906 70987 11109
rect 71842 11065 72042 11109
rect 71838 11031 71854 11065
rect 72030 11031 72046 11065
rect 71838 10913 71854 10947
rect 72030 10913 72046 10947
rect 68008 10890 68655 10898
rect 68008 10796 68012 10890
rect 68135 10796 68655 10890
rect 70505 10872 70521 10906
rect 70897 10872 70987 10906
rect 68008 10783 68655 10796
rect 67500 10753 67534 10769
rect 70430 10754 70521 10788
rect 70897 10754 70913 10788
rect 67307 10685 67323 10719
rect 67357 10685 67373 10719
rect 67425 10685 67441 10719
rect 67475 10685 67491 10719
rect 65778 10618 66587 10658
rect 65797 10617 66587 10618
rect 65675 10528 65742 10544
rect 65675 10494 65691 10528
rect 65725 10494 65742 10528
rect 65675 10478 65742 10494
rect 65506 10461 65540 10477
rect 65506 10411 65540 10427
rect 65852 10376 65886 10617
rect 67540 10614 67708 10632
rect 67540 10558 67556 10614
rect 67690 10558 67708 10614
rect 66322 10528 66389 10544
rect 67540 10542 67708 10558
rect 70430 10552 70469 10754
rect 70948 10670 70987 10872
rect 70505 10636 70521 10670
rect 70897 10636 70987 10670
rect 66322 10494 66339 10528
rect 66373 10494 66389 10528
rect 70430 10518 70521 10552
rect 70897 10518 70913 10552
rect 66322 10478 66389 10494
rect 66629 10460 66663 10476
rect 65941 10410 65957 10444
rect 65991 10410 66007 10444
rect 66059 10411 66075 10445
rect 66109 10411 66125 10445
rect 66629 10410 66663 10426
rect 70705 10399 70721 10433
rect 70897 10399 70990 10433
rect 65359 10360 65393 10376
rect 65359 10168 65393 10184
rect 65477 10360 65511 10376
rect 65477 10168 65511 10184
rect 65779 10360 65813 10376
rect 65852 10360 65931 10376
rect 65852 10330 65897 10360
rect 65779 9917 65814 9984
rect 65897 9968 65931 9984
rect 66015 10360 66049 10376
rect 66015 9968 66049 9984
rect 66133 10360 66167 10376
rect 66251 10360 66285 10376
rect 66657 10360 66691 10376
rect 66657 10168 66691 10184
rect 66775 10360 66809 10376
rect 66775 10168 66809 10184
rect 70634 10281 70721 10315
rect 70897 10281 70913 10315
rect 70634 10079 70671 10281
rect 70951 10197 70990 10399
rect 70705 10163 70721 10197
rect 70897 10163 70990 10197
rect 71071 10245 71105 10261
rect 71071 10195 71105 10211
rect 70634 10045 70721 10079
rect 70897 10045 70913 10079
rect 66133 9968 66167 9984
rect 66250 9917 66285 9984
rect 65779 9882 66285 9917
rect 65926 9813 66168 9825
rect 65926 9711 65973 9813
rect 66108 9711 66168 9813
rect 65926 9694 66168 9711
rect 68209 9613 71571 9700
rect 68209 9476 68338 9613
rect 71485 9578 71571 9613
rect 71485 9529 71499 9578
rect 71559 9529 71571 9578
rect 71485 9510 71571 9529
rect 65859 8232 66303 8238
rect 65859 8032 65870 8232
rect 66291 8032 66303 8232
rect 65859 8026 66303 8032
rect 66074 7747 66344 7782
rect 65720 7694 65754 7710
rect 65236 7548 65506 7583
rect 65236 7494 65270 7548
rect 65236 7302 65270 7318
rect 65354 7494 65388 7510
rect 65354 7302 65388 7318
rect 65472 7494 65506 7548
rect 65472 7302 65506 7318
rect 65590 7494 65624 7510
rect 65590 7302 65624 7318
rect 65720 7302 65754 7318
rect 65838 7694 65872 7710
rect 65838 7302 65872 7318
rect 65956 7694 65990 7710
rect 65956 7302 65990 7318
rect 66074 7694 66108 7747
rect 66074 7302 66108 7318
rect 66192 7694 66226 7710
rect 66192 7302 66226 7318
rect 66310 7694 66344 7747
rect 67318 7731 67486 7747
rect 66310 7302 66344 7318
rect 66428 7694 66462 7710
rect 67318 7661 67334 7731
rect 67470 7661 67486 7731
rect 67318 7645 67486 7661
rect 67855 7541 68125 7575
rect 66428 7302 66462 7318
rect 66557 7494 66591 7510
rect 66557 7302 66591 7318
rect 66675 7494 66709 7510
rect 66675 7302 66709 7318
rect 66793 7494 66827 7510
rect 66793 7302 66827 7318
rect 66911 7494 66945 7510
rect 66911 7302 66945 7318
rect 67029 7491 67063 7507
rect 67029 7299 67063 7315
rect 67147 7491 67181 7507
rect 67147 7299 67181 7315
rect 67265 7491 67299 7507
rect 67265 7299 67299 7315
rect 67383 7491 67417 7507
rect 67383 7299 67417 7315
rect 67501 7491 67535 7507
rect 67501 7299 67535 7315
rect 67619 7491 67653 7507
rect 67619 7299 67653 7315
rect 67737 7491 67771 7507
rect 67737 7299 67771 7315
rect 67855 7491 67889 7541
rect 67855 7299 67889 7315
rect 67973 7491 68007 7507
rect 67973 7299 68007 7315
rect 68091 7491 68125 7541
rect 68091 7299 68125 7315
rect 67780 7221 67796 7255
rect 67830 7221 67846 7255
rect 66888 7136 66922 7152
rect 67662 7104 67678 7138
rect 67712 7104 67728 7138
rect 66888 7086 66922 7102
rect 67266 7054 67300 7070
rect 65482 7017 65538 7034
rect 65482 6983 65488 7017
rect 65522 6983 65538 7017
rect 65482 6966 65538 6983
rect 65663 7001 65697 7017
rect 65781 7001 65815 7017
rect 65663 6609 65697 6625
rect 65780 6625 65781 6672
rect 65899 7001 65933 7017
rect 65815 6625 65816 6672
rect 65780 6567 65816 6625
rect 66017 7001 66051 7017
rect 65899 6609 65933 6625
rect 66015 6625 66017 6672
rect 66015 6567 66051 6625
rect 66135 7001 66169 7017
rect 66135 6609 66169 6625
rect 66253 7001 66287 7017
rect 66371 7001 66405 7017
rect 66287 6625 66289 6671
rect 66253 6567 66289 6625
rect 66533 6796 66603 6800
rect 66533 6705 66537 6796
rect 66599 6705 66603 6796
rect 66533 6700 66603 6705
rect 66371 6609 66405 6625
rect 66548 6567 66589 6700
rect 67266 6662 67300 6678
rect 67384 7054 67418 7070
rect 67384 6662 67418 6678
rect 67502 7054 67536 7070
rect 67619 7054 67653 7070
rect 67619 6862 67653 6878
rect 67737 7054 67771 7070
rect 67969 7044 68125 7050
rect 67969 6973 67984 7044
rect 68111 6973 68125 7044
rect 67969 6963 68125 6973
rect 67737 6862 67771 6878
rect 67502 6662 67536 6678
rect 67309 6594 67325 6628
rect 67359 6594 67375 6628
rect 67427 6594 67443 6628
rect 67477 6594 67493 6628
rect 65780 6527 66589 6567
rect 65799 6526 66589 6527
rect 65677 6437 65744 6453
rect 65677 6403 65693 6437
rect 65727 6403 65744 6437
rect 65677 6387 65744 6403
rect 65508 6370 65542 6386
rect 65508 6320 65542 6336
rect 65854 6285 65888 6526
rect 67542 6523 67710 6541
rect 67542 6467 67558 6523
rect 67692 6467 67710 6523
rect 66324 6437 66391 6453
rect 67542 6451 67710 6467
rect 66324 6403 66341 6437
rect 66375 6403 66391 6437
rect 66324 6387 66391 6403
rect 66631 6369 66665 6385
rect 65943 6319 65959 6353
rect 65993 6319 66009 6353
rect 66061 6320 66077 6354
rect 66111 6320 66127 6354
rect 66631 6319 66665 6335
rect 65361 6269 65395 6285
rect 65361 6077 65395 6093
rect 65479 6269 65513 6285
rect 65479 6077 65513 6093
rect 65781 6269 65815 6285
rect 65854 6269 65933 6285
rect 65854 6239 65899 6269
rect 65781 5826 65816 5893
rect 65899 5877 65933 5893
rect 66017 6269 66051 6285
rect 66017 5877 66051 5893
rect 66135 6269 66169 6285
rect 66253 6269 66287 6285
rect 66659 6269 66693 6285
rect 66659 6077 66693 6093
rect 66777 6269 66811 6285
rect 66777 6077 66811 6093
rect 66135 5877 66169 5893
rect 66252 5826 66287 5893
rect 65781 5791 66287 5826
rect 65928 5722 66170 5734
rect 65928 5620 65975 5722
rect 66110 5620 66170 5722
rect 65928 5603 66170 5620
rect 50163 5249 65082 5250
rect 47698 5248 65082 5249
rect 42943 5139 65082 5248
rect 42943 5137 53370 5139
rect 62421 5138 65082 5139
rect 42943 5136 49947 5137
rect 36898 4994 64923 4996
rect 68032 4994 68125 6963
rect 36898 4867 68125 4994
rect 48289 4865 68125 4867
rect 65859 4737 66303 4743
rect 38183 4605 38406 4680
rect 38183 4456 38259 4605
rect 38326 4604 38406 4605
rect 38183 4455 38262 4456
rect 38329 4455 38406 4604
rect 38183 4349 38406 4455
rect 40665 4660 40888 4734
rect 40665 4511 40739 4660
rect 40806 4658 40888 4660
rect 40665 4509 40744 4511
rect 40811 4509 40888 4658
rect 39998 4438 40032 4454
rect 39998 4388 40032 4404
rect 40665 4403 40888 4509
rect 41812 4658 42035 4734
rect 41812 4509 41891 4658
rect 41958 4657 42035 4658
rect 41812 4508 41895 4509
rect 41962 4508 42035 4657
rect 41128 4444 41162 4460
rect 41128 4394 41162 4410
rect 41812 4403 42035 4508
rect 44734 4603 44957 4678
rect 44734 4602 44814 4603
rect 44734 4453 44813 4602
rect 44881 4454 44957 4603
rect 44880 4453 44957 4454
rect 44734 4347 44957 4453
rect 47216 4656 47439 4732
rect 47216 4507 47295 4656
rect 47362 4507 47439 4656
rect 46549 4436 46583 4452
rect 46549 4386 46583 4402
rect 47216 4401 47439 4507
rect 48363 4656 48586 4732
rect 48363 4507 48442 4656
rect 48510 4507 48586 4656
rect 47679 4442 47713 4458
rect 47679 4392 47713 4408
rect 48363 4401 48586 4507
rect 50145 4661 50307 4677
rect 50145 4593 50188 4661
rect 50258 4593 50307 4661
rect 39998 4320 40032 4336
rect 38614 4240 38884 4274
rect 39998 4270 40032 4286
rect 41128 4324 41162 4340
rect 37788 4190 37822 4206
rect 37788 3998 37822 4014
rect 37906 4190 37940 4206
rect 37906 3998 37940 4014
rect 38024 4190 38058 4206
rect 38024 3998 38058 4014
rect 38142 4190 38176 4206
rect 38142 3998 38176 4014
rect 38260 4190 38294 4206
rect 38260 3998 38294 4014
rect 38378 4190 38412 4206
rect 38378 3998 38412 4014
rect 38496 4190 38530 4206
rect 38496 3998 38530 4014
rect 38614 4190 38648 4240
rect 38614 3998 38648 4014
rect 38732 4190 38766 4206
rect 38732 3998 38766 4014
rect 38850 4190 38884 4240
rect 38850 3998 38884 4014
rect 40113 4262 40147 4278
rect 38539 3920 38555 3954
rect 38589 3920 38605 3954
rect 40113 3870 40147 3886
rect 40231 4262 40265 4278
rect 40231 3870 40265 3886
rect 40349 4262 40383 4278
rect 40349 3870 40383 3886
rect 40467 4262 40501 4278
rect 40467 3870 40501 3886
rect 40585 4262 40619 4278
rect 40585 3870 40619 3886
rect 40703 4262 40737 4278
rect 40703 3870 40737 3886
rect 40821 4262 40855 4278
rect 41128 4274 41162 4290
rect 46549 4318 46583 4334
rect 40821 3870 40855 3886
rect 41255 4266 41289 4282
rect 41255 3874 41289 3890
rect 41373 4266 41407 4282
rect 41373 3874 41407 3890
rect 41491 4266 41525 4282
rect 41491 3874 41525 3890
rect 41609 4266 41643 4282
rect 41609 3874 41643 3890
rect 41727 4266 41761 4282
rect 41727 3874 41761 3890
rect 41845 4266 41879 4282
rect 41845 3874 41879 3890
rect 41963 4266 41997 4282
rect 45165 4238 45435 4272
rect 46549 4268 46583 4284
rect 47679 4322 47713 4338
rect 44339 4188 44373 4204
rect 44339 3996 44373 4012
rect 44457 4188 44491 4204
rect 44457 3996 44491 4012
rect 44575 4188 44609 4204
rect 44575 3996 44609 4012
rect 44693 4188 44727 4204
rect 44693 3996 44727 4012
rect 44811 4188 44845 4204
rect 44811 3996 44845 4012
rect 44929 4188 44963 4204
rect 44929 3996 44963 4012
rect 45047 4188 45081 4204
rect 45047 3996 45081 4012
rect 45165 4188 45199 4238
rect 45165 3996 45199 4012
rect 45283 4188 45317 4204
rect 45283 3996 45317 4012
rect 45401 4188 45435 4238
rect 45401 3996 45435 4012
rect 46664 4260 46698 4276
rect 45090 3918 45106 3952
rect 45140 3918 45156 3952
rect 41963 3874 41997 3890
rect 46664 3868 46698 3884
rect 46782 4260 46816 4276
rect 46782 3868 46816 3884
rect 46900 4260 46934 4276
rect 46900 3868 46934 3884
rect 47018 4260 47052 4276
rect 47018 3868 47052 3884
rect 47136 4260 47170 4276
rect 47136 3868 47170 3884
rect 47254 4260 47288 4276
rect 47254 3868 47288 3884
rect 47372 4260 47406 4276
rect 47679 4272 47713 4288
rect 47372 3868 47406 3884
rect 47806 4264 47840 4280
rect 47806 3872 47840 3888
rect 47924 4264 47958 4280
rect 47924 3872 47958 3888
rect 48042 4264 48076 4280
rect 48042 3872 48076 3888
rect 48160 4264 48194 4280
rect 48160 3872 48194 3888
rect 48278 4264 48312 4280
rect 48278 3872 48312 3888
rect 48396 4264 48430 4280
rect 48396 3872 48430 3888
rect 48514 4264 48548 4280
rect 50145 4075 50307 4593
rect 51389 4603 51612 4679
rect 51389 4600 51468 4603
rect 51389 4451 51465 4600
rect 51535 4454 51612 4603
rect 51532 4451 51612 4454
rect 53871 4660 54094 4733
rect 53871 4508 53950 4660
rect 54017 4508 54094 4660
rect 51389 4348 51612 4451
rect 53204 4437 53238 4453
rect 53204 4387 53238 4403
rect 53871 4402 54094 4508
rect 55018 4657 55241 4733
rect 55018 4508 55097 4657
rect 55166 4508 55241 4657
rect 54334 4443 54368 4459
rect 54334 4393 54368 4409
rect 55018 4402 55241 4508
rect 58011 4605 58234 4680
rect 58011 4456 58089 4605
rect 58156 4604 58234 4605
rect 58011 4455 58090 4456
rect 58157 4455 58234 4604
rect 58011 4349 58234 4455
rect 60493 4658 60716 4734
rect 60493 4653 60572 4658
rect 60493 4504 60568 4653
rect 60639 4509 60716 4658
rect 60635 4504 60716 4509
rect 59826 4438 59860 4454
rect 59826 4388 59860 4404
rect 60493 4403 60716 4504
rect 61640 4659 61863 4734
rect 61640 4510 61716 4659
rect 61783 4658 61863 4659
rect 61640 4509 61719 4510
rect 61786 4509 61863 4658
rect 63781 4706 63949 4722
rect 63781 4636 63797 4706
rect 63933 4636 63949 4706
rect 63781 4620 63949 4636
rect 60956 4444 60990 4460
rect 60956 4394 60990 4410
rect 61640 4403 61863 4509
rect 64318 4516 64588 4550
rect 65859 4537 65870 4737
rect 66291 4537 66303 4737
rect 65859 4531 66303 4537
rect 63492 4466 63526 4482
rect 53204 4319 53238 4335
rect 51820 4239 52090 4273
rect 53204 4269 53238 4285
rect 54334 4323 54368 4339
rect 50994 4189 51028 4205
rect 48514 3872 48548 3888
rect 38421 3803 38437 3837
rect 38471 3803 38487 3837
rect 44972 3801 44988 3835
rect 45022 3801 45038 3835
rect 38025 3753 38059 3769
rect 38025 3361 38059 3377
rect 38143 3753 38177 3769
rect 38143 3361 38177 3377
rect 38261 3753 38295 3769
rect 38378 3753 38412 3769
rect 38378 3561 38412 3577
rect 38496 3753 38530 3769
rect 38496 3561 38530 3577
rect 44576 3751 44610 3767
rect 40302 3530 40318 3564
rect 40352 3530 40368 3564
rect 41444 3534 41460 3568
rect 41494 3534 41510 3568
rect 40023 3479 40057 3495
rect 38261 3361 38295 3377
rect 38548 3427 38797 3470
rect 38548 3337 38595 3427
rect 38758 3337 38797 3427
rect 38068 3293 38084 3327
rect 38118 3293 38134 3327
rect 38186 3293 38202 3327
rect 38236 3293 38252 3327
rect 38548 3298 38797 3337
rect 40023 3287 40057 3303
rect 40141 3479 40175 3495
rect 40141 3287 40175 3303
rect 40259 3479 40293 3495
rect 40259 3287 40293 3303
rect 40377 3479 40411 3495
rect 40377 3287 40411 3303
rect 40542 3479 40576 3495
rect 40542 3287 40576 3303
rect 40660 3479 40694 3495
rect 40660 3287 40694 3303
rect 40778 3479 40812 3495
rect 40778 3287 40812 3303
rect 40896 3479 40930 3495
rect 40896 3287 40930 3303
rect 41165 3483 41199 3499
rect 41165 3291 41199 3307
rect 41283 3483 41317 3499
rect 41283 3291 41317 3307
rect 41401 3483 41435 3499
rect 41401 3291 41435 3307
rect 41519 3483 41553 3499
rect 41519 3291 41553 3307
rect 41684 3483 41718 3499
rect 41684 3291 41718 3307
rect 41802 3483 41836 3499
rect 41802 3291 41836 3307
rect 41920 3483 41954 3499
rect 41920 3291 41954 3307
rect 42038 3483 42072 3499
rect 44576 3359 44610 3375
rect 44694 3751 44728 3767
rect 44694 3359 44728 3375
rect 44812 3751 44846 3767
rect 44929 3751 44963 3767
rect 44929 3559 44963 3575
rect 45047 3751 45081 3767
rect 45047 3559 45081 3575
rect 46853 3528 46869 3562
rect 46903 3528 46919 3562
rect 47995 3532 48011 3566
rect 48045 3532 48061 3566
rect 46574 3477 46608 3493
rect 44812 3359 44846 3375
rect 45099 3425 45348 3468
rect 45099 3335 45146 3425
rect 45309 3335 45348 3425
rect 42038 3291 42072 3307
rect 44619 3291 44635 3325
rect 44669 3291 44685 3325
rect 44737 3291 44753 3325
rect 44787 3291 44803 3325
rect 45099 3296 45348 3335
rect 46574 3285 46608 3301
rect 46692 3477 46726 3493
rect 46692 3285 46726 3301
rect 46810 3477 46844 3493
rect 46810 3285 46844 3301
rect 46928 3477 46962 3493
rect 46928 3285 46962 3301
rect 47093 3477 47127 3493
rect 47093 3285 47127 3301
rect 47211 3477 47245 3493
rect 47211 3285 47245 3301
rect 47329 3477 47363 3493
rect 47329 3285 47363 3301
rect 47447 3477 47481 3493
rect 47447 3285 47481 3301
rect 47716 3481 47750 3497
rect 47716 3289 47750 3305
rect 47834 3481 47868 3497
rect 47834 3289 47868 3305
rect 47952 3481 47986 3497
rect 47952 3289 47986 3305
rect 48070 3481 48104 3497
rect 48070 3289 48104 3305
rect 48235 3481 48269 3497
rect 48235 3289 48269 3305
rect 48353 3481 48387 3497
rect 48353 3289 48387 3305
rect 48471 3481 48505 3497
rect 48471 3289 48505 3305
rect 48589 3481 48623 3497
rect 48589 3289 48623 3305
rect 40038 3056 40210 3103
rect 38197 2954 38420 3030
rect 38197 2805 38276 2954
rect 38343 2952 38420 2954
rect 38197 2803 38280 2805
rect 38347 2803 38420 2952
rect 40038 2893 40077 3056
rect 40167 2893 40210 3056
rect 40038 2854 40210 2893
rect 41180 3054 41352 3101
rect 41180 2891 41219 3054
rect 41309 2891 41352 3054
rect 46589 3054 46761 3101
rect 41180 2852 41352 2891
rect 44748 2959 44971 3028
rect 38197 2699 38420 2803
rect 44748 2810 44825 2959
rect 44892 2952 44971 2959
rect 44748 2803 44827 2810
rect 44894 2803 44971 2952
rect 46589 2891 46628 3054
rect 46718 2891 46761 3054
rect 46589 2852 46761 2891
rect 47731 3052 47903 3099
rect 47731 2889 47770 3052
rect 47860 2889 47903 3052
rect 47731 2885 47778 2889
rect 47845 2885 47903 2889
rect 47731 2850 47903 2885
rect 44748 2697 44971 2803
rect 38628 2590 38898 2624
rect 37802 2540 37836 2556
rect 37802 2348 37836 2364
rect 37920 2540 37954 2556
rect 37920 2348 37954 2364
rect 38038 2540 38072 2556
rect 38038 2348 38072 2364
rect 38156 2540 38190 2556
rect 38156 2348 38190 2364
rect 38274 2540 38308 2556
rect 38274 2348 38308 2364
rect 38392 2540 38426 2556
rect 38392 2348 38426 2364
rect 38510 2540 38544 2556
rect 38510 2348 38544 2364
rect 38628 2540 38662 2590
rect 38628 2348 38662 2364
rect 38746 2540 38780 2556
rect 38746 2348 38780 2364
rect 38864 2540 38898 2590
rect 38864 2348 38898 2364
rect 41908 2611 42133 2687
rect 41908 2462 41986 2611
rect 42054 2462 42133 2611
rect 45179 2588 45449 2622
rect 41908 2356 42133 2462
rect 44353 2538 44387 2554
rect 44353 2346 44387 2362
rect 44471 2538 44505 2554
rect 44471 2346 44505 2362
rect 44589 2538 44623 2554
rect 44589 2346 44623 2362
rect 44707 2538 44741 2554
rect 44707 2346 44741 2362
rect 44825 2538 44859 2554
rect 44825 2346 44859 2362
rect 44943 2538 44977 2554
rect 44943 2346 44977 2362
rect 45061 2538 45095 2554
rect 45061 2346 45095 2362
rect 45179 2538 45213 2588
rect 45179 2346 45213 2362
rect 45297 2538 45331 2554
rect 45297 2346 45331 2362
rect 45415 2538 45449 2588
rect 45415 2346 45449 2362
rect 48459 2610 48684 2685
rect 48459 2609 48542 2610
rect 48459 2460 48538 2609
rect 48609 2461 48684 2610
rect 48605 2460 48684 2461
rect 48459 2354 48684 2460
rect 38553 2270 38569 2304
rect 38603 2270 38619 2304
rect 45104 2268 45120 2302
rect 45154 2268 45170 2302
rect 38435 2153 38451 2187
rect 38485 2153 38501 2187
rect 40104 2176 40374 2211
rect 39750 2123 39784 2139
rect 38039 2103 38073 2119
rect 38039 1711 38073 1727
rect 38157 2103 38191 2119
rect 38157 1711 38191 1727
rect 38275 2103 38309 2119
rect 38392 2103 38426 2119
rect 38392 1911 38426 1927
rect 38510 2103 38544 2119
rect 38510 1911 38544 1927
rect 39266 1977 39536 2012
rect 39266 1923 39300 1977
rect 38275 1711 38309 1727
rect 38562 1777 38811 1820
rect 38562 1687 38609 1777
rect 38772 1687 38811 1777
rect 39266 1731 39300 1747
rect 39384 1923 39418 1939
rect 39384 1731 39418 1747
rect 39502 1923 39536 1977
rect 39502 1731 39536 1747
rect 39620 1923 39654 1939
rect 39620 1731 39654 1747
rect 39750 1731 39784 1747
rect 39868 2123 39902 2139
rect 39868 1731 39902 1747
rect 39986 2123 40020 2139
rect 39986 1731 40020 1747
rect 40104 2123 40138 2176
rect 40104 1731 40138 1747
rect 40222 2123 40256 2139
rect 40222 1731 40256 1747
rect 40340 2123 40374 2176
rect 42002 2176 42272 2211
rect 40340 1731 40374 1747
rect 40458 2123 40492 2139
rect 41648 2123 41682 2139
rect 41164 1977 41434 2012
rect 40458 1731 40492 1747
rect 40587 1923 40621 1939
rect 40587 1731 40621 1747
rect 40705 1923 40739 1939
rect 40705 1731 40739 1747
rect 40823 1923 40857 1939
rect 40823 1731 40857 1747
rect 40941 1923 40975 1939
rect 40941 1731 40975 1747
rect 41164 1923 41198 1977
rect 41164 1731 41198 1747
rect 41282 1923 41316 1939
rect 41282 1731 41316 1747
rect 41400 1923 41434 1977
rect 41400 1731 41434 1747
rect 41518 1923 41552 1939
rect 41518 1731 41552 1747
rect 41648 1731 41682 1747
rect 41766 2123 41800 2139
rect 41766 1731 41800 1747
rect 41884 2123 41918 2139
rect 41884 1731 41918 1747
rect 42002 2123 42036 2176
rect 42002 1731 42036 1747
rect 42120 2123 42154 2139
rect 42120 1731 42154 1747
rect 42238 2123 42272 2176
rect 44986 2151 45002 2185
rect 45036 2151 45052 2185
rect 46655 2174 46925 2209
rect 42238 1731 42272 1747
rect 42356 2123 42390 2139
rect 46301 2121 46335 2137
rect 44590 2101 44624 2117
rect 42356 1731 42390 1747
rect 42485 1923 42519 1939
rect 42485 1731 42519 1747
rect 42603 1923 42637 1939
rect 42603 1731 42637 1747
rect 42721 1923 42755 1939
rect 42721 1731 42755 1747
rect 42839 1923 42873 1939
rect 42839 1731 42873 1747
rect 44590 1709 44624 1725
rect 44708 2101 44742 2117
rect 44708 1709 44742 1725
rect 44826 2101 44860 2117
rect 44943 2101 44977 2117
rect 44943 1909 44977 1925
rect 45061 2101 45095 2117
rect 45061 1909 45095 1925
rect 45817 1975 46087 2010
rect 45817 1921 45851 1975
rect 44826 1709 44860 1725
rect 45113 1775 45362 1818
rect 38082 1643 38098 1677
rect 38132 1643 38148 1677
rect 38200 1643 38216 1677
rect 38250 1643 38266 1677
rect 38562 1648 38811 1687
rect 45113 1685 45160 1775
rect 45323 1685 45362 1775
rect 45817 1729 45851 1745
rect 45935 1921 45969 1937
rect 45935 1729 45969 1745
rect 46053 1921 46087 1975
rect 46053 1729 46087 1745
rect 46171 1921 46205 1937
rect 46171 1729 46205 1745
rect 46301 1729 46335 1745
rect 46419 2121 46453 2137
rect 46419 1729 46453 1745
rect 46537 2121 46571 2137
rect 46537 1729 46571 1745
rect 46655 2121 46689 2174
rect 46655 1729 46689 1745
rect 46773 2121 46807 2137
rect 46773 1729 46807 1745
rect 46891 2121 46925 2174
rect 48553 2174 48823 2209
rect 46891 1729 46925 1745
rect 47009 2121 47043 2137
rect 48199 2121 48233 2137
rect 47715 1975 47985 2010
rect 47009 1729 47043 1745
rect 47138 1921 47172 1937
rect 47138 1729 47172 1745
rect 47256 1921 47290 1937
rect 47256 1729 47290 1745
rect 47374 1921 47408 1937
rect 47374 1729 47408 1745
rect 47492 1921 47526 1937
rect 47492 1729 47526 1745
rect 47715 1921 47749 1975
rect 47715 1729 47749 1745
rect 47833 1921 47867 1937
rect 47833 1729 47867 1745
rect 47951 1921 47985 1975
rect 47951 1729 47985 1745
rect 48069 1921 48103 1937
rect 48069 1729 48103 1745
rect 48199 1729 48233 1745
rect 48317 2121 48351 2137
rect 48317 1729 48351 1745
rect 48435 2121 48469 2137
rect 48435 1729 48469 1745
rect 48553 2121 48587 2174
rect 48553 1729 48587 1745
rect 48671 2121 48705 2137
rect 48671 1729 48705 1745
rect 48789 2121 48823 2174
rect 48789 1729 48823 1745
rect 48907 2121 48941 2137
rect 48907 1729 48941 1745
rect 49036 1921 49070 1937
rect 49036 1729 49070 1745
rect 49154 1921 49188 1937
rect 49154 1729 49188 1745
rect 49272 1921 49306 1937
rect 49272 1729 49306 1745
rect 49390 1921 49424 1937
rect 49390 1729 49424 1745
rect 44633 1641 44649 1675
rect 44683 1641 44699 1675
rect 44751 1641 44767 1675
rect 44801 1641 44817 1675
rect 45113 1646 45362 1685
rect 40730 1509 40764 1525
rect 47281 1507 47315 1523
rect 40730 1459 40764 1475
rect 42820 1488 42887 1504
rect 42820 1454 42837 1488
rect 42871 1454 42887 1488
rect 47281 1457 47315 1473
rect 49371 1486 49438 1502
rect 39693 1430 39727 1446
rect 38192 1353 38415 1426
rect 38192 1204 38269 1353
rect 38336 1350 38415 1353
rect 38192 1201 38271 1204
rect 38338 1201 38415 1350
rect 38192 1095 38415 1201
rect 39811 1430 39845 1446
rect 39693 1038 39727 1054
rect 39810 1054 39811 1101
rect 39929 1430 39963 1446
rect 39845 1054 39846 1101
rect 38623 986 38893 1020
rect 37797 936 37831 952
rect 37797 744 37831 760
rect 37915 936 37949 952
rect 37915 744 37949 760
rect 38033 936 38067 952
rect 38033 744 38067 760
rect 38151 936 38185 952
rect 38151 744 38185 760
rect 38269 936 38303 952
rect 38269 744 38303 760
rect 38387 936 38421 952
rect 38387 744 38421 760
rect 38505 936 38539 952
rect 38505 744 38539 760
rect 38623 936 38657 986
rect 38623 744 38657 760
rect 38741 936 38775 952
rect 38741 744 38775 760
rect 38859 936 38893 986
rect 39810 996 39846 1054
rect 40047 1430 40081 1446
rect 39929 1038 39963 1054
rect 40045 1054 40047 1101
rect 40045 996 40081 1054
rect 40165 1430 40199 1446
rect 40165 1038 40199 1054
rect 40283 1430 40317 1446
rect 40401 1430 40435 1446
rect 40317 1054 40319 1100
rect 40283 996 40319 1054
rect 40401 1038 40435 1054
rect 41591 1430 41625 1446
rect 41709 1430 41743 1446
rect 41591 1038 41625 1054
rect 41708 1054 41709 1101
rect 41827 1430 41861 1446
rect 41743 1054 41744 1101
rect 40906 996 41403 1014
rect 39810 993 41403 996
rect 39810 959 41351 993
rect 41385 959 41403 993
rect 39810 956 41403 959
rect 41708 996 41744 1054
rect 41945 1430 41979 1446
rect 41827 1038 41861 1054
rect 41943 1054 41945 1101
rect 41943 996 41979 1054
rect 42063 1430 42097 1446
rect 42063 1038 42097 1054
rect 42181 1430 42215 1446
rect 42299 1430 42333 1446
rect 42820 1438 42887 1454
rect 49371 1452 49388 1486
rect 49422 1452 49438 1486
rect 42215 1054 42217 1100
rect 42181 996 42217 1054
rect 46244 1428 46278 1444
rect 44743 1348 44966 1424
rect 44743 1199 44822 1348
rect 44892 1199 44966 1348
rect 44743 1093 44966 1199
rect 42299 1038 42333 1054
rect 46362 1428 46396 1444
rect 46244 1036 46278 1052
rect 46361 1052 46362 1099
rect 46480 1428 46514 1444
rect 46396 1052 46397 1099
rect 42804 1025 42904 1026
rect 42804 996 42960 1025
rect 41708 956 42960 996
rect 39829 955 41403 956
rect 41727 955 42960 956
rect 39707 866 39774 882
rect 39707 832 39723 866
rect 39757 832 39774 866
rect 39707 816 39774 832
rect 38859 744 38893 760
rect 39538 799 39572 815
rect 39538 749 39572 765
rect 39884 714 39918 955
rect 40906 938 41403 955
rect 40354 866 40421 882
rect 40354 832 40371 866
rect 40405 832 40421 866
rect 40354 816 40421 832
rect 41605 866 41672 882
rect 41605 832 41621 866
rect 41655 832 41672 866
rect 41605 816 41672 832
rect 40661 798 40695 814
rect 39973 748 39989 782
rect 40023 748 40039 782
rect 40091 749 40107 783
rect 40141 749 40157 783
rect 40661 748 40695 764
rect 41436 799 41470 815
rect 41436 749 41470 765
rect 41782 714 41816 955
rect 42804 927 42960 955
rect 45174 984 45444 1018
rect 44348 934 44382 950
rect 42804 926 42904 927
rect 42250 867 42317 883
rect 42250 833 42267 867
rect 42301 833 42317 867
rect 42250 817 42317 833
rect 42559 798 42593 814
rect 41871 748 41887 782
rect 41921 748 41937 782
rect 41989 749 42005 783
rect 42039 749 42055 783
rect 42559 748 42593 764
rect 44348 742 44382 758
rect 44466 934 44500 950
rect 44466 742 44500 758
rect 44584 934 44618 950
rect 44584 742 44618 758
rect 44702 934 44736 950
rect 44702 742 44736 758
rect 44820 934 44854 950
rect 44820 742 44854 758
rect 44938 934 44972 950
rect 44938 742 44972 758
rect 45056 934 45090 950
rect 45056 742 45090 758
rect 45174 934 45208 984
rect 45174 742 45208 758
rect 45292 934 45326 950
rect 45292 742 45326 758
rect 45410 934 45444 984
rect 46361 994 46397 1052
rect 46598 1428 46632 1444
rect 46480 1036 46514 1052
rect 46596 1052 46598 1099
rect 46596 994 46632 1052
rect 46716 1428 46750 1444
rect 46716 1036 46750 1052
rect 46834 1428 46868 1444
rect 46952 1428 46986 1444
rect 46868 1052 46870 1098
rect 46834 994 46870 1052
rect 46952 1036 46986 1052
rect 48142 1428 48176 1444
rect 48260 1428 48294 1444
rect 48142 1036 48176 1052
rect 48259 1052 48260 1099
rect 48378 1428 48412 1444
rect 48294 1052 48295 1099
rect 47457 994 47954 1012
rect 46361 991 47954 994
rect 46361 957 47902 991
rect 47936 957 47954 991
rect 46361 954 47954 957
rect 48259 994 48295 1052
rect 48496 1428 48530 1444
rect 48378 1036 48412 1052
rect 48494 1052 48496 1099
rect 48494 994 48530 1052
rect 48614 1428 48648 1444
rect 48614 1036 48648 1052
rect 48732 1428 48766 1444
rect 48850 1428 48884 1444
rect 49371 1436 49438 1452
rect 48766 1052 48768 1098
rect 48732 994 48768 1052
rect 48850 1036 48884 1052
rect 49355 994 49662 1024
rect 48259 954 49662 994
rect 46380 953 47954 954
rect 48278 953 49662 954
rect 46258 864 46325 880
rect 46258 830 46274 864
rect 46308 830 46325 864
rect 46258 814 46325 830
rect 45410 742 45444 758
rect 46089 797 46123 813
rect 46089 747 46123 763
rect 38548 666 38564 700
rect 38598 666 38614 700
rect 39391 698 39425 714
rect 38430 549 38446 583
rect 38480 549 38496 583
rect 38034 499 38068 515
rect 38034 107 38068 123
rect 38152 499 38186 515
rect 38152 107 38186 123
rect 38270 499 38304 515
rect 38387 499 38421 515
rect 38387 307 38421 323
rect 38505 499 38539 515
rect 39391 506 39425 522
rect 39509 698 39543 714
rect 39509 506 39543 522
rect 39811 698 39845 714
rect 38505 307 38539 323
rect 39884 698 39963 714
rect 39884 668 39929 698
rect 39811 255 39846 322
rect 39929 306 39963 322
rect 40047 698 40081 714
rect 40047 306 40081 322
rect 40165 698 40199 714
rect 40283 698 40317 714
rect 40689 698 40723 714
rect 40689 506 40723 522
rect 40807 698 40841 714
rect 40807 506 40841 522
rect 41289 698 41323 714
rect 41289 506 41323 522
rect 41407 698 41441 714
rect 41407 506 41441 522
rect 41709 698 41743 714
rect 40165 306 40199 322
rect 40282 255 40317 322
rect 39811 220 40317 255
rect 41782 698 41861 714
rect 41782 668 41827 698
rect 41709 255 41744 322
rect 41827 306 41861 322
rect 41945 698 41979 714
rect 41945 306 41979 322
rect 42063 698 42097 714
rect 42181 698 42215 714
rect 42587 698 42621 714
rect 42587 506 42621 522
rect 42705 698 42739 714
rect 46435 712 46469 953
rect 47457 936 47954 953
rect 46905 864 46972 880
rect 46905 830 46922 864
rect 46956 830 46972 864
rect 46905 814 46972 830
rect 48156 864 48223 880
rect 48156 830 48172 864
rect 48206 830 48223 864
rect 48156 814 48223 830
rect 47212 796 47246 812
rect 46524 746 46540 780
rect 46574 746 46590 780
rect 46642 747 46658 781
rect 46692 747 46708 781
rect 47212 746 47246 762
rect 47987 797 48021 813
rect 47987 747 48021 763
rect 48333 712 48367 953
rect 49355 924 49662 953
rect 49427 923 49662 924
rect 48801 865 48868 881
rect 48801 831 48818 865
rect 48852 831 48868 865
rect 48801 815 48868 831
rect 49110 796 49144 812
rect 48422 746 48438 780
rect 48472 746 48488 780
rect 48540 747 48556 781
rect 48590 747 48606 781
rect 49110 746 49144 762
rect 45099 664 45115 698
rect 45149 664 45165 698
rect 45942 696 45976 712
rect 44981 547 44997 581
rect 45031 547 45047 581
rect 42705 506 42739 522
rect 42063 306 42097 322
rect 42180 255 42215 322
rect 41709 220 42215 255
rect 44585 497 44619 513
rect 38270 107 38304 123
rect 38557 173 38806 216
rect 38557 83 38604 173
rect 38767 83 38806 173
rect 44585 105 44619 121
rect 44703 497 44737 513
rect 44703 105 44737 121
rect 44821 497 44855 513
rect 44938 497 44972 513
rect 44938 305 44972 321
rect 45056 497 45090 513
rect 45942 504 45976 520
rect 46060 696 46094 712
rect 46060 504 46094 520
rect 46362 696 46396 712
rect 45056 305 45090 321
rect 46435 696 46514 712
rect 46435 666 46480 696
rect 46362 253 46397 320
rect 46480 304 46514 320
rect 46598 696 46632 712
rect 46598 304 46632 320
rect 46716 696 46750 712
rect 46834 696 46868 712
rect 47240 696 47274 712
rect 47240 504 47274 520
rect 47358 696 47392 712
rect 47358 504 47392 520
rect 47840 696 47874 712
rect 47840 504 47874 520
rect 47958 696 47992 712
rect 47958 504 47992 520
rect 48260 696 48294 712
rect 46716 304 46750 320
rect 46833 253 46868 320
rect 46362 218 46868 253
rect 48333 696 48412 712
rect 48333 666 48378 696
rect 48260 253 48295 320
rect 48378 304 48412 320
rect 48496 696 48530 712
rect 48496 304 48530 320
rect 48614 696 48648 712
rect 48732 696 48766 712
rect 49138 696 49172 712
rect 49138 504 49172 520
rect 49256 696 49290 712
rect 49256 504 49290 520
rect 48614 304 48648 320
rect 48731 253 48766 320
rect 48260 218 48766 253
rect 44821 105 44855 121
rect 45108 171 45357 214
rect 38077 39 38093 73
rect 38127 39 38143 73
rect 38195 39 38211 73
rect 38245 39 38261 73
rect 38557 44 38806 83
rect 45108 81 45155 171
rect 45318 81 45357 171
rect 39982 13 40154 60
rect 44628 37 44644 71
rect 44678 37 44694 71
rect 44746 37 44762 71
rect 44796 37 44812 71
rect 45108 42 45357 81
rect 39982 -150 40021 13
rect 40111 -150 40154 13
rect 39982 -190 40154 -150
rect 46533 11 46705 58
rect 46533 -152 46572 11
rect 46662 -152 46705 11
rect 46533 -192 46705 -152
rect 49528 -432 49662 923
rect 50142 -97 50310 4075
rect 50994 3997 51028 4013
rect 51112 4189 51146 4205
rect 51112 3997 51146 4013
rect 51230 4189 51264 4205
rect 51230 3997 51264 4013
rect 51348 4189 51382 4205
rect 51348 3997 51382 4013
rect 51466 4189 51500 4205
rect 51466 3997 51500 4013
rect 51584 4189 51618 4205
rect 51584 3997 51618 4013
rect 51702 4189 51736 4205
rect 51702 3997 51736 4013
rect 51820 4189 51854 4239
rect 51820 3997 51854 4013
rect 51938 4189 51972 4205
rect 51938 3997 51972 4013
rect 52056 4189 52090 4239
rect 52056 3997 52090 4013
rect 53319 4261 53353 4277
rect 51745 3919 51761 3953
rect 51795 3919 51811 3953
rect 53319 3869 53353 3885
rect 53437 4261 53471 4277
rect 53437 3869 53471 3885
rect 53555 4261 53589 4277
rect 53555 3869 53589 3885
rect 53673 4261 53707 4277
rect 53673 3869 53707 3885
rect 53791 4261 53825 4277
rect 53791 3869 53825 3885
rect 53909 4261 53943 4277
rect 53909 3869 53943 3885
rect 54027 4261 54061 4277
rect 54334 4273 54368 4289
rect 59826 4320 59860 4336
rect 54027 3869 54061 3885
rect 54461 4265 54495 4281
rect 54461 3873 54495 3889
rect 54579 4265 54613 4281
rect 54579 3873 54613 3889
rect 54697 4265 54731 4281
rect 54697 3873 54731 3889
rect 54815 4265 54849 4281
rect 54815 3873 54849 3889
rect 54933 4265 54967 4281
rect 54933 3873 54967 3889
rect 55051 4265 55085 4281
rect 55051 3873 55085 3889
rect 55169 4265 55203 4281
rect 58442 4240 58712 4274
rect 59826 4270 59860 4286
rect 60956 4324 60990 4340
rect 57616 4190 57650 4206
rect 57616 3998 57650 4014
rect 57734 4190 57768 4206
rect 57734 3998 57768 4014
rect 57852 4190 57886 4206
rect 57852 3998 57886 4014
rect 57970 4190 58004 4206
rect 57970 3998 58004 4014
rect 58088 4190 58122 4206
rect 58088 3998 58122 4014
rect 58206 4190 58240 4206
rect 58206 3998 58240 4014
rect 58324 4190 58358 4206
rect 58324 3998 58358 4014
rect 58442 4190 58476 4240
rect 58442 3998 58476 4014
rect 58560 4190 58594 4206
rect 58560 3998 58594 4014
rect 58678 4190 58712 4240
rect 58678 3998 58712 4014
rect 59941 4262 59975 4278
rect 58367 3920 58383 3954
rect 58417 3920 58433 3954
rect 55169 3873 55203 3889
rect 59941 3870 59975 3886
rect 60059 4262 60093 4278
rect 60059 3870 60093 3886
rect 60177 4262 60211 4278
rect 60177 3870 60211 3886
rect 60295 4262 60329 4278
rect 60295 3870 60329 3886
rect 60413 4262 60447 4278
rect 60413 3870 60447 3886
rect 60531 4262 60565 4278
rect 60531 3870 60565 3886
rect 60649 4262 60683 4278
rect 60956 4274 60990 4290
rect 60649 3870 60683 3886
rect 61083 4266 61117 4282
rect 61083 3874 61117 3890
rect 61201 4266 61235 4282
rect 61201 3874 61235 3890
rect 61319 4266 61353 4282
rect 61319 3874 61353 3890
rect 61437 4266 61471 4282
rect 61437 3874 61471 3890
rect 61555 4266 61589 4282
rect 61555 3874 61589 3890
rect 61673 4266 61707 4282
rect 61673 3874 61707 3890
rect 61791 4266 61825 4282
rect 63492 4274 63526 4290
rect 63610 4466 63644 4482
rect 63610 4274 63644 4290
rect 63728 4466 63762 4482
rect 63728 4274 63762 4290
rect 63846 4466 63880 4482
rect 63846 4274 63880 4290
rect 63964 4466 63998 4482
rect 63964 4274 63998 4290
rect 64082 4466 64116 4482
rect 64082 4274 64116 4290
rect 64200 4466 64234 4482
rect 64200 4274 64234 4290
rect 64318 4466 64352 4516
rect 64318 4274 64352 4290
rect 64436 4466 64470 4482
rect 64436 4274 64470 4290
rect 64554 4466 64588 4516
rect 64554 4274 64588 4290
rect 66074 4252 66344 4287
rect 64243 4196 64259 4230
rect 64293 4196 64309 4230
rect 65720 4199 65754 4215
rect 64125 4079 64141 4113
rect 64175 4079 64191 4113
rect 65236 4053 65506 4088
rect 61791 3874 61825 3890
rect 63729 4029 63763 4045
rect 51627 3802 51643 3836
rect 51677 3802 51693 3836
rect 58249 3803 58265 3837
rect 58299 3803 58315 3837
rect 51231 3752 51265 3768
rect 51231 3360 51265 3376
rect 51349 3752 51383 3768
rect 51349 3360 51383 3376
rect 51467 3752 51501 3768
rect 51584 3752 51618 3768
rect 51584 3560 51618 3576
rect 51702 3752 51736 3768
rect 51702 3560 51736 3576
rect 57853 3753 57887 3769
rect 53508 3529 53524 3563
rect 53558 3529 53574 3563
rect 54650 3533 54666 3567
rect 54700 3533 54716 3567
rect 53229 3478 53263 3494
rect 51467 3360 51501 3376
rect 51754 3426 52003 3469
rect 51754 3336 51801 3426
rect 51964 3336 52003 3426
rect 51274 3292 51290 3326
rect 51324 3292 51340 3326
rect 51392 3292 51408 3326
rect 51442 3292 51458 3326
rect 51754 3297 52003 3336
rect 53229 3286 53263 3302
rect 53347 3478 53381 3494
rect 53347 3286 53381 3302
rect 53465 3478 53499 3494
rect 53465 3286 53499 3302
rect 53583 3478 53617 3494
rect 53583 3286 53617 3302
rect 53748 3478 53782 3494
rect 53748 3286 53782 3302
rect 53866 3478 53900 3494
rect 53866 3286 53900 3302
rect 53984 3478 54018 3494
rect 53984 3286 54018 3302
rect 54102 3478 54136 3494
rect 54102 3286 54136 3302
rect 54371 3482 54405 3498
rect 54371 3290 54405 3306
rect 54489 3482 54523 3498
rect 54489 3290 54523 3306
rect 54607 3482 54641 3498
rect 54607 3290 54641 3306
rect 54725 3482 54759 3498
rect 54725 3290 54759 3306
rect 54890 3482 54924 3498
rect 54890 3290 54924 3306
rect 55008 3482 55042 3498
rect 55008 3290 55042 3306
rect 55126 3482 55160 3498
rect 55126 3290 55160 3306
rect 55244 3482 55278 3498
rect 57853 3361 57887 3377
rect 57971 3753 58005 3769
rect 57971 3361 58005 3377
rect 58089 3753 58123 3769
rect 58206 3753 58240 3769
rect 58206 3561 58240 3577
rect 58324 3753 58358 3769
rect 63729 3637 63763 3653
rect 63847 4029 63881 4045
rect 63847 3637 63881 3653
rect 63965 4029 63999 4045
rect 64082 4029 64116 4045
rect 64082 3837 64116 3853
rect 64200 4029 64234 4045
rect 64200 3837 64234 3853
rect 65236 3999 65270 4053
rect 65236 3807 65270 3823
rect 65354 3999 65388 4015
rect 65354 3807 65388 3823
rect 65472 3999 65506 4053
rect 65472 3807 65506 3823
rect 65590 3999 65624 4015
rect 65590 3807 65624 3823
rect 65720 3807 65754 3823
rect 65838 4199 65872 4215
rect 65838 3807 65872 3823
rect 65956 4199 65990 4215
rect 65956 3807 65990 3823
rect 66074 4199 66108 4252
rect 66074 3807 66108 3823
rect 66192 4199 66226 4215
rect 66192 3807 66226 3823
rect 66310 4199 66344 4252
rect 67318 4236 67486 4252
rect 66310 3807 66344 3823
rect 66428 4199 66462 4215
rect 67318 4166 67334 4236
rect 67470 4166 67486 4236
rect 67318 4150 67486 4166
rect 67855 4046 68125 4080
rect 66428 3807 66462 3823
rect 66557 3999 66591 4015
rect 66557 3807 66591 3823
rect 66675 3999 66709 4015
rect 66675 3807 66709 3823
rect 66793 3999 66827 4015
rect 66793 3807 66827 3823
rect 66911 3999 66945 4015
rect 66911 3807 66945 3823
rect 67029 3996 67063 4012
rect 67029 3804 67063 3820
rect 67147 3996 67181 4012
rect 67147 3804 67181 3820
rect 67265 3996 67299 4012
rect 67265 3804 67299 3820
rect 67383 3996 67417 4012
rect 67383 3804 67417 3820
rect 67501 3996 67535 4012
rect 67501 3804 67535 3820
rect 67619 3996 67653 4012
rect 67619 3804 67653 3820
rect 67737 3996 67771 4012
rect 67737 3804 67771 3820
rect 67855 3996 67889 4046
rect 67855 3804 67889 3820
rect 67973 3996 68007 4012
rect 67973 3804 68007 3820
rect 68091 3996 68125 4046
rect 68091 3804 68125 3820
rect 67780 3726 67796 3760
rect 67830 3726 67846 3760
rect 63965 3637 63999 3653
rect 66888 3641 66922 3657
rect 67662 3609 67678 3643
rect 67712 3609 67728 3643
rect 58324 3561 58358 3577
rect 63772 3569 63788 3603
rect 63822 3569 63838 3603
rect 63890 3569 63906 3603
rect 63940 3569 63956 3603
rect 66888 3591 66922 3607
rect 60130 3530 60146 3564
rect 60180 3530 60196 3564
rect 61272 3534 61288 3568
rect 61322 3534 61338 3568
rect 67266 3559 67300 3575
rect 65482 3522 65538 3539
rect 59851 3479 59885 3495
rect 58089 3361 58123 3377
rect 58376 3427 58625 3470
rect 58376 3337 58423 3427
rect 58586 3337 58625 3427
rect 55244 3290 55278 3306
rect 57896 3293 57912 3327
rect 57946 3293 57962 3327
rect 58014 3293 58030 3327
rect 58064 3293 58080 3327
rect 58376 3298 58625 3337
rect 59851 3287 59885 3303
rect 59969 3479 60003 3495
rect 59969 3287 60003 3303
rect 60087 3479 60121 3495
rect 60087 3287 60121 3303
rect 60205 3479 60239 3495
rect 60205 3287 60239 3303
rect 60370 3479 60404 3495
rect 60370 3287 60404 3303
rect 60488 3479 60522 3495
rect 60488 3287 60522 3303
rect 60606 3479 60640 3495
rect 60606 3287 60640 3303
rect 60724 3479 60758 3495
rect 60724 3287 60758 3303
rect 60993 3483 61027 3499
rect 60993 3291 61027 3307
rect 61111 3483 61145 3499
rect 61111 3291 61145 3307
rect 61229 3483 61263 3499
rect 61229 3291 61263 3307
rect 61347 3483 61381 3499
rect 61347 3291 61381 3307
rect 61512 3483 61546 3499
rect 61512 3291 61546 3307
rect 61630 3483 61664 3499
rect 61630 3291 61664 3307
rect 61748 3483 61782 3499
rect 61748 3291 61782 3307
rect 61866 3483 61900 3499
rect 64005 3498 64173 3516
rect 64005 3442 64021 3498
rect 64155 3442 64173 3498
rect 65482 3488 65488 3522
rect 65522 3488 65538 3522
rect 65482 3471 65538 3488
rect 65663 3506 65697 3522
rect 64005 3426 64173 3442
rect 61866 3291 61900 3307
rect 65781 3506 65815 3522
rect 65663 3114 65697 3130
rect 65780 3130 65781 3177
rect 65899 3506 65933 3522
rect 65815 3130 65816 3177
rect 53244 3055 53416 3102
rect 51403 2954 51626 3029
rect 51403 2953 51485 2954
rect 51403 2804 51482 2953
rect 51552 2805 51626 2954
rect 53244 2892 53283 3055
rect 53373 2892 53416 3055
rect 53244 2853 53416 2892
rect 54386 3053 54558 3100
rect 54386 2890 54425 3053
rect 54515 2890 54558 3053
rect 59866 3056 60038 3103
rect 54386 2851 54558 2890
rect 58025 2955 58248 3030
rect 51549 2804 51626 2805
rect 51403 2698 51626 2804
rect 58025 2805 58104 2955
rect 58171 2805 58248 2955
rect 59866 2893 59905 3056
rect 59995 2893 60038 3056
rect 59866 2854 60038 2893
rect 61008 3054 61180 3101
rect 61008 2891 61047 3054
rect 61137 2891 61180 3054
rect 65780 3072 65816 3130
rect 66017 3506 66051 3522
rect 65899 3114 65933 3130
rect 66015 3130 66017 3177
rect 66015 3072 66051 3130
rect 66135 3506 66169 3522
rect 66135 3114 66169 3130
rect 66253 3506 66287 3522
rect 66371 3506 66405 3522
rect 66287 3130 66289 3176
rect 66253 3072 66289 3130
rect 66533 3301 66603 3305
rect 66533 3210 66537 3301
rect 66599 3210 66603 3301
rect 66533 3205 66603 3210
rect 66371 3114 66405 3130
rect 66548 3072 66589 3205
rect 67266 3167 67300 3183
rect 67384 3559 67418 3575
rect 67384 3167 67418 3183
rect 67502 3559 67536 3575
rect 67619 3559 67653 3575
rect 67619 3367 67653 3383
rect 67737 3559 67771 3575
rect 67737 3367 67771 3383
rect 68209 3313 68339 9476
rect 70635 9405 70725 9439
rect 70901 9405 70917 9439
rect 70635 9203 70674 9405
rect 71199 9334 71284 9350
rect 70709 9287 70725 9321
rect 70901 9287 70991 9321
rect 70635 9169 70725 9203
rect 70901 9169 70917 9203
rect 70952 9085 70991 9287
rect 71199 9274 71216 9334
rect 71271 9274 71284 9334
rect 71199 9258 71284 9274
rect 70709 9051 70725 9085
rect 70901 9051 70991 9085
rect 70433 8964 70525 8998
rect 70901 8964 70917 8998
rect 70433 8762 70472 8964
rect 70509 8846 70525 8880
rect 70901 8846 70991 8880
rect 70433 8728 70525 8762
rect 70901 8728 70917 8762
rect 70952 8644 70991 8846
rect 70509 8610 70525 8644
rect 70901 8610 70991 8644
rect 70434 8497 70525 8531
rect 70901 8497 70917 8531
rect 70434 8295 70473 8497
rect 70952 8413 70991 8610
rect 71842 8571 71858 8605
rect 72034 8571 72050 8605
rect 71842 8453 71858 8487
rect 72034 8453 72050 8487
rect 71846 8413 72046 8453
rect 70509 8379 70525 8413
rect 70901 8379 70991 8413
rect 70237 8253 70347 8269
rect 70434 8261 70525 8295
rect 70901 8261 70917 8295
rect 70237 8057 70255 8253
rect 70331 8057 70347 8253
rect 70952 8177 70991 8379
rect 71487 8367 71572 8383
rect 71842 8379 71858 8413
rect 72234 8379 72250 8413
rect 71100 8319 71116 8353
rect 71150 8319 71166 8353
rect 71487 8307 71500 8367
rect 71555 8307 71572 8367
rect 71487 8291 71572 8307
rect 70509 8143 70525 8177
rect 70901 8143 70991 8177
rect 71202 8249 71287 8265
rect 71842 8261 71858 8295
rect 72234 8261 72250 8295
rect 71202 8189 71215 8249
rect 71270 8189 71287 8249
rect 72483 8195 72569 8211
rect 71202 8173 71287 8189
rect 71842 8143 71858 8177
rect 72234 8143 72250 8177
rect 72335 8176 72369 8192
rect 70237 8041 70347 8057
rect 70434 8025 70525 8059
rect 70901 8025 70917 8059
rect 70434 7823 70473 8025
rect 70952 7941 70991 8143
rect 72335 8126 72369 8142
rect 72483 8173 72501 8195
rect 71720 8084 71736 8118
rect 71770 8084 71786 8118
rect 72483 8115 72487 8173
rect 72483 8091 72501 8115
rect 72547 8091 72569 8195
rect 72483 8075 72569 8091
rect 71842 8025 71858 8059
rect 72234 8025 72250 8059
rect 71330 7965 71346 7999
rect 71380 7965 71396 7999
rect 70509 7907 70525 7941
rect 70901 7907 70991 7941
rect 71842 7907 71858 7941
rect 72234 7907 72250 7941
rect 70434 7789 70525 7823
rect 70901 7789 70917 7823
rect 70952 7704 70991 7907
rect 71846 7863 72046 7907
rect 71842 7829 71858 7863
rect 72034 7829 72050 7863
rect 71842 7711 71858 7745
rect 72034 7711 72050 7745
rect 70509 7670 70525 7704
rect 70901 7670 70991 7704
rect 70434 7552 70525 7586
rect 70901 7552 70917 7586
rect 70434 7350 70473 7552
rect 70952 7468 70991 7670
rect 70509 7434 70525 7468
rect 70901 7434 70991 7468
rect 70434 7316 70525 7350
rect 70901 7316 70917 7350
rect 70709 7197 70725 7231
rect 70901 7197 70994 7231
rect 70638 7079 70725 7113
rect 70901 7079 70917 7113
rect 70638 6877 70675 7079
rect 70955 6995 70994 7197
rect 70709 6961 70725 6995
rect 70901 6961 70994 6995
rect 71075 7043 71109 7059
rect 71075 6993 71109 7009
rect 70638 6843 70725 6877
rect 70901 6843 70917 6877
rect 70635 6261 70725 6295
rect 70901 6261 70917 6295
rect 70635 6059 70674 6261
rect 71199 6190 71284 6206
rect 70709 6143 70725 6177
rect 70901 6143 70991 6177
rect 70635 6025 70725 6059
rect 70901 6025 70917 6059
rect 70952 5941 70991 6143
rect 71199 6130 71216 6190
rect 71271 6130 71284 6190
rect 71199 6114 71284 6130
rect 70709 5907 70725 5941
rect 70901 5907 70991 5941
rect 70433 5820 70525 5854
rect 70901 5820 70917 5854
rect 70433 5618 70472 5820
rect 70509 5702 70525 5736
rect 70901 5702 70991 5736
rect 70433 5584 70525 5618
rect 70901 5584 70917 5618
rect 70952 5500 70991 5702
rect 70509 5466 70525 5500
rect 70901 5466 70991 5500
rect 70434 5353 70525 5387
rect 70901 5353 70917 5387
rect 70434 5151 70473 5353
rect 70952 5269 70991 5466
rect 71842 5427 71858 5461
rect 72034 5427 72050 5461
rect 71842 5309 71858 5343
rect 72034 5309 72050 5343
rect 71846 5269 72046 5309
rect 70509 5235 70525 5269
rect 70901 5235 70991 5269
rect 70237 5109 70347 5125
rect 70434 5117 70525 5151
rect 70901 5117 70917 5151
rect 70237 4913 70255 5109
rect 70331 4913 70347 5109
rect 70952 5033 70991 5235
rect 71487 5223 71572 5239
rect 71842 5235 71858 5269
rect 72234 5235 72250 5269
rect 71100 5175 71116 5209
rect 71150 5175 71166 5209
rect 71487 5163 71500 5223
rect 71555 5163 71572 5223
rect 71487 5147 71572 5163
rect 70509 4999 70525 5033
rect 70901 4999 70991 5033
rect 71202 5105 71287 5121
rect 71842 5117 71858 5151
rect 72234 5117 72250 5151
rect 71202 5045 71215 5105
rect 71270 5045 71287 5105
rect 72483 5051 72569 5067
rect 71202 5029 71287 5045
rect 71842 4999 71858 5033
rect 72234 4999 72250 5033
rect 72335 5032 72369 5048
rect 70237 4897 70347 4913
rect 70434 4881 70525 4915
rect 70901 4881 70917 4915
rect 70434 4679 70473 4881
rect 70952 4797 70991 4999
rect 72335 4982 72369 4998
rect 72483 5029 72501 5051
rect 71720 4940 71736 4974
rect 71770 4940 71786 4974
rect 72483 4971 72487 5029
rect 72483 4947 72501 4971
rect 72547 4947 72569 5051
rect 72483 4931 72569 4947
rect 71842 4881 71858 4915
rect 72234 4881 72250 4915
rect 71330 4821 71346 4855
rect 71380 4821 71396 4855
rect 70509 4763 70525 4797
rect 70901 4763 70991 4797
rect 71842 4763 71858 4797
rect 72234 4763 72250 4797
rect 70434 4645 70525 4679
rect 70901 4645 70917 4679
rect 70952 4560 70991 4763
rect 71846 4719 72046 4763
rect 71842 4685 71858 4719
rect 72034 4685 72050 4719
rect 71842 4567 71858 4601
rect 72034 4567 72050 4601
rect 70509 4526 70525 4560
rect 70901 4526 70991 4560
rect 70434 4408 70525 4442
rect 70901 4408 70917 4442
rect 70434 4206 70473 4408
rect 70952 4324 70991 4526
rect 70509 4290 70525 4324
rect 70901 4290 70991 4324
rect 70434 4172 70525 4206
rect 70901 4172 70917 4206
rect 70709 4053 70725 4087
rect 70901 4053 70994 4087
rect 70638 3935 70725 3969
rect 70901 3935 70917 3969
rect 70638 3733 70675 3935
rect 70955 3851 70994 4053
rect 70709 3817 70725 3851
rect 70901 3817 70994 3851
rect 71075 3899 71109 3915
rect 71075 3849 71109 3865
rect 70638 3699 70725 3733
rect 70901 3699 70917 3733
rect 68409 3399 71570 3416
rect 68409 3331 68420 3399
rect 68486 3331 71570 3399
rect 68409 3321 71570 3331
rect 68162 3288 68339 3313
rect 68162 3216 68192 3288
rect 68287 3216 68339 3288
rect 71481 3302 71570 3321
rect 71481 3253 71495 3302
rect 71555 3253 71570 3302
rect 71481 3233 71570 3253
rect 68162 3200 68339 3216
rect 67502 3167 67536 3183
rect 67309 3099 67325 3133
rect 67359 3099 67375 3133
rect 67427 3099 67443 3133
rect 67477 3099 67493 3133
rect 70631 3129 70721 3163
rect 70897 3129 70913 3163
rect 65780 3032 66589 3072
rect 65799 3031 66589 3032
rect 65677 2942 65744 2958
rect 65677 2908 65693 2942
rect 65727 2908 65744 2942
rect 65677 2892 65744 2908
rect 61008 2852 61180 2891
rect 65508 2875 65542 2891
rect 65508 2825 65542 2841
rect 58025 2699 58248 2805
rect 65854 2790 65888 3031
rect 67542 3028 67710 3046
rect 67542 2972 67558 3028
rect 67692 2972 67710 3028
rect 66324 2942 66391 2958
rect 67542 2956 67710 2972
rect 66324 2908 66341 2942
rect 66375 2908 66391 2942
rect 66324 2892 66391 2908
rect 70631 2927 70670 3129
rect 71195 3058 71280 3074
rect 70705 3011 70721 3045
rect 70897 3011 70987 3045
rect 70631 2893 70721 2927
rect 70897 2893 70913 2927
rect 66631 2874 66665 2890
rect 65943 2824 65959 2858
rect 65993 2824 66009 2858
rect 66061 2825 66077 2859
rect 66111 2825 66127 2859
rect 66631 2824 66665 2840
rect 70948 2809 70987 3011
rect 71195 2998 71212 3058
rect 71267 2998 71280 3058
rect 71195 2982 71280 2998
rect 65361 2774 65395 2790
rect 51834 2589 52104 2623
rect 51008 2539 51042 2555
rect 51008 2347 51042 2363
rect 51126 2539 51160 2555
rect 51126 2347 51160 2363
rect 51244 2539 51278 2555
rect 51244 2347 51278 2363
rect 51362 2539 51396 2555
rect 51362 2347 51396 2363
rect 51480 2539 51514 2555
rect 51480 2347 51514 2363
rect 51598 2539 51632 2555
rect 51598 2347 51632 2363
rect 51716 2539 51750 2555
rect 51716 2347 51750 2363
rect 51834 2539 51868 2589
rect 51834 2347 51868 2363
rect 51952 2539 51986 2555
rect 51952 2347 51986 2363
rect 52070 2539 52104 2589
rect 52070 2347 52104 2363
rect 55114 2612 55339 2686
rect 55114 2610 55196 2612
rect 55114 2461 55193 2610
rect 55263 2463 55339 2612
rect 58456 2590 58726 2624
rect 55260 2461 55339 2463
rect 55114 2355 55339 2461
rect 57630 2540 57664 2556
rect 57630 2348 57664 2364
rect 57748 2540 57782 2556
rect 57748 2348 57782 2364
rect 57866 2540 57900 2556
rect 57866 2348 57900 2364
rect 57984 2540 58018 2556
rect 57984 2348 58018 2364
rect 58102 2540 58136 2556
rect 58102 2348 58136 2364
rect 58220 2540 58254 2556
rect 58220 2348 58254 2364
rect 58338 2540 58372 2556
rect 58338 2348 58372 2364
rect 58456 2540 58490 2590
rect 58456 2348 58490 2364
rect 58574 2540 58608 2556
rect 58574 2348 58608 2364
rect 58692 2540 58726 2590
rect 58692 2348 58726 2364
rect 61736 2611 61961 2687
rect 61736 2462 61815 2611
rect 61882 2610 61961 2611
rect 61736 2461 61817 2462
rect 61884 2461 61961 2610
rect 65361 2582 65395 2598
rect 65479 2774 65513 2790
rect 65479 2582 65513 2598
rect 65781 2774 65815 2790
rect 61736 2356 61961 2461
rect 65854 2774 65933 2790
rect 65854 2744 65899 2774
rect 65781 2331 65816 2398
rect 65899 2382 65933 2398
rect 66017 2774 66051 2790
rect 66017 2382 66051 2398
rect 66135 2774 66169 2790
rect 66253 2774 66287 2790
rect 66659 2774 66693 2790
rect 66659 2582 66693 2598
rect 66777 2774 66811 2790
rect 70705 2775 70721 2809
rect 70897 2775 70987 2809
rect 66777 2582 66811 2598
rect 70429 2688 70521 2722
rect 70897 2688 70913 2722
rect 70429 2486 70468 2688
rect 70505 2570 70521 2604
rect 70897 2570 70987 2604
rect 70429 2452 70521 2486
rect 70897 2452 70913 2486
rect 66135 2382 66169 2398
rect 66252 2331 66287 2398
rect 70948 2368 70987 2570
rect 70505 2334 70521 2368
rect 70897 2334 70987 2368
rect 51759 2269 51775 2303
rect 51809 2269 51825 2303
rect 58381 2270 58397 2304
rect 58431 2270 58447 2304
rect 65781 2296 66287 2331
rect 65928 2227 66170 2239
rect 51641 2152 51657 2186
rect 51691 2152 51707 2186
rect 53310 2175 53580 2210
rect 52956 2122 52990 2138
rect 51245 2102 51279 2118
rect 51245 1710 51279 1726
rect 51363 2102 51397 2118
rect 51363 1710 51397 1726
rect 51481 2102 51515 2118
rect 51598 2102 51632 2118
rect 51598 1910 51632 1926
rect 51716 2102 51750 2118
rect 51716 1910 51750 1926
rect 52472 1976 52742 2011
rect 52472 1922 52506 1976
rect 51481 1710 51515 1726
rect 51768 1776 52017 1819
rect 51768 1686 51815 1776
rect 51978 1686 52017 1776
rect 52472 1730 52506 1746
rect 52590 1922 52624 1938
rect 52590 1730 52624 1746
rect 52708 1922 52742 1976
rect 52708 1730 52742 1746
rect 52826 1922 52860 1938
rect 52826 1730 52860 1746
rect 52956 1730 52990 1746
rect 53074 2122 53108 2138
rect 53074 1730 53108 1746
rect 53192 2122 53226 2138
rect 53192 1730 53226 1746
rect 53310 2122 53344 2175
rect 53310 1730 53344 1746
rect 53428 2122 53462 2138
rect 53428 1730 53462 1746
rect 53546 2122 53580 2175
rect 55208 2175 55478 2210
rect 53546 1730 53580 1746
rect 53664 2122 53698 2138
rect 54854 2122 54888 2138
rect 54370 1976 54640 2011
rect 53664 1730 53698 1746
rect 53793 1922 53827 1938
rect 53793 1730 53827 1746
rect 53911 1922 53945 1938
rect 53911 1730 53945 1746
rect 54029 1922 54063 1938
rect 54029 1730 54063 1746
rect 54147 1922 54181 1938
rect 54147 1730 54181 1746
rect 54370 1922 54404 1976
rect 54370 1730 54404 1746
rect 54488 1922 54522 1938
rect 54488 1730 54522 1746
rect 54606 1922 54640 1976
rect 54606 1730 54640 1746
rect 54724 1922 54758 1938
rect 54724 1730 54758 1746
rect 54854 1730 54888 1746
rect 54972 2122 55006 2138
rect 54972 1730 55006 1746
rect 55090 2122 55124 2138
rect 55090 1730 55124 1746
rect 55208 2122 55242 2175
rect 55208 1730 55242 1746
rect 55326 2122 55360 2138
rect 55326 1730 55360 1746
rect 55444 2122 55478 2175
rect 58263 2153 58279 2187
rect 58313 2153 58329 2187
rect 59932 2176 60202 2211
rect 55444 1730 55478 1746
rect 55562 2122 55596 2138
rect 59578 2123 59612 2139
rect 57867 2103 57901 2119
rect 55562 1730 55596 1746
rect 55691 1922 55725 1938
rect 55691 1730 55725 1746
rect 55809 1922 55843 1938
rect 55809 1730 55843 1746
rect 55927 1922 55961 1938
rect 55927 1730 55961 1746
rect 56045 1922 56079 1938
rect 56045 1730 56079 1746
rect 57867 1711 57901 1727
rect 57985 2103 58019 2119
rect 57985 1711 58019 1727
rect 58103 2103 58137 2119
rect 58220 2103 58254 2119
rect 58220 1911 58254 1927
rect 58338 2103 58372 2119
rect 58338 1911 58372 1927
rect 59094 1977 59364 2012
rect 59094 1923 59128 1977
rect 58103 1711 58137 1727
rect 58390 1777 58639 1820
rect 51288 1642 51304 1676
rect 51338 1642 51354 1676
rect 51406 1642 51422 1676
rect 51456 1642 51472 1676
rect 51768 1647 52017 1686
rect 58390 1687 58437 1777
rect 58600 1687 58639 1777
rect 59094 1731 59128 1747
rect 59212 1923 59246 1939
rect 59212 1731 59246 1747
rect 59330 1923 59364 1977
rect 59330 1731 59364 1747
rect 59448 1923 59482 1939
rect 59448 1731 59482 1747
rect 59578 1731 59612 1747
rect 59696 2123 59730 2139
rect 59696 1731 59730 1747
rect 59814 2123 59848 2139
rect 59814 1731 59848 1747
rect 59932 2123 59966 2176
rect 59932 1731 59966 1747
rect 60050 2123 60084 2139
rect 60050 1731 60084 1747
rect 60168 2123 60202 2176
rect 61830 2176 62100 2211
rect 60168 1731 60202 1747
rect 60286 2123 60320 2139
rect 61476 2123 61510 2139
rect 60992 1977 61262 2012
rect 60286 1731 60320 1747
rect 60415 1923 60449 1939
rect 60415 1731 60449 1747
rect 60533 1923 60567 1939
rect 60533 1731 60567 1747
rect 60651 1923 60685 1939
rect 60651 1731 60685 1747
rect 60769 1923 60803 1939
rect 60769 1731 60803 1747
rect 60992 1923 61026 1977
rect 60992 1731 61026 1747
rect 61110 1923 61144 1939
rect 61110 1731 61144 1747
rect 61228 1923 61262 1977
rect 61228 1731 61262 1747
rect 61346 1923 61380 1939
rect 61346 1731 61380 1747
rect 61476 1731 61510 1747
rect 61594 2123 61628 2139
rect 61594 1731 61628 1747
rect 61712 2123 61746 2139
rect 61712 1731 61746 1747
rect 61830 2123 61864 2176
rect 61830 1731 61864 1747
rect 61948 2123 61982 2139
rect 61948 1731 61982 1747
rect 62066 2123 62100 2176
rect 62066 1731 62100 1747
rect 62184 2123 62218 2139
rect 65928 2125 65975 2227
rect 66110 2125 66170 2227
rect 65928 2108 66170 2125
rect 70430 2221 70521 2255
rect 70897 2221 70913 2255
rect 70430 2019 70469 2221
rect 70948 2137 70987 2334
rect 71838 2295 71854 2329
rect 72030 2295 72046 2329
rect 71838 2177 71854 2211
rect 72030 2177 72046 2211
rect 71842 2137 72042 2177
rect 70505 2103 70521 2137
rect 70897 2103 70987 2137
rect 70233 1977 70343 1993
rect 70430 1985 70521 2019
rect 70897 1985 70913 2019
rect 62184 1731 62218 1747
rect 62313 1923 62347 1939
rect 62313 1731 62347 1747
rect 62431 1923 62465 1939
rect 62431 1731 62465 1747
rect 62549 1923 62583 1939
rect 62549 1731 62583 1747
rect 62667 1923 62701 1939
rect 70233 1781 70251 1977
rect 70327 1781 70343 1977
rect 70948 1901 70987 2103
rect 71483 2091 71568 2107
rect 71838 2103 71854 2137
rect 72230 2103 72246 2137
rect 71096 2043 71112 2077
rect 71146 2043 71162 2077
rect 71483 2031 71496 2091
rect 71551 2031 71568 2091
rect 71483 2015 71568 2031
rect 70505 1867 70521 1901
rect 70897 1867 70987 1901
rect 71198 1973 71283 1989
rect 71838 1985 71854 2019
rect 72230 1985 72246 2019
rect 71198 1913 71211 1973
rect 71266 1913 71283 1973
rect 72479 1919 72565 1935
rect 71198 1897 71283 1913
rect 71838 1867 71854 1901
rect 72230 1867 72246 1901
rect 72331 1900 72365 1916
rect 70233 1765 70343 1781
rect 62667 1731 62701 1747
rect 70430 1749 70521 1783
rect 70897 1749 70913 1783
rect 57910 1643 57926 1677
rect 57960 1643 57976 1677
rect 58028 1643 58044 1677
rect 58078 1643 58094 1677
rect 58390 1648 58639 1687
rect 63778 1636 63946 1652
rect 63778 1566 63794 1636
rect 63930 1566 63946 1636
rect 63778 1550 63946 1566
rect 70430 1547 70469 1749
rect 70948 1665 70987 1867
rect 72331 1850 72365 1866
rect 72479 1897 72497 1919
rect 71716 1808 71732 1842
rect 71766 1808 71782 1842
rect 72479 1839 72483 1897
rect 72479 1815 72497 1839
rect 72543 1815 72565 1919
rect 72479 1799 72565 1815
rect 71838 1749 71854 1783
rect 72230 1749 72246 1783
rect 71326 1689 71342 1723
rect 71376 1689 71392 1723
rect 70505 1631 70521 1665
rect 70897 1631 70987 1665
rect 71838 1631 71854 1665
rect 72230 1631 72246 1665
rect 53936 1508 53970 1524
rect 60558 1509 60592 1525
rect 70430 1513 70521 1547
rect 70897 1513 70913 1547
rect 53936 1458 53970 1474
rect 56026 1487 56093 1503
rect 56026 1453 56043 1487
rect 56077 1453 56093 1487
rect 60558 1459 60592 1475
rect 62648 1488 62715 1504
rect 52899 1429 52933 1445
rect 51398 1349 51621 1425
rect 51398 1200 51477 1349
rect 51544 1346 51621 1349
rect 51398 1197 51480 1200
rect 51547 1197 51621 1346
rect 51398 1094 51621 1197
rect 53017 1429 53051 1445
rect 52899 1037 52933 1053
rect 53016 1053 53017 1100
rect 53135 1429 53169 1445
rect 53051 1053 53052 1100
rect 51829 985 52099 1019
rect 51003 935 51037 951
rect 51003 743 51037 759
rect 51121 935 51155 951
rect 51121 743 51155 759
rect 51239 935 51273 951
rect 51239 743 51273 759
rect 51357 935 51391 951
rect 51357 743 51391 759
rect 51475 935 51509 951
rect 51475 743 51509 759
rect 51593 935 51627 951
rect 51593 743 51627 759
rect 51711 935 51745 951
rect 51711 743 51745 759
rect 51829 935 51863 985
rect 51829 743 51863 759
rect 51947 935 51981 951
rect 51947 743 51981 759
rect 52065 935 52099 985
rect 53016 995 53052 1053
rect 53253 1429 53287 1445
rect 53135 1037 53169 1053
rect 53251 1053 53253 1100
rect 53251 995 53287 1053
rect 53371 1429 53405 1445
rect 53371 1037 53405 1053
rect 53489 1429 53523 1445
rect 53607 1429 53641 1445
rect 53523 1053 53525 1099
rect 53489 995 53525 1053
rect 53607 1037 53641 1053
rect 54797 1429 54831 1445
rect 54915 1429 54949 1445
rect 54797 1037 54831 1053
rect 54914 1053 54915 1100
rect 55033 1429 55067 1445
rect 54949 1053 54950 1100
rect 54112 995 54609 1013
rect 53016 992 54609 995
rect 53016 958 54557 992
rect 54591 958 54609 992
rect 53016 955 54609 958
rect 54914 995 54950 1053
rect 55151 1429 55185 1445
rect 55033 1037 55067 1053
rect 55149 1053 55151 1100
rect 55149 995 55185 1053
rect 55269 1429 55303 1445
rect 55269 1037 55303 1053
rect 55387 1429 55421 1445
rect 55505 1429 55539 1445
rect 56026 1437 56093 1453
rect 62648 1454 62665 1488
rect 62699 1454 62715 1488
rect 55421 1053 55423 1099
rect 55387 995 55423 1053
rect 59521 1430 59555 1446
rect 58020 1350 58243 1426
rect 58020 1201 58099 1350
rect 58166 1346 58243 1350
rect 58020 1197 58101 1201
rect 58168 1197 58243 1346
rect 58020 1095 58243 1197
rect 55505 1037 55539 1053
rect 59639 1430 59673 1446
rect 59521 1038 59555 1054
rect 59638 1054 59639 1101
rect 59757 1430 59791 1446
rect 59673 1054 59674 1101
rect 56010 1024 56110 1025
rect 56010 995 56166 1024
rect 54914 955 56166 995
rect 53035 954 54609 955
rect 54933 954 56166 955
rect 52913 865 52980 881
rect 52913 831 52929 865
rect 52963 831 52980 865
rect 52913 815 52980 831
rect 52065 743 52099 759
rect 52744 798 52778 814
rect 52744 748 52778 764
rect 53090 713 53124 954
rect 54112 937 54609 954
rect 53560 865 53627 881
rect 53560 831 53577 865
rect 53611 831 53627 865
rect 53560 815 53627 831
rect 54811 865 54878 881
rect 54811 831 54827 865
rect 54861 831 54878 865
rect 54811 815 54878 831
rect 53867 797 53901 813
rect 53179 747 53195 781
rect 53229 747 53245 781
rect 53297 748 53313 782
rect 53347 748 53363 782
rect 53867 747 53901 763
rect 54642 798 54676 814
rect 54642 748 54676 764
rect 54988 713 55022 954
rect 56010 926 56166 954
rect 58451 986 58721 1020
rect 57625 936 57659 952
rect 56010 925 56110 926
rect 55456 866 55523 882
rect 55456 832 55473 866
rect 55507 832 55523 866
rect 55456 816 55523 832
rect 55765 797 55799 813
rect 55077 747 55093 781
rect 55127 747 55143 781
rect 55195 748 55211 782
rect 55245 748 55261 782
rect 55765 747 55799 763
rect 57625 744 57659 760
rect 57743 936 57777 952
rect 57743 744 57777 760
rect 57861 936 57895 952
rect 57861 744 57895 760
rect 57979 936 58013 952
rect 57979 744 58013 760
rect 58097 936 58131 952
rect 58097 744 58131 760
rect 58215 936 58249 952
rect 58215 744 58249 760
rect 58333 936 58367 952
rect 58333 744 58367 760
rect 58451 936 58485 986
rect 58451 744 58485 760
rect 58569 936 58603 952
rect 58569 744 58603 760
rect 58687 936 58721 986
rect 59638 996 59674 1054
rect 59875 1430 59909 1446
rect 59757 1038 59791 1054
rect 59873 1054 59875 1101
rect 59873 996 59909 1054
rect 59993 1430 60027 1446
rect 59993 1038 60027 1054
rect 60111 1430 60145 1446
rect 60229 1430 60263 1446
rect 60145 1054 60147 1100
rect 60111 996 60147 1054
rect 60229 1038 60263 1054
rect 61419 1430 61453 1446
rect 61537 1430 61571 1446
rect 61419 1038 61453 1054
rect 61536 1054 61537 1101
rect 61655 1430 61689 1446
rect 61571 1054 61572 1101
rect 60734 996 61231 1014
rect 59638 993 61231 996
rect 59638 959 61179 993
rect 61213 959 61231 993
rect 59638 956 61231 959
rect 61536 996 61572 1054
rect 61773 1430 61807 1446
rect 61655 1038 61689 1054
rect 61771 1054 61773 1101
rect 61771 996 61807 1054
rect 61891 1430 61925 1446
rect 61891 1038 61925 1054
rect 62009 1430 62043 1446
rect 62127 1430 62161 1446
rect 62648 1438 62715 1454
rect 64315 1446 64585 1480
rect 62043 1054 62045 1100
rect 62009 996 62045 1054
rect 63489 1396 63523 1412
rect 63489 1204 63523 1220
rect 63607 1396 63641 1412
rect 63607 1204 63641 1220
rect 63725 1396 63759 1412
rect 63725 1204 63759 1220
rect 63843 1396 63877 1412
rect 63843 1204 63877 1220
rect 63961 1396 63995 1412
rect 63961 1204 63995 1220
rect 64079 1396 64113 1412
rect 64079 1204 64113 1220
rect 64197 1396 64231 1412
rect 64197 1204 64231 1220
rect 64315 1396 64349 1446
rect 64315 1204 64349 1220
rect 64433 1396 64467 1412
rect 64433 1204 64467 1220
rect 64551 1396 64585 1446
rect 70948 1428 70987 1631
rect 71842 1587 72042 1631
rect 71838 1553 71854 1587
rect 72030 1553 72046 1587
rect 71838 1435 71854 1469
rect 72030 1435 72046 1469
rect 70505 1394 70521 1428
rect 70897 1394 70987 1428
rect 64551 1204 64585 1220
rect 70430 1276 70521 1310
rect 70897 1276 70913 1310
rect 64240 1126 64256 1160
rect 64290 1126 64306 1160
rect 62127 1038 62161 1054
rect 70430 1074 70469 1276
rect 70948 1192 70987 1394
rect 70505 1158 70521 1192
rect 70897 1158 70987 1192
rect 62632 1025 62732 1026
rect 62632 996 62788 1025
rect 61536 956 62788 996
rect 59657 955 61231 956
rect 61555 955 62788 956
rect 59535 866 59602 882
rect 59535 832 59551 866
rect 59585 832 59602 866
rect 59535 816 59602 832
rect 58687 744 58721 760
rect 59366 799 59400 815
rect 59366 749 59400 765
rect 59712 714 59746 955
rect 60734 938 61231 955
rect 60182 866 60249 882
rect 60182 832 60199 866
rect 60233 832 60249 866
rect 60182 816 60249 832
rect 61433 866 61500 882
rect 61433 832 61449 866
rect 61483 832 61500 866
rect 61433 816 61500 832
rect 60489 798 60523 814
rect 59801 748 59817 782
rect 59851 748 59867 782
rect 59919 749 59935 783
rect 59969 749 59985 783
rect 60489 748 60523 764
rect 61264 799 61298 815
rect 61264 749 61298 765
rect 61610 714 61644 955
rect 62632 927 62788 955
rect 64122 1009 64138 1043
rect 64172 1009 64188 1043
rect 70430 1040 70521 1074
rect 70897 1040 70913 1074
rect 63726 959 63760 975
rect 62632 926 62732 927
rect 62078 867 62145 883
rect 62078 833 62095 867
rect 62129 833 62145 867
rect 62078 817 62145 833
rect 62387 798 62421 814
rect 61699 748 61715 782
rect 61749 748 61765 782
rect 61817 749 61833 783
rect 61867 749 61883 783
rect 62387 748 62421 764
rect 51754 665 51770 699
rect 51804 665 51820 699
rect 52597 697 52631 713
rect 51636 548 51652 582
rect 51686 548 51702 582
rect 51240 498 51274 514
rect 51240 106 51274 122
rect 51358 498 51392 514
rect 51358 106 51392 122
rect 51476 498 51510 514
rect 51593 498 51627 514
rect 51593 306 51627 322
rect 51711 498 51745 514
rect 52597 505 52631 521
rect 52715 697 52749 713
rect 52715 505 52749 521
rect 53017 697 53051 713
rect 51711 306 51745 322
rect 53090 697 53169 713
rect 53090 667 53135 697
rect 53017 254 53052 321
rect 53135 305 53169 321
rect 53253 697 53287 713
rect 53253 305 53287 321
rect 53371 697 53405 713
rect 53489 697 53523 713
rect 53895 697 53929 713
rect 53895 505 53929 521
rect 54013 697 54047 713
rect 54013 505 54047 521
rect 54495 697 54529 713
rect 54495 505 54529 521
rect 54613 697 54647 713
rect 54613 505 54647 521
rect 54915 697 54949 713
rect 53371 305 53405 321
rect 53488 254 53523 321
rect 53017 219 53523 254
rect 54988 697 55067 713
rect 54988 667 55033 697
rect 54915 254 54950 321
rect 55033 305 55067 321
rect 55151 697 55185 713
rect 55151 305 55185 321
rect 55269 697 55303 713
rect 55387 697 55421 713
rect 55793 697 55827 713
rect 55793 505 55827 521
rect 55911 697 55945 713
rect 58376 666 58392 700
rect 58426 666 58442 700
rect 59219 698 59253 714
rect 58258 549 58274 583
rect 58308 549 58324 583
rect 55911 505 55945 521
rect 55269 305 55303 321
rect 55386 254 55421 321
rect 54915 219 55421 254
rect 57862 499 57896 515
rect 51476 106 51510 122
rect 51763 172 52012 215
rect 51763 82 51810 172
rect 51973 152 52012 172
rect 51976 85 52012 152
rect 57862 107 57896 123
rect 57980 499 58014 515
rect 57980 107 58014 123
rect 58098 499 58132 515
rect 58215 499 58249 515
rect 58215 307 58249 323
rect 58333 499 58367 515
rect 59219 506 59253 522
rect 59337 698 59371 714
rect 59337 506 59371 522
rect 59639 698 59673 714
rect 58333 307 58367 323
rect 59712 698 59791 714
rect 59712 668 59757 698
rect 59639 255 59674 322
rect 59757 306 59791 322
rect 59875 698 59909 714
rect 59875 306 59909 322
rect 59993 698 60027 714
rect 60111 698 60145 714
rect 60517 698 60551 714
rect 60517 506 60551 522
rect 60635 698 60669 714
rect 60635 506 60669 522
rect 61117 698 61151 714
rect 61117 506 61151 522
rect 61235 698 61269 714
rect 61235 506 61269 522
rect 61537 698 61571 714
rect 59993 306 60027 322
rect 60110 255 60145 322
rect 59639 220 60145 255
rect 61610 698 61689 714
rect 61610 668 61655 698
rect 61537 255 61572 322
rect 61655 306 61689 322
rect 61773 698 61807 714
rect 61773 306 61807 322
rect 61891 698 61925 714
rect 62009 698 62043 714
rect 62415 698 62449 714
rect 62415 506 62449 522
rect 62533 698 62567 714
rect 63726 567 63760 583
rect 63844 959 63878 975
rect 63844 567 63878 583
rect 63962 959 63996 975
rect 64079 959 64113 975
rect 64079 767 64113 783
rect 64197 959 64231 975
rect 70705 921 70721 955
rect 70897 921 70990 955
rect 64197 767 64231 783
rect 70634 803 70721 837
rect 70897 803 70913 837
rect 63962 567 63996 583
rect 70634 601 70671 803
rect 70951 719 70990 921
rect 70705 685 70721 719
rect 70897 685 70990 719
rect 71071 767 71105 783
rect 71071 717 71105 733
rect 70634 567 70721 601
rect 70897 567 70913 601
rect 62533 506 62567 522
rect 63769 499 63785 533
rect 63819 499 63835 533
rect 63887 499 63903 533
rect 63937 499 63953 533
rect 64002 428 64170 446
rect 64002 372 64018 428
rect 64152 372 64170 428
rect 64002 356 64170 372
rect 65859 389 66303 395
rect 61891 306 61925 322
rect 62008 255 62043 322
rect 61537 220 62043 255
rect 58098 107 58132 123
rect 58385 173 58634 216
rect 65859 189 65870 389
rect 66291 189 66303 389
rect 65859 183 66303 189
rect 68537 262 68655 274
rect 68537 254 71567 262
rect 68537 188 68555 254
rect 68648 210 71567 254
rect 68648 188 71568 210
rect 68537 181 71568 188
rect 51973 82 52012 85
rect 51283 38 51299 72
rect 51333 38 51349 72
rect 51401 38 51417 72
rect 51451 38 51467 72
rect 51763 43 52012 82
rect 58385 83 58432 173
rect 58595 83 58634 173
rect 50142 -165 50188 -97
rect 50258 -165 50310 -97
rect 50142 -178 50310 -165
rect 53188 12 53360 59
rect 57905 39 57921 73
rect 57955 39 57971 73
rect 58023 39 58039 73
rect 58073 39 58089 73
rect 58385 44 58634 83
rect 71482 158 71568 181
rect 71482 109 71495 158
rect 71555 109 71568 158
rect 71482 78 71568 109
rect 53188 -151 53227 12
rect 53317 -151 53360 12
rect 53188 -191 53360 -151
rect 59810 13 59982 60
rect 59810 -150 59849 13
rect 59939 -150 59982 13
rect 70631 -15 70721 19
rect 70897 -15 70913 19
rect 66074 -96 66344 -61
rect 59810 -190 59982 -150
rect 65720 -149 65754 -133
rect 65236 -295 65506 -260
rect 65236 -349 65270 -295
rect 49528 -584 64874 -432
rect 65236 -541 65270 -525
rect 65354 -349 65388 -333
rect 65354 -541 65388 -525
rect 65472 -349 65506 -295
rect 65472 -541 65506 -525
rect 65590 -349 65624 -333
rect 65590 -541 65624 -525
rect 65720 -541 65754 -525
rect 65838 -149 65872 -133
rect 65838 -541 65872 -525
rect 65956 -149 65990 -133
rect 65956 -541 65990 -525
rect 66074 -149 66108 -96
rect 66074 -541 66108 -525
rect 66192 -149 66226 -133
rect 66192 -541 66226 -525
rect 66310 -149 66344 -96
rect 67318 -112 67486 -96
rect 66310 -541 66344 -525
rect 66428 -149 66462 -133
rect 67318 -182 67334 -112
rect 67470 -182 67486 -112
rect 67318 -198 67486 -182
rect 70631 -217 70670 -15
rect 71195 -86 71280 -70
rect 70705 -133 70721 -99
rect 70897 -133 70987 -99
rect 70631 -251 70721 -217
rect 70897 -251 70913 -217
rect 67855 -302 68125 -268
rect 66428 -541 66462 -525
rect 66557 -349 66591 -333
rect 66557 -541 66591 -525
rect 66675 -349 66709 -333
rect 66675 -541 66709 -525
rect 66793 -349 66827 -333
rect 66793 -541 66827 -525
rect 66911 -349 66945 -333
rect 66911 -541 66945 -525
rect 67029 -352 67063 -336
rect 67029 -544 67063 -528
rect 67147 -352 67181 -336
rect 67147 -544 67181 -528
rect 67265 -352 67299 -336
rect 67265 -544 67299 -528
rect 67383 -352 67417 -336
rect 67383 -544 67417 -528
rect 67501 -352 67535 -336
rect 67501 -544 67535 -528
rect 67619 -352 67653 -336
rect 67619 -544 67653 -528
rect 67737 -352 67771 -336
rect 67737 -544 67771 -528
rect 67855 -352 67889 -302
rect 67855 -544 67889 -528
rect 67973 -352 68007 -336
rect 67973 -544 68007 -528
rect 68091 -352 68125 -302
rect 70948 -335 70987 -133
rect 71195 -146 71212 -86
rect 71267 -146 71280 -86
rect 71195 -162 71280 -146
rect 70705 -369 70721 -335
rect 70897 -369 70987 -335
rect 68091 -544 68125 -528
rect 70429 -456 70521 -422
rect 70897 -456 70913 -422
rect 64782 -681 64874 -584
rect 67780 -622 67796 -588
rect 67830 -622 67846 -588
rect 70429 -658 70468 -456
rect 70505 -574 70521 -540
rect 70897 -574 70987 -540
rect 64782 -687 65302 -681
rect 42118 -719 42286 -703
rect 42118 -775 42134 -719
rect 42268 -775 42286 -719
rect 42118 -793 42286 -775
rect 48672 -714 48840 -698
rect 48672 -770 48688 -714
rect 48822 -770 48840 -714
rect 48672 -788 48840 -770
rect 55321 -726 55489 -710
rect 55321 -782 55337 -726
rect 55471 -782 55489 -726
rect 64782 -757 65216 -687
rect 64783 -758 65216 -757
rect 65289 -758 65302 -687
rect 66888 -707 66922 -691
rect 70429 -692 70521 -658
rect 70897 -692 70913 -658
rect 67662 -739 67678 -705
rect 67712 -739 67728 -705
rect 66888 -757 66922 -741
rect 64783 -765 65302 -758
rect 55321 -800 55489 -782
rect 67266 -789 67300 -773
rect 65482 -826 65538 -809
rect 41885 -880 41901 -846
rect 41935 -880 41951 -846
rect 42003 -880 42019 -846
rect 42053 -880 42069 -846
rect 48439 -875 48455 -841
rect 48489 -875 48505 -841
rect 48557 -875 48573 -841
rect 48607 -875 48623 -841
rect 55088 -887 55104 -853
rect 55138 -887 55154 -853
rect 55206 -887 55222 -853
rect 55256 -887 55272 -853
rect 65482 -860 65488 -826
rect 65522 -860 65538 -826
rect 65482 -877 65538 -860
rect 65663 -842 65697 -826
rect 41842 -930 41876 -914
rect 41842 -1322 41876 -1306
rect 41960 -930 41994 -914
rect 41960 -1322 41994 -1306
rect 42078 -930 42112 -914
rect 48396 -925 48430 -909
rect 42078 -1322 42112 -1306
rect 42195 -1130 42229 -1114
rect 42195 -1322 42229 -1306
rect 42313 -1130 42347 -1114
rect 42313 -1322 42347 -1306
rect 48396 -1317 48430 -1301
rect 48514 -925 48548 -909
rect 48514 -1317 48548 -1301
rect 48632 -925 48666 -909
rect 55045 -937 55079 -921
rect 48632 -1317 48666 -1301
rect 48749 -1125 48783 -1109
rect 48749 -1317 48783 -1301
rect 48867 -1125 48901 -1109
rect 48867 -1317 48901 -1301
rect 55045 -1329 55079 -1313
rect 55163 -937 55197 -921
rect 55163 -1329 55197 -1313
rect 55281 -937 55315 -921
rect 55281 -1329 55315 -1313
rect 55398 -1137 55432 -1121
rect 55398 -1329 55432 -1313
rect 55516 -1137 55550 -1121
rect 63785 -1209 63953 -1193
rect 63785 -1279 63801 -1209
rect 63937 -1279 63953 -1209
rect 65781 -842 65815 -826
rect 65663 -1234 65697 -1218
rect 65780 -1218 65781 -1171
rect 65899 -842 65933 -826
rect 65815 -1218 65816 -1171
rect 63785 -1295 63953 -1279
rect 65780 -1276 65816 -1218
rect 66017 -842 66051 -826
rect 65899 -1234 65933 -1218
rect 66015 -1218 66017 -1171
rect 66015 -1276 66051 -1218
rect 66135 -842 66169 -826
rect 66135 -1234 66169 -1218
rect 66253 -842 66287 -826
rect 66371 -842 66405 -826
rect 66287 -1218 66289 -1172
rect 66253 -1276 66289 -1218
rect 66533 -1047 66603 -1043
rect 66533 -1138 66537 -1047
rect 66599 -1138 66603 -1047
rect 66533 -1143 66603 -1138
rect 66371 -1234 66405 -1218
rect 66548 -1276 66589 -1143
rect 67266 -1181 67300 -1165
rect 67384 -789 67418 -773
rect 67384 -1181 67418 -1165
rect 67502 -789 67536 -773
rect 67619 -789 67653 -773
rect 67619 -981 67653 -965
rect 67737 -789 67771 -773
rect 70948 -776 70987 -574
rect 70505 -810 70521 -776
rect 70897 -810 70987 -776
rect 67737 -981 67771 -965
rect 70430 -923 70521 -889
rect 70897 -923 70913 -889
rect 70430 -1125 70469 -923
rect 70948 -1007 70987 -810
rect 71838 -849 71854 -815
rect 72030 -849 72046 -815
rect 71838 -967 71854 -933
rect 72030 -967 72046 -933
rect 71842 -1007 72042 -967
rect 70505 -1041 70521 -1007
rect 70897 -1041 70987 -1007
rect 67502 -1181 67536 -1165
rect 70233 -1167 70343 -1151
rect 70430 -1159 70521 -1125
rect 70897 -1159 70913 -1125
rect 67309 -1249 67325 -1215
rect 67359 -1249 67375 -1215
rect 67427 -1249 67443 -1215
rect 67477 -1249 67493 -1215
rect 55516 -1329 55550 -1313
rect 65780 -1316 66589 -1276
rect 65799 -1317 66589 -1316
rect 42238 -1390 42254 -1356
rect 42288 -1390 42304 -1356
rect 48792 -1385 48808 -1351
rect 48842 -1385 48858 -1351
rect 55441 -1397 55457 -1363
rect 55491 -1397 55507 -1363
rect 64322 -1399 64592 -1365
rect 63496 -1449 63530 -1433
rect 42356 -1507 42372 -1473
rect 42406 -1507 42422 -1473
rect 48910 -1502 48926 -1468
rect 48960 -1502 48976 -1468
rect 55559 -1514 55575 -1480
rect 55609 -1514 55625 -1480
rect 41605 -1567 41639 -1551
rect 41605 -1759 41639 -1743
rect 41723 -1567 41757 -1551
rect 41723 -1759 41757 -1743
rect 41841 -1567 41875 -1551
rect 41841 -1759 41875 -1743
rect 41959 -1567 41993 -1551
rect 41959 -1759 41993 -1743
rect 42077 -1567 42111 -1551
rect 42077 -1759 42111 -1743
rect 42195 -1567 42229 -1551
rect 42195 -1759 42229 -1743
rect 42313 -1567 42347 -1551
rect 42313 -1759 42347 -1743
rect 42431 -1567 42465 -1551
rect 42431 -1793 42465 -1743
rect 42549 -1567 42583 -1551
rect 42549 -1759 42583 -1743
rect 42667 -1567 42701 -1551
rect 42667 -1793 42701 -1743
rect 48159 -1562 48193 -1546
rect 48159 -1754 48193 -1738
rect 48277 -1562 48311 -1546
rect 48277 -1754 48311 -1738
rect 48395 -1562 48429 -1546
rect 48395 -1754 48429 -1738
rect 48513 -1562 48547 -1546
rect 48513 -1754 48547 -1738
rect 48631 -1562 48665 -1546
rect 48631 -1754 48665 -1738
rect 48749 -1562 48783 -1546
rect 48749 -1754 48783 -1738
rect 48867 -1562 48901 -1546
rect 48867 -1754 48901 -1738
rect 48985 -1562 49019 -1546
rect 42431 -1827 42701 -1793
rect 48985 -1788 49019 -1738
rect 49103 -1562 49137 -1546
rect 49103 -1754 49137 -1738
rect 49221 -1562 49255 -1546
rect 49221 -1788 49255 -1738
rect 54808 -1574 54842 -1558
rect 54808 -1766 54842 -1750
rect 54926 -1574 54960 -1558
rect 54926 -1766 54960 -1750
rect 55044 -1574 55078 -1558
rect 55044 -1766 55078 -1750
rect 55162 -1574 55196 -1558
rect 55162 -1766 55196 -1750
rect 55280 -1574 55314 -1558
rect 55280 -1766 55314 -1750
rect 55398 -1574 55432 -1558
rect 55398 -1766 55432 -1750
rect 55516 -1574 55550 -1558
rect 55516 -1766 55550 -1750
rect 55634 -1574 55668 -1558
rect 48985 -1822 49255 -1788
rect 55634 -1800 55668 -1750
rect 55752 -1574 55786 -1558
rect 55752 -1766 55786 -1750
rect 55870 -1574 55904 -1558
rect 63496 -1641 63530 -1625
rect 63614 -1449 63648 -1433
rect 63614 -1641 63648 -1625
rect 63732 -1449 63766 -1433
rect 63732 -1641 63766 -1625
rect 63850 -1449 63884 -1433
rect 63850 -1641 63884 -1625
rect 63968 -1449 64002 -1433
rect 63968 -1641 64002 -1625
rect 64086 -1449 64120 -1433
rect 64086 -1641 64120 -1625
rect 64204 -1449 64238 -1433
rect 64204 -1641 64238 -1625
rect 64322 -1449 64356 -1399
rect 64322 -1641 64356 -1625
rect 64440 -1449 64474 -1433
rect 64440 -1641 64474 -1625
rect 64558 -1449 64592 -1399
rect 65677 -1406 65744 -1390
rect 65677 -1440 65693 -1406
rect 65727 -1440 65744 -1406
rect 65677 -1456 65744 -1440
rect 65508 -1473 65542 -1457
rect 65508 -1523 65542 -1507
rect 65854 -1558 65888 -1317
rect 67542 -1320 67710 -1302
rect 67542 -1376 67558 -1320
rect 67692 -1376 67710 -1320
rect 66324 -1406 66391 -1390
rect 67542 -1392 67710 -1376
rect 70233 -1363 70251 -1167
rect 70327 -1363 70343 -1167
rect 70948 -1243 70987 -1041
rect 71483 -1053 71568 -1037
rect 71838 -1041 71854 -1007
rect 72230 -1041 72246 -1007
rect 71096 -1101 71112 -1067
rect 71146 -1101 71162 -1067
rect 71483 -1113 71496 -1053
rect 71551 -1113 71568 -1053
rect 71483 -1129 71568 -1113
rect 70505 -1277 70521 -1243
rect 70897 -1277 70987 -1243
rect 71198 -1171 71283 -1155
rect 71838 -1159 71854 -1125
rect 72230 -1159 72246 -1125
rect 71198 -1231 71211 -1171
rect 71266 -1231 71283 -1171
rect 72479 -1225 72565 -1209
rect 71198 -1247 71283 -1231
rect 71838 -1277 71854 -1243
rect 72230 -1277 72246 -1243
rect 72331 -1244 72365 -1228
rect 70233 -1379 70343 -1363
rect 66324 -1440 66341 -1406
rect 66375 -1440 66391 -1406
rect 66324 -1456 66391 -1440
rect 70430 -1395 70521 -1361
rect 70897 -1395 70913 -1361
rect 66631 -1474 66665 -1458
rect 65943 -1524 65959 -1490
rect 65993 -1524 66009 -1490
rect 66061 -1523 66077 -1489
rect 66111 -1523 66127 -1489
rect 66631 -1524 66665 -1508
rect 64558 -1641 64592 -1625
rect 65361 -1574 65395 -1558
rect 64247 -1719 64263 -1685
rect 64297 -1719 64313 -1685
rect 55870 -1800 55904 -1750
rect 65361 -1766 65395 -1750
rect 65479 -1574 65513 -1558
rect 65479 -1766 65513 -1750
rect 65781 -1574 65815 -1558
rect 55634 -1834 55904 -1800
rect 64129 -1836 64145 -1802
rect 64179 -1836 64195 -1802
rect 63733 -1886 63767 -1870
rect 41894 -1913 42062 -1897
rect 41894 -1983 41910 -1913
rect 42046 -1983 42062 -1913
rect 41894 -1999 42062 -1983
rect 48448 -1908 48616 -1892
rect 48448 -1978 48464 -1908
rect 48600 -1978 48616 -1908
rect 48448 -1994 48616 -1978
rect 55097 -1920 55265 -1904
rect 55097 -1990 55113 -1920
rect 55249 -1990 55265 -1920
rect 55097 -2006 55265 -1990
rect 63733 -2278 63767 -2262
rect 63851 -1886 63885 -1870
rect 63851 -2278 63885 -2262
rect 63969 -1886 64003 -1870
rect 64086 -1886 64120 -1870
rect 64086 -2078 64120 -2062
rect 64204 -1886 64238 -1870
rect 65854 -1574 65933 -1558
rect 65854 -1604 65899 -1574
rect 65781 -2017 65816 -1950
rect 65899 -1966 65933 -1950
rect 66017 -1574 66051 -1558
rect 66017 -1966 66051 -1950
rect 66135 -1574 66169 -1558
rect 66253 -1574 66287 -1558
rect 66659 -1574 66693 -1558
rect 66659 -1766 66693 -1750
rect 66777 -1574 66811 -1558
rect 70430 -1597 70469 -1395
rect 70948 -1479 70987 -1277
rect 72331 -1294 72365 -1278
rect 72479 -1247 72497 -1225
rect 71716 -1336 71732 -1302
rect 71766 -1336 71782 -1302
rect 72479 -1305 72483 -1247
rect 72479 -1329 72497 -1305
rect 72543 -1329 72565 -1225
rect 72479 -1345 72565 -1329
rect 71838 -1395 71854 -1361
rect 72230 -1395 72246 -1361
rect 71326 -1455 71342 -1421
rect 71376 -1455 71392 -1421
rect 70505 -1513 70521 -1479
rect 70897 -1513 70987 -1479
rect 71838 -1513 71854 -1479
rect 72230 -1513 72246 -1479
rect 70430 -1631 70521 -1597
rect 70897 -1631 70913 -1597
rect 70948 -1716 70987 -1513
rect 71842 -1557 72042 -1513
rect 71838 -1591 71854 -1557
rect 72030 -1591 72046 -1557
rect 71838 -1709 71854 -1675
rect 72030 -1709 72046 -1675
rect 70505 -1750 70521 -1716
rect 70897 -1750 70987 -1716
rect 66777 -1766 66811 -1750
rect 66135 -1966 66169 -1950
rect 66252 -2017 66287 -1950
rect 65781 -2052 66287 -2017
rect 70430 -1868 70521 -1834
rect 70897 -1868 70913 -1834
rect 64204 -2078 64238 -2062
rect 70430 -2070 70469 -1868
rect 70948 -1952 70987 -1750
rect 70505 -1986 70521 -1952
rect 70897 -1986 70987 -1952
rect 70430 -2104 70521 -2070
rect 70897 -2104 70913 -2070
rect 65928 -2121 66170 -2109
rect 65928 -2223 65975 -2121
rect 66110 -2223 66170 -2121
rect 70705 -2223 70721 -2189
rect 70897 -2223 70990 -2189
rect 65928 -2240 66170 -2223
rect 63969 -2278 64003 -2262
rect 63776 -2346 63792 -2312
rect 63826 -2346 63842 -2312
rect 63894 -2346 63910 -2312
rect 63944 -2346 63960 -2312
rect 70634 -2341 70721 -2307
rect 70897 -2341 70913 -2307
rect 64009 -2417 64177 -2399
rect 64009 -2473 64025 -2417
rect 64159 -2473 64177 -2417
rect 64009 -2489 64177 -2473
rect 70634 -2543 70671 -2341
rect 70951 -2425 70990 -2223
rect 70705 -2459 70721 -2425
rect 70897 -2459 70990 -2425
rect 71071 -2377 71105 -2361
rect 71071 -2427 71105 -2411
rect 70634 -2577 70721 -2543
rect 70897 -2577 70913 -2543
rect 31371 -2768 31387 -2734
rect 31563 -2768 31579 -2734
rect 32528 -2809 33773 -2726
rect 33880 -2809 33894 -2726
rect 32528 -2822 33894 -2809
rect 36481 -2732 36672 -2717
rect 36481 -2798 36506 -2732
rect 36650 -2798 36672 -2732
rect 36481 -2819 36672 -2798
rect 31371 -2886 31387 -2852
rect 31563 -2886 31579 -2852
rect 1613 -2975 1647 -2959
rect 1613 -3025 1647 -3009
rect 4757 -2975 4791 -2959
rect 4757 -3025 4791 -3009
rect 7889 -2971 7923 -2955
rect 7889 -3021 7923 -3005
rect 11033 -2971 11067 -2955
rect 11033 -3021 11067 -3005
rect 14235 -2975 14269 -2959
rect 14235 -3025 14269 -3009
rect 17379 -2975 17413 -2959
rect 17379 -3025 17413 -3009
rect 20511 -2971 20545 -2955
rect 20511 -3021 20545 -3005
rect 23655 -2971 23689 -2955
rect 23655 -3021 23689 -3005
rect 30146 -3020 30162 -2986
rect 30338 -3020 30354 -2986
rect 1126 -3097 1160 -3081
rect 1126 -3289 1160 -3273
rect 1244 -3085 1278 -3081
rect 1318 -3085 1352 -3081
rect 1244 -3097 1352 -3085
rect 1278 -3273 1318 -3097
rect 1244 -3285 1318 -3273
rect 1244 -3289 1278 -3285
rect 1318 -3489 1352 -3473
rect 1436 -3097 1470 -3081
rect 1436 -3489 1470 -3473
rect 1554 -3097 1588 -3081
rect 1554 -3489 1588 -3473
rect 1672 -3097 1706 -3081
rect 1672 -3489 1706 -3473
rect 1790 -3085 1824 -3081
rect 1868 -3085 1902 -3081
rect 1790 -3097 1902 -3085
rect 1824 -3273 1868 -3097
rect 1824 -3285 1902 -3273
rect 1868 -3289 1902 -3285
rect 1986 -3097 2020 -3081
rect 1986 -3289 2020 -3273
rect 4270 -3097 4304 -3081
rect 4270 -3289 4304 -3273
rect 4388 -3085 4422 -3081
rect 4462 -3085 4496 -3081
rect 4388 -3097 4496 -3085
rect 4422 -3273 4462 -3097
rect 4388 -3285 4462 -3273
rect 4388 -3289 4422 -3285
rect 1790 -3489 1824 -3473
rect 4462 -3489 4496 -3473
rect 4580 -3097 4614 -3081
rect 4580 -3489 4614 -3473
rect 4698 -3097 4732 -3081
rect 4698 -3489 4732 -3473
rect 4816 -3097 4850 -3081
rect 4816 -3489 4850 -3473
rect 4934 -3085 4968 -3081
rect 5012 -3085 5046 -3081
rect 4934 -3097 5046 -3085
rect 4968 -3273 5012 -3097
rect 4968 -3285 5046 -3273
rect 5012 -3289 5046 -3285
rect 5130 -3097 5164 -3081
rect 5130 -3289 5164 -3273
rect 7402 -3093 7436 -3077
rect 7402 -3285 7436 -3269
rect 7520 -3081 7554 -3077
rect 7594 -3081 7628 -3077
rect 7520 -3093 7628 -3081
rect 7554 -3269 7594 -3093
rect 7520 -3281 7594 -3269
rect 7520 -3285 7554 -3281
rect 4934 -3489 4968 -3473
rect 7594 -3485 7628 -3469
rect 7712 -3093 7746 -3077
rect 7712 -3485 7746 -3469
rect 7830 -3093 7864 -3077
rect 7830 -3485 7864 -3469
rect 7948 -3093 7982 -3077
rect 7948 -3485 7982 -3469
rect 8066 -3081 8100 -3077
rect 8144 -3081 8178 -3077
rect 8066 -3093 8178 -3081
rect 8100 -3269 8144 -3093
rect 8100 -3281 8178 -3269
rect 8144 -3285 8178 -3281
rect 8262 -3093 8296 -3077
rect 8262 -3285 8296 -3269
rect 10546 -3093 10580 -3077
rect 10546 -3285 10580 -3269
rect 10664 -3081 10698 -3077
rect 10738 -3081 10772 -3077
rect 10664 -3093 10772 -3081
rect 10698 -3269 10738 -3093
rect 10664 -3281 10738 -3269
rect 10664 -3285 10698 -3281
rect 8066 -3485 8100 -3469
rect 10738 -3485 10772 -3469
rect 10856 -3093 10890 -3077
rect 10856 -3485 10890 -3469
rect 10974 -3093 11008 -3077
rect 10974 -3485 11008 -3469
rect 11092 -3093 11126 -3077
rect 11092 -3485 11126 -3469
rect 11210 -3081 11244 -3077
rect 11288 -3081 11322 -3077
rect 11210 -3093 11322 -3081
rect 11244 -3269 11288 -3093
rect 11244 -3281 11322 -3269
rect 11288 -3285 11322 -3281
rect 11406 -3093 11440 -3077
rect 11406 -3285 11440 -3269
rect 13748 -3097 13782 -3081
rect 13748 -3289 13782 -3273
rect 13866 -3085 13900 -3081
rect 13940 -3085 13974 -3081
rect 13866 -3097 13974 -3085
rect 13900 -3273 13940 -3097
rect 13866 -3285 13940 -3273
rect 13866 -3289 13900 -3285
rect 11210 -3485 11244 -3469
rect 13940 -3489 13974 -3473
rect 14058 -3097 14092 -3081
rect 14058 -3489 14092 -3473
rect 14176 -3097 14210 -3081
rect 14176 -3489 14210 -3473
rect 14294 -3097 14328 -3081
rect 14294 -3489 14328 -3473
rect 14412 -3085 14446 -3081
rect 14490 -3085 14524 -3081
rect 14412 -3097 14524 -3085
rect 14446 -3273 14490 -3097
rect 14446 -3285 14524 -3273
rect 14490 -3289 14524 -3285
rect 14608 -3097 14642 -3081
rect 14608 -3289 14642 -3273
rect 16892 -3097 16926 -3081
rect 16892 -3289 16926 -3273
rect 17010 -3085 17044 -3081
rect 17084 -3085 17118 -3081
rect 17010 -3097 17118 -3085
rect 17044 -3273 17084 -3097
rect 17010 -3285 17084 -3273
rect 17010 -3289 17044 -3285
rect 14412 -3489 14446 -3473
rect 17084 -3489 17118 -3473
rect 17202 -3097 17236 -3081
rect 17202 -3489 17236 -3473
rect 17320 -3097 17354 -3081
rect 17320 -3489 17354 -3473
rect 17438 -3097 17472 -3081
rect 17438 -3489 17472 -3473
rect 17556 -3085 17590 -3081
rect 17634 -3085 17668 -3081
rect 17556 -3097 17668 -3085
rect 17590 -3273 17634 -3097
rect 17590 -3285 17668 -3273
rect 17634 -3289 17668 -3285
rect 17752 -3097 17786 -3081
rect 17752 -3289 17786 -3273
rect 20024 -3093 20058 -3077
rect 20024 -3285 20058 -3269
rect 20142 -3081 20176 -3077
rect 20216 -3081 20250 -3077
rect 20142 -3093 20250 -3081
rect 20176 -3269 20216 -3093
rect 20142 -3281 20216 -3269
rect 20142 -3285 20176 -3281
rect 17556 -3489 17590 -3473
rect 20216 -3485 20250 -3469
rect 20334 -3093 20368 -3077
rect 20334 -3485 20368 -3469
rect 20452 -3093 20486 -3077
rect 20452 -3485 20486 -3469
rect 20570 -3093 20604 -3077
rect 20570 -3485 20604 -3469
rect 20688 -3081 20722 -3077
rect 20766 -3081 20800 -3077
rect 20688 -3093 20800 -3081
rect 20722 -3269 20766 -3093
rect 20722 -3281 20800 -3269
rect 20766 -3285 20800 -3281
rect 20884 -3093 20918 -3077
rect 20884 -3285 20918 -3269
rect 23168 -3093 23202 -3077
rect 23168 -3285 23202 -3269
rect 23286 -3081 23320 -3077
rect 23360 -3081 23394 -3077
rect 23286 -3093 23394 -3081
rect 23320 -3269 23360 -3093
rect 23286 -3281 23360 -3269
rect 23286 -3285 23320 -3281
rect 20688 -3485 20722 -3469
rect 23360 -3485 23394 -3469
rect 23478 -3093 23512 -3077
rect 23478 -3485 23512 -3469
rect 23596 -3093 23630 -3077
rect 23596 -3485 23630 -3469
rect 23714 -3093 23748 -3077
rect 23714 -3485 23748 -3469
rect 23832 -3081 23866 -3077
rect 23910 -3081 23944 -3077
rect 23832 -3093 23944 -3081
rect 23866 -3269 23910 -3093
rect 23866 -3281 23944 -3269
rect 23910 -3285 23944 -3281
rect 24028 -3093 24062 -3077
rect 24028 -3285 24062 -3269
rect 23832 -3485 23866 -3469
rect 1539 -3608 1555 -3574
rect 1589 -3608 1605 -3574
rect 4683 -3608 4699 -3574
rect 4733 -3608 4749 -3574
rect 7815 -3604 7831 -3570
rect 7865 -3604 7881 -3570
rect 10959 -3604 10975 -3570
rect 11009 -3604 11025 -3570
rect 14161 -3608 14177 -3574
rect 14211 -3608 14227 -3574
rect 17305 -3608 17321 -3574
rect 17355 -3608 17371 -3574
rect 20437 -3604 20453 -3570
rect 20487 -3604 20503 -3570
rect 23581 -3604 23597 -3570
rect 23631 -3604 23647 -3570
rect 7796 -3722 7932 -3718
rect 1520 -3726 1656 -3722
rect 1520 -3740 1558 -3726
rect 1616 -3740 1656 -3726
rect 1520 -3786 1536 -3740
rect 1640 -3786 1656 -3740
rect 1520 -3808 1656 -3786
rect 4664 -3726 4800 -3722
rect 4664 -3740 4702 -3726
rect 4760 -3740 4800 -3726
rect 4664 -3786 4680 -3740
rect 4784 -3786 4800 -3740
rect 4664 -3808 4800 -3786
rect 7796 -3736 7834 -3722
rect 7892 -3736 7932 -3722
rect 7796 -3782 7812 -3736
rect 7916 -3782 7932 -3736
rect 7796 -3804 7932 -3782
rect 10940 -3722 11076 -3718
rect 20418 -3722 20554 -3718
rect 10940 -3736 10978 -3722
rect 11036 -3736 11076 -3722
rect 10940 -3782 10956 -3736
rect 11060 -3782 11076 -3736
rect 10940 -3804 11076 -3782
rect 14142 -3726 14278 -3722
rect 14142 -3740 14180 -3726
rect 14238 -3740 14278 -3726
rect 14142 -3786 14158 -3740
rect 14262 -3786 14278 -3740
rect 14142 -3808 14278 -3786
rect 17286 -3726 17422 -3722
rect 17286 -3740 17324 -3726
rect 17382 -3740 17422 -3726
rect 17286 -3786 17302 -3740
rect 17406 -3786 17422 -3740
rect 17286 -3808 17422 -3786
rect 20418 -3736 20456 -3722
rect 20514 -3736 20554 -3722
rect 20418 -3782 20434 -3736
rect 20538 -3782 20554 -3736
rect 20418 -3804 20554 -3782
rect 23562 -3722 23698 -3718
rect 23562 -3736 23600 -3722
rect 23658 -3736 23698 -3722
rect 23562 -3782 23578 -3736
rect 23682 -3782 23698 -3736
rect 23562 -3804 23698 -3782
<< viali >>
rect 41810 24735 41844 24769
rect 42940 24741 42974 24775
rect 48323 24732 48357 24766
rect 49453 24738 49487 24772
rect 54857 24727 54891 24761
rect 55987 24733 56021 24767
rect 61415 24731 61449 24765
rect 62545 24737 62579 24771
rect 41810 24617 41844 24651
rect 42940 24621 42974 24655
rect 39600 24345 39634 24521
rect 39718 24345 39752 24521
rect 39836 24345 39870 24521
rect 39954 24345 39988 24521
rect 40072 24345 40106 24521
rect 40190 24345 40224 24521
rect 40308 24345 40342 24521
rect 40426 24345 40460 24521
rect 40544 24345 40578 24521
rect 40662 24345 40696 24521
rect 40367 24251 40401 24285
rect 41925 24217 41959 24593
rect 42043 24217 42077 24593
rect 42161 24217 42195 24593
rect 42279 24217 42313 24593
rect 42397 24217 42431 24593
rect 42515 24217 42549 24593
rect 48323 24614 48357 24648
rect 42633 24217 42667 24593
rect 43067 24221 43101 24597
rect 43185 24221 43219 24597
rect 43303 24221 43337 24597
rect 43421 24221 43455 24597
rect 43539 24221 43573 24597
rect 43657 24221 43691 24597
rect 43775 24221 43809 24597
rect 49453 24618 49487 24652
rect 46113 24342 46147 24518
rect 46231 24342 46265 24518
rect 46349 24342 46383 24518
rect 46467 24342 46501 24518
rect 46585 24342 46619 24518
rect 46703 24342 46737 24518
rect 46821 24342 46855 24518
rect 46939 24342 46973 24518
rect 47057 24342 47091 24518
rect 47175 24342 47209 24518
rect 46880 24248 46914 24282
rect 48438 24214 48472 24590
rect 48556 24214 48590 24590
rect 48674 24214 48708 24590
rect 48792 24214 48826 24590
rect 48910 24214 48944 24590
rect 49028 24214 49062 24590
rect 49146 24214 49180 24590
rect 49580 24218 49614 24594
rect 49698 24218 49732 24594
rect 49816 24218 49850 24594
rect 49934 24218 49968 24594
rect 50052 24218 50086 24594
rect 50170 24218 50204 24594
rect 54857 24609 54891 24643
rect 50288 24218 50322 24594
rect 55987 24613 56021 24647
rect 52647 24337 52681 24513
rect 52765 24337 52799 24513
rect 52883 24337 52917 24513
rect 53001 24337 53035 24513
rect 53119 24337 53153 24513
rect 53237 24337 53271 24513
rect 53355 24337 53389 24513
rect 53473 24337 53507 24513
rect 53591 24337 53625 24513
rect 53709 24337 53743 24513
rect 53414 24243 53448 24277
rect 54972 24209 55006 24585
rect 55090 24209 55124 24585
rect 55208 24209 55242 24585
rect 55326 24209 55360 24585
rect 55444 24209 55478 24585
rect 55562 24209 55596 24585
rect 61415 24613 61449 24647
rect 55680 24209 55714 24585
rect 56114 24213 56148 24589
rect 56232 24213 56266 24589
rect 56350 24213 56384 24589
rect 56468 24213 56502 24589
rect 56586 24213 56620 24589
rect 56704 24213 56738 24589
rect 56822 24213 56856 24589
rect 62545 24617 62579 24651
rect 59205 24341 59239 24517
rect 59323 24341 59357 24517
rect 59441 24341 59475 24517
rect 59559 24341 59593 24517
rect 59677 24341 59711 24517
rect 59795 24341 59829 24517
rect 59913 24341 59947 24517
rect 60031 24341 60065 24517
rect 60149 24341 60183 24517
rect 60267 24341 60301 24517
rect 59972 24247 60006 24281
rect 61530 24213 61564 24589
rect 61648 24213 61682 24589
rect 61766 24213 61800 24589
rect 61884 24213 61918 24589
rect 62002 24213 62036 24589
rect 62120 24213 62154 24589
rect 62238 24213 62272 24589
rect 62672 24217 62706 24593
rect 62790 24217 62824 24593
rect 62908 24217 62942 24593
rect 63026 24217 63060 24593
rect 63144 24217 63178 24593
rect 63262 24217 63296 24593
rect 63380 24217 63414 24593
rect 28285 24096 28342 24163
rect 40249 24134 40283 24168
rect 46762 24131 46796 24165
rect 53296 24126 53330 24160
rect 59854 24130 59888 24164
rect 4284 22180 4356 22234
rect 7428 22180 7500 22234
rect 10560 22176 10632 22230
rect 13704 22176 13776 22230
rect 16906 22180 16978 22234
rect 20050 22180 20122 22234
rect 23182 22176 23254 22230
rect 26326 22176 26398 22230
rect 3012 21608 3046 21784
rect 3130 21608 3164 21784
rect 3248 21608 3282 21784
rect 3366 21608 3400 21784
rect 3485 21608 3519 21984
rect 3603 21608 3637 21984
rect 3721 21608 3755 21984
rect 3839 21608 3873 21984
rect 3958 21608 3992 21984
rect 4076 21608 4110 21984
rect 4194 21608 4228 21984
rect 4312 21608 4346 21984
rect 4430 21608 4464 21984
rect 4548 21608 4582 21984
rect 4666 21608 4700 21984
rect 4779 21608 4813 21984
rect 4897 21608 4931 21984
rect 5015 21608 5049 21984
rect 5133 21608 5167 21984
rect 5220 21608 5254 21784
rect 5338 21608 5372 21784
rect 5456 21608 5490 21784
rect 5574 21608 5608 21784
rect 6156 21608 6190 21784
rect 6274 21608 6308 21784
rect 6392 21608 6426 21784
rect 6510 21608 6544 21784
rect 6629 21608 6663 21984
rect 6747 21608 6781 21984
rect 6865 21608 6899 21984
rect 6983 21608 7017 21984
rect 7102 21608 7136 21984
rect 7220 21608 7254 21984
rect 7338 21608 7372 21984
rect 7456 21608 7490 21984
rect 7574 21608 7608 21984
rect 7692 21608 7726 21984
rect 7810 21608 7844 21984
rect 7923 21608 7957 21984
rect 8041 21608 8075 21984
rect 8159 21608 8193 21984
rect 8277 21608 8311 21984
rect 8364 21608 8398 21784
rect 8482 21608 8516 21784
rect 8600 21608 8634 21784
rect 8718 21608 8752 21784
rect 9288 21604 9322 21780
rect 9406 21604 9440 21780
rect 9524 21604 9558 21780
rect 9642 21604 9676 21780
rect 9761 21604 9795 21980
rect 9879 21604 9913 21980
rect 9997 21604 10031 21980
rect 10115 21604 10149 21980
rect 10234 21604 10268 21980
rect 10352 21604 10386 21980
rect 10470 21604 10504 21980
rect 10588 21604 10622 21980
rect 10706 21604 10740 21980
rect 10824 21604 10858 21980
rect 10942 21604 10976 21980
rect 11055 21604 11089 21980
rect 11173 21604 11207 21980
rect 11291 21604 11325 21980
rect 11409 21604 11443 21980
rect 11496 21604 11530 21780
rect 11614 21604 11648 21780
rect 11732 21604 11766 21780
rect 11850 21604 11884 21780
rect 12432 21604 12466 21780
rect 12550 21604 12584 21780
rect 12668 21604 12702 21780
rect 12786 21604 12820 21780
rect 12905 21604 12939 21980
rect 13023 21604 13057 21980
rect 13141 21604 13175 21980
rect 13259 21604 13293 21980
rect 13378 21604 13412 21980
rect 13496 21604 13530 21980
rect 13614 21604 13648 21980
rect 13732 21604 13766 21980
rect 13850 21604 13884 21980
rect 13968 21604 14002 21980
rect 14086 21604 14120 21980
rect 14199 21604 14233 21980
rect 14317 21604 14351 21980
rect 14435 21604 14469 21980
rect 14553 21604 14587 21980
rect 14640 21604 14674 21780
rect 14758 21604 14792 21780
rect 14876 21604 14910 21780
rect 14994 21604 15028 21780
rect 15634 21608 15668 21784
rect 15752 21608 15786 21784
rect 15870 21608 15904 21784
rect 15988 21608 16022 21784
rect 16107 21608 16141 21984
rect 16225 21608 16259 21984
rect 16343 21608 16377 21984
rect 16461 21608 16495 21984
rect 16580 21608 16614 21984
rect 16698 21608 16732 21984
rect 16816 21608 16850 21984
rect 16934 21608 16968 21984
rect 17052 21608 17086 21984
rect 17170 21608 17204 21984
rect 17288 21608 17322 21984
rect 17401 21608 17435 21984
rect 17519 21608 17553 21984
rect 17637 21608 17671 21984
rect 17755 21608 17789 21984
rect 17842 21608 17876 21784
rect 17960 21608 17994 21784
rect 18078 21608 18112 21784
rect 18196 21608 18230 21784
rect 18778 21608 18812 21784
rect 18896 21608 18930 21784
rect 19014 21608 19048 21784
rect 19132 21608 19166 21784
rect 19251 21608 19285 21984
rect 19369 21608 19403 21984
rect 19487 21608 19521 21984
rect 19605 21608 19639 21984
rect 19724 21608 19758 21984
rect 19842 21608 19876 21984
rect 19960 21608 19994 21984
rect 20078 21608 20112 21984
rect 20196 21608 20230 21984
rect 20314 21608 20348 21984
rect 20432 21608 20466 21984
rect 20545 21608 20579 21984
rect 20663 21608 20697 21984
rect 20781 21608 20815 21984
rect 20899 21608 20933 21984
rect 20986 21608 21020 21784
rect 21104 21608 21138 21784
rect 21222 21608 21256 21784
rect 21340 21608 21374 21784
rect 21910 21604 21944 21780
rect 22028 21604 22062 21780
rect 22146 21604 22180 21780
rect 22264 21604 22298 21780
rect 22383 21604 22417 21980
rect 22501 21604 22535 21980
rect 22619 21604 22653 21980
rect 22737 21604 22771 21980
rect 22856 21604 22890 21980
rect 22974 21604 23008 21980
rect 23092 21604 23126 21980
rect 23210 21604 23244 21980
rect 23328 21604 23362 21980
rect 23446 21604 23480 21980
rect 23564 21604 23598 21980
rect 23677 21604 23711 21980
rect 23795 21604 23829 21980
rect 23913 21604 23947 21980
rect 24031 21604 24065 21980
rect 24118 21604 24152 21780
rect 24236 21604 24270 21780
rect 24354 21604 24388 21780
rect 24472 21604 24506 21780
rect 25054 21604 25088 21780
rect 25172 21604 25206 21780
rect 25290 21604 25324 21780
rect 25408 21604 25442 21780
rect 25527 21604 25561 21980
rect 25645 21604 25679 21980
rect 25763 21604 25797 21980
rect 25881 21604 25915 21980
rect 26000 21604 26034 21980
rect 26118 21604 26152 21980
rect 26236 21604 26270 21980
rect 26354 21604 26388 21980
rect 26472 21604 26506 21980
rect 26590 21604 26624 21980
rect 26708 21604 26742 21980
rect 26821 21604 26855 21980
rect 26939 21604 26973 21980
rect 27057 21604 27091 21980
rect 27175 21604 27209 21980
rect 27262 21604 27296 21780
rect 27380 21604 27414 21780
rect 27498 21604 27532 21780
rect 27616 21604 27650 21780
rect 3178 21400 3212 21434
rect 6322 21400 6356 21434
rect 4488 21359 4522 21393
rect 9454 21396 9488 21430
rect 7632 21359 7666 21393
rect 12598 21396 12632 21430
rect 10764 21355 10798 21389
rect 15800 21400 15834 21434
rect 13908 21355 13942 21389
rect 18944 21400 18978 21434
rect 17110 21359 17144 21393
rect 22076 21396 22110 21430
rect 20254 21359 20288 21393
rect 25220 21396 25254 21430
rect 23386 21355 23420 21389
rect 26530 21355 26564 21389
rect 27950 21392 28042 21436
rect 28412 23975 28469 24042
rect 4358 21239 4416 21294
rect 4416 21239 4418 21294
rect 5443 21238 5445 21293
rect 5445 21238 5503 21293
rect 7502 21239 7560 21294
rect 7560 21239 7562 21294
rect 8587 21238 8589 21293
rect 8589 21238 8647 21293
rect 10634 21235 10692 21290
rect 10692 21235 10694 21290
rect 11719 21234 11721 21289
rect 11721 21234 11779 21289
rect 13778 21235 13836 21290
rect 13836 21235 13838 21290
rect 14863 21234 14865 21289
rect 14865 21234 14923 21289
rect 16980 21239 17038 21294
rect 17038 21239 17040 21294
rect 18065 21238 18067 21293
rect 18067 21238 18125 21293
rect 20124 21239 20182 21294
rect 20182 21239 20184 21294
rect 21209 21238 21211 21293
rect 21211 21238 21269 21293
rect 23256 21235 23314 21290
rect 23314 21235 23316 21290
rect 24341 21234 24343 21289
rect 24343 21234 24401 21289
rect 26400 21235 26458 21290
rect 26458 21235 26460 21290
rect 27485 21234 27487 21289
rect 27487 21234 27545 21289
rect 27740 21230 27789 21290
rect 4134 21129 4168 21163
rect 5698 21118 5747 21178
rect 4476 20954 4534 21009
rect 4534 20954 4536 21009
rect 7278 21129 7312 21163
rect 8842 21118 8891 21178
rect 10410 21125 10444 21159
rect 11974 21114 12023 21174
rect 7620 20954 7678 21009
rect 7678 20954 7680 21009
rect 8842 20950 8891 21010
rect 10752 20950 10810 21005
rect 10810 20950 10812 21005
rect 11974 20946 12023 21006
rect 13554 21125 13588 21159
rect 16756 21129 16790 21163
rect 18320 21118 18369 21178
rect 19900 21129 19934 21163
rect 23032 21125 23066 21159
rect 24596 21114 24645 21174
rect 26176 21125 26210 21159
rect 13896 20950 13954 21005
rect 13954 20950 13956 21005
rect 15118 20946 15167 21006
rect 17098 20954 17156 21009
rect 17156 20954 17158 21009
rect 18320 20950 18369 21010
rect 20242 20954 20300 21009
rect 20300 20954 20302 21009
rect 21464 20950 21513 21010
rect 23374 20950 23432 21005
rect 23432 20950 23434 21005
rect 24596 20946 24645 21006
rect 26518 20950 26576 21005
rect 26576 20950 26578 21005
rect 27740 20946 27789 21006
rect 27950 20954 28042 20998
rect 28534 23857 28591 23924
rect 28541 20820 28591 20861
rect 4253 20739 4287 20773
rect 7397 20739 7431 20773
rect 10529 20735 10563 20769
rect 13673 20735 13707 20769
rect 16875 20739 16909 20773
rect 20019 20739 20053 20773
rect 23151 20735 23185 20769
rect 28658 23735 28715 23802
rect 26295 20735 26329 20769
rect 27950 20714 28042 20758
rect 3880 20475 3914 20651
rect 3998 20475 4032 20651
rect 4076 20275 4110 20651
rect 4194 20275 4228 20651
rect 4312 20275 4346 20651
rect 4430 20275 4464 20651
rect 4548 20275 4582 20651
rect 4622 20475 4656 20651
rect 4740 20475 4774 20651
rect 7024 20475 7058 20651
rect 7142 20475 7176 20651
rect 7220 20275 7254 20651
rect 7338 20275 7372 20651
rect 7456 20275 7490 20651
rect 7574 20275 7608 20651
rect 7692 20275 7726 20651
rect 7766 20475 7800 20651
rect 7884 20475 7918 20651
rect 10156 20471 10190 20647
rect 10274 20471 10308 20647
rect 10352 20271 10386 20647
rect 10470 20271 10504 20647
rect 10588 20271 10622 20647
rect 10706 20271 10740 20647
rect 10824 20271 10858 20647
rect 10898 20471 10932 20647
rect 11016 20471 11050 20647
rect 13300 20471 13334 20647
rect 13418 20471 13452 20647
rect 13496 20271 13530 20647
rect 13614 20271 13648 20647
rect 13732 20271 13766 20647
rect 13850 20271 13884 20647
rect 13968 20271 14002 20647
rect 14042 20471 14076 20647
rect 14160 20471 14194 20647
rect 16502 20475 16536 20651
rect 16620 20475 16654 20651
rect 16698 20275 16732 20651
rect 16816 20275 16850 20651
rect 16934 20275 16968 20651
rect 17052 20275 17086 20651
rect 17170 20275 17204 20651
rect 17244 20475 17278 20651
rect 17362 20475 17396 20651
rect 19646 20475 19680 20651
rect 19764 20475 19798 20651
rect 19842 20275 19876 20651
rect 19960 20275 19994 20651
rect 20078 20275 20112 20651
rect 20196 20275 20230 20651
rect 20314 20275 20348 20651
rect 20388 20475 20422 20651
rect 20506 20475 20540 20651
rect 22778 20471 22812 20647
rect 22896 20471 22930 20647
rect 22974 20271 23008 20647
rect 23092 20271 23126 20647
rect 23210 20271 23244 20647
rect 23328 20271 23362 20647
rect 23446 20271 23480 20647
rect 23520 20471 23554 20647
rect 23638 20471 23672 20647
rect 25922 20471 25956 20647
rect 26040 20471 26074 20647
rect 26118 20271 26152 20647
rect 26236 20271 26270 20647
rect 26354 20271 26388 20647
rect 26472 20271 26506 20647
rect 26590 20271 26624 20647
rect 26664 20471 26698 20647
rect 26782 20471 26816 20647
rect 39837 23708 39871 24084
rect 39955 23708 39989 24084
rect 40073 23708 40107 24084
rect 40190 23908 40224 24084
rect 40308 23908 40342 24084
rect 42130 23861 42164 23895
rect 43272 23865 43306 23899
rect 28780 23616 28837 23683
rect 39896 23624 39930 23658
rect 40014 23624 40048 23658
rect 41835 23634 41869 23810
rect 41953 23634 41987 23810
rect 42071 23634 42105 23810
rect 42189 23634 42223 23810
rect 42354 23634 42388 23810
rect 42472 23634 42506 23810
rect 42590 23634 42624 23810
rect 42708 23634 42742 23810
rect 42977 23638 43011 23814
rect 43095 23638 43129 23814
rect 43213 23638 43247 23814
rect 43331 23638 43365 23814
rect 43496 23638 43530 23814
rect 43614 23638 43648 23814
rect 43732 23638 43766 23814
rect 43850 23638 43884 23814
rect 46350 23705 46384 24081
rect 46468 23705 46502 24081
rect 46586 23705 46620 24081
rect 46703 23905 46737 24081
rect 46821 23905 46855 24081
rect 48643 23858 48677 23892
rect 49785 23862 49819 23896
rect 46409 23621 46443 23655
rect 46527 23621 46561 23655
rect 48348 23631 48382 23807
rect 48466 23631 48500 23807
rect 48584 23631 48618 23807
rect 48702 23631 48736 23807
rect 48867 23631 48901 23807
rect 48985 23631 49019 23807
rect 49103 23631 49137 23807
rect 49221 23631 49255 23807
rect 49490 23635 49524 23811
rect 49608 23635 49642 23811
rect 49726 23635 49760 23811
rect 49844 23635 49878 23811
rect 50009 23635 50043 23811
rect 50127 23635 50161 23811
rect 50245 23635 50279 23811
rect 50363 23635 50397 23811
rect 52884 23700 52918 24076
rect 53002 23700 53036 24076
rect 53120 23700 53154 24076
rect 53237 23900 53271 24076
rect 53355 23900 53389 24076
rect 55177 23853 55211 23887
rect 56319 23857 56353 23891
rect 52943 23616 52977 23650
rect 53061 23616 53095 23650
rect 54882 23626 54916 23802
rect 55000 23626 55034 23802
rect 55118 23626 55152 23802
rect 55236 23626 55270 23802
rect 55401 23626 55435 23802
rect 55519 23626 55553 23802
rect 55637 23626 55671 23802
rect 55755 23626 55789 23802
rect 56024 23630 56058 23806
rect 56142 23630 56176 23806
rect 56260 23630 56294 23806
rect 56378 23630 56412 23806
rect 56543 23630 56577 23806
rect 56661 23630 56695 23806
rect 56779 23630 56813 23806
rect 56897 23630 56931 23806
rect 59442 23704 59476 24080
rect 59560 23704 59594 24080
rect 59678 23704 59712 24080
rect 59795 23904 59829 24080
rect 59913 23904 59947 24080
rect 61735 23857 61769 23891
rect 62877 23861 62911 23895
rect 59501 23620 59535 23654
rect 59619 23620 59653 23654
rect 61440 23630 61474 23806
rect 61558 23630 61592 23806
rect 61676 23630 61710 23806
rect 61794 23630 61828 23806
rect 61959 23630 61993 23806
rect 62077 23630 62111 23806
rect 62195 23630 62229 23806
rect 62313 23630 62347 23806
rect 62582 23634 62616 23810
rect 62700 23634 62734 23810
rect 62818 23634 62852 23810
rect 62936 23634 62970 23810
rect 63101 23634 63135 23810
rect 63219 23634 63253 23810
rect 63337 23634 63371 23810
rect 63455 23634 63489 23810
rect 27951 20578 28043 20622
rect 33822 22803 33876 22852
rect 33666 22360 33735 22431
rect 28910 21963 28970 22039
rect 27950 20468 28042 20512
rect 33519 21936 33590 22007
rect 27949 20341 28042 20385
rect 29049 21508 29109 21584
rect 4311 20140 4345 20174
rect 7455 20140 7489 20174
rect 10587 20136 10621 20170
rect 13731 20136 13765 20170
rect 16933 20140 16967 20174
rect 20077 20140 20111 20174
rect 23209 20136 23243 20170
rect 26353 20136 26387 20170
rect 33376 21486 33447 21547
rect 27949 20103 28042 20147
rect 29192 21089 29252 21165
rect 4284 20008 4342 20022
rect 4284 19976 4342 20008
rect 7428 20008 7486 20022
rect 7428 19976 7486 20008
rect 10560 20004 10618 20018
rect 10560 19972 10618 20004
rect 13704 20004 13762 20018
rect 13704 19972 13762 20004
rect 16906 20008 16964 20022
rect 16906 19976 16964 20008
rect 20050 20008 20108 20022
rect 20050 19976 20108 20008
rect 23182 20004 23240 20018
rect 23182 19972 23240 20004
rect 26326 20004 26384 20018
rect 26326 19972 26384 20004
rect 27948 19879 28041 19923
rect 4624 16976 4704 17046
rect 4624 16974 4704 16976
rect 5792 16976 5872 17046
rect 5792 16974 5872 16976
rect 5318 16936 5352 16970
rect 6960 16976 7040 17046
rect 6960 16974 7040 16976
rect 6486 16936 6520 16970
rect 8128 16976 8208 17046
rect 8128 16974 8208 16976
rect 7654 16936 7688 16970
rect 9302 16974 9382 17044
rect 9302 16972 9382 16974
rect 8822 16936 8856 16970
rect 10470 16974 10550 17044
rect 10470 16972 10550 16974
rect 9996 16934 10030 16968
rect 11638 16974 11718 17044
rect 11638 16972 11718 16974
rect 11164 16934 11198 16968
rect 12806 16974 12886 17044
rect 12806 16972 12886 16974
rect 12332 16934 12366 16968
rect 13500 16934 13534 16968
rect 5318 16828 5352 16862
rect 6486 16828 6520 16862
rect 7654 16828 7688 16862
rect 8822 16828 8856 16862
rect 9996 16826 10030 16860
rect 11164 16826 11198 16860
rect 12332 16826 12366 16860
rect 13500 16826 13534 16860
rect 4520 16420 4554 16796
rect 4638 16420 4672 16796
rect 4756 16420 4790 16796
rect 4874 16420 4908 16796
rect 4992 16420 5026 16796
rect 5110 16420 5144 16796
rect 5228 16420 5262 16796
rect 5688 16422 5722 16798
rect 5806 16422 5840 16798
rect 5924 16422 5958 16798
rect 6042 16422 6076 16798
rect 6160 16422 6194 16798
rect 6278 16422 6312 16798
rect 6396 16422 6430 16798
rect 6856 16420 6890 16796
rect 6974 16420 7008 16796
rect 7092 16420 7126 16796
rect 7210 16420 7244 16796
rect 7328 16420 7362 16796
rect 7446 16420 7480 16796
rect 7564 16420 7598 16796
rect 8024 16422 8058 16798
rect 8142 16422 8176 16798
rect 8260 16422 8294 16798
rect 8378 16422 8412 16798
rect 8496 16422 8530 16798
rect 8614 16422 8648 16798
rect 8732 16422 8766 16798
rect 9198 16420 9232 16796
rect 9316 16420 9350 16796
rect 9434 16420 9468 16796
rect 9552 16420 9586 16796
rect 9670 16420 9704 16796
rect 9788 16420 9822 16796
rect 9906 16420 9940 16796
rect 10366 16418 10400 16794
rect 10484 16418 10518 16794
rect 10602 16418 10636 16794
rect 10720 16418 10754 16794
rect 10838 16418 10872 16794
rect 10956 16418 10990 16794
rect 11074 16418 11108 16794
rect 11534 16420 11568 16796
rect 11652 16420 11686 16796
rect 11770 16420 11804 16796
rect 11888 16420 11922 16796
rect 12006 16420 12040 16796
rect 12124 16420 12158 16796
rect 12242 16420 12276 16796
rect 12702 16420 12736 16796
rect 12820 16420 12854 16796
rect 12938 16420 12972 16796
rect 13056 16420 13090 16796
rect 13174 16420 13208 16796
rect 13292 16420 13326 16796
rect 13410 16420 13444 16796
rect 14498 16777 14558 16839
rect 15946 16777 16006 16839
rect 17444 16775 17504 16837
rect 18892 16775 18952 16837
rect 20412 16777 20472 16839
rect 21860 16777 21920 16839
rect 23358 16775 23418 16837
rect 24806 16775 24866 16837
rect 13803 16425 13837 16601
rect 13921 16425 13955 16601
rect 14039 16425 14073 16601
rect 14157 16425 14191 16601
rect 14275 16425 14309 16601
rect 14393 16425 14427 16601
rect 14511 16425 14545 16601
rect 14629 16425 14663 16601
rect 14747 16425 14781 16601
rect 14865 16425 14899 16601
rect 15251 16425 15285 16601
rect 15369 16425 15403 16601
rect 15487 16425 15521 16601
rect 15605 16425 15639 16601
rect 15723 16425 15757 16601
rect 15841 16425 15875 16601
rect 15959 16425 15993 16601
rect 16077 16425 16111 16601
rect 16195 16425 16229 16601
rect 16313 16425 16347 16601
rect 16749 16423 16783 16599
rect 16867 16423 16901 16599
rect 16985 16423 17019 16599
rect 17103 16423 17137 16599
rect 17221 16423 17255 16599
rect 17339 16423 17373 16599
rect 17457 16423 17491 16599
rect 17575 16423 17609 16599
rect 17693 16423 17727 16599
rect 17811 16423 17845 16599
rect 18197 16423 18231 16599
rect 18315 16423 18349 16599
rect 18433 16423 18467 16599
rect 18551 16423 18585 16599
rect 18669 16423 18703 16599
rect 18787 16423 18821 16599
rect 18905 16423 18939 16599
rect 19023 16423 19057 16599
rect 19141 16423 19175 16599
rect 19259 16423 19293 16599
rect 19717 16425 19751 16601
rect 19835 16425 19869 16601
rect 19953 16425 19987 16601
rect 20071 16425 20105 16601
rect 20189 16425 20223 16601
rect 20307 16425 20341 16601
rect 20425 16425 20459 16601
rect 20543 16425 20577 16601
rect 20661 16425 20695 16601
rect 20779 16425 20813 16601
rect 21165 16425 21199 16601
rect 21283 16425 21317 16601
rect 21401 16425 21435 16601
rect 21519 16425 21553 16601
rect 21637 16425 21671 16601
rect 21755 16425 21789 16601
rect 21873 16425 21907 16601
rect 21991 16425 22025 16601
rect 22109 16425 22143 16601
rect 22227 16425 22261 16601
rect 22663 16423 22697 16599
rect 22781 16423 22815 16599
rect 22899 16423 22933 16599
rect 23017 16423 23051 16599
rect 23135 16423 23169 16599
rect 23253 16423 23287 16599
rect 23371 16423 23405 16599
rect 23489 16423 23523 16599
rect 23607 16423 23641 16599
rect 23725 16423 23759 16599
rect 24111 16423 24145 16599
rect 24229 16423 24263 16599
rect 24347 16423 24381 16599
rect 24465 16423 24499 16599
rect 24583 16423 24617 16599
rect 24701 16423 24735 16599
rect 24819 16423 24853 16599
rect 24937 16423 24971 16599
rect 25055 16423 25089 16599
rect 25173 16423 25207 16599
rect 14098 16331 14132 16365
rect 15546 16331 15580 16365
rect 17044 16329 17078 16363
rect 18492 16329 18526 16363
rect 20012 16331 20046 16365
rect 21460 16331 21494 16365
rect 22958 16329 22992 16363
rect 24406 16329 24440 16363
rect 14216 16214 14250 16248
rect 15664 16214 15698 16248
rect 17162 16212 17196 16246
rect 18610 16212 18644 16246
rect 20130 16214 20164 16248
rect 21578 16214 21612 16248
rect 23076 16212 23110 16246
rect 24524 16212 24558 16246
rect 5023 16065 5057 16099
rect 6191 16065 6225 16099
rect 7359 16065 7393 16099
rect 8527 16065 8561 16099
rect 9701 16063 9735 16097
rect 4445 15832 4479 16008
rect 4563 15832 4597 16008
rect 4681 15832 4715 16008
rect 4799 15832 4833 16008
rect 4964 15838 4998 16014
rect 5082 15838 5116 16014
rect 5200 15838 5234 16014
rect 5318 15838 5352 16014
rect 5613 15831 5647 16007
rect 5731 15831 5765 16007
rect 5849 15831 5883 16007
rect 5967 15831 6001 16007
rect 6132 15838 6166 16014
rect 6250 15838 6284 16014
rect 6368 15838 6402 16014
rect 6486 15838 6520 16014
rect 6781 15831 6815 16007
rect 6899 15831 6933 16007
rect 7017 15831 7051 16007
rect 7135 15831 7169 16007
rect 7300 15836 7334 16012
rect 7418 15836 7452 16012
rect 7536 15836 7570 16012
rect 7654 15836 7688 16012
rect 7950 15832 7984 16008
rect 8068 15832 8102 16008
rect 5102 15704 5168 15708
rect 1782 15042 1854 15096
rect 510 14470 544 14646
rect 628 14470 662 14646
rect 746 14470 780 14646
rect 864 14470 898 14646
rect 983 14470 1017 14846
rect 1101 14470 1135 14846
rect 1219 14470 1253 14846
rect 1337 14470 1371 14846
rect 1456 14470 1490 14846
rect 1574 14470 1608 14846
rect 1692 14470 1726 14846
rect 1810 14470 1844 14846
rect 1928 14470 1962 14846
rect 2046 14470 2080 14846
rect 2164 14470 2198 14846
rect 2277 14470 2311 14846
rect 2395 14470 2429 14846
rect 2513 14470 2547 14846
rect 2631 14470 2665 14846
rect 2718 14470 2752 14646
rect 2836 14470 2870 14646
rect 2954 14470 2988 14646
rect 3072 14470 3106 14646
rect 676 14262 710 14296
rect 1986 14221 2020 14255
rect 1856 14101 1914 14156
rect 1914 14101 1916 14156
rect 2941 14100 2943 14155
rect 2943 14100 3001 14155
rect 1632 13991 1666 14025
rect 3196 13980 3245 14040
rect 5102 15638 5168 15704
rect 8186 15832 8220 16008
rect 8304 15832 8338 16008
rect 8468 15836 8502 16012
rect 8586 15836 8620 16012
rect 8704 15836 8738 16012
rect 8822 15836 8856 16012
rect 9122 15836 9156 16012
rect 9240 15836 9274 16012
rect 9358 15836 9392 16012
rect 9476 15836 9510 16012
rect 9642 15836 9676 16012
rect 9760 15836 9794 16012
rect 9878 15836 9912 16012
rect 9996 15836 10030 16012
rect 6270 15704 6336 15708
rect 6270 15638 6336 15704
rect 7438 15704 7504 15708
rect 7438 15638 7504 15704
rect 8606 15704 8672 15708
rect 8606 15638 8672 15704
rect 9780 15702 9846 15706
rect 9780 15636 9846 15702
rect 4926 15042 4998 15096
rect 3654 14470 3688 14646
rect 3772 14470 3806 14646
rect 3890 14470 3924 14646
rect 4008 14470 4042 14646
rect 4127 14470 4161 14846
rect 4245 14470 4279 14846
rect 4363 14470 4397 14846
rect 4481 14470 4515 14846
rect 4600 14470 4634 14846
rect 4718 14470 4752 14846
rect 4836 14470 4870 14846
rect 4954 14470 4988 14846
rect 5072 14470 5106 14846
rect 5190 14470 5224 14846
rect 5308 14470 5342 14846
rect 5421 14470 5455 14846
rect 5539 14470 5573 14846
rect 5657 14470 5691 14846
rect 5775 14470 5809 14846
rect 5862 14470 5896 14646
rect 5980 14470 6014 14646
rect 6098 14470 6132 14646
rect 6216 14470 6250 14646
rect 3820 14262 3854 14296
rect 5130 14221 5164 14255
rect 8058 15038 8130 15092
rect 6786 14466 6820 14642
rect 6904 14466 6938 14642
rect 7022 14466 7056 14642
rect 7140 14466 7174 14642
rect 7259 14466 7293 14842
rect 7377 14466 7411 14842
rect 7495 14466 7529 14842
rect 7613 14466 7647 14842
rect 7732 14466 7766 14842
rect 7850 14466 7884 14842
rect 7968 14466 8002 14842
rect 8086 14466 8120 14842
rect 8204 14466 8238 14842
rect 8322 14466 8356 14842
rect 8440 14466 8474 14842
rect 8553 14466 8587 14842
rect 8671 14466 8705 14842
rect 8789 14466 8823 14842
rect 8907 14466 8941 14842
rect 8994 14466 9028 14642
rect 9112 14466 9146 14642
rect 9230 14466 9264 14642
rect 9348 14466 9382 14642
rect 6952 14258 6986 14292
rect 5000 14101 5058 14156
rect 5058 14101 5060 14156
rect 6085 14100 6087 14155
rect 6087 14100 6145 14155
rect 4776 13991 4810 14025
rect 6340 13980 6389 14040
rect 1974 13816 2032 13871
rect 2032 13816 2034 13871
rect 3196 13812 3245 13872
rect 5118 13816 5176 13871
rect 5176 13816 5178 13871
rect 8262 14217 8296 14251
rect 8132 14097 8190 14152
rect 8190 14097 8192 14152
rect 9217 14096 9219 14151
rect 9219 14096 9277 14151
rect 7908 13987 7942 14021
rect 9472 13976 9521 14036
rect 6340 13812 6389 13872
rect 8250 13812 8308 13867
rect 8308 13812 8310 13867
rect 9472 13808 9521 13868
rect 10869 16063 10903 16097
rect 12037 16063 12071 16097
rect 13205 16063 13239 16097
rect 10291 15836 10325 16012
rect 10409 15836 10443 16012
rect 10527 15836 10561 16012
rect 10645 15836 10679 16012
rect 10810 15836 10844 16012
rect 10928 15836 10962 16012
rect 11046 15836 11080 16012
rect 11164 15836 11198 16012
rect 11459 15836 11493 16012
rect 11577 15836 11611 16012
rect 11695 15836 11729 16012
rect 11813 15836 11847 16012
rect 11978 15836 12012 16012
rect 12096 15836 12130 16012
rect 12214 15836 12248 16012
rect 12332 15836 12366 16012
rect 12626 15830 12660 16006
rect 12744 15830 12778 16006
rect 12862 15830 12896 16006
rect 12980 15830 13014 16006
rect 13146 15834 13180 16010
rect 13264 15834 13298 16010
rect 13382 15834 13416 16010
rect 13500 15834 13534 16010
rect 14157 15988 14191 16164
rect 14275 15988 14309 16164
rect 14392 15788 14426 16164
rect 14510 15788 14544 16164
rect 14628 15788 14662 16164
rect 15605 15988 15639 16164
rect 15723 15988 15757 16164
rect 15840 15788 15874 16164
rect 15958 15788 15992 16164
rect 16076 15788 16110 16164
rect 17103 15986 17137 16162
rect 17221 15986 17255 16162
rect 17338 15786 17372 16162
rect 17456 15786 17490 16162
rect 17574 15786 17608 16162
rect 18551 15986 18585 16162
rect 18669 15986 18703 16162
rect 18786 15786 18820 16162
rect 18904 15786 18938 16162
rect 19022 15786 19056 16162
rect 20071 15988 20105 16164
rect 20189 15988 20223 16164
rect 20306 15788 20340 16164
rect 20424 15788 20458 16164
rect 20542 15788 20576 16164
rect 21519 15988 21553 16164
rect 21637 15988 21671 16164
rect 21754 15788 21788 16164
rect 21872 15788 21906 16164
rect 21990 15788 22024 16164
rect 23017 15986 23051 16162
rect 23135 15986 23169 16162
rect 23252 15786 23286 16162
rect 23370 15786 23404 16162
rect 23488 15786 23522 16162
rect 24465 15986 24499 16162
rect 24583 15986 24617 16162
rect 24700 15786 24734 16162
rect 24818 15786 24852 16162
rect 24936 15786 24970 16162
rect 10948 15702 11014 15706
rect 10948 15636 11014 15702
rect 12116 15702 12182 15706
rect 12116 15636 12182 15702
rect 13284 15702 13350 15706
rect 14451 15704 14485 15738
rect 14569 15704 14603 15738
rect 15899 15704 15933 15738
rect 16017 15704 16051 15738
rect 17397 15702 17431 15736
rect 17515 15702 17549 15736
rect 18845 15702 18879 15736
rect 18963 15702 18997 15736
rect 20365 15704 20399 15738
rect 20483 15704 20517 15738
rect 21813 15704 21847 15738
rect 21931 15704 21965 15738
rect 23311 15702 23345 15736
rect 23429 15702 23463 15736
rect 24759 15702 24793 15736
rect 24877 15702 24911 15736
rect 13284 15636 13350 15702
rect 14278 15581 14330 15627
rect 15726 15581 15778 15627
rect 17224 15579 17276 15625
rect 18672 15579 18724 15625
rect 20192 15581 20244 15627
rect 21640 15581 21692 15627
rect 23138 15579 23190 15625
rect 24586 15579 24638 15625
rect 11202 15038 11274 15092
rect 9930 14466 9964 14642
rect 10048 14466 10082 14642
rect 10166 14466 10200 14642
rect 10284 14466 10318 14642
rect 10403 14466 10437 14842
rect 10521 14466 10555 14842
rect 10639 14466 10673 14842
rect 10757 14466 10791 14842
rect 10876 14466 10910 14842
rect 10994 14466 11028 14842
rect 11112 14466 11146 14842
rect 11230 14466 11264 14842
rect 11348 14466 11382 14842
rect 11466 14466 11500 14842
rect 11584 14466 11618 14842
rect 11697 14466 11731 14842
rect 11815 14466 11849 14842
rect 11933 14466 11967 14842
rect 12051 14466 12085 14842
rect 12138 14466 12172 14642
rect 12256 14466 12290 14642
rect 12374 14466 12408 14642
rect 12492 14466 12526 14642
rect 10096 14258 10130 14292
rect 11406 14217 11440 14251
rect 11276 14097 11334 14152
rect 11334 14097 11336 14152
rect 12361 14096 12363 14151
rect 12363 14096 12421 14151
rect 11052 13987 11086 14021
rect 12616 13976 12665 14036
rect 14404 15042 14476 15096
rect 17548 15042 17620 15096
rect 13132 14470 13166 14646
rect 13250 14470 13284 14646
rect 13368 14470 13402 14646
rect 13486 14470 13520 14646
rect 13605 14470 13639 14846
rect 13723 14470 13757 14846
rect 13841 14470 13875 14846
rect 13959 14470 13993 14846
rect 14078 14470 14112 14846
rect 14196 14470 14230 14846
rect 14314 14470 14348 14846
rect 14432 14470 14466 14846
rect 14550 14470 14584 14846
rect 14668 14470 14702 14846
rect 14786 14470 14820 14846
rect 14899 14470 14933 14846
rect 15017 14470 15051 14846
rect 15135 14470 15169 14846
rect 15253 14470 15287 14846
rect 15340 14470 15374 14646
rect 15458 14470 15492 14646
rect 15576 14470 15610 14646
rect 15694 14470 15728 14646
rect 16276 14470 16310 14646
rect 16394 14470 16428 14646
rect 16512 14470 16546 14646
rect 16630 14470 16664 14646
rect 16749 14470 16783 14846
rect 16867 14470 16901 14846
rect 16985 14470 17019 14846
rect 17103 14470 17137 14846
rect 17222 14470 17256 14846
rect 17340 14470 17374 14846
rect 17458 14470 17492 14846
rect 17576 14470 17610 14846
rect 17694 14470 17728 14846
rect 17812 14470 17846 14846
rect 17930 14470 17964 14846
rect 18043 14470 18077 14846
rect 18161 14470 18195 14846
rect 18279 14470 18313 14846
rect 18397 14470 18431 14846
rect 18484 14470 18518 14646
rect 18602 14470 18636 14646
rect 18720 14470 18754 14646
rect 18838 14470 18872 14646
rect 13298 14262 13332 14296
rect 16442 14262 16476 14296
rect 14608 14221 14642 14255
rect 17752 14221 17786 14255
rect 14478 14101 14536 14156
rect 14536 14101 14538 14156
rect 15563 14100 15565 14155
rect 15565 14100 15623 14155
rect 17622 14101 17680 14156
rect 17680 14101 17682 14156
rect 18707 14100 18709 14155
rect 18709 14100 18767 14155
rect 14254 13991 14288 14025
rect 15818 13980 15867 14040
rect 17398 13991 17432 14025
rect 18962 13980 19011 14040
rect 20680 15038 20752 15092
rect 19408 14466 19442 14642
rect 19526 14466 19560 14642
rect 19644 14466 19678 14642
rect 19762 14466 19796 14642
rect 19881 14466 19915 14842
rect 19999 14466 20033 14842
rect 20117 14466 20151 14842
rect 20235 14466 20269 14842
rect 20354 14466 20388 14842
rect 20472 14466 20506 14842
rect 20590 14466 20624 14842
rect 20708 14466 20742 14842
rect 20826 14466 20860 14842
rect 20944 14466 20978 14842
rect 21062 14466 21096 14842
rect 21175 14466 21209 14842
rect 21293 14466 21327 14842
rect 21411 14466 21445 14842
rect 21529 14466 21563 14842
rect 21616 14466 21650 14642
rect 21734 14466 21768 14642
rect 21852 14466 21886 14642
rect 21970 14466 22004 14642
rect 19574 14258 19608 14292
rect 20884 14217 20918 14251
rect 20754 14097 20812 14152
rect 20812 14097 20814 14152
rect 21839 14096 21841 14151
rect 21841 14096 21899 14151
rect 20530 13987 20564 14021
rect 22094 13976 22143 14036
rect 17740 13816 17798 13871
rect 17798 13816 17800 13871
rect 18962 13812 19011 13872
rect 23824 15038 23896 15092
rect 22552 14466 22586 14642
rect 22670 14466 22704 14642
rect 22788 14466 22822 14642
rect 22906 14466 22940 14642
rect 23025 14466 23059 14842
rect 23143 14466 23177 14842
rect 23261 14466 23295 14842
rect 23379 14466 23413 14842
rect 23498 14466 23532 14842
rect 23616 14466 23650 14842
rect 23734 14466 23768 14842
rect 23852 14466 23886 14842
rect 23970 14466 24004 14842
rect 24088 14466 24122 14842
rect 24206 14466 24240 14842
rect 24319 14466 24353 14842
rect 24437 14466 24471 14842
rect 24555 14466 24589 14842
rect 24673 14466 24707 14842
rect 24760 14466 24794 14642
rect 24878 14466 24912 14642
rect 24996 14466 25030 14642
rect 25114 14466 25148 14642
rect 22718 14258 22752 14292
rect 24028 14217 24062 14251
rect 23898 14097 23956 14152
rect 23956 14097 23958 14152
rect 24983 14096 24985 14151
rect 24985 14096 25043 14151
rect 23674 13987 23708 14021
rect 25238 13976 25287 14036
rect 20872 13812 20930 13867
rect 20930 13812 20932 13867
rect 22094 13808 22143 13868
rect 24016 13812 24074 13867
rect 24074 13812 24076 13867
rect 25238 13808 25287 13868
rect 1751 13601 1785 13635
rect 4895 13601 4929 13635
rect 8027 13597 8061 13631
rect 11171 13597 11205 13631
rect 14373 13601 14407 13635
rect 17517 13601 17551 13635
rect 20649 13597 20683 13631
rect 23793 13597 23827 13631
rect 1378 13337 1412 13513
rect 1496 13337 1530 13513
rect 1574 13137 1608 13513
rect 1692 13137 1726 13513
rect 1810 13137 1844 13513
rect 1928 13137 1962 13513
rect 2046 13137 2080 13513
rect 2120 13337 2154 13513
rect 2238 13337 2272 13513
rect 4522 13337 4556 13513
rect 4640 13337 4674 13513
rect 4718 13137 4752 13513
rect 4836 13137 4870 13513
rect 4954 13137 4988 13513
rect 5072 13137 5106 13513
rect 5190 13137 5224 13513
rect 5264 13337 5298 13513
rect 5382 13337 5416 13513
rect 7654 13333 7688 13509
rect 7772 13333 7806 13509
rect 7850 13133 7884 13509
rect 7968 13133 8002 13509
rect 8086 13133 8120 13509
rect 8204 13133 8238 13509
rect 8322 13133 8356 13509
rect 8396 13333 8430 13509
rect 8514 13333 8548 13509
rect 10798 13333 10832 13509
rect 10916 13333 10950 13509
rect 10994 13133 11028 13509
rect 11112 13133 11146 13509
rect 11230 13133 11264 13509
rect 11348 13133 11382 13509
rect 11466 13133 11500 13509
rect 11540 13333 11574 13509
rect 11658 13333 11692 13509
rect 14000 13337 14034 13513
rect 14118 13337 14152 13513
rect 14196 13137 14230 13513
rect 14314 13137 14348 13513
rect 14432 13137 14466 13513
rect 14550 13137 14584 13513
rect 14668 13137 14702 13513
rect 14742 13337 14776 13513
rect 14860 13337 14894 13513
rect 17144 13337 17178 13513
rect 17262 13337 17296 13513
rect 17340 13137 17374 13513
rect 17458 13137 17492 13513
rect 17576 13137 17610 13513
rect 17694 13137 17728 13513
rect 17812 13137 17846 13513
rect 17886 13337 17920 13513
rect 18004 13337 18038 13513
rect 20276 13333 20310 13509
rect 20394 13333 20428 13509
rect 20472 13133 20506 13509
rect 20590 13133 20624 13509
rect 20708 13133 20742 13509
rect 20826 13133 20860 13509
rect 20944 13133 20978 13509
rect 21018 13333 21052 13509
rect 21136 13333 21170 13509
rect 23420 13333 23454 13509
rect 23538 13333 23572 13509
rect 23616 13133 23650 13509
rect 23734 13133 23768 13509
rect 23852 13133 23886 13509
rect 23970 13133 24004 13509
rect 24088 13133 24122 13509
rect 24162 13333 24196 13509
rect 24280 13333 24314 13509
rect 30166 13134 30342 13168
rect 30701 13145 30761 13161
rect 1809 13002 1843 13036
rect 4953 13002 4987 13036
rect 8085 12998 8119 13032
rect 11229 12998 11263 13032
rect 14431 13002 14465 13036
rect 17575 13002 17609 13036
rect 20707 12998 20741 13032
rect 23851 12998 23885 13032
rect 30701 13111 30715 13145
rect 30715 13111 30749 13145
rect 30749 13111 30761 13145
rect 30701 13095 30761 13111
rect 30166 13016 30342 13050
rect 31391 13009 31567 13043
rect 30166 12898 30342 12932
rect 1782 12870 1840 12884
rect 1782 12838 1840 12870
rect 4926 12870 4984 12884
rect 4926 12838 4984 12870
rect 8058 12866 8116 12880
rect 8058 12834 8116 12866
rect 11202 12866 11260 12880
rect 11202 12834 11260 12866
rect 14404 12870 14462 12884
rect 14404 12838 14462 12870
rect 17548 12870 17606 12884
rect 17548 12838 17606 12870
rect 20680 12866 20738 12880
rect 20680 12834 20738 12866
rect 23824 12866 23882 12880
rect 23824 12834 23882 12866
rect 31290 12862 31324 12896
rect 31391 12891 31567 12925
rect 30166 12780 30342 12814
rect 30659 12707 31035 12741
rect 29966 12650 30342 12684
rect 31223 12677 31257 12711
rect 30659 12589 31035 12623
rect 31391 12589 31767 12623
rect 29966 12532 30342 12566
rect 30659 12471 31035 12505
rect 1782 12308 1854 12362
rect 4926 12308 4998 12362
rect 8058 12304 8130 12358
rect 11202 12304 11274 12358
rect 14404 12308 14476 12362
rect 17548 12308 17620 12362
rect 20680 12304 20752 12358
rect 23824 12304 23896 12358
rect 29966 12414 30342 12448
rect 31391 12471 31767 12505
rect 31307 12411 31341 12445
rect 30659 12353 31035 12387
rect 31391 12353 31767 12387
rect 29711 12293 29739 12331
rect 29739 12293 29749 12331
rect 29966 12296 30342 12330
rect 510 11736 544 11912
rect 628 11736 662 11912
rect 746 11736 780 11912
rect 864 11736 898 11912
rect 983 11736 1017 12112
rect 1101 11736 1135 12112
rect 1219 11736 1253 12112
rect 1337 11736 1371 12112
rect 1456 11736 1490 12112
rect 1574 11736 1608 12112
rect 1692 11736 1726 12112
rect 1810 11736 1844 12112
rect 1928 11736 1962 12112
rect 2046 11736 2080 12112
rect 2164 11736 2198 12112
rect 2277 11736 2311 12112
rect 2395 11736 2429 12112
rect 2513 11736 2547 12112
rect 2631 11736 2665 12112
rect 2718 11736 2752 11912
rect 2836 11736 2870 11912
rect 2954 11736 2988 11912
rect 3072 11736 3106 11912
rect 3654 11736 3688 11912
rect 3772 11736 3806 11912
rect 3890 11736 3924 11912
rect 4008 11736 4042 11912
rect 4127 11736 4161 12112
rect 4245 11736 4279 12112
rect 4363 11736 4397 12112
rect 4481 11736 4515 12112
rect 4600 11736 4634 12112
rect 4718 11736 4752 12112
rect 4836 11736 4870 12112
rect 4954 11736 4988 12112
rect 5072 11736 5106 12112
rect 5190 11736 5224 12112
rect 5308 11736 5342 12112
rect 5421 11736 5455 12112
rect 5539 11736 5573 12112
rect 5657 11736 5691 12112
rect 5775 11736 5809 12112
rect 5862 11736 5896 11912
rect 5980 11736 6014 11912
rect 6098 11736 6132 11912
rect 6216 11736 6250 11912
rect 6786 11732 6820 11908
rect 6904 11732 6938 11908
rect 7022 11732 7056 11908
rect 7140 11732 7174 11908
rect 7259 11732 7293 12108
rect 7377 11732 7411 12108
rect 7495 11732 7529 12108
rect 7613 11732 7647 12108
rect 7732 11732 7766 12108
rect 7850 11732 7884 12108
rect 7968 11732 8002 12108
rect 8086 11732 8120 12108
rect 8204 11732 8238 12108
rect 8322 11732 8356 12108
rect 8440 11732 8474 12108
rect 8553 11732 8587 12108
rect 8671 11732 8705 12108
rect 8789 11732 8823 12108
rect 8907 11732 8941 12108
rect 8994 11732 9028 11908
rect 9112 11732 9146 11908
rect 9230 11732 9264 11908
rect 9348 11732 9382 11908
rect 9930 11732 9964 11908
rect 10048 11732 10082 11908
rect 10166 11732 10200 11908
rect 10284 11732 10318 11908
rect 10403 11732 10437 12108
rect 10521 11732 10555 12108
rect 10639 11732 10673 12108
rect 10757 11732 10791 12108
rect 10876 11732 10910 12108
rect 10994 11732 11028 12108
rect 11112 11732 11146 12108
rect 11230 11732 11264 12108
rect 11348 11732 11382 12108
rect 11466 11732 11500 12108
rect 11584 11732 11618 12108
rect 11697 11732 11731 12108
rect 11815 11732 11849 12108
rect 11933 11732 11967 12108
rect 12051 11732 12085 12108
rect 12138 11732 12172 11908
rect 12256 11732 12290 11908
rect 12374 11732 12408 11908
rect 12492 11732 12526 11908
rect 13132 11736 13166 11912
rect 13250 11736 13284 11912
rect 13368 11736 13402 11912
rect 13486 11736 13520 11912
rect 13605 11736 13639 12112
rect 13723 11736 13757 12112
rect 13841 11736 13875 12112
rect 13959 11736 13993 12112
rect 14078 11736 14112 12112
rect 14196 11736 14230 12112
rect 14314 11736 14348 12112
rect 14432 11736 14466 12112
rect 14550 11736 14584 12112
rect 14668 11736 14702 12112
rect 14786 11736 14820 12112
rect 14899 11736 14933 12112
rect 15017 11736 15051 12112
rect 15135 11736 15169 12112
rect 15253 11736 15287 12112
rect 15340 11736 15374 11912
rect 15458 11736 15492 11912
rect 15576 11736 15610 11912
rect 15694 11736 15728 11912
rect 16276 11736 16310 11912
rect 16394 11736 16428 11912
rect 16512 11736 16546 11912
rect 16630 11736 16664 11912
rect 16749 11736 16783 12112
rect 16867 11736 16901 12112
rect 16985 11736 17019 12112
rect 17103 11736 17137 12112
rect 17222 11736 17256 12112
rect 17340 11736 17374 12112
rect 17458 11736 17492 12112
rect 17576 11736 17610 12112
rect 17694 11736 17728 12112
rect 17812 11736 17846 12112
rect 17930 11736 17964 12112
rect 18043 11736 18077 12112
rect 18161 11736 18195 12112
rect 18279 11736 18313 12112
rect 18397 11736 18431 12112
rect 18484 11736 18518 11912
rect 18602 11736 18636 11912
rect 18720 11736 18754 11912
rect 18838 11736 18872 11912
rect 19408 11732 19442 11908
rect 19526 11732 19560 11908
rect 19644 11732 19678 11908
rect 19762 11732 19796 11908
rect 19881 11732 19915 12108
rect 19999 11732 20033 12108
rect 20117 11732 20151 12108
rect 20235 11732 20269 12108
rect 20354 11732 20388 12108
rect 20472 11732 20506 12108
rect 20590 11732 20624 12108
rect 20708 11732 20742 12108
rect 20826 11732 20860 12108
rect 20944 11732 20978 12108
rect 21062 11732 21096 12108
rect 21175 11732 21209 12108
rect 21293 11732 21327 12108
rect 21411 11732 21445 12108
rect 21529 11732 21563 12108
rect 21616 11732 21650 11908
rect 21734 11732 21768 11908
rect 21852 11732 21886 11908
rect 21970 11732 22004 11908
rect 22552 11732 22586 11908
rect 22670 11732 22704 11908
rect 22788 11732 22822 11908
rect 22906 11732 22940 11908
rect 23025 11732 23059 12108
rect 23143 11732 23177 12108
rect 23261 11732 23295 12108
rect 23379 11732 23413 12108
rect 23498 11732 23532 12108
rect 23616 11732 23650 12108
rect 23734 11732 23768 12108
rect 23852 11732 23886 12108
rect 23970 11732 24004 12108
rect 24088 11732 24122 12108
rect 24206 11732 24240 12108
rect 24319 11732 24353 12108
rect 24437 11732 24471 12108
rect 24555 11732 24589 12108
rect 24673 11732 24707 12108
rect 30659 12235 31035 12269
rect 29966 12178 30342 12212
rect 31306 12293 31340 12327
rect 31391 12235 31767 12269
rect 31933 12343 31955 12393
rect 31955 12343 31975 12393
rect 30659 12117 31035 12151
rect 31391 12117 31767 12151
rect 29966 12060 30342 12094
rect 30659 11999 31035 12033
rect 24760 11732 24794 11908
rect 24878 11732 24912 11908
rect 24996 11732 25030 11908
rect 29966 11942 30342 11976
rect 25114 11732 25148 11908
rect 30166 11813 30342 11847
rect 30511 11751 30565 11761
rect 30166 11695 30342 11729
rect 30511 11717 30521 11751
rect 30521 11717 30555 11751
rect 30555 11717 30565 11751
rect 30511 11707 30565 11717
rect 30166 11577 30342 11611
rect 676 11528 710 11562
rect 3820 11528 3854 11562
rect 1986 11487 2020 11521
rect 6952 11524 6986 11558
rect 5130 11487 5164 11521
rect 10096 11524 10130 11558
rect 8262 11483 8296 11517
rect 13298 11528 13332 11562
rect 11406 11483 11440 11517
rect 16442 11528 16476 11562
rect 14608 11487 14642 11521
rect 19574 11524 19608 11558
rect 17752 11487 17786 11521
rect 22718 11524 22752 11558
rect 20884 11483 20918 11517
rect 31223 12029 31257 12063
rect 31291 11739 31325 11773
rect 31391 11711 31567 11745
rect 31391 11593 31567 11627
rect 24028 11483 24062 11517
rect 30166 11459 30342 11493
rect 1856 11367 1914 11422
rect 1914 11367 1916 11422
rect 2941 11366 2943 11421
rect 2943 11366 3001 11421
rect 5000 11367 5058 11422
rect 5058 11367 5060 11422
rect 6085 11366 6087 11421
rect 6087 11366 6145 11421
rect 8132 11363 8190 11418
rect 8190 11363 8192 11418
rect 9217 11362 9219 11417
rect 9219 11362 9277 11417
rect 9472 11358 9521 11418
rect 11276 11363 11334 11418
rect 11334 11363 11336 11418
rect 12361 11362 12363 11417
rect 12363 11362 12421 11417
rect 14478 11367 14536 11422
rect 14536 11367 14538 11422
rect 15563 11366 15565 11421
rect 15565 11366 15623 11421
rect 17622 11367 17680 11422
rect 17680 11367 17682 11422
rect 18707 11366 18709 11421
rect 18709 11366 18767 11421
rect 20754 11363 20812 11418
rect 20812 11363 20814 11418
rect 21839 11362 21841 11417
rect 21841 11362 21899 11417
rect 23898 11363 23956 11418
rect 23956 11363 23958 11418
rect 31063 11427 31165 11529
rect 24983 11362 24985 11417
rect 24985 11362 25043 11417
rect 1632 11257 1666 11291
rect 3196 11246 3245 11306
rect 4776 11257 4810 11291
rect 6340 11246 6389 11306
rect 7908 11253 7942 11287
rect 9472 11242 9521 11302
rect 11052 11253 11086 11287
rect 12616 11242 12665 11302
rect 14254 11257 14288 11291
rect 15818 11246 15867 11306
rect 17398 11257 17432 11291
rect 18962 11246 19011 11306
rect 20530 11253 20564 11287
rect 22094 11242 22143 11302
rect 23674 11253 23708 11287
rect 25238 11242 25287 11302
rect 1974 11082 2032 11137
rect 2032 11082 2034 11137
rect 3196 11078 3245 11138
rect 5118 11082 5176 11137
rect 5176 11082 5178 11137
rect 6340 11078 6389 11138
rect 8250 11078 8308 11133
rect 8308 11078 8310 11133
rect 9472 11074 9521 11134
rect 11394 11078 11452 11133
rect 11452 11078 11454 11133
rect 12616 11074 12665 11134
rect 14596 11082 14654 11137
rect 14654 11082 14656 11137
rect 15818 11078 15867 11138
rect 17740 11082 17798 11137
rect 17798 11082 17800 11137
rect 18962 11078 19011 11138
rect 20872 11078 20930 11133
rect 20930 11078 20932 11133
rect 22094 11074 22143 11134
rect 24016 11078 24074 11133
rect 24074 11078 24076 11133
rect 25238 11074 25287 11134
rect 30164 11066 30340 11100
rect 30699 11077 30759 11093
rect 1751 10867 1785 10901
rect 4895 10867 4929 10901
rect 8027 10863 8061 10897
rect 11171 10863 11205 10897
rect 14373 10867 14407 10901
rect 17517 10867 17551 10901
rect 20649 10863 20683 10897
rect 23793 10863 23827 10897
rect 30699 11043 30713 11077
rect 30713 11043 30747 11077
rect 30747 11043 30759 11077
rect 30699 11027 30759 11043
rect 30164 10948 30340 10982
rect 31389 10941 31565 10975
rect 30164 10830 30340 10864
rect 1378 10603 1412 10779
rect 1496 10603 1530 10779
rect 1574 10403 1608 10779
rect 1692 10403 1726 10779
rect 1810 10403 1844 10779
rect 1928 10403 1962 10779
rect 2046 10403 2080 10779
rect 2120 10603 2154 10779
rect 2238 10603 2272 10779
rect 4522 10603 4556 10779
rect 4640 10603 4674 10779
rect 4718 10403 4752 10779
rect 4836 10403 4870 10779
rect 4954 10403 4988 10779
rect 5072 10403 5106 10779
rect 5190 10403 5224 10779
rect 5264 10603 5298 10779
rect 5382 10603 5416 10779
rect 7654 10599 7688 10775
rect 7772 10599 7806 10775
rect 7850 10399 7884 10775
rect 7968 10399 8002 10775
rect 8086 10399 8120 10775
rect 8204 10399 8238 10775
rect 8322 10399 8356 10775
rect 8396 10599 8430 10775
rect 8514 10599 8548 10775
rect 10798 10599 10832 10775
rect 10916 10599 10950 10775
rect 10994 10399 11028 10775
rect 11112 10399 11146 10775
rect 11230 10399 11264 10775
rect 11348 10399 11382 10775
rect 11466 10399 11500 10775
rect 11540 10599 11574 10775
rect 11658 10599 11692 10775
rect 14000 10603 14034 10779
rect 14118 10603 14152 10779
rect 14196 10403 14230 10779
rect 14314 10403 14348 10779
rect 14432 10403 14466 10779
rect 14550 10403 14584 10779
rect 14668 10403 14702 10779
rect 14742 10603 14776 10779
rect 14860 10603 14894 10779
rect 17144 10603 17178 10779
rect 17262 10603 17296 10779
rect 17340 10403 17374 10779
rect 17458 10403 17492 10779
rect 17576 10403 17610 10779
rect 17694 10403 17728 10779
rect 17812 10403 17846 10779
rect 17886 10603 17920 10779
rect 31288 10794 31322 10828
rect 31389 10823 31565 10857
rect 18004 10603 18038 10779
rect 20276 10599 20310 10775
rect 20394 10599 20428 10775
rect 20472 10399 20506 10775
rect 20590 10399 20624 10775
rect 20708 10399 20742 10775
rect 20826 10399 20860 10775
rect 20944 10399 20978 10775
rect 21018 10599 21052 10775
rect 21136 10599 21170 10775
rect 23420 10599 23454 10775
rect 23538 10599 23572 10775
rect 23616 10399 23650 10775
rect 23734 10399 23768 10775
rect 23852 10399 23886 10775
rect 23970 10399 24004 10775
rect 24088 10399 24122 10775
rect 24162 10599 24196 10775
rect 24280 10599 24314 10775
rect 30164 10712 30340 10746
rect 30657 10639 31033 10673
rect 29964 10582 30340 10616
rect 31221 10609 31255 10643
rect 30657 10521 31033 10555
rect 31389 10521 31765 10555
rect 29964 10464 30340 10498
rect 30657 10403 31033 10437
rect 29964 10346 30340 10380
rect 31389 10403 31765 10437
rect 31305 10343 31339 10377
rect 1809 10268 1843 10302
rect 4953 10268 4987 10302
rect 8085 10264 8119 10298
rect 11229 10264 11263 10298
rect 14431 10268 14465 10302
rect 17575 10268 17609 10302
rect 20707 10264 20741 10298
rect 23851 10264 23885 10298
rect 30657 10285 31033 10319
rect 31389 10285 31765 10319
rect 29709 10225 29737 10263
rect 29737 10225 29747 10263
rect 1782 10136 1840 10150
rect 1782 10104 1840 10136
rect 4926 10136 4984 10150
rect 4926 10104 4984 10136
rect 8058 10132 8116 10146
rect 8058 10100 8116 10132
rect 11202 10132 11260 10146
rect 11202 10100 11260 10132
rect 14404 10136 14462 10150
rect 14404 10104 14462 10136
rect 17548 10136 17606 10150
rect 17548 10104 17606 10136
rect 20680 10132 20738 10146
rect 20680 10100 20738 10132
rect 29964 10228 30340 10262
rect 23824 10132 23882 10146
rect 23824 10100 23882 10132
rect 30657 10167 31033 10201
rect 29964 10110 30340 10144
rect 31304 10225 31338 10259
rect 31389 10167 31765 10201
rect 31931 10275 31953 10325
rect 31953 10275 31973 10325
rect 30657 10049 31033 10083
rect 31389 10049 31765 10083
rect 29964 9992 30340 10026
rect 30657 9931 31033 9965
rect 29964 9874 30340 9908
rect 30164 9745 30340 9779
rect 30509 9683 30563 9693
rect 1792 9576 1864 9630
rect 4936 9576 5008 9630
rect 8068 9572 8140 9626
rect 11212 9572 11284 9626
rect 14414 9576 14486 9630
rect 17558 9576 17630 9630
rect 20690 9572 20762 9626
rect 23834 9572 23906 9626
rect 30164 9627 30340 9661
rect 30509 9649 30519 9683
rect 30519 9649 30553 9683
rect 30553 9649 30563 9683
rect 30509 9639 30563 9649
rect 30164 9509 30340 9543
rect 520 9004 554 9180
rect 638 9004 672 9180
rect 756 9004 790 9180
rect 874 9004 908 9180
rect 993 9004 1027 9380
rect 1111 9004 1145 9380
rect 1229 9004 1263 9380
rect 1347 9004 1381 9380
rect 1466 9004 1500 9380
rect 1584 9004 1618 9380
rect 1702 9004 1736 9380
rect 1820 9004 1854 9380
rect 1938 9004 1972 9380
rect 2056 9004 2090 9380
rect 2174 9004 2208 9380
rect 2287 9004 2321 9380
rect 2405 9004 2439 9380
rect 2523 9004 2557 9380
rect 2641 9004 2675 9380
rect 2728 9004 2762 9180
rect 2846 9004 2880 9180
rect 2964 9004 2998 9180
rect 3082 9004 3116 9180
rect 3664 9004 3698 9180
rect 3782 9004 3816 9180
rect 3900 9004 3934 9180
rect 4018 9004 4052 9180
rect 4137 9004 4171 9380
rect 4255 9004 4289 9380
rect 4373 9004 4407 9380
rect 4491 9004 4525 9380
rect 4610 9004 4644 9380
rect 4728 9004 4762 9380
rect 4846 9004 4880 9380
rect 4964 9004 4998 9380
rect 5082 9004 5116 9380
rect 5200 9004 5234 9380
rect 5318 9004 5352 9380
rect 5431 9004 5465 9380
rect 5549 9004 5583 9380
rect 5667 9004 5701 9380
rect 5785 9004 5819 9380
rect 5872 9004 5906 9180
rect 5990 9004 6024 9180
rect 6108 9004 6142 9180
rect 6226 9004 6260 9180
rect 6796 9000 6830 9176
rect 6914 9000 6948 9176
rect 7032 9000 7066 9176
rect 7150 9000 7184 9176
rect 7269 9000 7303 9376
rect 7387 9000 7421 9376
rect 7505 9000 7539 9376
rect 7623 9000 7657 9376
rect 7742 9000 7776 9376
rect 7860 9000 7894 9376
rect 7978 9000 8012 9376
rect 8096 9000 8130 9376
rect 8214 9000 8248 9376
rect 8332 9000 8366 9376
rect 8450 9000 8484 9376
rect 8563 9000 8597 9376
rect 8681 9000 8715 9376
rect 8799 9000 8833 9376
rect 8917 9000 8951 9376
rect 9004 9000 9038 9176
rect 9122 9000 9156 9176
rect 9240 9000 9274 9176
rect 9358 9000 9392 9176
rect 9940 9000 9974 9176
rect 10058 9000 10092 9176
rect 10176 9000 10210 9176
rect 10294 9000 10328 9176
rect 10413 9000 10447 9376
rect 10531 9000 10565 9376
rect 10649 9000 10683 9376
rect 10767 9000 10801 9376
rect 10886 9000 10920 9376
rect 11004 9000 11038 9376
rect 11122 9000 11156 9376
rect 11240 9000 11274 9376
rect 11358 9000 11392 9376
rect 11476 9000 11510 9376
rect 11594 9000 11628 9376
rect 11707 9000 11741 9376
rect 11825 9000 11859 9376
rect 11943 9000 11977 9376
rect 12061 9000 12095 9376
rect 12148 9000 12182 9176
rect 12266 9000 12300 9176
rect 12384 9000 12418 9176
rect 12502 9000 12536 9176
rect 13142 9004 13176 9180
rect 13260 9004 13294 9180
rect 13378 9004 13412 9180
rect 13496 9004 13530 9180
rect 13615 9004 13649 9380
rect 13733 9004 13767 9380
rect 13851 9004 13885 9380
rect 13969 9004 14003 9380
rect 14088 9004 14122 9380
rect 14206 9004 14240 9380
rect 14324 9004 14358 9380
rect 14442 9004 14476 9380
rect 14560 9004 14594 9380
rect 14678 9004 14712 9380
rect 14796 9004 14830 9380
rect 14909 9004 14943 9380
rect 15027 9004 15061 9380
rect 15145 9004 15179 9380
rect 15263 9004 15297 9380
rect 15350 9004 15384 9180
rect 15468 9004 15502 9180
rect 15586 9004 15620 9180
rect 15704 9004 15738 9180
rect 16286 9004 16320 9180
rect 16404 9004 16438 9180
rect 16522 9004 16556 9180
rect 16640 9004 16674 9180
rect 16759 9004 16793 9380
rect 16877 9004 16911 9380
rect 16995 9004 17029 9380
rect 17113 9004 17147 9380
rect 17232 9004 17266 9380
rect 17350 9004 17384 9380
rect 17468 9004 17502 9380
rect 17586 9004 17620 9380
rect 17704 9004 17738 9380
rect 17822 9004 17856 9380
rect 17940 9004 17974 9380
rect 18053 9004 18087 9380
rect 18171 9004 18205 9380
rect 18289 9004 18323 9380
rect 18407 9004 18441 9380
rect 18494 9004 18528 9180
rect 18612 9004 18646 9180
rect 18730 9004 18764 9180
rect 18848 9004 18882 9180
rect 19418 9000 19452 9176
rect 19536 9000 19570 9176
rect 19654 9000 19688 9176
rect 19772 9000 19806 9176
rect 19891 9000 19925 9376
rect 20009 9000 20043 9376
rect 20127 9000 20161 9376
rect 20245 9000 20279 9376
rect 20364 9000 20398 9376
rect 20482 9000 20516 9376
rect 20600 9000 20634 9376
rect 20718 9000 20752 9376
rect 20836 9000 20870 9376
rect 20954 9000 20988 9376
rect 21072 9000 21106 9376
rect 21185 9000 21219 9376
rect 21303 9000 21337 9376
rect 21421 9000 21455 9376
rect 21539 9000 21573 9376
rect 21626 9000 21660 9176
rect 21744 9000 21778 9176
rect 21862 9000 21896 9176
rect 21980 9000 22014 9176
rect 22562 9000 22596 9176
rect 22680 9000 22714 9176
rect 22798 9000 22832 9176
rect 22916 9000 22950 9176
rect 23035 9000 23069 9376
rect 23153 9000 23187 9376
rect 23271 9000 23305 9376
rect 23389 9000 23423 9376
rect 23508 9000 23542 9376
rect 23626 9000 23660 9376
rect 23744 9000 23778 9376
rect 23862 9000 23896 9376
rect 23980 9000 24014 9376
rect 24098 9000 24132 9376
rect 31221 9961 31255 9995
rect 31289 9671 31323 9705
rect 31389 9643 31565 9677
rect 31389 9525 31565 9559
rect 24216 9000 24250 9376
rect 24329 9000 24363 9376
rect 24447 9000 24481 9376
rect 24565 9000 24599 9376
rect 30164 9391 30340 9425
rect 24683 9000 24717 9376
rect 31061 9359 31163 9461
rect 24770 9000 24804 9176
rect 24888 9000 24922 9176
rect 25006 9000 25040 9176
rect 25124 9000 25158 9176
rect 30166 8997 30342 9031
rect 30701 9008 30761 9024
rect 686 8796 720 8830
rect 3830 8796 3864 8830
rect 1996 8755 2030 8789
rect 6962 8792 6996 8826
rect 5140 8755 5174 8789
rect 10106 8792 10140 8826
rect 8272 8751 8306 8785
rect 13308 8796 13342 8830
rect 11416 8751 11450 8785
rect 16452 8796 16486 8830
rect 14618 8755 14652 8789
rect 19584 8792 19618 8826
rect 17762 8755 17796 8789
rect 22728 8792 22762 8826
rect 20894 8751 20928 8785
rect 24038 8751 24072 8785
rect 30701 8974 30715 9008
rect 30715 8974 30749 9008
rect 30749 8974 30761 9008
rect 30701 8958 30761 8974
rect 30166 8879 30342 8913
rect 31391 8872 31567 8906
rect 30166 8761 30342 8795
rect 31290 8725 31324 8759
rect 31391 8754 31567 8788
rect 1866 8635 1924 8690
rect 1924 8635 1926 8690
rect 2951 8634 2953 8689
rect 2953 8634 3011 8689
rect 3206 8630 3255 8690
rect 5010 8635 5068 8690
rect 5068 8635 5070 8690
rect 6095 8634 6097 8689
rect 6097 8634 6155 8689
rect 6350 8630 6399 8690
rect 8142 8631 8200 8686
rect 8200 8631 8202 8686
rect 9227 8630 9229 8685
rect 9229 8630 9287 8685
rect 9482 8626 9531 8686
rect 11286 8631 11344 8686
rect 11344 8631 11346 8686
rect 12371 8630 12373 8685
rect 12373 8630 12431 8685
rect 12626 8626 12675 8686
rect 14488 8635 14546 8690
rect 14546 8635 14548 8690
rect 15573 8634 15575 8689
rect 15575 8634 15633 8689
rect 15828 8630 15877 8690
rect 17632 8635 17690 8690
rect 17690 8635 17692 8690
rect 18717 8634 18719 8689
rect 18719 8634 18777 8689
rect 18972 8630 19021 8690
rect 20764 8631 20822 8686
rect 20822 8631 20824 8686
rect 21849 8630 21851 8685
rect 21851 8630 21909 8685
rect 22104 8626 22153 8686
rect 23908 8631 23966 8686
rect 23966 8631 23968 8686
rect 24993 8630 24995 8685
rect 24995 8630 25053 8685
rect 25248 8626 25297 8686
rect 30166 8643 30342 8677
rect 1642 8525 1676 8559
rect 3206 8514 3255 8574
rect 1984 8350 2042 8405
rect 2042 8350 2044 8405
rect 3206 8346 3255 8406
rect 1761 8135 1795 8169
rect 1388 7871 1422 8047
rect 1506 7871 1540 8047
rect 1584 7671 1618 8047
rect 1702 7671 1736 8047
rect 1820 7671 1854 8047
rect 1938 7671 1972 8047
rect 2056 7671 2090 8047
rect 2130 7871 2164 8047
rect 2248 7871 2282 8047
rect 1819 7536 1853 7570
rect 1792 7404 1850 7418
rect 1792 7372 1850 7404
rect 4786 8525 4820 8559
rect 6350 8514 6399 8574
rect 5128 8350 5186 8405
rect 5186 8350 5188 8405
rect 6350 8346 6399 8406
rect 4905 8135 4939 8169
rect 4532 7871 4566 8047
rect 4650 7871 4684 8047
rect 4728 7671 4762 8047
rect 4846 7671 4880 8047
rect 4964 7671 4998 8047
rect 5082 7671 5116 8047
rect 5200 7671 5234 8047
rect 5274 7871 5308 8047
rect 5392 7871 5426 8047
rect 4963 7536 4997 7570
rect 4936 7404 4994 7418
rect 4936 7372 4994 7404
rect 7918 8521 7952 8555
rect 9482 8510 9531 8570
rect 8260 8346 8318 8401
rect 8318 8346 8320 8401
rect 9482 8342 9531 8402
rect 8037 8131 8071 8165
rect 7664 7867 7698 8043
rect 7782 7867 7816 8043
rect 7860 7667 7894 8043
rect 7978 7667 8012 8043
rect 8096 7667 8130 8043
rect 8214 7667 8248 8043
rect 8332 7667 8366 8043
rect 8406 7867 8440 8043
rect 8524 7867 8558 8043
rect 8095 7532 8129 7566
rect 8068 7400 8126 7414
rect 8068 7368 8126 7400
rect 11062 8521 11096 8555
rect 12626 8510 12675 8570
rect 14264 8525 14298 8559
rect 15828 8514 15877 8574
rect 11404 8346 11462 8401
rect 11462 8346 11464 8401
rect 12626 8342 12675 8402
rect 11181 8131 11215 8165
rect 10808 7867 10842 8043
rect 10926 7867 10960 8043
rect 11004 7667 11038 8043
rect 11122 7667 11156 8043
rect 11240 7667 11274 8043
rect 11358 7667 11392 8043
rect 11476 7667 11510 8043
rect 11550 7867 11584 8043
rect 11668 7867 11702 8043
rect 11239 7532 11273 7566
rect 11212 7400 11270 7414
rect 11212 7368 11270 7400
rect 14606 8350 14664 8405
rect 14664 8350 14666 8405
rect 15828 8346 15877 8406
rect 14383 8135 14417 8169
rect 14010 7871 14044 8047
rect 14128 7871 14162 8047
rect 14206 7671 14240 8047
rect 14324 7671 14358 8047
rect 14442 7671 14476 8047
rect 14560 7671 14594 8047
rect 14678 7671 14712 8047
rect 14752 7871 14786 8047
rect 14870 7871 14904 8047
rect 14441 7536 14475 7570
rect 14414 7404 14472 7418
rect 14414 7372 14472 7404
rect 3277 6695 3373 6731
rect 4015 6695 4111 6731
rect 4753 6695 4849 6731
rect 5491 6695 5587 6731
rect 6231 6695 6327 6731
rect 6973 6695 7069 6731
rect 7711 6695 7807 6731
rect 8449 6697 8545 6733
rect 3129 6369 3163 6545
rect 3247 6369 3281 6545
rect 3365 6369 3399 6545
rect 3483 6369 3517 6545
rect 3867 6369 3901 6545
rect 3985 6369 4019 6545
rect 4103 6369 4137 6545
rect 4221 6369 4255 6545
rect 4605 6369 4639 6545
rect 4723 6369 4757 6545
rect 4841 6369 4875 6545
rect 4959 6369 4993 6545
rect 5343 6369 5377 6545
rect 5461 6369 5495 6545
rect 5579 6369 5613 6545
rect 5697 6369 5731 6545
rect 6083 6369 6117 6545
rect 6201 6369 6235 6545
rect 6319 6369 6353 6545
rect 6437 6369 6471 6545
rect 6825 6371 6859 6547
rect 6943 6371 6977 6547
rect 7061 6371 7095 6547
rect 7179 6371 7213 6547
rect 7563 6375 7597 6551
rect 7681 6375 7715 6551
rect 7799 6375 7833 6551
rect 7917 6375 7951 6551
rect 8301 6371 8335 6547
rect 8419 6371 8453 6547
rect 8537 6371 8571 6547
rect 8655 6371 8689 6547
rect 3307 6229 3341 6263
rect 3487 6223 3525 6269
rect 4045 6229 4079 6263
rect 4226 6223 4262 6269
rect 4783 6229 4817 6263
rect 5521 6229 5555 6263
rect 6261 6229 6295 6263
rect 7003 6229 7037 6263
rect 7741 6229 7775 6263
rect 8479 6231 8513 6265
rect 3247 5987 3281 6163
rect 3365 5987 3399 6163
rect 3345 5809 3423 5863
rect 3985 5987 4019 6163
rect 4103 5987 4137 6163
rect 4083 5809 4161 5863
rect -1976 3361 -1883 3398
rect 151 3354 205 3398
rect 4723 5983 4757 6159
rect 4841 5983 4875 6159
rect 4821 5809 4899 5863
rect 5461 5983 5495 6159
rect 5579 5983 5613 6159
rect 5559 5809 5637 5863
rect 6201 5983 6235 6159
rect 6319 5983 6353 6159
rect 6299 5809 6377 5863
rect 6943 5983 6977 6159
rect 7061 5983 7095 6159
rect 7041 5809 7119 5863
rect 7681 5987 7715 6163
rect 7799 5987 7833 6163
rect 7779 5809 7857 5863
rect 8419 5985 8453 6161
rect 8537 5985 8571 6161
rect 8517 5811 8595 5865
rect 10067 6662 10105 6690
rect 10067 6652 10105 6662
rect 9233 6059 9267 6235
rect 9351 6059 9385 6235
rect 9469 6059 9503 6235
rect 9587 6059 9621 6235
rect 9716 6059 9750 6435
rect 9834 6059 9868 6435
rect 9952 6059 9986 6435
rect 10070 6059 10104 6435
rect 10188 6059 10222 6435
rect 10306 6059 10340 6435
rect 10424 6059 10458 6435
rect 10554 6059 10588 6235
rect 10672 6059 10706 6235
rect 10790 6059 10824 6235
rect 10908 6059 10942 6235
rect 9481 5880 9535 5890
rect 9481 5846 9491 5880
rect 9491 5846 9525 5880
rect 9525 5846 9535 5880
rect 9481 5836 9535 5846
rect 9773 5366 9807 5742
rect 9891 5366 9925 5742
rect 9201 5236 9303 5338
rect 10009 5366 10043 5742
rect 10127 5366 10161 5742
rect 10245 5366 10279 5742
rect 10363 5366 10397 5742
rect 10481 5366 10515 5742
rect 10869 5686 10935 5700
rect 10869 5652 10885 5686
rect 10885 5652 10919 5686
rect 10919 5652 10935 5686
rect 10869 5640 10935 5652
rect 12135 6660 12173 6688
rect 12135 6650 12173 6660
rect 11301 6057 11335 6233
rect 11419 6057 11453 6233
rect 11537 6057 11571 6233
rect 11655 6057 11689 6233
rect 11784 6057 11818 6433
rect 11902 6057 11936 6433
rect 12020 6057 12054 6433
rect 12138 6057 12172 6433
rect 12256 6057 12290 6433
rect 12374 6057 12408 6433
rect 12492 6057 12526 6433
rect 12622 6057 12656 6233
rect 12740 6057 12774 6233
rect 12858 6057 12892 6233
rect 12976 6057 13010 6233
rect 11549 5878 11603 5888
rect 11549 5844 11559 5878
rect 11559 5844 11593 5878
rect 11593 5844 11603 5878
rect 11549 5834 11603 5844
rect 11841 5364 11875 5740
rect 11959 5364 11993 5740
rect 9803 5144 9837 5178
rect 9513 5076 9547 5110
rect 10067 5061 10101 5095
rect 10185 5060 10219 5094
rect 11269 5234 11371 5336
rect 12077 5364 12111 5740
rect 12195 5364 12229 5740
rect 12313 5364 12347 5740
rect 12431 5364 12465 5740
rect 12549 5364 12583 5740
rect 12937 5684 13003 5698
rect 12937 5650 12953 5684
rect 12953 5650 12987 5684
rect 12987 5650 13003 5684
rect 12937 5638 13003 5650
rect 14204 6662 14242 6690
rect 14204 6652 14242 6662
rect 13370 6059 13404 6235
rect 13488 6059 13522 6235
rect 13606 6059 13640 6235
rect 13724 6059 13758 6235
rect 13853 6059 13887 6435
rect 13971 6059 14005 6435
rect 14089 6059 14123 6435
rect 14207 6059 14241 6435
rect 14325 6059 14359 6435
rect 14443 6059 14477 6435
rect 14561 6059 14595 6435
rect 14691 6059 14725 6235
rect 14809 6059 14843 6235
rect 14927 6059 14961 6235
rect 15045 6059 15079 6235
rect 13618 5880 13672 5890
rect 13618 5846 13628 5880
rect 13628 5846 13662 5880
rect 13662 5846 13672 5880
rect 13618 5836 13672 5846
rect 13910 5366 13944 5742
rect 14028 5366 14062 5742
rect 10451 5144 10485 5178
rect 11871 5142 11905 5176
rect 10636 5077 10670 5111
rect 11581 5074 11615 5108
rect 12135 5059 12169 5093
rect 12253 5058 12287 5092
rect 9367 4834 9401 5010
rect 9485 4834 9519 5010
rect 9891 4634 9925 5010
rect 10009 4634 10043 5010
rect 10127 4634 10161 5010
rect 10245 4634 10279 5010
rect 10363 4634 10397 5010
rect 10665 4834 10699 5010
rect 13338 5236 13440 5338
rect 14146 5366 14180 5742
rect 14264 5366 14298 5742
rect 14382 5366 14416 5742
rect 14500 5366 14534 5742
rect 14618 5366 14652 5742
rect 15006 5686 15072 5700
rect 15006 5652 15022 5686
rect 15022 5652 15056 5686
rect 15056 5652 15072 5686
rect 15006 5640 15072 5652
rect 17408 8525 17442 8559
rect 18972 8514 19021 8574
rect 17750 8350 17808 8405
rect 17808 8350 17810 8405
rect 18972 8346 19021 8406
rect 17527 8135 17561 8169
rect 20540 8521 20574 8555
rect 22104 8510 22153 8570
rect 20882 8346 20940 8401
rect 20940 8346 20942 8401
rect 22104 8342 22153 8402
rect 20659 8131 20693 8165
rect 17154 7871 17188 8047
rect 17272 7871 17306 8047
rect 17350 7671 17384 8047
rect 17468 7671 17502 8047
rect 17586 7671 17620 8047
rect 17704 7671 17738 8047
rect 17822 7671 17856 8047
rect 17896 7871 17930 8047
rect 18014 7871 18048 8047
rect 17585 7536 17619 7570
rect 17558 7404 17616 7418
rect 17558 7372 17616 7404
rect 16272 6660 16310 6688
rect 16272 6650 16310 6660
rect 15438 6057 15472 6233
rect 15556 6057 15590 6233
rect 15674 6057 15708 6233
rect 15792 6057 15826 6233
rect 15921 6057 15955 6433
rect 16039 6057 16073 6433
rect 16157 6057 16191 6433
rect 16275 6057 16309 6433
rect 16393 6057 16427 6433
rect 16511 6057 16545 6433
rect 16629 6057 16663 6433
rect 16759 6057 16793 6233
rect 16877 6057 16911 6233
rect 16995 6057 17029 6233
rect 17113 6057 17147 6233
rect 15686 5878 15740 5888
rect 15686 5844 15696 5878
rect 15696 5844 15730 5878
rect 15730 5844 15740 5878
rect 15686 5834 15740 5844
rect 15978 5364 16012 5740
rect 16096 5364 16130 5740
rect 12519 5142 12553 5176
rect 13940 5144 13974 5178
rect 12704 5075 12738 5109
rect 13650 5076 13684 5110
rect 14204 5061 14238 5095
rect 14322 5060 14356 5094
rect 15406 5234 15508 5336
rect 16214 5364 16248 5740
rect 16332 5364 16366 5740
rect 16450 5364 16484 5740
rect 16568 5364 16602 5740
rect 16686 5364 16720 5740
rect 17074 5684 17140 5698
rect 17074 5650 17090 5684
rect 17090 5650 17124 5684
rect 17124 5650 17140 5684
rect 17074 5638 17140 5650
rect 18341 6660 18379 6688
rect 18341 6650 18379 6660
rect 17507 6057 17541 6233
rect 17625 6057 17659 6233
rect 17743 6057 17777 6233
rect 17861 6057 17895 6233
rect 17990 6057 18024 6433
rect 18108 6057 18142 6433
rect 18226 6057 18260 6433
rect 18344 6057 18378 6433
rect 18462 6057 18496 6433
rect 18580 6057 18614 6433
rect 18698 6057 18732 6433
rect 18828 6057 18862 6233
rect 18946 6057 18980 6233
rect 19064 6057 19098 6233
rect 19182 6057 19216 6233
rect 17755 5878 17809 5888
rect 17755 5844 17765 5878
rect 17765 5844 17799 5878
rect 17799 5844 17809 5878
rect 17755 5834 17809 5844
rect 18047 5364 18081 5740
rect 18165 5364 18199 5740
rect 14588 5144 14622 5178
rect 16008 5142 16042 5176
rect 14773 5077 14807 5111
rect 15718 5074 15752 5108
rect 16272 5059 16306 5093
rect 16390 5058 16424 5092
rect 10783 4834 10817 5010
rect 11435 4832 11469 5008
rect 11553 4832 11587 5008
rect 11959 4632 11993 5008
rect 12077 4632 12111 5008
rect 12195 4632 12229 5008
rect 12313 4632 12347 5008
rect 12431 4632 12465 5008
rect 12733 4832 12767 5008
rect 12851 4832 12885 5008
rect 13504 4834 13538 5010
rect 13622 4834 13656 5010
rect 14028 4634 14062 5010
rect 14146 4634 14180 5010
rect 14264 4634 14298 5010
rect 14382 4634 14416 5010
rect 14500 4634 14534 5010
rect 14802 4834 14836 5010
rect 17475 5234 17577 5336
rect 18283 5364 18317 5740
rect 18401 5364 18435 5740
rect 18519 5364 18553 5740
rect 18637 5364 18671 5740
rect 18755 5364 18789 5740
rect 19143 5684 19209 5698
rect 19143 5650 19159 5684
rect 19159 5650 19193 5684
rect 19193 5650 19209 5684
rect 19143 5638 19209 5650
rect 20286 7867 20320 8043
rect 20404 7867 20438 8043
rect 20482 7667 20516 8043
rect 20600 7667 20634 8043
rect 20718 7667 20752 8043
rect 20836 7667 20870 8043
rect 20954 7667 20988 8043
rect 21028 7867 21062 8043
rect 21146 7867 21180 8043
rect 20717 7532 20751 7566
rect 20690 7400 20748 7414
rect 20690 7368 20748 7400
rect 23684 8521 23718 8555
rect 30659 8570 31035 8604
rect 25248 8510 25297 8570
rect 29966 8513 30342 8547
rect 31223 8540 31257 8574
rect 24026 8346 24084 8401
rect 24084 8346 24086 8401
rect 25248 8342 25297 8402
rect 23803 8131 23837 8165
rect 23430 7867 23464 8043
rect 23548 7867 23582 8043
rect 23626 7667 23660 8043
rect 23744 7667 23778 8043
rect 23862 7667 23896 8043
rect 23980 7667 24014 8043
rect 24098 7667 24132 8043
rect 24172 7867 24206 8043
rect 24290 7867 24324 8043
rect 23861 7532 23895 7566
rect 23834 7400 23892 7414
rect 23834 7368 23892 7400
rect 30659 8452 31035 8486
rect 31391 8452 31767 8486
rect 29966 8395 30342 8429
rect 30659 8334 31035 8368
rect 29966 8277 30342 8311
rect 31391 8334 31767 8368
rect 31307 8274 31341 8308
rect 30659 8216 31035 8250
rect 31391 8216 31767 8250
rect 29711 8156 29739 8194
rect 29739 8156 29749 8194
rect 29966 8159 30342 8193
rect 30659 8098 31035 8132
rect 29966 8041 30342 8075
rect 31306 8156 31340 8190
rect 31391 8098 31767 8132
rect 31933 8206 31955 8256
rect 31955 8206 31975 8256
rect 30659 7980 31035 8014
rect 31391 7980 31767 8014
rect 29966 7923 30342 7957
rect 30659 7862 31035 7896
rect 29966 7805 30342 7839
rect 30166 7676 30342 7710
rect 30511 7614 30565 7624
rect 30166 7558 30342 7592
rect 30511 7580 30521 7614
rect 30521 7580 30555 7614
rect 30555 7580 30565 7614
rect 30511 7570 30565 7580
rect 30166 7440 30342 7474
rect 31223 7892 31257 7926
rect 31291 7602 31325 7636
rect 31391 7574 31567 7608
rect 31391 7456 31567 7490
rect 30166 7322 30342 7356
rect 31063 7290 31165 7392
rect 30164 6929 30340 6963
rect 30699 6940 30759 6956
rect 20409 6658 20447 6686
rect 20409 6648 20447 6658
rect 19575 6055 19609 6231
rect 19693 6055 19727 6231
rect 19811 6055 19845 6231
rect 19929 6055 19963 6231
rect 20058 6055 20092 6431
rect 20176 6055 20210 6431
rect 20294 6055 20328 6431
rect 20412 6055 20446 6431
rect 20530 6055 20564 6431
rect 20648 6055 20682 6431
rect 20766 6055 20800 6431
rect 20896 6055 20930 6231
rect 21014 6055 21048 6231
rect 21132 6055 21166 6231
rect 21250 6055 21284 6231
rect 19823 5876 19877 5886
rect 19823 5842 19833 5876
rect 19833 5842 19867 5876
rect 19867 5842 19877 5876
rect 19823 5832 19877 5842
rect 20115 5362 20149 5738
rect 20233 5362 20267 5738
rect 16656 5142 16690 5176
rect 18077 5142 18111 5176
rect 16841 5075 16875 5109
rect 17787 5074 17821 5108
rect 18341 5059 18375 5093
rect 18459 5058 18493 5092
rect 19543 5232 19645 5334
rect 20351 5362 20385 5738
rect 20469 5362 20503 5738
rect 20587 5362 20621 5738
rect 20705 5362 20739 5738
rect 20823 5362 20857 5738
rect 21211 5682 21277 5696
rect 21211 5648 21227 5682
rect 21227 5648 21261 5682
rect 21261 5648 21277 5682
rect 21211 5636 21277 5648
rect 22478 6660 22516 6688
rect 22478 6650 22516 6660
rect 21644 6057 21678 6233
rect 21762 6057 21796 6233
rect 21880 6057 21914 6233
rect 21998 6057 22032 6233
rect 22127 6057 22161 6433
rect 22245 6057 22279 6433
rect 22363 6057 22397 6433
rect 22481 6057 22515 6433
rect 22599 6057 22633 6433
rect 22717 6057 22751 6433
rect 22835 6057 22869 6433
rect 22965 6057 22999 6233
rect 23083 6057 23117 6233
rect 23201 6057 23235 6233
rect 23319 6057 23353 6233
rect 21892 5878 21946 5888
rect 21892 5844 21902 5878
rect 21902 5844 21936 5878
rect 21936 5844 21946 5878
rect 21892 5834 21946 5844
rect 22184 5364 22218 5740
rect 22302 5364 22336 5740
rect 18725 5142 18759 5176
rect 20145 5140 20179 5174
rect 18910 5075 18944 5109
rect 19855 5072 19889 5106
rect 20409 5057 20443 5091
rect 20527 5056 20561 5090
rect 14920 4834 14954 5010
rect 15572 4832 15606 5008
rect 15690 4832 15724 5008
rect 16096 4632 16130 5008
rect 16214 4632 16248 5008
rect 16332 4632 16366 5008
rect 16450 4632 16484 5008
rect 16568 4632 16602 5008
rect 16870 4832 16904 5008
rect 16988 4832 17022 5008
rect 17641 4832 17675 5008
rect 17759 4832 17793 5008
rect 18165 4632 18199 5008
rect 18283 4632 18317 5008
rect 18401 4632 18435 5008
rect 18519 4632 18553 5008
rect 18637 4632 18671 5008
rect 18939 4832 18973 5008
rect 21612 5234 21714 5336
rect 22420 5364 22454 5740
rect 22538 5364 22572 5740
rect 22656 5364 22690 5740
rect 22774 5364 22808 5740
rect 22892 5364 22926 5740
rect 23280 5684 23346 5698
rect 23280 5650 23296 5684
rect 23296 5650 23330 5684
rect 23330 5650 23346 5684
rect 23280 5638 23346 5650
rect 30699 6906 30713 6940
rect 30713 6906 30747 6940
rect 30747 6906 30759 6940
rect 30699 6890 30759 6906
rect 30164 6811 30340 6845
rect 31389 6804 31565 6838
rect 24546 6658 24584 6686
rect 30164 6693 30340 6727
rect 24546 6648 24584 6658
rect 31288 6657 31322 6691
rect 31389 6686 31565 6720
rect 30164 6575 30340 6609
rect 30657 6502 31033 6536
rect 23712 6055 23746 6231
rect 23830 6055 23864 6231
rect 23948 6055 23982 6231
rect 24066 6055 24100 6231
rect 24195 6055 24229 6431
rect 24313 6055 24347 6431
rect 24431 6055 24465 6431
rect 24549 6055 24583 6431
rect 24667 6055 24701 6431
rect 24785 6055 24819 6431
rect 29964 6445 30340 6479
rect 31221 6472 31255 6506
rect 24903 6055 24937 6431
rect 30657 6384 31033 6418
rect 31389 6384 31765 6418
rect 29964 6327 30340 6361
rect 25033 6055 25067 6231
rect 25151 6055 25185 6231
rect 25269 6055 25303 6231
rect 30657 6266 31033 6300
rect 25387 6055 25421 6231
rect 29964 6209 30340 6243
rect 31389 6266 31765 6300
rect 31305 6206 31339 6240
rect 30657 6148 31033 6182
rect 31389 6148 31765 6182
rect 29709 6088 29737 6126
rect 29737 6088 29747 6126
rect 29964 6091 30340 6125
rect 30657 6030 31033 6064
rect 29964 5973 30340 6007
rect 31304 6088 31338 6122
rect 31389 6030 31765 6064
rect 31931 6138 31953 6188
rect 31953 6138 31973 6188
rect 30657 5912 31033 5946
rect 31389 5912 31765 5946
rect 23960 5876 24014 5886
rect 23960 5842 23970 5876
rect 23970 5842 24004 5876
rect 24004 5842 24014 5876
rect 29964 5855 30340 5889
rect 23960 5832 24014 5842
rect 30657 5794 31033 5828
rect 24252 5362 24286 5738
rect 24370 5362 24404 5738
rect 20793 5140 20827 5174
rect 22214 5142 22248 5176
rect 20978 5073 21012 5107
rect 21924 5074 21958 5108
rect 22478 5059 22512 5093
rect 22596 5058 22630 5092
rect 23680 5232 23782 5334
rect 24488 5362 24522 5738
rect 24606 5362 24640 5738
rect 24724 5362 24758 5738
rect 24842 5362 24876 5738
rect 24960 5362 24994 5738
rect 29964 5737 30340 5771
rect 25348 5682 25414 5696
rect 25348 5648 25364 5682
rect 25364 5648 25398 5682
rect 25398 5648 25414 5682
rect 25348 5636 25414 5648
rect 30164 5608 30340 5642
rect 22862 5142 22896 5176
rect 24282 5140 24316 5174
rect 23047 5075 23081 5109
rect 23992 5072 24026 5106
rect 24546 5057 24580 5091
rect 24664 5056 24698 5090
rect 19057 4832 19091 5008
rect 19709 4830 19743 5006
rect 19827 4830 19861 5006
rect 20233 4630 20267 5006
rect 20351 4630 20385 5006
rect 20469 4630 20503 5006
rect 20587 4630 20621 5006
rect 20705 4630 20739 5006
rect 21007 4830 21041 5006
rect 21125 4830 21159 5006
rect 21778 4832 21812 5008
rect 21896 4832 21930 5008
rect 22302 4632 22336 5008
rect 22420 4632 22454 5008
rect 22538 4632 22572 5008
rect 22656 4632 22690 5008
rect 22774 4632 22808 5008
rect 23076 4832 23110 5008
rect 24930 5140 24964 5174
rect 25115 5073 25149 5107
rect 23194 4832 23228 5008
rect 23846 4830 23880 5006
rect 23964 4830 23998 5006
rect 24370 4630 24404 5006
rect 24488 4630 24522 5006
rect 24606 4630 24640 5006
rect 24724 4630 24758 5006
rect 24842 4630 24876 5006
rect 25144 4830 25178 5006
rect 25262 4830 25296 5006
rect 10117 4446 10167 4468
rect 10117 4426 10167 4446
rect 12185 4444 12235 4466
rect 12185 4424 12235 4444
rect 14254 4446 14304 4468
rect 14254 4426 14304 4446
rect 16322 4444 16372 4466
rect 16322 4424 16372 4444
rect 18391 4444 18441 4466
rect 18391 4424 18441 4444
rect 20459 4442 20509 4464
rect 20459 4422 20509 4442
rect 22528 4444 22578 4466
rect 22528 4424 22578 4444
rect 24596 4442 24646 4464
rect 24596 4422 24646 4442
rect 30509 5546 30563 5556
rect 30164 5490 30340 5524
rect 30509 5512 30519 5546
rect 30519 5512 30553 5546
rect 30553 5512 30563 5546
rect 30509 5502 30563 5512
rect 30164 5372 30340 5406
rect 31221 5824 31255 5858
rect 31289 5534 31323 5568
rect 31389 5506 31565 5540
rect 31389 5388 31565 5422
rect 30164 5254 30340 5288
rect 31061 5222 31163 5324
rect 30164 4860 30340 4894
rect 30699 4871 30759 4887
rect 30699 4837 30713 4871
rect 30713 4837 30747 4871
rect 30747 4837 30759 4871
rect 30699 4821 30759 4837
rect 30164 4742 30340 4776
rect 31389 4735 31565 4769
rect 30164 4624 30340 4658
rect 31288 4588 31322 4622
rect 31389 4617 31565 4651
rect 30164 4506 30340 4540
rect 30657 4433 31033 4467
rect 29964 4376 30340 4410
rect 31221 4403 31255 4437
rect 30657 4315 31033 4349
rect 31389 4315 31765 4349
rect 29964 4258 30340 4292
rect 30657 4197 31033 4231
rect 29964 4140 30340 4174
rect 31389 4197 31765 4231
rect 31305 4137 31339 4171
rect 23350 4004 23401 4055
rect 30657 4079 31033 4113
rect 31389 4079 31765 4113
rect 29709 4019 29737 4057
rect 29737 4019 29747 4057
rect 21319 3896 21366 3950
rect 29964 4022 30340 4056
rect 19272 3793 19319 3847
rect 30657 3961 31033 3995
rect 29964 3904 30340 3938
rect 31304 4019 31338 4053
rect 31389 3961 31765 3995
rect 31931 4069 31953 4119
rect 31953 4069 31973 4119
rect 30657 3843 31033 3877
rect 31389 3843 31765 3877
rect 29964 3786 30340 3820
rect 17179 3686 17229 3737
rect 30657 3725 31033 3759
rect 29964 3668 30340 3702
rect 15107 3589 15158 3642
rect 30164 3539 30340 3573
rect 13011 3447 13055 3498
rect 30509 3477 30563 3487
rect 30164 3421 30340 3455
rect 30509 3443 30519 3477
rect 30519 3443 30553 3477
rect 30553 3443 30563 3477
rect 30509 3433 30563 3443
rect 10934 3349 10987 3403
rect 30164 3303 30340 3337
rect 31221 3755 31255 3789
rect 31289 3465 31323 3499
rect 31389 3437 31565 3471
rect 31389 3319 31565 3353
rect 30164 3185 30340 3219
rect -1506 3122 -1414 3158
rect 31061 3153 31163 3255
rect 150 3106 204 3150
rect -1246 3001 -1166 3044
rect 149 2990 203 3034
rect 32681 2938 32747 3000
rect -1030 2876 -952 2933
rect 149 2866 203 2910
rect 30162 2792 30338 2826
rect 30697 2803 30757 2819
rect 1512 2324 1584 2378
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 2656 1544 2690 1578
rect 1346 1503 1380 1537
rect 121 1378 170 1438
rect 4656 2324 4728 2378
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 5800 1544 5834 1578
rect 4490 1503 4524 1537
rect 7788 2328 7860 2382
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 8932 1548 8966 1582
rect 7622 1507 7656 1541
rect 365 1382 423 1437
rect 423 1382 425 1437
rect 1450 1383 1452 1438
rect 1452 1383 1510 1438
rect 3265 1378 3314 1438
rect 3509 1382 3567 1437
rect 3567 1382 3569 1437
rect 4594 1383 4596 1438
rect 4596 1383 4654 1438
rect 6397 1382 6446 1442
rect 10932 2328 11004 2382
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 12076 1548 12110 1582
rect 10766 1507 10800 1541
rect 6641 1386 6699 1441
rect 6699 1386 6701 1441
rect 7726 1387 7728 1442
rect 7728 1387 7786 1442
rect 9541 1382 9590 1442
rect 9785 1386 9843 1441
rect 9843 1386 9845 1441
rect 10870 1387 10872 1442
rect 10872 1387 10930 1442
rect 14134 2324 14206 2378
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 15278 1544 15312 1578
rect 13968 1503 14002 1537
rect 12743 1378 12792 1438
rect 17278 2324 17350 2378
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 18422 1544 18456 1578
rect 17112 1503 17146 1537
rect 20410 2328 20482 2382
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 21554 1548 21588 1582
rect 20244 1507 20278 1541
rect 12987 1382 13045 1437
rect 13045 1382 13047 1437
rect 14072 1383 14074 1438
rect 14074 1383 14132 1438
rect 15887 1378 15936 1438
rect 16131 1382 16189 1437
rect 16189 1382 16191 1437
rect 17216 1383 17218 1438
rect 17218 1383 17276 1438
rect 19019 1382 19068 1442
rect 30697 2769 30711 2803
rect 30711 2769 30745 2803
rect 30745 2769 30757 2803
rect 30697 2753 30757 2769
rect 30162 2674 30338 2708
rect 31387 2667 31563 2701
rect 30162 2556 30338 2590
rect 31286 2520 31320 2554
rect 31387 2549 31563 2583
rect 30162 2438 30338 2472
rect 23554 2328 23626 2382
rect 30655 2365 31031 2399
rect 29962 2308 30338 2342
rect 31219 2335 31253 2369
rect 30655 2247 31031 2281
rect 31387 2247 31763 2281
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 29962 2190 30338 2224
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 30655 2129 31031 2163
rect 29962 2072 30338 2106
rect 31387 2129 31763 2163
rect 31303 2069 31337 2103
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 30655 2011 31031 2045
rect 31387 2011 31763 2045
rect 29707 1951 29735 1989
rect 29735 1951 29745 1989
rect 29962 1954 30338 1988
rect 30655 1893 31031 1927
rect 29962 1836 30338 1870
rect 31302 1951 31336 1985
rect 31387 1893 31763 1927
rect 31929 2001 31951 2051
rect 31951 2001 31971 2051
rect 30655 1775 31031 1809
rect 31387 1775 31763 1809
rect 29962 1718 30338 1752
rect 30655 1657 31031 1691
rect 29962 1600 30338 1634
rect 24698 1548 24732 1582
rect 23388 1507 23422 1541
rect 30162 1471 30338 1505
rect 19263 1386 19321 1441
rect 19321 1386 19323 1441
rect 20348 1387 20350 1442
rect 20350 1387 20408 1442
rect 22163 1382 22212 1442
rect 22407 1386 22465 1441
rect 22465 1386 22467 1441
rect 23492 1387 23494 1442
rect 23494 1387 23552 1442
rect 30507 1409 30561 1419
rect 30162 1353 30338 1387
rect 30507 1375 30517 1409
rect 30517 1375 30551 1409
rect 30551 1375 30561 1409
rect 30507 1365 30561 1375
rect 121 1262 170 1322
rect 1700 1273 1734 1307
rect 3265 1262 3314 1322
rect 4844 1273 4878 1307
rect 6397 1266 6446 1326
rect 7976 1277 8010 1311
rect 9541 1266 9590 1326
rect 11120 1277 11154 1311
rect 12743 1262 12792 1322
rect 14322 1273 14356 1307
rect 15887 1262 15936 1322
rect 17466 1273 17500 1307
rect 19019 1266 19068 1326
rect 20598 1277 20632 1311
rect 22163 1266 22212 1326
rect 23742 1277 23776 1311
rect 30162 1235 30338 1269
rect 31219 1687 31253 1721
rect 31287 1397 31321 1431
rect 31387 1369 31563 1403
rect 31387 1251 31563 1285
rect 1332 1098 1334 1153
rect 1334 1098 1392 1153
rect 4476 1098 4478 1153
rect 4478 1098 4536 1153
rect 7608 1102 7610 1157
rect 7610 1102 7668 1157
rect 10752 1102 10754 1157
rect 10754 1102 10812 1157
rect 13954 1098 13956 1153
rect 13956 1098 14014 1153
rect 17098 1098 17100 1153
rect 17100 1098 17158 1153
rect 20230 1102 20232 1157
rect 20232 1102 20290 1157
rect 23374 1102 23376 1157
rect 23376 1102 23434 1157
rect 30162 1117 30338 1151
rect 31059 1085 31161 1187
rect 1581 883 1615 917
rect 4725 883 4759 917
rect 7857 887 7891 921
rect 11001 887 11035 921
rect 14203 883 14237 917
rect 17347 883 17381 917
rect 20479 887 20513 921
rect 23623 887 23657 921
rect 32534 866 32604 921
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 30164 723 30340 757
rect 30699 734 30759 750
rect 30699 700 30713 734
rect 30713 700 30747 734
rect 30747 700 30759 734
rect 30699 684 30759 700
rect 30164 605 30340 639
rect 31389 598 31565 632
rect 30164 487 30340 521
rect 31288 451 31322 485
rect 31389 480 31565 514
rect 30164 369 30340 403
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 23565 288 23599 322
rect 30657 296 31033 330
rect 29964 239 30340 273
rect 31221 266 31255 300
rect 30657 178 31033 212
rect 31389 178 31765 212
rect 1526 152 1584 166
rect 1526 120 1584 152
rect 4670 152 4728 166
rect 4670 120 4728 152
rect 7802 156 7860 170
rect 7802 124 7860 156
rect 10946 156 11004 170
rect 10946 124 11004 156
rect 14148 152 14206 166
rect 14148 120 14206 152
rect 17292 152 17350 166
rect 17292 120 17350 152
rect 20424 156 20482 170
rect 20424 124 20482 156
rect 23568 156 23626 170
rect 23568 124 23626 156
rect 29964 121 30340 155
rect 30657 60 31033 94
rect 29964 3 30340 37
rect 31389 60 31765 94
rect 31305 0 31339 34
rect 30657 -58 31033 -24
rect 31389 -58 31765 -24
rect 29709 -118 29737 -80
rect 29737 -118 29747 -80
rect 29964 -115 30340 -81
rect 30657 -176 31033 -142
rect 29964 -233 30340 -199
rect 31304 -118 31338 -84
rect 31389 -176 31765 -142
rect 31931 -68 31953 -18
rect 31953 -68 31973 -18
rect 30657 -294 31033 -260
rect 31389 -294 31765 -260
rect 29964 -351 30340 -317
rect 30657 -412 31033 -378
rect 29964 -469 30340 -435
rect 30164 -598 30340 -564
rect 30509 -660 30563 -650
rect 30164 -716 30340 -682
rect 30509 -694 30519 -660
rect 30519 -694 30553 -660
rect 30553 -694 30563 -660
rect 30509 -704 30563 -694
rect 30164 -834 30340 -800
rect 31221 -382 31255 -348
rect 31289 -672 31323 -638
rect 31389 -700 31565 -666
rect 31389 -818 31565 -784
rect 30164 -952 30340 -918
rect 31061 -984 31163 -882
rect 1544 -1568 1616 -1514
rect 292 -2140 326 -1964
rect 410 -2140 444 -1964
rect 528 -2140 562 -1964
rect 646 -2140 680 -1964
rect 733 -2140 767 -1764
rect 851 -2140 885 -1764
rect 969 -2140 1003 -1764
rect 1087 -2140 1121 -1764
rect 1200 -2140 1234 -1764
rect 1318 -2140 1352 -1764
rect 1436 -2140 1470 -1764
rect 1554 -2140 1588 -1764
rect 1672 -2140 1706 -1764
rect 1790 -2140 1824 -1764
rect 1908 -2140 1942 -1764
rect 2027 -2140 2061 -1764
rect 2145 -2140 2179 -1764
rect 2263 -2140 2297 -1764
rect 2381 -2140 2415 -1764
rect 2500 -2140 2534 -1964
rect 2618 -2140 2652 -1964
rect 2736 -2140 2770 -1964
rect 2854 -2140 2888 -1964
rect 2688 -2348 2722 -2314
rect 1378 -2389 1412 -2355
rect 4688 -1568 4760 -1514
rect 3436 -2140 3470 -1964
rect 3554 -2140 3588 -1964
rect 3672 -2140 3706 -1964
rect 3790 -2140 3824 -1964
rect 3877 -2140 3911 -1764
rect 3995 -2140 4029 -1764
rect 4113 -2140 4147 -1764
rect 4231 -2140 4265 -1764
rect 4344 -2140 4378 -1764
rect 4462 -2140 4496 -1764
rect 4580 -2140 4614 -1764
rect 4698 -2140 4732 -1764
rect 4816 -2140 4850 -1764
rect 4934 -2140 4968 -1764
rect 5052 -2140 5086 -1764
rect 5171 -2140 5205 -1764
rect 5289 -2140 5323 -1764
rect 5407 -2140 5441 -1764
rect 5525 -2140 5559 -1764
rect 5644 -2140 5678 -1964
rect 5762 -2140 5796 -1964
rect 5880 -2140 5914 -1964
rect 5998 -2140 6032 -1964
rect 5832 -2348 5866 -2314
rect 4522 -2389 4556 -2355
rect 7820 -1564 7892 -1510
rect 6568 -2136 6602 -1960
rect 6686 -2136 6720 -1960
rect 6804 -2136 6838 -1960
rect 6922 -2136 6956 -1960
rect 7009 -2136 7043 -1760
rect 7127 -2136 7161 -1760
rect 7245 -2136 7279 -1760
rect 7363 -2136 7397 -1760
rect 7476 -2136 7510 -1760
rect 7594 -2136 7628 -1760
rect 7712 -2136 7746 -1760
rect 7830 -2136 7864 -1760
rect 7948 -2136 7982 -1760
rect 8066 -2136 8100 -1760
rect 8184 -2136 8218 -1760
rect 8303 -2136 8337 -1760
rect 8421 -2136 8455 -1760
rect 8539 -2136 8573 -1760
rect 8657 -2136 8691 -1760
rect 8776 -2136 8810 -1960
rect 8894 -2136 8928 -1960
rect 9012 -2136 9046 -1960
rect 9130 -2136 9164 -1960
rect 8964 -2344 8998 -2310
rect 7654 -2385 7688 -2351
rect 153 -2514 202 -2454
rect 397 -2510 455 -2455
rect 455 -2510 457 -2455
rect 1482 -2509 1484 -2454
rect 1484 -2509 1542 -2454
rect 3297 -2514 3346 -2454
rect 3541 -2510 3599 -2455
rect 3599 -2510 3601 -2455
rect 4626 -2509 4628 -2454
rect 4628 -2509 4686 -2454
rect 10964 -1564 11036 -1510
rect 9712 -2136 9746 -1960
rect 9830 -2136 9864 -1960
rect 9948 -2136 9982 -1960
rect 10066 -2136 10100 -1960
rect 10153 -2136 10187 -1760
rect 10271 -2136 10305 -1760
rect 10389 -2136 10423 -1760
rect 10507 -2136 10541 -1760
rect 10620 -2136 10654 -1760
rect 10738 -2136 10772 -1760
rect 10856 -2136 10890 -1760
rect 10974 -2136 11008 -1760
rect 11092 -2136 11126 -1760
rect 11210 -2136 11244 -1760
rect 11328 -2136 11362 -1760
rect 11447 -2136 11481 -1760
rect 11565 -2136 11599 -1760
rect 11683 -2136 11717 -1760
rect 11801 -2136 11835 -1760
rect 11920 -2136 11954 -1960
rect 12038 -2136 12072 -1960
rect 12156 -2136 12190 -1960
rect 12274 -2136 12308 -1960
rect 12108 -2344 12142 -2310
rect 10798 -2385 10832 -2351
rect 14166 -1568 14238 -1514
rect 12914 -2140 12948 -1964
rect 13032 -2140 13066 -1964
rect 13150 -2140 13184 -1964
rect 13268 -2140 13302 -1964
rect 13355 -2140 13389 -1764
rect 13473 -2140 13507 -1764
rect 13591 -2140 13625 -1764
rect 13709 -2140 13743 -1764
rect 13822 -2140 13856 -1764
rect 13940 -2140 13974 -1764
rect 14058 -2140 14092 -1764
rect 14176 -2140 14210 -1764
rect 14294 -2140 14328 -1764
rect 14412 -2140 14446 -1764
rect 14530 -2140 14564 -1764
rect 14649 -2140 14683 -1764
rect 14767 -2140 14801 -1764
rect 14885 -2140 14919 -1764
rect 15003 -2140 15037 -1764
rect 15122 -2140 15156 -1964
rect 15240 -2140 15274 -1964
rect 15358 -2140 15392 -1964
rect 15476 -2140 15510 -1964
rect 15310 -2348 15344 -2314
rect 14000 -2389 14034 -2355
rect 17310 -1568 17382 -1514
rect 16058 -2140 16092 -1964
rect 16176 -2140 16210 -1964
rect 16294 -2140 16328 -1964
rect 16412 -2140 16446 -1964
rect 16499 -2140 16533 -1764
rect 16617 -2140 16651 -1764
rect 16735 -2140 16769 -1764
rect 16853 -2140 16887 -1764
rect 16966 -2140 17000 -1764
rect 17084 -2140 17118 -1764
rect 17202 -2140 17236 -1764
rect 17320 -2140 17354 -1764
rect 17438 -2140 17472 -1764
rect 17556 -2140 17590 -1764
rect 17674 -2140 17708 -1764
rect 17793 -2140 17827 -1764
rect 17911 -2140 17945 -1764
rect 18029 -2140 18063 -1764
rect 18147 -2140 18181 -1764
rect 18266 -2140 18300 -1964
rect 18384 -2140 18418 -1964
rect 18502 -2140 18536 -1964
rect 18620 -2140 18654 -1964
rect 18454 -2348 18488 -2314
rect 17144 -2389 17178 -2355
rect 20442 -1564 20514 -1510
rect 19190 -2136 19224 -1960
rect 19308 -2136 19342 -1960
rect 19426 -2136 19460 -1960
rect 19544 -2136 19578 -1960
rect 19631 -2136 19665 -1760
rect 19749 -2136 19783 -1760
rect 19867 -2136 19901 -1760
rect 19985 -2136 20019 -1760
rect 20098 -2136 20132 -1760
rect 20216 -2136 20250 -1760
rect 20334 -2136 20368 -1760
rect 20452 -2136 20486 -1760
rect 20570 -2136 20604 -1760
rect 20688 -2136 20722 -1760
rect 20806 -2136 20840 -1760
rect 20925 -2136 20959 -1760
rect 21043 -2136 21077 -1760
rect 21161 -2136 21195 -1760
rect 21279 -2136 21313 -1760
rect 21398 -2136 21432 -1960
rect 21516 -2136 21550 -1960
rect 21634 -2136 21668 -1960
rect 21752 -2136 21786 -1960
rect 21586 -2344 21620 -2310
rect 20276 -2385 20310 -2351
rect 6429 -2510 6478 -2450
rect 6673 -2506 6731 -2451
rect 6731 -2506 6733 -2451
rect 7758 -2505 7760 -2450
rect 7760 -2505 7818 -2450
rect 9573 -2510 9622 -2450
rect 9817 -2506 9875 -2451
rect 9875 -2506 9877 -2451
rect 10902 -2505 10904 -2450
rect 10904 -2505 10962 -2450
rect 12775 -2514 12824 -2454
rect 13019 -2510 13077 -2455
rect 13077 -2510 13079 -2455
rect 14104 -2509 14106 -2454
rect 14106 -2509 14164 -2454
rect 15919 -2514 15968 -2454
rect 16163 -2510 16221 -2455
rect 16221 -2510 16223 -2455
rect 17248 -2509 17250 -2454
rect 17250 -2509 17308 -2454
rect 30162 -1345 30338 -1311
rect 30697 -1334 30757 -1318
rect 23586 -1564 23658 -1510
rect 30697 -1368 30711 -1334
rect 30711 -1368 30745 -1334
rect 30745 -1368 30757 -1334
rect 30697 -1384 30757 -1368
rect 30162 -1463 30338 -1429
rect 31387 -1470 31563 -1436
rect 30162 -1581 30338 -1547
rect 31286 -1617 31320 -1583
rect 31387 -1588 31563 -1554
rect 22334 -2136 22368 -1960
rect 22452 -2136 22486 -1960
rect 22570 -2136 22604 -1960
rect 22688 -2136 22722 -1960
rect 22775 -2136 22809 -1760
rect 22893 -2136 22927 -1760
rect 23011 -2136 23045 -1760
rect 23129 -2136 23163 -1760
rect 23242 -2136 23276 -1760
rect 23360 -2136 23394 -1760
rect 23478 -2136 23512 -1760
rect 23596 -2136 23630 -1760
rect 23714 -2136 23748 -1760
rect 23832 -2136 23866 -1760
rect 30162 -1699 30338 -1665
rect 23950 -2136 23984 -1760
rect 24069 -2136 24103 -1760
rect 24187 -2136 24221 -1760
rect 24305 -2136 24339 -1760
rect 24423 -2136 24457 -1760
rect 30655 -1772 31031 -1738
rect 29962 -1829 30338 -1795
rect 31219 -1802 31253 -1768
rect 30655 -1890 31031 -1856
rect 31387 -1890 31763 -1856
rect 24542 -2136 24576 -1960
rect 24660 -2136 24694 -1960
rect 24778 -2136 24812 -1960
rect 29962 -1947 30338 -1913
rect 24896 -2136 24930 -1960
rect 30655 -2008 31031 -1974
rect 29962 -2065 30338 -2031
rect 31387 -2008 31763 -1974
rect 31303 -2068 31337 -2034
rect 30655 -2126 31031 -2092
rect 31387 -2126 31763 -2092
rect 29707 -2186 29735 -2148
rect 29735 -2186 29745 -2148
rect 29962 -2183 30338 -2149
rect 24730 -2344 24764 -2310
rect 23420 -2385 23454 -2351
rect 30655 -2244 31031 -2210
rect 29962 -2301 30338 -2267
rect 31302 -2186 31336 -2152
rect 31387 -2244 31763 -2210
rect 31929 -2136 31951 -2086
rect 31951 -2136 31971 -2086
rect 30655 -2362 31031 -2328
rect 31387 -2362 31763 -2328
rect 29962 -2419 30338 -2385
rect 19051 -2510 19100 -2450
rect 19295 -2506 19353 -2451
rect 19353 -2506 19355 -2451
rect 20380 -2505 20382 -2450
rect 20382 -2505 20440 -2450
rect 22195 -2510 22244 -2450
rect 22439 -2506 22497 -2451
rect 22497 -2506 22499 -2451
rect 23524 -2505 23526 -2450
rect 23526 -2505 23584 -2450
rect 30655 -2480 31031 -2446
rect 29962 -2537 30338 -2503
rect 1732 -2619 1766 -2585
rect 4876 -2619 4910 -2585
rect 8008 -2615 8042 -2581
rect 11152 -2615 11186 -2581
rect 14354 -2619 14388 -2585
rect 17498 -2619 17532 -2585
rect 20630 -2615 20664 -2581
rect 23774 -2615 23808 -2581
rect 30162 -2666 30338 -2632
rect 1364 -2794 1366 -2739
rect 1366 -2794 1424 -2739
rect 4508 -2794 4510 -2739
rect 4510 -2794 4568 -2739
rect 7640 -2790 7642 -2735
rect 7642 -2790 7700 -2735
rect 10784 -2790 10786 -2735
rect 10786 -2790 10844 -2735
rect 13986 -2794 13988 -2739
rect 13988 -2794 14046 -2739
rect 17130 -2794 17132 -2739
rect 17132 -2794 17190 -2739
rect 20262 -2790 20264 -2735
rect 20264 -2790 20322 -2735
rect 23406 -2790 23408 -2735
rect 23408 -2790 23466 -2735
rect 30507 -2728 30561 -2718
rect 30162 -2784 30338 -2750
rect 30507 -2762 30517 -2728
rect 30517 -2762 30551 -2728
rect 30551 -2762 30561 -2728
rect 30507 -2772 30561 -2762
rect 30162 -2902 30338 -2868
rect 31219 -2450 31253 -2416
rect 31287 -2740 31321 -2706
rect 39614 22695 39648 22871
rect 39732 22695 39766 22871
rect 39850 22695 39884 22871
rect 39968 22695 40002 22871
rect 40086 22695 40120 22871
rect 40204 22695 40238 22871
rect 40322 22695 40356 22871
rect 40440 22695 40474 22871
rect 40558 22695 40592 22871
rect 40676 22695 40710 22871
rect 46127 22692 46161 22868
rect 46245 22692 46279 22868
rect 46363 22692 46397 22868
rect 46481 22692 46515 22868
rect 46599 22692 46633 22868
rect 46717 22692 46751 22868
rect 46835 22692 46869 22868
rect 46953 22692 46987 22868
rect 47071 22692 47105 22868
rect 47189 22692 47223 22868
rect 52661 22687 52695 22863
rect 52779 22687 52813 22863
rect 52897 22687 52931 22863
rect 53015 22687 53049 22863
rect 53133 22687 53167 22863
rect 53251 22687 53285 22863
rect 53369 22687 53403 22863
rect 53487 22687 53521 22863
rect 53605 22687 53639 22863
rect 53723 22687 53757 22863
rect 59219 22691 59253 22867
rect 59337 22691 59371 22867
rect 59455 22691 59489 22867
rect 59573 22691 59607 22867
rect 59691 22691 59725 22867
rect 59809 22691 59843 22867
rect 59927 22691 59961 22867
rect 60045 22691 60079 22867
rect 60163 22691 60197 22867
rect 60281 22691 60315 22867
rect 40381 22601 40415 22635
rect 46894 22598 46928 22632
rect 53428 22593 53462 22627
rect 59986 22597 60020 22631
rect 40263 22484 40297 22518
rect 39851 22058 39885 22434
rect 39969 22058 40003 22434
rect 40087 22058 40121 22434
rect 40204 22258 40238 22434
rect 40322 22258 40356 22434
rect 41078 22078 41112 22254
rect 41196 22078 41230 22254
rect 41314 22078 41348 22254
rect 41432 22078 41466 22254
rect 41562 22078 41596 22454
rect 41680 22078 41714 22454
rect 41798 22078 41832 22454
rect 41916 22078 41950 22454
rect 42034 22078 42068 22454
rect 42152 22078 42186 22454
rect 42270 22078 42304 22454
rect 42399 22078 42433 22254
rect 42517 22078 42551 22254
rect 42635 22078 42669 22254
rect 42753 22078 42787 22254
rect 42976 22078 43010 22254
rect 43094 22078 43128 22254
rect 43212 22078 43246 22254
rect 43330 22078 43364 22254
rect 43460 22078 43494 22454
rect 43578 22078 43612 22454
rect 43696 22078 43730 22454
rect 43814 22078 43848 22454
rect 43932 22078 43966 22454
rect 46776 22481 46810 22515
rect 44050 22078 44084 22454
rect 44168 22078 44202 22454
rect 44297 22078 44331 22254
rect 44415 22078 44449 22254
rect 44533 22078 44567 22254
rect 44651 22078 44685 22254
rect 46364 22055 46398 22431
rect 46482 22055 46516 22431
rect 46600 22055 46634 22431
rect 46717 22255 46751 22431
rect 46835 22255 46869 22431
rect 39910 21974 39944 22008
rect 40028 21974 40062 22008
rect 47591 22075 47625 22251
rect 47709 22075 47743 22251
rect 47827 22075 47861 22251
rect 47945 22075 47979 22251
rect 48075 22075 48109 22451
rect 48193 22075 48227 22451
rect 48311 22075 48345 22451
rect 48429 22075 48463 22451
rect 48547 22075 48581 22451
rect 48665 22075 48699 22451
rect 48783 22075 48817 22451
rect 48912 22075 48946 22251
rect 49030 22075 49064 22251
rect 49148 22075 49182 22251
rect 49266 22075 49300 22251
rect 49489 22075 49523 22251
rect 49607 22075 49641 22251
rect 49725 22075 49759 22251
rect 49843 22075 49877 22251
rect 49973 22075 50007 22451
rect 50091 22075 50125 22451
rect 50209 22075 50243 22451
rect 50327 22075 50361 22451
rect 50445 22075 50479 22451
rect 53310 22476 53344 22510
rect 50563 22075 50597 22451
rect 50681 22075 50715 22451
rect 50810 22075 50844 22251
rect 50928 22075 50962 22251
rect 51046 22075 51080 22251
rect 51164 22075 51198 22251
rect 52898 22050 52932 22426
rect 53016 22050 53050 22426
rect 53134 22050 53168 22426
rect 53251 22250 53285 22426
rect 53369 22250 53403 22426
rect 46423 21971 46457 22005
rect 46541 21971 46575 22005
rect 54125 22070 54159 22246
rect 54243 22070 54277 22246
rect 54361 22070 54395 22246
rect 54479 22070 54513 22246
rect 54609 22070 54643 22446
rect 54727 22070 54761 22446
rect 54845 22070 54879 22446
rect 54963 22070 54997 22446
rect 55081 22070 55115 22446
rect 55199 22070 55233 22446
rect 55317 22070 55351 22446
rect 55446 22070 55480 22246
rect 55564 22070 55598 22246
rect 55682 22070 55716 22246
rect 55800 22070 55834 22246
rect 56023 22070 56057 22246
rect 56141 22070 56175 22246
rect 56259 22070 56293 22246
rect 56377 22070 56411 22246
rect 56507 22070 56541 22446
rect 56625 22070 56659 22446
rect 56743 22070 56777 22446
rect 56861 22070 56895 22446
rect 56979 22070 57013 22446
rect 59868 22480 59902 22514
rect 57097 22070 57131 22446
rect 57215 22070 57249 22446
rect 57344 22070 57378 22246
rect 57462 22070 57496 22246
rect 57580 22070 57614 22246
rect 57698 22070 57732 22246
rect 59456 22054 59490 22430
rect 59574 22054 59608 22430
rect 59692 22054 59726 22430
rect 59809 22254 59843 22430
rect 59927 22254 59961 22430
rect 52957 21966 52991 22000
rect 53075 21966 53109 22000
rect 60683 22074 60717 22250
rect 60801 22074 60835 22250
rect 60919 22074 60953 22250
rect 61037 22074 61071 22250
rect 61167 22074 61201 22450
rect 61285 22074 61319 22450
rect 61403 22074 61437 22450
rect 61521 22074 61555 22450
rect 61639 22074 61673 22450
rect 61757 22074 61791 22450
rect 61875 22074 61909 22450
rect 62004 22074 62038 22250
rect 62122 22074 62156 22250
rect 62240 22074 62274 22250
rect 62358 22074 62392 22250
rect 62581 22074 62615 22250
rect 62699 22074 62733 22250
rect 62817 22074 62851 22250
rect 62935 22074 62969 22250
rect 63065 22074 63099 22450
rect 63183 22074 63217 22450
rect 63301 22074 63335 22450
rect 63419 22074 63453 22450
rect 63537 22074 63571 22450
rect 63655 22074 63689 22450
rect 63773 22074 63807 22450
rect 63902 22074 63936 22250
rect 64020 22074 64054 22250
rect 64138 22074 64172 22250
rect 64256 22074 64290 22250
rect 68618 22235 68701 22300
rect 59515 21970 59549 22004
rect 59633 21970 59667 22004
rect 42542 21806 42576 21840
rect 44649 21785 44683 21819
rect 49055 21803 49089 21837
rect 41505 21385 41539 21761
rect 41623 21385 41657 21761
rect 39609 21091 39643 21267
rect 39727 21091 39761 21267
rect 39845 21091 39879 21267
rect 39963 21091 39997 21267
rect 40081 21091 40115 21267
rect 40199 21091 40233 21267
rect 40317 21091 40351 21267
rect 40435 21091 40469 21267
rect 40553 21091 40587 21267
rect 41741 21385 41775 21761
rect 41859 21385 41893 21761
rect 41977 21385 42011 21761
rect 42095 21385 42129 21761
rect 42213 21385 42247 21761
rect 43403 21385 43437 21761
rect 43521 21385 43555 21761
rect 43639 21385 43673 21761
rect 43757 21385 43791 21761
rect 43875 21385 43909 21761
rect 43993 21385 44027 21761
rect 51162 21782 51196 21816
rect 55589 21798 55623 21832
rect 44111 21385 44145 21761
rect 48018 21382 48052 21758
rect 48136 21382 48170 21758
rect 40671 21091 40705 21267
rect 41535 21163 41569 21197
rect 41350 21096 41384 21130
rect 42183 21163 42217 21197
rect 43433 21163 43467 21197
rect 41801 21079 41835 21113
rect 41919 21080 41953 21114
rect 42473 21095 42507 21129
rect 43248 21096 43282 21130
rect 44079 21164 44113 21198
rect 43699 21079 43733 21113
rect 43817 21080 43851 21114
rect 44371 21095 44405 21129
rect 40376 20997 40410 21031
rect 40258 20880 40292 20914
rect 41203 20853 41237 21029
rect 39846 20454 39880 20830
rect 39964 20454 39998 20830
rect 40082 20454 40116 20830
rect 40199 20654 40233 20830
rect 41321 20853 41355 21029
rect 40317 20654 40351 20830
rect 41623 20653 41657 21029
rect 41741 20653 41775 21029
rect 41859 20653 41893 21029
rect 41977 20653 42011 21029
rect 42095 20653 42129 21029
rect 42501 20853 42535 21029
rect 42619 20853 42653 21029
rect 43101 20853 43135 21029
rect 43219 20853 43253 21029
rect 43521 20653 43555 21029
rect 43639 20653 43673 21029
rect 43757 20653 43791 21029
rect 43875 20653 43909 21029
rect 43993 20653 44027 21029
rect 44399 20853 44433 21029
rect 44517 20853 44551 21029
rect 39905 20370 39939 20404
rect 40023 20370 40057 20404
rect 46122 21088 46156 21264
rect 46240 21088 46274 21264
rect 46358 21088 46392 21264
rect 46476 21088 46510 21264
rect 46594 21088 46628 21264
rect 46712 21088 46746 21264
rect 46830 21088 46864 21264
rect 46948 21088 46982 21264
rect 47066 21088 47100 21264
rect 48254 21382 48288 21758
rect 48372 21382 48406 21758
rect 48490 21382 48524 21758
rect 48608 21382 48642 21758
rect 48726 21382 48760 21758
rect 49916 21382 49950 21758
rect 50034 21382 50068 21758
rect 50152 21382 50186 21758
rect 50270 21382 50304 21758
rect 50388 21382 50422 21758
rect 50506 21382 50540 21758
rect 57696 21777 57730 21811
rect 62147 21802 62181 21836
rect 50624 21382 50658 21758
rect 54552 21377 54586 21753
rect 54670 21377 54704 21753
rect 47184 21088 47218 21264
rect 48048 21160 48082 21194
rect 47863 21093 47897 21127
rect 48696 21160 48730 21194
rect 49946 21160 49980 21194
rect 48314 21076 48348 21110
rect 48432 21077 48466 21111
rect 48986 21092 49020 21126
rect 49761 21093 49795 21127
rect 50592 21161 50626 21195
rect 50212 21076 50246 21110
rect 50330 21077 50364 21111
rect 50884 21092 50918 21126
rect 46889 20994 46923 21028
rect 46771 20877 46805 20911
rect 47716 20850 47750 21026
rect 46359 20451 46393 20827
rect 46477 20451 46511 20827
rect 46595 20451 46629 20827
rect 46712 20651 46746 20827
rect 47834 20850 47868 21026
rect 46830 20651 46864 20827
rect 48136 20650 48170 21026
rect 48254 20650 48288 21026
rect 48372 20650 48406 21026
rect 48490 20650 48524 21026
rect 48608 20650 48642 21026
rect 49014 20850 49048 21026
rect 49132 20850 49166 21026
rect 49614 20850 49648 21026
rect 49732 20850 49766 21026
rect 50034 20650 50068 21026
rect 50152 20650 50186 21026
rect 50270 20650 50304 21026
rect 50388 20650 50422 21026
rect 50506 20650 50540 21026
rect 50912 20850 50946 21026
rect 51030 20850 51064 21026
rect 46418 20367 46452 20401
rect 46536 20367 46570 20401
rect 52656 21083 52690 21259
rect 52774 21083 52808 21259
rect 52892 21083 52926 21259
rect 53010 21083 53044 21259
rect 53128 21083 53162 21259
rect 53246 21083 53280 21259
rect 53364 21083 53398 21259
rect 53482 21083 53516 21259
rect 53600 21083 53634 21259
rect 54788 21377 54822 21753
rect 54906 21377 54940 21753
rect 55024 21377 55058 21753
rect 55142 21377 55176 21753
rect 55260 21377 55294 21753
rect 56450 21377 56484 21753
rect 56568 21377 56602 21753
rect 56686 21377 56720 21753
rect 56804 21377 56838 21753
rect 56922 21377 56956 21753
rect 57040 21377 57074 21753
rect 64254 21781 64288 21815
rect 57158 21377 57192 21753
rect 61110 21381 61144 21757
rect 61228 21381 61262 21757
rect 53718 21083 53752 21259
rect 54582 21155 54616 21189
rect 54397 21088 54431 21122
rect 55230 21155 55264 21189
rect 56480 21155 56514 21189
rect 54848 21071 54882 21105
rect 54966 21072 55000 21106
rect 55520 21087 55554 21121
rect 56295 21088 56329 21122
rect 57126 21156 57160 21190
rect 56746 21071 56780 21105
rect 56864 21072 56898 21106
rect 57418 21087 57452 21121
rect 53423 20989 53457 21023
rect 53305 20872 53339 20906
rect 54250 20845 54284 21021
rect 52893 20446 52927 20822
rect 53011 20446 53045 20822
rect 53129 20446 53163 20822
rect 53246 20646 53280 20822
rect 54368 20845 54402 21021
rect 53364 20646 53398 20822
rect 54670 20645 54704 21021
rect 54788 20645 54822 21021
rect 54906 20645 54940 21021
rect 55024 20645 55058 21021
rect 55142 20645 55176 21021
rect 55548 20845 55582 21021
rect 55666 20845 55700 21021
rect 56148 20845 56182 21021
rect 56266 20845 56300 21021
rect 56568 20645 56602 21021
rect 56686 20645 56720 21021
rect 56804 20645 56838 21021
rect 56922 20645 56956 21021
rect 57040 20645 57074 21021
rect 57446 20845 57480 21021
rect 57564 20845 57598 21021
rect 52952 20362 52986 20396
rect 53070 20362 53104 20396
rect 59214 21087 59248 21263
rect 59332 21087 59366 21263
rect 59450 21087 59484 21263
rect 59568 21087 59602 21263
rect 59686 21087 59720 21263
rect 59804 21087 59838 21263
rect 59922 21087 59956 21263
rect 60040 21087 60074 21263
rect 60158 21087 60192 21263
rect 61346 21381 61380 21757
rect 61464 21381 61498 21757
rect 61582 21381 61616 21757
rect 61700 21381 61734 21757
rect 61818 21381 61852 21757
rect 63008 21381 63042 21757
rect 63126 21381 63160 21757
rect 63244 21381 63278 21757
rect 63362 21381 63396 21757
rect 63480 21381 63514 21757
rect 63598 21381 63632 21757
rect 63716 21381 63750 21757
rect 60276 21087 60310 21263
rect 61140 21159 61174 21193
rect 60955 21092 60989 21126
rect 61788 21159 61822 21193
rect 63038 21159 63072 21193
rect 61406 21075 61440 21109
rect 61524 21076 61558 21110
rect 62078 21091 62112 21125
rect 62853 21092 62887 21126
rect 65917 21264 66062 21342
rect 63684 21160 63718 21194
rect 63304 21075 63338 21109
rect 63422 21076 63456 21110
rect 63976 21091 64010 21125
rect 59981 20993 60015 21027
rect 59863 20876 59897 20910
rect 60808 20849 60842 21025
rect 59451 20450 59485 20826
rect 59569 20450 59603 20826
rect 59687 20450 59721 20826
rect 59804 20650 59838 20826
rect 60926 20849 60960 21025
rect 59922 20650 59956 20826
rect 61228 20649 61262 21025
rect 61346 20649 61380 21025
rect 61464 20649 61498 21025
rect 61582 20649 61616 21025
rect 61700 20649 61734 21025
rect 62106 20849 62140 21025
rect 62224 20849 62258 21025
rect 62706 20849 62740 21025
rect 62824 20849 62858 21025
rect 63126 20649 63160 21025
rect 63244 20649 63278 21025
rect 63362 20649 63396 21025
rect 63480 20649 63514 21025
rect 63598 20649 63632 21025
rect 64004 20849 64038 21025
rect 64122 20849 64156 21025
rect 59510 20366 59544 20400
rect 59628 20366 59662 20400
rect 66434 19890 66569 19962
rect 67002 19722 67132 19812
rect 71499 22151 71559 22200
rect 70725 22027 70901 22061
rect 70725 21909 70901 21943
rect 70725 21791 70901 21825
rect 71216 21898 71271 21956
rect 71216 21896 71271 21898
rect 70725 21673 70901 21707
rect 70525 21586 70901 21620
rect 70525 21468 70901 21502
rect 70525 21350 70901 21384
rect 70525 21232 70901 21266
rect 70525 21119 70901 21153
rect 71858 21193 72034 21227
rect 71858 21075 72034 21109
rect 70525 21001 70901 21035
rect 70525 20883 70901 20917
rect 70275 20737 70329 20809
rect 71858 21001 72234 21035
rect 71116 20941 71150 20975
rect 71500 20987 71555 20989
rect 71500 20929 71555 20987
rect 70525 20765 70901 20799
rect 71858 20883 72234 20917
rect 71215 20869 71270 20871
rect 71215 20811 71270 20869
rect 71858 20765 72234 20799
rect 70525 20647 70901 20681
rect 72335 20764 72369 20798
rect 71736 20706 71770 20740
rect 72487 20737 72501 20795
rect 72501 20737 72533 20795
rect 71858 20647 72234 20681
rect 71346 20587 71380 20621
rect 70525 20529 70901 20563
rect 71858 20529 72234 20563
rect 70525 20411 70901 20445
rect 71858 20451 72034 20485
rect 71858 20333 72034 20367
rect 70525 20292 70901 20326
rect 70525 20174 70901 20208
rect 70525 20056 70901 20090
rect 70525 19938 70901 19972
rect 70725 19819 70901 19853
rect 40446 19133 40480 19167
rect 41576 19127 41610 19161
rect 47004 19129 47038 19163
rect 48134 19123 48168 19157
rect 53538 19134 53572 19168
rect 54668 19128 54702 19162
rect 70725 19701 70901 19735
rect 70725 19583 70901 19617
rect 71075 19631 71109 19665
rect 70725 19465 70901 19499
rect 60051 19137 60085 19171
rect 61181 19131 61215 19165
rect 40446 19013 40480 19047
rect 39611 18613 39645 18989
rect 39729 18613 39763 18989
rect 39847 18613 39881 18989
rect 39965 18613 39999 18989
rect 40083 18613 40117 18989
rect 40201 18613 40235 18989
rect 41576 19009 41610 19043
rect 40319 18613 40353 18989
rect 40753 18609 40787 18985
rect 40871 18609 40905 18985
rect 40989 18609 41023 18985
rect 41107 18609 41141 18985
rect 41225 18609 41259 18985
rect 41343 18609 41377 18985
rect 47004 19009 47038 19043
rect 41461 18609 41495 18985
rect 42724 18737 42758 18913
rect 42842 18737 42876 18913
rect 42960 18737 42994 18913
rect 43078 18737 43112 18913
rect 43196 18737 43230 18913
rect 43314 18737 43348 18913
rect 43432 18737 43466 18913
rect 43550 18737 43584 18913
rect 43668 18737 43702 18913
rect 43786 18737 43820 18913
rect 43019 18643 43053 18677
rect 46169 18609 46203 18985
rect 46287 18609 46321 18985
rect 46405 18609 46439 18985
rect 46523 18609 46557 18985
rect 46641 18609 46675 18985
rect 46759 18609 46793 18985
rect 48134 19005 48168 19039
rect 53538 19014 53572 19048
rect 46877 18609 46911 18985
rect 47311 18605 47345 18981
rect 47429 18605 47463 18981
rect 47547 18605 47581 18981
rect 47665 18605 47699 18981
rect 47783 18605 47817 18981
rect 47901 18605 47935 18981
rect 48019 18605 48053 18981
rect 49282 18733 49316 18909
rect 49400 18733 49434 18909
rect 49518 18733 49552 18909
rect 49636 18733 49670 18909
rect 49754 18733 49788 18909
rect 49872 18733 49906 18909
rect 49990 18733 50024 18909
rect 50108 18733 50142 18909
rect 50226 18733 50260 18909
rect 50344 18733 50378 18909
rect 49577 18639 49611 18673
rect 52703 18614 52737 18990
rect 52821 18614 52855 18990
rect 52939 18614 52973 18990
rect 53057 18614 53091 18990
rect 53175 18614 53209 18990
rect 53293 18614 53327 18990
rect 54668 19010 54702 19044
rect 53411 18614 53445 18990
rect 53845 18610 53879 18986
rect 53963 18610 53997 18986
rect 54081 18610 54115 18986
rect 54199 18610 54233 18986
rect 54317 18610 54351 18986
rect 54435 18610 54469 18986
rect 60051 19017 60085 19051
rect 54553 18610 54587 18986
rect 55816 18738 55850 18914
rect 55934 18738 55968 18914
rect 56052 18738 56086 18914
rect 56170 18738 56204 18914
rect 56288 18738 56322 18914
rect 56406 18738 56440 18914
rect 56524 18738 56558 18914
rect 56642 18738 56676 18914
rect 56760 18738 56794 18914
rect 56878 18738 56912 18914
rect 56111 18644 56145 18678
rect 59216 18617 59250 18993
rect 59334 18617 59368 18993
rect 59452 18617 59486 18993
rect 59570 18617 59604 18993
rect 59688 18617 59722 18993
rect 59806 18617 59840 18993
rect 61181 19013 61215 19047
rect 59924 18617 59958 18993
rect 60358 18613 60392 18989
rect 60476 18613 60510 18989
rect 60594 18613 60628 18989
rect 60712 18613 60746 18989
rect 60830 18613 60864 18989
rect 60948 18613 60982 18989
rect 61066 18613 61100 18989
rect 62329 18741 62363 18917
rect 62447 18741 62481 18917
rect 62565 18741 62599 18917
rect 62683 18741 62717 18917
rect 62801 18741 62835 18917
rect 62919 18741 62953 18917
rect 63037 18741 63071 18917
rect 63155 18741 63189 18917
rect 63273 18741 63307 18917
rect 63391 18741 63425 18917
rect 62624 18647 62658 18681
rect 43137 18526 43171 18560
rect 49695 18522 49729 18556
rect 56229 18527 56263 18561
rect 62742 18530 62776 18564
rect 43078 18300 43112 18476
rect 40114 18257 40148 18291
rect 41256 18253 41290 18287
rect 43196 18300 43230 18476
rect 39536 18030 39570 18206
rect 39654 18030 39688 18206
rect 39772 18030 39806 18206
rect 39890 18030 39924 18206
rect 40055 18030 40089 18206
rect 40173 18030 40207 18206
rect 40291 18030 40325 18206
rect 40409 18030 40443 18206
rect 40678 18026 40712 18202
rect 40796 18026 40830 18202
rect 40914 18026 40948 18202
rect 41032 18026 41066 18202
rect 41197 18026 41231 18202
rect 41315 18026 41349 18202
rect 41433 18026 41467 18202
rect 41551 18026 41585 18202
rect 43313 18100 43347 18476
rect 43431 18100 43465 18476
rect 43549 18100 43583 18476
rect 49636 18296 49670 18472
rect 46672 18253 46706 18287
rect 47814 18249 47848 18283
rect 49754 18296 49788 18472
rect 43372 18016 43406 18050
rect 43490 18016 43524 18050
rect 46094 18026 46128 18202
rect 46212 18026 46246 18202
rect 46330 18026 46364 18202
rect 46448 18026 46482 18202
rect 46613 18026 46647 18202
rect 46731 18026 46765 18202
rect 46849 18026 46883 18202
rect 46967 18026 47001 18202
rect 47236 18022 47270 18198
rect 47354 18022 47388 18198
rect 47472 18022 47506 18198
rect 47590 18022 47624 18198
rect 47755 18022 47789 18198
rect 47873 18022 47907 18198
rect 47991 18022 48025 18198
rect 48109 18022 48143 18198
rect 49871 18096 49905 18472
rect 49989 18096 50023 18472
rect 50107 18096 50141 18472
rect 56170 18301 56204 18477
rect 53206 18258 53240 18292
rect 54348 18254 54382 18288
rect 56288 18301 56322 18477
rect 49930 18012 49964 18046
rect 50048 18012 50082 18046
rect 52628 18031 52662 18207
rect 52746 18031 52780 18207
rect 52864 18031 52898 18207
rect 52982 18031 53016 18207
rect 53147 18031 53181 18207
rect 53265 18031 53299 18207
rect 53383 18031 53417 18207
rect 53501 18031 53535 18207
rect 53770 18027 53804 18203
rect 53888 18027 53922 18203
rect 54006 18027 54040 18203
rect 54124 18027 54158 18203
rect 54289 18027 54323 18203
rect 54407 18027 54441 18203
rect 54525 18027 54559 18203
rect 54643 18027 54677 18203
rect 56405 18101 56439 18477
rect 56523 18101 56557 18477
rect 56641 18101 56675 18477
rect 62683 18304 62717 18480
rect 59719 18261 59753 18295
rect 60861 18257 60895 18291
rect 62801 18304 62835 18480
rect 56464 18017 56498 18051
rect 56582 18017 56616 18051
rect 59141 18034 59175 18210
rect 59259 18034 59293 18210
rect 59377 18034 59411 18210
rect 59495 18034 59529 18210
rect 59660 18034 59694 18210
rect 59778 18034 59812 18210
rect 59896 18034 59930 18210
rect 60014 18034 60048 18210
rect 60283 18030 60317 18206
rect 60401 18030 60435 18206
rect 60519 18030 60553 18206
rect 60637 18030 60671 18206
rect 60802 18030 60836 18206
rect 60920 18030 60954 18206
rect 61038 18030 61072 18206
rect 61156 18030 61190 18206
rect 62918 18104 62952 18480
rect 63036 18104 63070 18480
rect 63154 18104 63188 18480
rect 62977 18020 63011 18054
rect 63095 18020 63129 18054
rect 44496 17462 44607 17571
rect 42710 17087 42744 17263
rect 42828 17087 42862 17263
rect 42946 17087 42980 17263
rect 43064 17087 43098 17263
rect 43182 17087 43216 17263
rect 43300 17087 43334 17263
rect 43418 17087 43452 17263
rect 43536 17087 43570 17263
rect 43654 17087 43688 17263
rect 43772 17087 43806 17263
rect 43005 16993 43039 17027
rect 38735 16470 38769 16646
rect 38853 16470 38887 16646
rect 38971 16470 39005 16646
rect 39089 16470 39123 16646
rect 39218 16470 39252 16846
rect 39336 16470 39370 16846
rect 39454 16470 39488 16846
rect 39572 16470 39606 16846
rect 39690 16470 39724 16846
rect 39808 16470 39842 16846
rect 39926 16470 39960 16846
rect 40056 16470 40090 16646
rect 40174 16470 40208 16646
rect 40292 16470 40326 16646
rect 40410 16470 40444 16646
rect 40633 16470 40667 16646
rect 40751 16470 40785 16646
rect 40869 16470 40903 16646
rect 40987 16470 41021 16646
rect 41116 16470 41150 16846
rect 41234 16470 41268 16846
rect 41352 16470 41386 16846
rect 43123 16876 43157 16910
rect 41470 16470 41504 16846
rect 41588 16470 41622 16846
rect 41706 16470 41740 16846
rect 41824 16470 41858 16846
rect 41954 16470 41988 16646
rect 42072 16470 42106 16646
rect 42190 16470 42224 16646
rect 42308 16470 42342 16646
rect 43064 16650 43098 16826
rect 43182 16650 43216 16826
rect 43299 16450 43333 16826
rect 43417 16450 43451 16826
rect 43535 16450 43569 16826
rect 43358 16366 43392 16400
rect 43476 16366 43510 16400
rect 38737 16177 38771 16211
rect 40844 16198 40878 16232
rect 39275 15777 39309 16153
rect 39393 15777 39427 16153
rect 38516 15650 38648 15748
rect 39511 15777 39545 16153
rect 39629 15777 39663 16153
rect 39747 15777 39781 16153
rect 39865 15777 39899 16153
rect 39983 15777 40017 16153
rect 41173 15777 41207 16153
rect 41291 15777 41325 16153
rect 41409 15777 41443 16153
rect 41527 15777 41561 16153
rect 41645 15777 41679 16153
rect 41763 15777 41797 16153
rect 41881 15777 41915 16153
rect 39307 15556 39341 15590
rect 39015 15487 39049 15521
rect 39569 15472 39603 15506
rect 39687 15471 39721 15505
rect 39953 15555 39987 15589
rect 41203 15555 41237 15589
rect 40138 15488 40172 15522
rect 40913 15487 40947 15521
rect 41467 15472 41501 15506
rect 41585 15471 41619 15505
rect 41851 15555 41885 15589
rect 42036 15488 42070 15522
rect 42715 15483 42749 15659
rect 42833 15483 42867 15659
rect 42951 15483 42985 15659
rect 43069 15483 43103 15659
rect 43187 15483 43221 15659
rect 43305 15483 43339 15659
rect 43423 15483 43457 15659
rect 43541 15483 43575 15659
rect 43659 15483 43693 15659
rect 43777 15483 43811 15659
rect 38869 15245 38903 15421
rect 38987 15245 39021 15421
rect 39393 15045 39427 15421
rect 39511 15045 39545 15421
rect 39629 15045 39663 15421
rect 39747 15045 39781 15421
rect 39865 15045 39899 15421
rect 40167 15245 40201 15421
rect 40285 15245 40319 15421
rect 40767 15245 40801 15421
rect 40885 15245 40919 15421
rect 41291 15045 41325 15421
rect 41409 15045 41443 15421
rect 41527 15045 41561 15421
rect 41645 15045 41679 15421
rect 41763 15045 41797 15421
rect 42065 15245 42099 15421
rect 42183 15245 42217 15421
rect 43010 15389 43044 15423
rect 43128 15272 43162 15306
rect 43069 15046 43103 15222
rect 43187 15046 43221 15222
rect 43304 14846 43338 15222
rect 43422 14846 43456 15222
rect 43540 14846 43574 15222
rect 43363 14762 43397 14796
rect 43481 14762 43515 14796
rect 51059 17462 51162 17559
rect 49268 17083 49302 17259
rect 49386 17083 49420 17259
rect 49504 17083 49538 17259
rect 49622 17083 49656 17259
rect 49740 17083 49774 17259
rect 49858 17083 49892 17259
rect 49976 17083 50010 17259
rect 50094 17083 50128 17259
rect 50212 17083 50246 17259
rect 50330 17083 50364 17259
rect 49563 16989 49597 17023
rect 45293 16466 45327 16642
rect 45411 16466 45445 16642
rect 45529 16466 45563 16642
rect 45647 16466 45681 16642
rect 45776 16466 45810 16842
rect 45894 16466 45928 16842
rect 46012 16466 46046 16842
rect 46130 16466 46164 16842
rect 46248 16466 46282 16842
rect 46366 16466 46400 16842
rect 46484 16466 46518 16842
rect 46614 16466 46648 16642
rect 46732 16466 46766 16642
rect 46850 16466 46884 16642
rect 46968 16466 47002 16642
rect 47191 16466 47225 16642
rect 47309 16466 47343 16642
rect 47427 16466 47461 16642
rect 47545 16466 47579 16642
rect 47674 16466 47708 16842
rect 47792 16466 47826 16842
rect 47910 16466 47944 16842
rect 49681 16872 49715 16906
rect 48028 16466 48062 16842
rect 48146 16466 48180 16842
rect 48264 16466 48298 16842
rect 48382 16466 48416 16842
rect 48512 16466 48546 16642
rect 48630 16466 48664 16642
rect 48748 16466 48782 16642
rect 48866 16466 48900 16642
rect 49622 16646 49656 16822
rect 49740 16646 49774 16822
rect 49857 16446 49891 16822
rect 49975 16446 50009 16822
rect 50093 16446 50127 16822
rect 49916 16362 49950 16396
rect 50034 16362 50068 16396
rect 45295 16173 45329 16207
rect 47402 16194 47436 16228
rect 45833 15773 45867 16149
rect 45951 15773 45985 16149
rect 45074 15646 45206 15744
rect 46069 15773 46103 16149
rect 46187 15773 46221 16149
rect 46305 15773 46339 16149
rect 46423 15773 46457 16149
rect 46541 15773 46575 16149
rect 47731 15773 47765 16149
rect 47849 15773 47883 16149
rect 47967 15773 48001 16149
rect 48085 15773 48119 16149
rect 48203 15773 48237 16149
rect 48321 15773 48355 16149
rect 48439 15773 48473 16149
rect 45865 15552 45899 15586
rect 45573 15483 45607 15517
rect 46127 15468 46161 15502
rect 46245 15467 46279 15501
rect 46511 15551 46545 15585
rect 47761 15551 47795 15585
rect 46696 15484 46730 15518
rect 47471 15483 47505 15517
rect 48025 15468 48059 15502
rect 48143 15467 48177 15501
rect 48409 15551 48443 15585
rect 48594 15484 48628 15518
rect 49273 15479 49307 15655
rect 49391 15479 49425 15655
rect 49509 15479 49543 15655
rect 49627 15479 49661 15655
rect 49745 15479 49779 15655
rect 49863 15479 49897 15655
rect 49981 15479 50015 15655
rect 50099 15479 50133 15655
rect 50217 15479 50251 15655
rect 50335 15479 50369 15655
rect 45427 15241 45461 15417
rect 45545 15241 45579 15417
rect 45951 15041 45985 15417
rect 46069 15041 46103 15417
rect 46187 15041 46221 15417
rect 46305 15041 46339 15417
rect 46423 15041 46457 15417
rect 46725 15241 46759 15417
rect 46843 15241 46877 15417
rect 47325 15241 47359 15417
rect 47443 15241 47477 15417
rect 47849 15041 47883 15417
rect 47967 15041 48001 15417
rect 48085 15041 48119 15417
rect 48203 15041 48237 15417
rect 48321 15041 48355 15417
rect 48623 15241 48657 15417
rect 48741 15241 48775 15417
rect 49568 15385 49602 15419
rect 49686 15268 49720 15302
rect 49627 15042 49661 15218
rect 49745 15042 49779 15218
rect 49862 14842 49896 15218
rect 49980 14842 50014 15218
rect 50098 14842 50132 15218
rect 49921 14758 49955 14792
rect 50039 14758 50073 14792
rect 57595 17471 57693 17563
rect 55802 17088 55836 17264
rect 55920 17088 55954 17264
rect 56038 17088 56072 17264
rect 56156 17088 56190 17264
rect 56274 17088 56308 17264
rect 56392 17088 56426 17264
rect 56510 17088 56544 17264
rect 56628 17088 56662 17264
rect 56746 17088 56780 17264
rect 56864 17088 56898 17264
rect 56097 16994 56131 17028
rect 51827 16471 51861 16647
rect 51945 16471 51979 16647
rect 52063 16471 52097 16647
rect 52181 16471 52215 16647
rect 52310 16471 52344 16847
rect 52428 16471 52462 16847
rect 52546 16471 52580 16847
rect 52664 16471 52698 16847
rect 52782 16471 52816 16847
rect 52900 16471 52934 16847
rect 53018 16471 53052 16847
rect 53148 16471 53182 16647
rect 53266 16471 53300 16647
rect 53384 16471 53418 16647
rect 53502 16471 53536 16647
rect 53725 16471 53759 16647
rect 53843 16471 53877 16647
rect 53961 16471 53995 16647
rect 54079 16471 54113 16647
rect 54208 16471 54242 16847
rect 54326 16471 54360 16847
rect 54444 16471 54478 16847
rect 56215 16877 56249 16911
rect 54562 16471 54596 16847
rect 54680 16471 54714 16847
rect 54798 16471 54832 16847
rect 54916 16471 54950 16847
rect 55046 16471 55080 16647
rect 55164 16471 55198 16647
rect 55282 16471 55316 16647
rect 55400 16471 55434 16647
rect 56156 16651 56190 16827
rect 56274 16651 56308 16827
rect 56391 16451 56425 16827
rect 56509 16451 56543 16827
rect 56627 16451 56661 16827
rect 56450 16367 56484 16401
rect 56568 16367 56602 16401
rect 51829 16178 51863 16212
rect 53936 16199 53970 16233
rect 52367 15778 52401 16154
rect 52485 15778 52519 16154
rect 51608 15651 51740 15749
rect 52603 15778 52637 16154
rect 52721 15778 52755 16154
rect 52839 15778 52873 16154
rect 52957 15778 52991 16154
rect 53075 15778 53109 16154
rect 54265 15778 54299 16154
rect 54383 15778 54417 16154
rect 54501 15778 54535 16154
rect 54619 15778 54653 16154
rect 54737 15778 54771 16154
rect 54855 15778 54889 16154
rect 54973 15778 55007 16154
rect 52399 15557 52433 15591
rect 52107 15488 52141 15522
rect 52661 15473 52695 15507
rect 52779 15472 52813 15506
rect 53045 15556 53079 15590
rect 54295 15556 54329 15590
rect 53230 15489 53264 15523
rect 54005 15488 54039 15522
rect 54559 15473 54593 15507
rect 54677 15472 54711 15506
rect 54943 15556 54977 15590
rect 55128 15489 55162 15523
rect 55807 15484 55841 15660
rect 55925 15484 55959 15660
rect 56043 15484 56077 15660
rect 56161 15484 56195 15660
rect 56279 15484 56313 15660
rect 56397 15484 56431 15660
rect 56515 15484 56549 15660
rect 56633 15484 56667 15660
rect 56751 15484 56785 15660
rect 56869 15484 56903 15660
rect 51961 15246 51995 15422
rect 52079 15246 52113 15422
rect 52485 15046 52519 15422
rect 52603 15046 52637 15422
rect 52721 15046 52755 15422
rect 52839 15046 52873 15422
rect 52957 15046 52991 15422
rect 53259 15246 53293 15422
rect 53377 15246 53411 15422
rect 53859 15246 53893 15422
rect 53977 15246 54011 15422
rect 54383 15046 54417 15422
rect 54501 15046 54535 15422
rect 54619 15046 54653 15422
rect 54737 15046 54771 15422
rect 54855 15046 54889 15422
rect 55157 15246 55191 15422
rect 55275 15246 55309 15422
rect 56102 15390 56136 15424
rect 56220 15273 56254 15307
rect 56161 15047 56195 15223
rect 56279 15047 56313 15223
rect 56396 14847 56430 15223
rect 56514 14847 56548 15223
rect 56632 14847 56666 15223
rect 56455 14763 56489 14797
rect 56573 14763 56607 14797
rect 62315 17091 62349 17267
rect 62433 17091 62467 17267
rect 62551 17091 62585 17267
rect 62669 17091 62703 17267
rect 62787 17091 62821 17267
rect 62905 17091 62939 17267
rect 63023 17091 63057 17267
rect 63141 17091 63175 17267
rect 63259 17091 63293 17267
rect 63377 17091 63411 17267
rect 62610 16997 62644 17031
rect 58340 16474 58374 16650
rect 58458 16474 58492 16650
rect 58576 16474 58610 16650
rect 58694 16474 58728 16650
rect 58823 16474 58857 16850
rect 58941 16474 58975 16850
rect 59059 16474 59093 16850
rect 59177 16474 59211 16850
rect 59295 16474 59329 16850
rect 59413 16474 59447 16850
rect 59531 16474 59565 16850
rect 59661 16474 59695 16650
rect 59779 16474 59813 16650
rect 59897 16474 59931 16650
rect 60015 16474 60049 16650
rect 60238 16474 60272 16650
rect 60356 16474 60390 16650
rect 60474 16474 60508 16650
rect 60592 16474 60626 16650
rect 60721 16474 60755 16850
rect 60839 16474 60873 16850
rect 60957 16474 60991 16850
rect 62728 16880 62762 16914
rect 61075 16474 61109 16850
rect 61193 16474 61227 16850
rect 61311 16474 61345 16850
rect 61429 16474 61463 16850
rect 61559 16474 61593 16650
rect 61677 16474 61711 16650
rect 61795 16474 61829 16650
rect 61913 16474 61947 16650
rect 62669 16654 62703 16830
rect 62787 16654 62821 16830
rect 62904 16454 62938 16830
rect 63022 16454 63056 16830
rect 63140 16454 63174 16830
rect 62963 16370 62997 16404
rect 63081 16370 63115 16404
rect 58342 16181 58376 16215
rect 60449 16202 60483 16236
rect 58880 15781 58914 16157
rect 58998 15781 59032 16157
rect 58121 15654 58253 15752
rect 59116 15781 59150 16157
rect 59234 15781 59268 16157
rect 59352 15781 59386 16157
rect 59470 15781 59504 16157
rect 59588 15781 59622 16157
rect 60778 15781 60812 16157
rect 60896 15781 60930 16157
rect 61014 15781 61048 16157
rect 61132 15781 61166 16157
rect 61250 15781 61284 16157
rect 61368 15781 61402 16157
rect 61486 15781 61520 16157
rect 58912 15560 58946 15594
rect 58620 15491 58654 15525
rect 59174 15476 59208 15510
rect 59292 15475 59326 15509
rect 59558 15559 59592 15593
rect 60808 15559 60842 15593
rect 59743 15492 59777 15526
rect 60518 15491 60552 15525
rect 61072 15476 61106 15510
rect 61190 15475 61224 15509
rect 61456 15559 61490 15593
rect 61641 15492 61675 15526
rect 62320 15487 62354 15663
rect 62438 15487 62472 15663
rect 62556 15487 62590 15663
rect 62674 15487 62708 15663
rect 62792 15487 62826 15663
rect 62910 15487 62944 15663
rect 63028 15487 63062 15663
rect 63146 15487 63180 15663
rect 63264 15487 63298 15663
rect 63382 15487 63416 15663
rect 58474 15249 58508 15425
rect 58592 15249 58626 15425
rect 58998 15049 59032 15425
rect 59116 15049 59150 15425
rect 59234 15049 59268 15425
rect 59352 15049 59386 15425
rect 59470 15049 59504 15425
rect 59772 15249 59806 15425
rect 59890 15249 59924 15425
rect 60372 15249 60406 15425
rect 60490 15249 60524 15425
rect 60896 15049 60930 15425
rect 61014 15049 61048 15425
rect 61132 15049 61166 15425
rect 61250 15049 61284 15425
rect 61368 15049 61402 15425
rect 61670 15249 61704 15425
rect 61788 15249 61822 15425
rect 62615 15393 62649 15427
rect 62733 15276 62767 15310
rect 62674 15050 62708 15226
rect 62792 15050 62826 15226
rect 62909 14850 62943 15226
rect 63027 14850 63061 15226
rect 63145 14850 63179 15226
rect 62968 14766 63002 14800
rect 63086 14766 63120 14800
rect 57742 13097 57810 13155
rect 51217 12980 51288 13036
rect 68260 19086 68309 19149
rect 71499 19007 71559 19056
rect 70725 18883 70901 18917
rect 70725 18765 70901 18799
rect 70725 18647 70901 18681
rect 71216 18754 71271 18812
rect 71216 18752 71271 18754
rect 70725 18529 70901 18563
rect 70525 18442 70901 18476
rect 70525 18324 70901 18358
rect 70525 18206 70901 18240
rect 70525 18088 70901 18122
rect 70525 17975 70901 18009
rect 71858 18049 72034 18083
rect 71858 17931 72034 17965
rect 70525 17857 70901 17891
rect 70525 17739 70901 17773
rect 70275 17593 70329 17665
rect 71858 17857 72234 17891
rect 71116 17797 71150 17831
rect 71500 17843 71555 17845
rect 71500 17785 71555 17843
rect 70525 17621 70901 17655
rect 71858 17739 72234 17773
rect 71215 17725 71270 17727
rect 71215 17667 71270 17725
rect 71858 17621 72234 17655
rect 70525 17503 70901 17537
rect 72335 17620 72369 17654
rect 71736 17562 71770 17596
rect 72487 17593 72501 17651
rect 72501 17593 72533 17651
rect 71858 17503 72234 17537
rect 71346 17443 71380 17477
rect 70525 17385 70901 17419
rect 71858 17385 72234 17419
rect 70525 17267 70901 17301
rect 71858 17307 72034 17341
rect 71858 17189 72034 17223
rect 70525 17148 70901 17182
rect 70525 17030 70901 17064
rect 70525 16912 70901 16946
rect 70525 16794 70901 16828
rect 70725 16675 70901 16709
rect 70725 16557 70901 16591
rect 70725 16439 70901 16473
rect 71075 16487 71109 16521
rect 70725 16321 70901 16355
rect 44641 12658 44720 12703
rect 41911 12313 41971 12375
rect 48460 12312 48520 12374
rect 55114 12333 55174 12395
rect 64610 12293 64688 12365
rect 41570 11961 41604 12137
rect 41688 11961 41722 12137
rect 41806 11961 41840 12137
rect 41924 11961 41958 12137
rect 42042 11961 42076 12137
rect 42160 11961 42194 12137
rect 42278 11961 42312 12137
rect 42396 11961 42430 12137
rect 42514 11961 42548 12137
rect 42632 11961 42666 12137
rect 48119 11960 48153 12136
rect 48237 11960 48271 12136
rect 48355 11960 48389 12136
rect 48473 11960 48507 12136
rect 48591 11960 48625 12136
rect 48709 11960 48743 12136
rect 48827 11960 48861 12136
rect 48945 11960 48979 12136
rect 49063 11960 49097 12136
rect 49181 11960 49215 12136
rect 54773 11981 54807 12157
rect 54891 11981 54925 12157
rect 55009 11981 55043 12157
rect 55127 11981 55161 12157
rect 55245 11981 55279 12157
rect 55363 11981 55397 12157
rect 55481 11981 55515 12157
rect 55599 11981 55633 12157
rect 55717 11981 55751 12157
rect 55835 11981 55869 12157
rect 63767 12166 63827 12228
rect 65868 12289 66289 12323
rect 65868 12144 65931 12289
rect 65931 12144 66240 12289
rect 66240 12144 66289 12289
rect 65868 12123 66289 12144
rect 42337 11867 42371 11901
rect 48886 11866 48920 11900
rect 55540 11887 55574 11921
rect 63426 11814 63460 11990
rect 42219 11750 42253 11784
rect 48768 11749 48802 11783
rect 55422 11770 55456 11804
rect 63544 11814 63578 11990
rect 63662 11814 63696 11990
rect 63780 11814 63814 11990
rect 63898 11814 63932 11990
rect 64016 11814 64050 11990
rect 64134 11814 64168 11990
rect 64252 11814 64286 11990
rect 64370 11814 64404 11990
rect 64488 11814 64522 11990
rect 41807 11324 41841 11700
rect 41925 11324 41959 11700
rect 42043 11324 42077 11700
rect 42160 11524 42194 11700
rect 42278 11524 42312 11700
rect 48356 11323 48390 11699
rect 48474 11323 48508 11699
rect 48592 11323 48626 11699
rect 48709 11523 48743 11699
rect 48827 11523 48861 11699
rect 55010 11344 55044 11720
rect 55128 11344 55162 11720
rect 55246 11344 55280 11720
rect 55363 11544 55397 11720
rect 64193 11720 64227 11754
rect 55481 11544 55515 11720
rect 64075 11603 64109 11637
rect 41866 11240 41900 11274
rect 41984 11240 42018 11274
rect 48269 11228 48318 11274
rect 48415 11239 48449 11273
rect 48533 11239 48567 11273
rect 54876 11248 54937 11296
rect 55069 11260 55103 11294
rect 55187 11260 55221 11294
rect 42139 11117 42191 11163
rect 33824 10784 33883 10840
rect 33985 10972 34046 11022
rect 33781 9425 33855 9495
rect 48688 11116 48740 11162
rect 41688 10795 41737 10849
rect 54978 11168 55023 11206
rect 55342 11137 55394 11183
rect 63663 11177 63697 11553
rect 63781 11177 63815 11553
rect 63899 11177 63933 11553
rect 64016 11377 64050 11553
rect 64134 11377 64168 11553
rect 65234 11409 65268 11585
rect 65352 11409 65386 11585
rect 65470 11409 65504 11585
rect 65588 11409 65622 11585
rect 65718 11409 65752 11785
rect 65836 11409 65870 11785
rect 65954 11409 65988 11785
rect 66072 11409 66106 11785
rect 66190 11409 66224 11785
rect 66308 11409 66342 11785
rect 66426 11409 66460 11785
rect 67368 11758 67428 11820
rect 66555 11409 66589 11585
rect 66673 11409 66707 11585
rect 66791 11409 66825 11585
rect 66909 11409 66943 11585
rect 67027 11406 67061 11582
rect 67145 11406 67179 11582
rect 67263 11406 67297 11582
rect 67381 11406 67415 11582
rect 67499 11406 67533 11582
rect 67617 11406 67651 11582
rect 67735 11406 67769 11582
rect 67853 11406 67887 11582
rect 67971 11406 68005 11582
rect 68089 11406 68123 11582
rect 67794 11312 67828 11346
rect 66886 11193 66920 11227
rect 67676 11195 67710 11229
rect 63722 11093 63756 11127
rect 63840 11093 63874 11127
rect 65213 11053 65293 11121
rect 65486 11074 65520 11108
rect 63995 10970 64047 11016
rect 34138 10404 34195 10449
rect 33965 9231 34078 9315
rect 33778 6607 33872 6688
rect 33779 832 33861 914
rect 33773 -2266 33867 -2190
rect 35247 10413 35307 10475
rect 34906 10061 34940 10237
rect 35024 10061 35058 10237
rect 35142 10061 35176 10237
rect 35260 10061 35294 10237
rect 35378 10061 35412 10237
rect 35496 10061 35530 10237
rect 35614 10061 35648 10237
rect 35732 10061 35766 10237
rect 35850 10061 35884 10237
rect 35968 10061 36002 10237
rect 35673 9967 35707 10001
rect 35555 9850 35589 9884
rect 34257 832 34359 913
rect 34403 9417 34492 9493
rect 35143 9424 35177 9800
rect 35261 9424 35295 9800
rect 35379 9424 35413 9800
rect 35496 9624 35530 9800
rect 35614 9624 35648 9800
rect 35202 9340 35236 9374
rect 35320 9340 35354 9374
rect 34897 9255 34953 9299
rect 35475 9217 35527 9263
rect 35239 7828 35299 7890
rect 34898 7476 34932 7652
rect 35016 7476 35050 7652
rect 35134 7476 35168 7652
rect 35252 7476 35286 7652
rect 35370 7476 35404 7652
rect 35488 7476 35522 7652
rect 35606 7476 35640 7652
rect 35724 7476 35758 7652
rect 35842 7476 35876 7652
rect 35960 7476 35994 7652
rect 35665 7382 35699 7416
rect 35547 7265 35581 7299
rect 35135 6839 35169 7215
rect 35253 6839 35287 7215
rect 35371 6839 35405 7215
rect 35488 7039 35522 7215
rect 35606 7039 35640 7215
rect 35194 6755 35228 6789
rect 35312 6755 35346 6789
rect 35467 6632 35519 6678
rect 35220 4550 35280 4612
rect 34879 4198 34913 4374
rect 34997 4198 35031 4374
rect 35115 4198 35149 4374
rect 35233 4198 35267 4374
rect 35351 4198 35385 4374
rect 35469 4198 35503 4374
rect 35587 4198 35621 4374
rect 35705 4198 35739 4374
rect 35823 4198 35857 4374
rect 35941 4198 35975 4374
rect 35646 4104 35680 4138
rect 35528 3987 35562 4021
rect 35116 3561 35150 3937
rect 35234 3561 35268 3937
rect 35352 3561 35386 3937
rect 35469 3761 35503 3937
rect 35587 3761 35621 3937
rect 35175 3477 35209 3511
rect 35293 3477 35327 3511
rect 34841 3387 34901 3440
rect 35448 3354 35500 3400
rect 35236 1790 35296 1852
rect 34895 1438 34929 1614
rect 35013 1438 35047 1614
rect 35131 1438 35165 1614
rect 35249 1438 35283 1614
rect 35367 1438 35401 1614
rect 35485 1438 35519 1614
rect 35603 1438 35637 1614
rect 35721 1438 35755 1614
rect 35839 1438 35873 1614
rect 35957 1438 35991 1614
rect 35662 1344 35696 1378
rect 35544 1227 35578 1261
rect 35132 801 35166 1177
rect 35250 801 35284 1177
rect 35368 801 35402 1177
rect 35485 1001 35519 1177
rect 35603 1001 35637 1177
rect 35191 717 35225 751
rect 35309 717 35343 751
rect 35464 594 35516 640
rect 34377 -2520 34521 -2454
rect 33962 -2665 34076 -2594
rect 38271 10384 38338 10385
rect 38271 10236 38337 10384
rect 38337 10236 38338 10384
rect 40753 10289 40819 10435
rect 40819 10289 40820 10435
rect 40753 10286 40820 10289
rect 40006 10184 40040 10218
rect 41895 10289 41899 10437
rect 41899 10289 41962 10437
rect 41895 10288 41962 10289
rect 41136 10190 41170 10224
rect 44820 10472 44887 10473
rect 44820 10324 44886 10472
rect 44886 10324 44887 10472
rect 47303 10377 47368 10524
rect 47368 10377 47370 10524
rect 47303 10375 47370 10377
rect 46555 10272 46589 10306
rect 48447 10377 48448 10526
rect 48448 10377 48514 10526
rect 47685 10278 47719 10312
rect 51473 10255 51540 10403
rect 51473 10254 51540 10255
rect 53954 10458 54021 10459
rect 53954 10310 53955 10458
rect 53955 10310 54021 10458
rect 46555 10154 46589 10188
rect 40006 10066 40040 10100
rect 41136 10070 41170 10104
rect 47685 10158 47719 10192
rect 37796 9794 37830 9970
rect 37914 9794 37948 9970
rect 38032 9794 38066 9970
rect 38150 9794 38184 9970
rect 38268 9794 38302 9970
rect 38386 9794 38420 9970
rect 38504 9794 38538 9970
rect 38622 9794 38656 9970
rect 38740 9794 38774 9970
rect 38858 9794 38892 9970
rect 38563 9700 38597 9734
rect 40121 9666 40155 10042
rect 40239 9666 40273 10042
rect 40357 9666 40391 10042
rect 40475 9666 40509 10042
rect 40593 9666 40627 10042
rect 40711 9666 40745 10042
rect 40829 9666 40863 10042
rect 41263 9670 41297 10046
rect 41381 9670 41415 10046
rect 41499 9670 41533 10046
rect 41617 9670 41651 10046
rect 41735 9670 41769 10046
rect 41853 9670 41887 10046
rect 41971 9670 42005 10046
rect 44345 9882 44379 10058
rect 44463 9882 44497 10058
rect 44581 9882 44615 10058
rect 44699 9882 44733 10058
rect 44817 9882 44851 10058
rect 44935 9882 44969 10058
rect 45053 9882 45087 10058
rect 45171 9882 45205 10058
rect 45289 9882 45323 10058
rect 45407 9882 45441 10058
rect 45112 9788 45146 9822
rect 46670 9754 46704 10130
rect 46788 9754 46822 10130
rect 46906 9754 46940 10130
rect 47024 9754 47058 10130
rect 47142 9754 47176 10130
rect 47260 9754 47294 10130
rect 47378 9754 47412 10130
rect 47812 9758 47846 10134
rect 47930 9758 47964 10134
rect 48048 9758 48082 10134
rect 48166 9758 48200 10134
rect 48284 9758 48318 10134
rect 48402 9758 48436 10134
rect 53209 10204 53243 10238
rect 55101 10309 55102 10458
rect 55102 10309 55168 10458
rect 54339 10210 54373 10244
rect 58093 10323 58098 10472
rect 58098 10323 58160 10472
rect 60577 10377 60580 10524
rect 60580 10377 60644 10524
rect 60577 10375 60644 10377
rect 59834 10272 59868 10306
rect 61726 10526 61793 10530
rect 61726 10381 61727 10526
rect 61727 10381 61793 10526
rect 60964 10278 60998 10312
rect 59834 10154 59868 10188
rect 48520 9758 48554 10134
rect 53209 10086 53243 10120
rect 54339 10090 54373 10124
rect 50999 9814 51033 9990
rect 51117 9814 51151 9990
rect 51235 9814 51269 9990
rect 51353 9814 51387 9990
rect 51471 9814 51505 9990
rect 51589 9814 51623 9990
rect 51707 9814 51741 9990
rect 51825 9814 51859 9990
rect 51943 9814 51977 9990
rect 52061 9814 52095 9990
rect 51766 9720 51800 9754
rect 44994 9671 45028 9705
rect 53324 9686 53358 10062
rect 53442 9686 53476 10062
rect 53560 9686 53594 10062
rect 53678 9686 53712 10062
rect 53796 9686 53830 10062
rect 53914 9686 53948 10062
rect 60964 10158 60998 10192
rect 54032 9686 54066 10062
rect 54466 9690 54500 10066
rect 54584 9690 54618 10066
rect 54702 9690 54736 10066
rect 54820 9690 54854 10066
rect 54938 9690 54972 10066
rect 55056 9690 55090 10066
rect 55174 9690 55208 10066
rect 57624 9882 57658 10058
rect 57742 9882 57776 10058
rect 57860 9882 57894 10058
rect 57978 9882 58012 10058
rect 58096 9882 58130 10058
rect 58214 9882 58248 10058
rect 58332 9882 58366 10058
rect 58450 9882 58484 10058
rect 58568 9882 58602 10058
rect 58686 9882 58720 10058
rect 58391 9788 58425 9822
rect 59949 9754 59983 10130
rect 60067 9754 60101 10130
rect 60185 9754 60219 10130
rect 60303 9754 60337 10130
rect 60421 9754 60455 10130
rect 60539 9754 60573 10130
rect 60657 9754 60691 10130
rect 61091 9758 61125 10134
rect 61209 9758 61243 10134
rect 61327 9758 61361 10134
rect 61445 9758 61479 10134
rect 61563 9758 61597 10134
rect 61681 9758 61715 10134
rect 61799 9758 61833 10134
rect 58273 9671 58307 9705
rect 38445 9583 38479 9617
rect 38033 9157 38067 9533
rect 38151 9157 38185 9533
rect 38269 9157 38303 9533
rect 38386 9357 38420 9533
rect 38504 9357 38538 9533
rect 40326 9310 40360 9344
rect 41468 9314 41502 9348
rect 38612 9129 38761 9196
rect 38092 9073 38126 9107
rect 38210 9073 38244 9107
rect 40031 9083 40065 9259
rect 40149 9083 40183 9259
rect 40267 9083 40301 9259
rect 40385 9083 40419 9259
rect 40550 9083 40584 9259
rect 40668 9083 40702 9259
rect 40786 9083 40820 9259
rect 40904 9083 40938 9259
rect 41173 9087 41207 9263
rect 41291 9087 41325 9263
rect 41409 9087 41443 9263
rect 41527 9087 41561 9263
rect 41692 9087 41726 9263
rect 41810 9087 41844 9263
rect 41928 9087 41962 9263
rect 42046 9087 42080 9263
rect 44582 9245 44616 9621
rect 44700 9245 44734 9621
rect 44818 9245 44852 9621
rect 44935 9445 44969 9621
rect 45053 9445 45087 9621
rect 51648 9603 51682 9637
rect 46875 9398 46909 9432
rect 48017 9402 48051 9436
rect 45158 9211 45307 9278
rect 44641 9161 44675 9195
rect 44759 9161 44793 9195
rect 46580 9171 46614 9347
rect 46698 9171 46732 9347
rect 46816 9171 46850 9347
rect 46934 9171 46968 9347
rect 47099 9171 47133 9347
rect 47217 9171 47251 9347
rect 47335 9171 47369 9347
rect 47453 9171 47487 9347
rect 47722 9175 47756 9351
rect 47840 9175 47874 9351
rect 47958 9175 47992 9351
rect 48076 9175 48110 9351
rect 48241 9175 48275 9351
rect 48359 9175 48393 9351
rect 48477 9175 48511 9351
rect 48595 9175 48629 9351
rect 51236 9177 51270 9553
rect 51354 9177 51388 9553
rect 51472 9177 51506 9553
rect 51589 9377 51623 9553
rect 51707 9377 51741 9553
rect 53529 9330 53563 9364
rect 54671 9334 54705 9368
rect 51808 9145 51957 9212
rect 51295 9093 51329 9127
rect 51413 9093 51447 9127
rect 53234 9103 53268 9279
rect 53352 9103 53386 9279
rect 53470 9103 53504 9279
rect 53588 9103 53622 9279
rect 53753 9103 53787 9279
rect 53871 9103 53905 9279
rect 53989 9103 54023 9279
rect 54107 9103 54141 9279
rect 54376 9107 54410 9283
rect 54494 9107 54528 9283
rect 54612 9107 54646 9283
rect 54730 9107 54764 9283
rect 54895 9107 54929 9283
rect 55013 9107 55047 9283
rect 55131 9107 55165 9283
rect 55249 9107 55283 9283
rect 57861 9245 57895 9621
rect 57979 9245 58013 9621
rect 58097 9245 58131 9621
rect 58214 9445 58248 9621
rect 58332 9445 58366 9621
rect 63762 9595 63822 9657
rect 60154 9398 60188 9432
rect 61296 9402 61330 9436
rect 58440 9221 58589 9288
rect 57920 9161 57954 9195
rect 58038 9161 58072 9195
rect 59859 9171 59893 9347
rect 59977 9171 60011 9347
rect 60095 9171 60129 9347
rect 60213 9171 60247 9347
rect 60378 9171 60412 9347
rect 60496 9171 60530 9347
rect 60614 9171 60648 9347
rect 60732 9171 60766 9347
rect 61001 9175 61035 9351
rect 61119 9175 61153 9351
rect 61237 9175 61271 9351
rect 61355 9175 61389 9351
rect 61520 9175 61554 9351
rect 61638 9175 61672 9351
rect 61756 9175 61790 9351
rect 61874 9175 61908 9351
rect 63421 9243 63455 9419
rect 63539 9243 63573 9419
rect 63657 9243 63691 9419
rect 63775 9243 63809 9419
rect 63893 9243 63927 9419
rect 64011 9243 64045 9419
rect 64129 9243 64163 9419
rect 64247 9243 64281 9419
rect 64365 9243 64399 9419
rect 64483 9243 64517 9419
rect 64188 9149 64222 9183
rect 64070 9032 64104 9066
rect 38283 8585 38284 8734
rect 38284 8585 38350 8734
rect 40098 8676 40165 8825
rect 41236 8678 41303 8827
rect 44834 8673 44900 8821
rect 44900 8673 44901 8821
rect 44834 8672 44901 8673
rect 46643 8772 46710 8921
rect 47782 8764 47849 8913
rect 51488 8754 51555 8755
rect 51488 8606 51554 8754
rect 51554 8606 51555 8754
rect 53296 8700 53363 8849
rect 54442 8703 54509 8852
rect 58116 8673 58179 8821
rect 58179 8673 58183 8821
rect 58116 8672 58183 8673
rect 59917 8761 59984 8908
rect 59917 8759 59984 8761
rect 61060 8761 61127 8910
rect 37810 8144 37844 8320
rect 37928 8144 37962 8320
rect 38046 8144 38080 8320
rect 38164 8144 38198 8320
rect 38282 8144 38316 8320
rect 38400 8144 38434 8320
rect 38518 8144 38552 8320
rect 38636 8144 38670 8320
rect 38754 8144 38788 8320
rect 38872 8144 38906 8320
rect 41995 8391 42062 8392
rect 41995 8243 42062 8391
rect 44359 8232 44393 8408
rect 44477 8232 44511 8408
rect 44595 8232 44629 8408
rect 44713 8232 44747 8408
rect 44831 8232 44865 8408
rect 44949 8232 44983 8408
rect 45067 8232 45101 8408
rect 45185 8232 45219 8408
rect 45303 8232 45337 8408
rect 45421 8232 45455 8408
rect 63658 8606 63692 8982
rect 63776 8606 63810 8982
rect 63894 8606 63928 8982
rect 64011 8806 64045 8982
rect 64129 8806 64163 8982
rect 48549 8330 48611 8479
rect 48611 8330 48616 8479
rect 45126 8138 45160 8172
rect 51013 8164 51047 8340
rect 51131 8164 51165 8340
rect 51249 8164 51283 8340
rect 51367 8164 51401 8340
rect 51485 8164 51519 8340
rect 51603 8164 51637 8340
rect 51721 8164 51755 8340
rect 51839 8164 51873 8340
rect 51957 8164 51991 8340
rect 52075 8164 52109 8340
rect 55195 8262 55198 8407
rect 55198 8262 55262 8407
rect 55195 8258 55262 8262
rect 57638 8232 57672 8408
rect 57756 8232 57790 8408
rect 57874 8232 57908 8408
rect 57992 8232 58026 8408
rect 58110 8232 58144 8408
rect 58228 8232 58262 8408
rect 58346 8232 58380 8408
rect 58464 8232 58498 8408
rect 58582 8232 58616 8408
rect 58700 8232 58734 8408
rect 63717 8522 63751 8556
rect 63835 8522 63869 8556
rect 61823 8330 61890 8476
rect 61823 8327 61890 8330
rect 63990 8399 64042 8445
rect 58405 8138 58439 8172
rect 38577 8050 38611 8084
rect 45008 8021 45042 8055
rect 38459 7933 38493 7967
rect 37008 7404 37126 7514
rect 38047 7507 38081 7883
rect 38165 7507 38199 7883
rect 38283 7507 38317 7883
rect 38400 7707 38434 7883
rect 38518 7707 38552 7883
rect 38627 7479 38776 7546
rect 39274 7527 39308 7703
rect 39392 7527 39426 7703
rect 39510 7527 39544 7703
rect 39628 7527 39662 7703
rect 39758 7527 39792 7903
rect 39876 7527 39910 7903
rect 39994 7527 40028 7903
rect 40112 7527 40146 7903
rect 40230 7527 40264 7903
rect 40348 7527 40382 7903
rect 40466 7527 40500 7903
rect 40595 7527 40629 7703
rect 40713 7527 40747 7703
rect 40831 7527 40865 7703
rect 40949 7527 40983 7703
rect 41172 7527 41206 7703
rect 41290 7527 41324 7703
rect 41408 7527 41442 7703
rect 41526 7527 41560 7703
rect 41656 7527 41690 7903
rect 41774 7527 41808 7903
rect 41892 7527 41926 7903
rect 42010 7527 42044 7903
rect 42128 7527 42162 7903
rect 42246 7527 42280 7903
rect 42364 7527 42398 7903
rect 42493 7527 42527 7703
rect 42611 7527 42645 7703
rect 42729 7527 42763 7703
rect 42847 7527 42881 7703
rect 44596 7595 44630 7971
rect 44714 7595 44748 7971
rect 44832 7595 44866 7971
rect 44949 7795 44983 7971
rect 45067 7795 45101 7971
rect 45176 7561 45325 7628
rect 45823 7615 45857 7791
rect 45941 7615 45975 7791
rect 46059 7615 46093 7791
rect 46177 7615 46211 7791
rect 46307 7615 46341 7991
rect 46425 7615 46459 7991
rect 46543 7615 46577 7991
rect 46661 7615 46695 7991
rect 46779 7615 46813 7991
rect 51780 8070 51814 8104
rect 46897 7615 46931 7991
rect 47015 7615 47049 7991
rect 47144 7615 47178 7791
rect 47262 7615 47296 7791
rect 47380 7615 47414 7791
rect 47498 7615 47532 7791
rect 47721 7615 47755 7791
rect 47839 7615 47873 7791
rect 47957 7615 47991 7791
rect 48075 7615 48109 7791
rect 48205 7615 48239 7991
rect 48323 7615 48357 7991
rect 48441 7615 48475 7991
rect 48559 7615 48593 7991
rect 48677 7615 48711 7991
rect 58287 8021 58321 8055
rect 48795 7615 48829 7991
rect 48913 7615 48947 7991
rect 51662 7953 51696 7987
rect 49042 7615 49076 7791
rect 49160 7615 49194 7791
rect 49278 7615 49312 7791
rect 49396 7615 49430 7791
rect 44655 7511 44689 7545
rect 44773 7511 44807 7545
rect 38106 7423 38140 7457
rect 38224 7423 38258 7457
rect 50210 7426 50349 7543
rect 51250 7527 51284 7903
rect 51368 7527 51402 7903
rect 51486 7527 51520 7903
rect 51603 7727 51637 7903
rect 51721 7727 51755 7903
rect 51825 7494 51974 7561
rect 52477 7547 52511 7723
rect 52595 7547 52629 7723
rect 52713 7547 52747 7723
rect 52831 7547 52865 7723
rect 52961 7547 52995 7923
rect 53079 7547 53113 7923
rect 53197 7547 53231 7923
rect 53315 7547 53349 7923
rect 53433 7547 53467 7923
rect 53551 7547 53585 7923
rect 53669 7547 53703 7923
rect 53798 7547 53832 7723
rect 53916 7547 53950 7723
rect 54034 7547 54068 7723
rect 54152 7547 54186 7723
rect 54375 7547 54409 7723
rect 54493 7547 54527 7723
rect 54611 7547 54645 7723
rect 54729 7547 54763 7723
rect 54859 7547 54893 7923
rect 54977 7547 55011 7923
rect 55095 7547 55129 7923
rect 55213 7547 55247 7923
rect 55331 7547 55365 7923
rect 55449 7547 55483 7923
rect 55567 7547 55601 7923
rect 55696 7547 55730 7723
rect 55814 7547 55848 7723
rect 55932 7547 55966 7723
rect 56050 7547 56084 7723
rect 57875 7595 57909 7971
rect 57993 7595 58027 7971
rect 58111 7595 58145 7971
rect 58228 7795 58262 7971
rect 58346 7795 58380 7971
rect 58445 7560 58594 7627
rect 59102 7615 59136 7791
rect 59220 7615 59254 7791
rect 59338 7615 59372 7791
rect 59456 7615 59490 7791
rect 59586 7615 59620 7991
rect 59704 7615 59738 7991
rect 59822 7615 59856 7991
rect 59940 7615 59974 7991
rect 60058 7615 60092 7991
rect 60176 7615 60210 7991
rect 60294 7615 60328 7991
rect 60423 7615 60457 7791
rect 60541 7615 60575 7791
rect 60659 7615 60693 7791
rect 60777 7615 60811 7791
rect 61000 7615 61034 7791
rect 61118 7615 61152 7791
rect 61236 7615 61270 7791
rect 61354 7615 61388 7791
rect 61484 7615 61518 7991
rect 61602 7615 61636 7991
rect 61720 7615 61754 7991
rect 61838 7615 61872 7991
rect 61956 7615 61990 7991
rect 62074 7615 62108 7991
rect 62192 7615 62226 7991
rect 62321 7615 62355 7791
rect 62439 7615 62473 7791
rect 62557 7615 62591 7791
rect 62675 7615 62709 7791
rect 57934 7511 57968 7545
rect 58052 7511 58086 7545
rect 51309 7443 51343 7477
rect 51427 7443 51461 7477
rect 47287 7343 47321 7377
rect 49394 7322 49428 7356
rect 40738 7255 40772 7289
rect 42845 7234 42879 7268
rect 38281 6981 38346 7128
rect 38346 6981 38348 7128
rect 38281 6979 38348 6981
rect 39701 6834 39735 7210
rect 39819 6834 39853 7210
rect 37805 6540 37839 6716
rect 37923 6540 37957 6716
rect 38041 6540 38075 6716
rect 38159 6540 38193 6716
rect 38277 6540 38311 6716
rect 38395 6540 38429 6716
rect 38513 6540 38547 6716
rect 38631 6540 38665 6716
rect 38749 6540 38783 6716
rect 39937 6834 39971 7210
rect 40055 6834 40089 7210
rect 40173 6834 40207 7210
rect 40291 6834 40325 7210
rect 40409 6834 40443 7210
rect 41599 6834 41633 7210
rect 41717 6834 41751 7210
rect 41835 6834 41869 7210
rect 41953 6834 41987 7210
rect 42071 6834 42105 7210
rect 42189 6834 42223 7210
rect 42307 6834 42341 7210
rect 44826 7218 44893 7221
rect 44826 7072 44828 7218
rect 44828 7072 44893 7218
rect 46250 6922 46284 7298
rect 46368 6922 46402 7298
rect 38867 6540 38901 6716
rect 39731 6612 39765 6646
rect 39546 6545 39580 6579
rect 40379 6612 40413 6646
rect 41629 6612 41663 6646
rect 39997 6528 40031 6562
rect 40115 6529 40149 6563
rect 40669 6544 40703 6578
rect 41444 6545 41478 6579
rect 42275 6613 42309 6647
rect 41895 6528 41929 6562
rect 42013 6529 42047 6563
rect 42567 6544 42601 6578
rect 38572 6446 38606 6480
rect 38454 6329 38488 6363
rect 39399 6302 39433 6478
rect 38042 5903 38076 6279
rect 38160 5903 38194 6279
rect 38278 5903 38312 6279
rect 38395 6103 38429 6279
rect 39517 6302 39551 6478
rect 38513 6103 38547 6279
rect 39819 6102 39853 6478
rect 39937 6102 39971 6478
rect 40055 6102 40089 6478
rect 40173 6102 40207 6478
rect 40291 6102 40325 6478
rect 40697 6302 40731 6478
rect 40815 6302 40849 6478
rect 41297 6302 41331 6478
rect 41415 6302 41449 6478
rect 41717 6102 41751 6478
rect 41835 6102 41869 6478
rect 41953 6102 41987 6478
rect 42071 6102 42105 6478
rect 42189 6102 42223 6478
rect 42595 6302 42629 6478
rect 42713 6302 42747 6478
rect 38625 5871 38774 5938
rect 38101 5819 38135 5853
rect 38219 5819 38253 5853
rect 40038 5636 40105 5785
rect 44354 6628 44388 6804
rect 44472 6628 44506 6804
rect 44590 6628 44624 6804
rect 44708 6628 44742 6804
rect 44826 6628 44860 6804
rect 44944 6628 44978 6804
rect 45062 6628 45096 6804
rect 45180 6628 45214 6804
rect 45298 6628 45332 6804
rect 46486 6922 46520 7298
rect 46604 6922 46638 7298
rect 46722 6922 46756 7298
rect 46840 6922 46874 7298
rect 46958 6922 46992 7298
rect 48148 6922 48182 7298
rect 48266 6922 48300 7298
rect 48384 6922 48418 7298
rect 48502 6922 48536 7298
rect 48620 6922 48654 7298
rect 48738 6922 48772 7298
rect 48856 6922 48890 7298
rect 45416 6628 45450 6804
rect 46280 6700 46314 6734
rect 46095 6633 46129 6667
rect 46928 6700 46962 6734
rect 48178 6700 48212 6734
rect 46546 6616 46580 6650
rect 46664 6617 46698 6651
rect 47218 6632 47252 6666
rect 47993 6633 48027 6667
rect 49517 6795 49649 6893
rect 48824 6701 48858 6735
rect 48444 6616 48478 6650
rect 48562 6617 48596 6651
rect 49116 6632 49150 6666
rect 45121 6534 45155 6568
rect 45003 6417 45037 6451
rect 45948 6390 45982 6566
rect 44591 5991 44625 6367
rect 44709 5991 44743 6367
rect 44827 5991 44861 6367
rect 44944 6191 44978 6367
rect 46066 6390 46100 6566
rect 45062 6191 45096 6367
rect 46368 6190 46402 6566
rect 46486 6190 46520 6566
rect 46604 6190 46638 6566
rect 46722 6190 46756 6566
rect 46840 6190 46874 6566
rect 47246 6390 47280 6566
rect 47364 6390 47398 6566
rect 47846 6390 47880 6566
rect 47964 6390 47998 6566
rect 48266 6190 48300 6566
rect 48384 6190 48418 6566
rect 48502 6190 48536 6566
rect 48620 6190 48654 6566
rect 48738 6190 48772 6566
rect 49144 6390 49178 6566
rect 49262 6390 49296 6566
rect 45173 5960 45322 6027
rect 44650 5907 44684 5941
rect 44768 5907 44802 5941
rect 46587 5721 46654 5870
rect 60566 7343 60600 7377
rect 62673 7322 62707 7356
rect 53941 7275 53975 7309
rect 56048 7254 56082 7288
rect 51483 7150 51550 7152
rect 51483 7003 51549 7150
rect 51549 7003 51550 7150
rect 52904 6854 52938 7230
rect 53022 6854 53056 7230
rect 51008 6560 51042 6736
rect 51126 6560 51160 6736
rect 51244 6560 51278 6736
rect 51362 6560 51396 6736
rect 51480 6560 51514 6736
rect 51598 6560 51632 6736
rect 51716 6560 51750 6736
rect 51834 6560 51868 6736
rect 51952 6560 51986 6736
rect 53140 6854 53174 7230
rect 53258 6854 53292 7230
rect 53376 6854 53410 7230
rect 53494 6854 53528 7230
rect 53612 6854 53646 7230
rect 54802 6854 54836 7230
rect 54920 6854 54954 7230
rect 55038 6854 55072 7230
rect 55156 6854 55190 7230
rect 55274 6854 55308 7230
rect 55392 6854 55426 7230
rect 55510 6854 55544 7230
rect 58108 7069 58174 7213
rect 58174 7069 58175 7213
rect 58108 7064 58175 7069
rect 59529 6922 59563 7298
rect 59647 6922 59681 7298
rect 52070 6560 52104 6736
rect 52934 6632 52968 6666
rect 52749 6565 52783 6599
rect 53582 6632 53616 6666
rect 54832 6632 54866 6666
rect 53200 6548 53234 6582
rect 53318 6549 53352 6583
rect 53872 6564 53906 6598
rect 54647 6565 54681 6599
rect 56632 6724 56728 6824
rect 55478 6633 55512 6667
rect 57633 6628 57667 6804
rect 57751 6628 57785 6804
rect 57869 6628 57903 6804
rect 57987 6628 58021 6804
rect 58105 6628 58139 6804
rect 58223 6628 58257 6804
rect 58341 6628 58375 6804
rect 58459 6628 58493 6804
rect 58577 6628 58611 6804
rect 59765 6922 59799 7298
rect 59883 6922 59917 7298
rect 60001 6922 60035 7298
rect 60119 6922 60153 7298
rect 60237 6922 60271 7298
rect 61427 6922 61461 7298
rect 61545 6922 61579 7298
rect 61663 6922 61697 7298
rect 61781 6922 61815 7298
rect 61899 6922 61933 7298
rect 62017 6922 62051 7298
rect 62135 6922 62169 7298
rect 58695 6628 58729 6804
rect 59559 6700 59593 6734
rect 59374 6633 59408 6667
rect 55098 6548 55132 6582
rect 55216 6549 55250 6583
rect 55770 6564 55804 6598
rect 60207 6700 60241 6734
rect 61457 6700 61491 6734
rect 59825 6616 59859 6650
rect 59943 6617 59977 6651
rect 60497 6632 60531 6666
rect 61272 6633 61306 6667
rect 62796 6795 62928 6893
rect 62103 6701 62137 6735
rect 61723 6616 61757 6650
rect 61841 6617 61875 6651
rect 62395 6632 62429 6666
rect 58400 6534 58434 6568
rect 51775 6466 51809 6500
rect 51657 6349 51691 6383
rect 52602 6322 52636 6498
rect 51245 5923 51279 6299
rect 51363 5923 51397 6299
rect 51481 5923 51515 6299
rect 51598 6123 51632 6299
rect 52720 6322 52754 6498
rect 51716 6123 51750 6299
rect 53022 6122 53056 6498
rect 53140 6122 53174 6498
rect 53258 6122 53292 6498
rect 53376 6122 53410 6498
rect 53494 6122 53528 6498
rect 53900 6322 53934 6498
rect 54018 6322 54052 6498
rect 54500 6322 54534 6498
rect 54618 6322 54652 6498
rect 54920 6122 54954 6498
rect 55038 6122 55072 6498
rect 55156 6122 55190 6498
rect 55274 6122 55308 6498
rect 55392 6122 55426 6498
rect 55798 6322 55832 6498
rect 55916 6322 55950 6498
rect 58282 6417 58316 6451
rect 59227 6390 59261 6566
rect 57870 5991 57904 6367
rect 57988 5991 58022 6367
rect 58106 5991 58140 6367
rect 58223 6191 58257 6367
rect 59345 6390 59379 6566
rect 58341 6191 58375 6367
rect 59647 6190 59681 6566
rect 59765 6190 59799 6566
rect 59883 6190 59917 6566
rect 60001 6190 60035 6566
rect 60119 6190 60153 6566
rect 60525 6390 60559 6566
rect 60643 6390 60677 6566
rect 61125 6390 61159 6566
rect 61243 6390 61277 6566
rect 61545 6190 61579 6566
rect 61663 6190 61697 6566
rect 61781 6190 61815 6566
rect 61899 6190 61933 6566
rect 62017 6190 62051 6566
rect 62423 6390 62457 6566
rect 62541 6390 62575 6566
rect 63762 6562 63822 6624
rect 63421 6210 63455 6386
rect 63539 6210 63573 6386
rect 63657 6210 63691 6386
rect 63775 6210 63809 6386
rect 63893 6210 63927 6386
rect 64011 6210 64045 6386
rect 64129 6210 64163 6386
rect 64247 6210 64281 6386
rect 64365 6210 64399 6386
rect 64483 6210 64517 6386
rect 64188 6116 64222 6150
rect 51827 5889 51976 5956
rect 58451 5955 58600 6022
rect 64070 5999 64104 6033
rect 57929 5907 57963 5941
rect 58047 5907 58081 5941
rect 51304 5839 51338 5873
rect 51422 5839 51456 5873
rect 53236 5655 53303 5804
rect 59867 5721 59934 5870
rect 63658 5573 63692 5949
rect 63776 5573 63810 5949
rect 63894 5573 63928 5949
rect 64011 5773 64045 5949
rect 64129 5773 64163 5949
rect 50189 5410 50259 5478
rect 56172 5404 56278 5503
rect 57281 5404 57387 5503
rect 63717 5489 63751 5523
rect 63835 5489 63869 5523
rect 63990 5366 64042 5412
rect 65661 10716 65695 11092
rect 65779 10716 65813 11092
rect 65897 10716 65931 11092
rect 66015 10716 66049 11092
rect 66133 10716 66167 11092
rect 66251 10716 66285 11092
rect 66369 10716 66403 11092
rect 66535 10796 66597 10887
rect 67264 10769 67298 11145
rect 67382 10769 67416 11145
rect 67500 10769 67534 11145
rect 67617 10969 67651 11145
rect 67735 10969 67769 11145
rect 71495 15875 71555 15924
rect 70721 15751 70897 15785
rect 70721 15633 70897 15667
rect 70721 15515 70897 15549
rect 71212 15622 71267 15680
rect 71212 15620 71267 15622
rect 70721 15397 70897 15431
rect 70521 15310 70897 15344
rect 70521 15192 70897 15226
rect 70521 15074 70897 15108
rect 70521 14956 70897 14990
rect 70521 14843 70897 14877
rect 71854 14917 72030 14951
rect 71854 14799 72030 14833
rect 70521 14725 70897 14759
rect 70521 14607 70897 14641
rect 70271 14461 70325 14533
rect 71854 14725 72230 14759
rect 71112 14665 71146 14699
rect 71496 14711 71551 14713
rect 71496 14653 71551 14711
rect 70521 14489 70897 14523
rect 71854 14607 72230 14641
rect 71211 14593 71266 14595
rect 71211 14535 71266 14593
rect 71854 14489 72230 14523
rect 70521 14371 70897 14405
rect 72331 14488 72365 14522
rect 71732 14430 71766 14464
rect 72483 14461 72497 14519
rect 72497 14461 72529 14519
rect 71854 14371 72230 14405
rect 71342 14311 71376 14345
rect 70521 14253 70897 14287
rect 71854 14253 72230 14287
rect 70521 14135 70897 14169
rect 71854 14175 72030 14209
rect 71854 14057 72030 14091
rect 70521 14016 70897 14050
rect 70521 13898 70897 13932
rect 70521 13780 70897 13814
rect 70521 13662 70897 13696
rect 70721 13543 70897 13577
rect 70721 13425 70897 13459
rect 70721 13307 70897 13341
rect 71071 13355 71105 13389
rect 70721 13189 70897 13223
rect 70721 12607 70897 12641
rect 70721 12489 70897 12523
rect 70721 12371 70897 12405
rect 71212 12478 71267 12536
rect 71212 12476 71267 12478
rect 70721 12253 70897 12287
rect 70521 12166 70897 12200
rect 70521 12048 70897 12082
rect 70521 11930 70897 11964
rect 70521 11812 70897 11846
rect 70521 11699 70897 11733
rect 71854 11773 72030 11807
rect 71854 11655 72030 11689
rect 70521 11581 70897 11615
rect 70521 11463 70897 11497
rect 70271 11317 70325 11389
rect 71854 11581 72230 11615
rect 71112 11521 71146 11555
rect 71496 11567 71551 11569
rect 71496 11509 71551 11567
rect 70521 11345 70897 11379
rect 71854 11463 72230 11497
rect 71211 11449 71266 11451
rect 71211 11391 71266 11449
rect 71854 11345 72230 11379
rect 70521 11227 70897 11261
rect 72331 11344 72365 11378
rect 71732 11286 71766 11320
rect 72483 11317 72497 11375
rect 72497 11317 72529 11375
rect 71854 11227 72230 11261
rect 71342 11167 71376 11201
rect 70521 11109 70897 11143
rect 71854 11109 72230 11143
rect 70521 10991 70897 11025
rect 71854 11031 72030 11065
rect 71854 10913 72030 10947
rect 68012 10796 68135 10890
rect 70521 10872 70897 10906
rect 70521 10754 70897 10788
rect 67323 10685 67357 10719
rect 67441 10685 67475 10719
rect 65691 10494 65725 10528
rect 65506 10427 65540 10461
rect 67596 10562 67648 10608
rect 70521 10636 70897 10670
rect 66339 10494 66373 10528
rect 70521 10518 70897 10552
rect 65957 10410 65991 10444
rect 66075 10411 66109 10445
rect 66629 10426 66663 10460
rect 70721 10399 70897 10433
rect 65359 10184 65393 10360
rect 65477 10184 65511 10360
rect 65779 9984 65813 10360
rect 65897 9984 65931 10360
rect 66015 9984 66049 10360
rect 66133 9984 66167 10360
rect 66251 9984 66285 10360
rect 66657 10184 66691 10360
rect 66775 10184 66809 10360
rect 70721 10281 70897 10315
rect 70721 10163 70897 10197
rect 71071 10211 71105 10245
rect 70721 10045 70897 10079
rect 65973 9711 66108 9813
rect 71499 9529 71559 9578
rect 65870 8198 66291 8232
rect 65870 8053 65933 8198
rect 65933 8053 66242 8198
rect 66242 8053 66291 8198
rect 65870 8032 66291 8053
rect 65236 7318 65270 7494
rect 65354 7318 65388 7494
rect 65472 7318 65506 7494
rect 65590 7318 65624 7494
rect 65720 7318 65754 7694
rect 65838 7318 65872 7694
rect 65956 7318 65990 7694
rect 66074 7318 66108 7694
rect 66192 7318 66226 7694
rect 66310 7318 66344 7694
rect 66428 7318 66462 7694
rect 67370 7667 67430 7729
rect 66557 7318 66591 7494
rect 66675 7318 66709 7494
rect 66793 7318 66827 7494
rect 66911 7318 66945 7494
rect 67029 7315 67063 7491
rect 67147 7315 67181 7491
rect 67265 7315 67299 7491
rect 67383 7315 67417 7491
rect 67501 7315 67535 7491
rect 67619 7315 67653 7491
rect 67737 7315 67771 7491
rect 67855 7315 67889 7491
rect 67973 7315 68007 7491
rect 68091 7315 68125 7491
rect 67796 7221 67830 7255
rect 66888 7102 66922 7136
rect 67678 7104 67712 7138
rect 65488 6983 65522 7017
rect 65663 6625 65697 7001
rect 65781 6625 65815 7001
rect 65899 6625 65933 7001
rect 66017 6625 66051 7001
rect 66135 6625 66169 7001
rect 66253 6625 66287 7001
rect 66371 6625 66405 7001
rect 66537 6705 66599 6796
rect 67266 6678 67300 7054
rect 67384 6678 67418 7054
rect 67502 6678 67536 7054
rect 67619 6878 67653 7054
rect 67737 6878 67771 7054
rect 67984 6973 68111 7044
rect 67325 6594 67359 6628
rect 67443 6594 67477 6628
rect 65693 6403 65727 6437
rect 65508 6336 65542 6370
rect 67598 6471 67650 6517
rect 66341 6403 66375 6437
rect 65959 6319 65993 6353
rect 66077 6320 66111 6354
rect 66631 6335 66665 6369
rect 65361 6093 65395 6269
rect 65479 6093 65513 6269
rect 65781 5893 65815 6269
rect 65899 5893 65933 6269
rect 66017 5893 66051 6269
rect 66135 5893 66169 6269
rect 66253 5893 66287 6269
rect 66659 6093 66693 6269
rect 66777 6093 66811 6269
rect 65975 5620 66110 5722
rect 38259 4604 38326 4605
rect 38259 4456 38262 4604
rect 38262 4456 38326 4604
rect 40739 4658 40806 4660
rect 40739 4511 40744 4658
rect 40744 4511 40806 4658
rect 39998 4404 40032 4438
rect 41895 4509 41958 4657
rect 41958 4509 41962 4657
rect 41895 4508 41962 4509
rect 41128 4410 41162 4444
rect 44814 4602 44881 4603
rect 44814 4454 44880 4602
rect 44880 4454 44881 4602
rect 47295 4507 47362 4656
rect 46549 4402 46583 4436
rect 48443 4507 48509 4656
rect 48509 4507 48510 4656
rect 47679 4408 47713 4442
rect 50188 4593 50258 4661
rect 39998 4286 40032 4320
rect 41128 4290 41162 4324
rect 37788 4014 37822 4190
rect 37906 4014 37940 4190
rect 38024 4014 38058 4190
rect 38142 4014 38176 4190
rect 38260 4014 38294 4190
rect 38378 4014 38412 4190
rect 38496 4014 38530 4190
rect 38614 4014 38648 4190
rect 38732 4014 38766 4190
rect 38850 4014 38884 4190
rect 38555 3920 38589 3954
rect 40113 3886 40147 4262
rect 40231 3886 40265 4262
rect 40349 3886 40383 4262
rect 40467 3886 40501 4262
rect 40585 3886 40619 4262
rect 40703 3886 40737 4262
rect 46549 4284 46583 4318
rect 40821 3886 40855 4262
rect 41255 3890 41289 4266
rect 41373 3890 41407 4266
rect 41491 3890 41525 4266
rect 41609 3890 41643 4266
rect 41727 3890 41761 4266
rect 41845 3890 41879 4266
rect 41963 3890 41997 4266
rect 47679 4288 47713 4322
rect 44339 4012 44373 4188
rect 44457 4012 44491 4188
rect 44575 4012 44609 4188
rect 44693 4012 44727 4188
rect 44811 4012 44845 4188
rect 44929 4012 44963 4188
rect 45047 4012 45081 4188
rect 45165 4012 45199 4188
rect 45283 4012 45317 4188
rect 45401 4012 45435 4188
rect 45106 3918 45140 3952
rect 46664 3884 46698 4260
rect 46782 3884 46816 4260
rect 46900 3884 46934 4260
rect 47018 3884 47052 4260
rect 47136 3884 47170 4260
rect 47254 3884 47288 4260
rect 47372 3884 47406 4260
rect 47806 3888 47840 4264
rect 47924 3888 47958 4264
rect 48042 3888 48076 4264
rect 48160 3888 48194 4264
rect 48278 3888 48312 4264
rect 48396 3888 48430 4264
rect 48514 3888 48548 4264
rect 51465 4454 51468 4600
rect 51468 4454 51532 4600
rect 51465 4451 51532 4454
rect 53950 4657 54017 4660
rect 53950 4511 54017 4657
rect 53204 4403 53238 4437
rect 55099 4508 55164 4657
rect 55164 4508 55166 4657
rect 54334 4409 54368 4443
rect 58089 4604 58156 4605
rect 58089 4456 58090 4604
rect 58090 4456 58156 4604
rect 60568 4509 60572 4653
rect 60572 4509 60635 4653
rect 60568 4504 60635 4509
rect 59826 4404 59860 4438
rect 61716 4658 61783 4659
rect 61716 4510 61719 4658
rect 61719 4510 61783 4658
rect 63833 4642 63893 4704
rect 60956 4410 60990 4444
rect 65870 4703 66291 4737
rect 65870 4558 65933 4703
rect 65933 4558 66242 4703
rect 66242 4558 66291 4703
rect 65870 4537 66291 4558
rect 53204 4285 53238 4319
rect 54334 4289 54368 4323
rect 38437 3803 38471 3837
rect 44988 3801 45022 3835
rect 38025 3377 38059 3753
rect 38143 3377 38177 3753
rect 38261 3377 38295 3753
rect 38378 3577 38412 3753
rect 38496 3577 38530 3753
rect 40318 3530 40352 3564
rect 41460 3534 41494 3568
rect 38602 3342 38751 3409
rect 38084 3293 38118 3327
rect 38202 3293 38236 3327
rect 40023 3303 40057 3479
rect 40141 3303 40175 3479
rect 40259 3303 40293 3479
rect 40377 3303 40411 3479
rect 40542 3303 40576 3479
rect 40660 3303 40694 3479
rect 40778 3303 40812 3479
rect 40896 3303 40930 3479
rect 41165 3307 41199 3483
rect 41283 3307 41317 3483
rect 41401 3307 41435 3483
rect 41519 3307 41553 3483
rect 41684 3307 41718 3483
rect 41802 3307 41836 3483
rect 41920 3307 41954 3483
rect 42038 3307 42072 3483
rect 44576 3375 44610 3751
rect 44694 3375 44728 3751
rect 44812 3375 44846 3751
rect 44929 3575 44963 3751
rect 45047 3575 45081 3751
rect 46869 3528 46903 3562
rect 48011 3532 48045 3566
rect 45152 3336 45301 3403
rect 44635 3291 44669 3325
rect 44753 3291 44787 3325
rect 46574 3301 46608 3477
rect 46692 3301 46726 3477
rect 46810 3301 46844 3477
rect 46928 3301 46962 3477
rect 47093 3301 47127 3477
rect 47211 3301 47245 3477
rect 47329 3301 47363 3477
rect 47447 3301 47481 3477
rect 47716 3305 47750 3481
rect 47834 3305 47868 3481
rect 47952 3305 47986 3481
rect 48070 3305 48104 3481
rect 48235 3305 48269 3481
rect 48353 3305 48387 3481
rect 48471 3305 48505 3481
rect 48589 3305 48623 3481
rect 38280 2805 38343 2952
rect 38343 2805 38347 2952
rect 38280 2803 38347 2805
rect 40079 2899 40146 3048
rect 41232 2894 41299 3043
rect 44825 2952 44892 2959
rect 44825 2810 44827 2952
rect 44827 2810 44892 2952
rect 46637 2896 46704 3045
rect 47778 2889 47845 3034
rect 47778 2885 47845 2889
rect 37802 2364 37836 2540
rect 37920 2364 37954 2540
rect 38038 2364 38072 2540
rect 38156 2364 38190 2540
rect 38274 2364 38308 2540
rect 38392 2364 38426 2540
rect 38510 2364 38544 2540
rect 38628 2364 38662 2540
rect 38746 2364 38780 2540
rect 38864 2364 38898 2540
rect 41986 2462 41987 2611
rect 41987 2462 42053 2611
rect 44353 2362 44387 2538
rect 44471 2362 44505 2538
rect 44589 2362 44623 2538
rect 44707 2362 44741 2538
rect 44825 2362 44859 2538
rect 44943 2362 44977 2538
rect 45061 2362 45095 2538
rect 45179 2362 45213 2538
rect 45297 2362 45331 2538
rect 45415 2362 45449 2538
rect 48542 2609 48609 2610
rect 48542 2461 48605 2609
rect 48605 2461 48609 2609
rect 38569 2270 38603 2304
rect 45120 2268 45154 2302
rect 38451 2153 38485 2187
rect 38039 1727 38073 2103
rect 38157 1727 38191 2103
rect 38275 1727 38309 2103
rect 38392 1927 38426 2103
rect 38510 1927 38544 2103
rect 38610 1692 38759 1759
rect 39266 1747 39300 1923
rect 39384 1747 39418 1923
rect 39502 1747 39536 1923
rect 39620 1747 39654 1923
rect 39750 1747 39784 2123
rect 39868 1747 39902 2123
rect 39986 1747 40020 2123
rect 40104 1747 40138 2123
rect 40222 1747 40256 2123
rect 40340 1747 40374 2123
rect 40458 1747 40492 2123
rect 40587 1747 40621 1923
rect 40705 1747 40739 1923
rect 40823 1747 40857 1923
rect 40941 1747 40975 1923
rect 41164 1747 41198 1923
rect 41282 1747 41316 1923
rect 41400 1747 41434 1923
rect 41518 1747 41552 1923
rect 41648 1747 41682 2123
rect 41766 1747 41800 2123
rect 41884 1747 41918 2123
rect 42002 1747 42036 2123
rect 42120 1747 42154 2123
rect 45002 2151 45036 2185
rect 42238 1747 42272 2123
rect 42356 1747 42390 2123
rect 42485 1747 42519 1923
rect 42603 1747 42637 1923
rect 42721 1747 42755 1923
rect 42839 1747 42873 1923
rect 44590 1725 44624 2101
rect 44708 1725 44742 2101
rect 44826 1725 44860 2101
rect 44943 1925 44977 2101
rect 45061 1925 45095 2101
rect 38098 1643 38132 1677
rect 38216 1643 38250 1677
rect 45168 1691 45317 1758
rect 45817 1745 45851 1921
rect 45935 1745 45969 1921
rect 46053 1745 46087 1921
rect 46171 1745 46205 1921
rect 46301 1745 46335 2121
rect 46419 1745 46453 2121
rect 46537 1745 46571 2121
rect 46655 1745 46689 2121
rect 46773 1745 46807 2121
rect 46891 1745 46925 2121
rect 47009 1745 47043 2121
rect 47138 1745 47172 1921
rect 47256 1745 47290 1921
rect 47374 1745 47408 1921
rect 47492 1745 47526 1921
rect 47715 1745 47749 1921
rect 47833 1745 47867 1921
rect 47951 1745 47985 1921
rect 48069 1745 48103 1921
rect 48199 1745 48233 2121
rect 48317 1745 48351 2121
rect 48435 1745 48469 2121
rect 48553 1745 48587 2121
rect 48671 1745 48705 2121
rect 48789 1745 48823 2121
rect 48907 1745 48941 2121
rect 49036 1745 49070 1921
rect 49154 1745 49188 1921
rect 49272 1745 49306 1921
rect 49390 1745 49424 1921
rect 44649 1641 44683 1675
rect 44767 1641 44801 1675
rect 40730 1475 40764 1509
rect 42837 1454 42871 1488
rect 47281 1473 47315 1507
rect 38269 1350 38336 1353
rect 38269 1204 38271 1350
rect 38271 1204 38336 1350
rect 39693 1054 39727 1430
rect 39811 1054 39845 1430
rect 37797 760 37831 936
rect 37915 760 37949 936
rect 38033 760 38067 936
rect 38151 760 38185 936
rect 38269 760 38303 936
rect 38387 760 38421 936
rect 38505 760 38539 936
rect 38623 760 38657 936
rect 38741 760 38775 936
rect 39929 1054 39963 1430
rect 40047 1054 40081 1430
rect 40165 1054 40199 1430
rect 40283 1054 40317 1430
rect 40401 1054 40435 1430
rect 41591 1054 41625 1430
rect 41709 1054 41743 1430
rect 41827 1054 41861 1430
rect 41945 1054 41979 1430
rect 42063 1054 42097 1430
rect 42181 1054 42215 1430
rect 49388 1452 49422 1486
rect 42299 1054 42333 1430
rect 44825 1199 44889 1348
rect 44889 1199 44892 1348
rect 46244 1052 46278 1428
rect 46362 1052 46396 1428
rect 38859 760 38893 936
rect 39723 832 39757 866
rect 39538 765 39572 799
rect 40371 832 40405 866
rect 41621 832 41655 866
rect 39989 748 40023 782
rect 40107 749 40141 783
rect 40661 764 40695 798
rect 41436 765 41470 799
rect 42960 927 43092 1025
rect 42267 833 42301 867
rect 41887 748 41921 782
rect 42005 749 42039 783
rect 42559 764 42593 798
rect 44348 758 44382 934
rect 44466 758 44500 934
rect 44584 758 44618 934
rect 44702 758 44736 934
rect 44820 758 44854 934
rect 44938 758 44972 934
rect 45056 758 45090 934
rect 45174 758 45208 934
rect 45292 758 45326 934
rect 46480 1052 46514 1428
rect 46598 1052 46632 1428
rect 46716 1052 46750 1428
rect 46834 1052 46868 1428
rect 46952 1052 46986 1428
rect 48142 1052 48176 1428
rect 48260 1052 48294 1428
rect 48378 1052 48412 1428
rect 48496 1052 48530 1428
rect 48614 1052 48648 1428
rect 48732 1052 48766 1428
rect 48850 1052 48884 1428
rect 45410 758 45444 934
rect 46274 830 46308 864
rect 46089 763 46123 797
rect 38564 666 38598 700
rect 38446 549 38480 583
rect 39391 522 39425 698
rect 38034 123 38068 499
rect 38152 123 38186 499
rect 38270 123 38304 499
rect 38387 323 38421 499
rect 39509 522 39543 698
rect 38505 323 38539 499
rect 39811 322 39845 698
rect 39929 322 39963 698
rect 40047 322 40081 698
rect 40165 322 40199 698
rect 40283 322 40317 698
rect 40689 522 40723 698
rect 40807 522 40841 698
rect 41289 522 41323 698
rect 41407 522 41441 698
rect 41709 322 41743 698
rect 41827 322 41861 698
rect 41945 322 41979 698
rect 42063 322 42097 698
rect 42181 322 42215 698
rect 42587 522 42621 698
rect 46922 830 46956 864
rect 48172 830 48206 864
rect 46540 746 46574 780
rect 46658 747 46692 781
rect 47212 762 47246 796
rect 47987 763 48021 797
rect 48818 831 48852 865
rect 48438 746 48472 780
rect 48556 747 48590 781
rect 49110 762 49144 796
rect 42705 522 42739 698
rect 45115 664 45149 698
rect 44997 547 45031 581
rect 45942 520 45976 696
rect 38610 100 38759 167
rect 44585 121 44619 497
rect 44703 121 44737 497
rect 44821 121 44855 497
rect 44938 321 44972 497
rect 46060 520 46094 696
rect 45056 321 45090 497
rect 46362 320 46396 696
rect 46480 320 46514 696
rect 46598 320 46632 696
rect 46716 320 46750 696
rect 46834 320 46868 696
rect 47240 520 47274 696
rect 47358 520 47392 696
rect 47840 520 47874 696
rect 47958 520 47992 696
rect 48260 320 48294 696
rect 48378 320 48412 696
rect 48496 320 48530 696
rect 48614 320 48648 696
rect 48732 320 48766 696
rect 49138 520 49172 696
rect 49256 520 49290 696
rect 38093 39 38127 73
rect 38211 39 38245 73
rect 45157 91 45306 158
rect 44644 37 44678 71
rect 44762 37 44796 71
rect 40031 -150 40098 -1
rect 46579 -151 46646 -2
rect 50994 4013 51028 4189
rect 51112 4013 51146 4189
rect 51230 4013 51264 4189
rect 51348 4013 51382 4189
rect 51466 4013 51500 4189
rect 51584 4013 51618 4189
rect 51702 4013 51736 4189
rect 51820 4013 51854 4189
rect 51938 4013 51972 4189
rect 52056 4013 52090 4189
rect 51761 3919 51795 3953
rect 53319 3885 53353 4261
rect 53437 3885 53471 4261
rect 53555 3885 53589 4261
rect 53673 3885 53707 4261
rect 53791 3885 53825 4261
rect 53909 3885 53943 4261
rect 59826 4286 59860 4320
rect 54027 3885 54061 4261
rect 54461 3889 54495 4265
rect 54579 3889 54613 4265
rect 54697 3889 54731 4265
rect 54815 3889 54849 4265
rect 54933 3889 54967 4265
rect 55051 3889 55085 4265
rect 55169 3889 55203 4265
rect 60956 4290 60990 4324
rect 57616 4014 57650 4190
rect 57734 4014 57768 4190
rect 57852 4014 57886 4190
rect 57970 4014 58004 4190
rect 58088 4014 58122 4190
rect 58206 4014 58240 4190
rect 58324 4014 58358 4190
rect 58442 4014 58476 4190
rect 58560 4014 58594 4190
rect 58678 4014 58712 4190
rect 58383 3920 58417 3954
rect 59941 3886 59975 4262
rect 60059 3886 60093 4262
rect 60177 3886 60211 4262
rect 60295 3886 60329 4262
rect 60413 3886 60447 4262
rect 60531 3886 60565 4262
rect 63492 4290 63526 4466
rect 60649 3886 60683 4262
rect 61083 3890 61117 4266
rect 61201 3890 61235 4266
rect 61319 3890 61353 4266
rect 61437 3890 61471 4266
rect 61555 3890 61589 4266
rect 61673 3890 61707 4266
rect 63610 4290 63644 4466
rect 63728 4290 63762 4466
rect 63846 4290 63880 4466
rect 63964 4290 63998 4466
rect 64082 4290 64116 4466
rect 64200 4290 64234 4466
rect 64318 4290 64352 4466
rect 64436 4290 64470 4466
rect 64554 4290 64588 4466
rect 61791 3890 61825 4266
rect 64259 4196 64293 4230
rect 64141 4079 64175 4113
rect 51643 3802 51677 3836
rect 58265 3803 58299 3837
rect 51231 3376 51265 3752
rect 51349 3376 51383 3752
rect 51467 3376 51501 3752
rect 51584 3576 51618 3752
rect 51702 3576 51736 3752
rect 53524 3529 53558 3563
rect 54666 3533 54700 3567
rect 51813 3345 51962 3412
rect 51290 3292 51324 3326
rect 51408 3292 51442 3326
rect 53229 3302 53263 3478
rect 53347 3302 53381 3478
rect 53465 3302 53499 3478
rect 53583 3302 53617 3478
rect 53748 3302 53782 3478
rect 53866 3302 53900 3478
rect 53984 3302 54018 3478
rect 54102 3302 54136 3478
rect 54371 3306 54405 3482
rect 54489 3306 54523 3482
rect 54607 3306 54641 3482
rect 54725 3306 54759 3482
rect 54890 3306 54924 3482
rect 55008 3306 55042 3482
rect 55126 3306 55160 3482
rect 55244 3306 55278 3482
rect 57853 3377 57887 3753
rect 57971 3377 58005 3753
rect 58089 3377 58123 3753
rect 58206 3577 58240 3753
rect 58324 3577 58358 3753
rect 63729 3653 63763 4029
rect 63847 3653 63881 4029
rect 63965 3653 63999 4029
rect 64082 3853 64116 4029
rect 64200 3853 64234 4029
rect 65236 3823 65270 3999
rect 65354 3823 65388 3999
rect 65472 3823 65506 3999
rect 65590 3823 65624 3999
rect 65720 3823 65754 4199
rect 65838 3823 65872 4199
rect 65956 3823 65990 4199
rect 66074 3823 66108 4199
rect 66192 3823 66226 4199
rect 66310 3823 66344 4199
rect 66428 3823 66462 4199
rect 67370 4172 67430 4234
rect 66557 3823 66591 3999
rect 66675 3823 66709 3999
rect 66793 3823 66827 3999
rect 66911 3823 66945 3999
rect 67029 3820 67063 3996
rect 67147 3820 67181 3996
rect 67265 3820 67299 3996
rect 67383 3820 67417 3996
rect 67501 3820 67535 3996
rect 67619 3820 67653 3996
rect 67737 3820 67771 3996
rect 67855 3820 67889 3996
rect 67973 3820 68007 3996
rect 68091 3820 68125 3996
rect 67796 3726 67830 3760
rect 66888 3607 66922 3641
rect 67678 3609 67712 3643
rect 63788 3569 63822 3603
rect 63906 3569 63940 3603
rect 60146 3530 60180 3564
rect 61288 3534 61322 3568
rect 58429 3350 58578 3417
rect 57912 3293 57946 3327
rect 58030 3293 58064 3327
rect 59851 3303 59885 3479
rect 59969 3303 60003 3479
rect 60087 3303 60121 3479
rect 60205 3303 60239 3479
rect 60370 3303 60404 3479
rect 60488 3303 60522 3479
rect 60606 3303 60640 3479
rect 60724 3303 60758 3479
rect 60993 3307 61027 3483
rect 61111 3307 61145 3483
rect 61229 3307 61263 3483
rect 61347 3307 61381 3483
rect 61512 3307 61546 3483
rect 61630 3307 61664 3483
rect 61748 3307 61782 3483
rect 61866 3307 61900 3483
rect 64061 3446 64113 3492
rect 65488 3488 65522 3522
rect 65663 3130 65697 3506
rect 65781 3130 65815 3506
rect 51485 2953 51552 2954
rect 51485 2805 51549 2953
rect 51549 2805 51552 2953
rect 53289 2900 53356 3049
rect 54435 2903 54502 3052
rect 58104 2954 58171 2955
rect 58104 2806 58171 2954
rect 59920 2904 59987 3053
rect 61054 2895 61121 3044
rect 65899 3130 65933 3506
rect 66017 3130 66051 3506
rect 66135 3130 66169 3506
rect 66253 3130 66287 3506
rect 66371 3130 66405 3506
rect 66537 3210 66599 3301
rect 67266 3183 67300 3559
rect 67384 3183 67418 3559
rect 67502 3183 67536 3559
rect 67619 3383 67653 3559
rect 67737 3383 67771 3559
rect 70725 9405 70901 9439
rect 70725 9287 70901 9321
rect 70725 9169 70901 9203
rect 71216 9276 71271 9334
rect 71216 9274 71271 9276
rect 70725 9051 70901 9085
rect 70525 8964 70901 8998
rect 70525 8846 70901 8880
rect 70525 8728 70901 8762
rect 70525 8610 70901 8644
rect 70525 8497 70901 8531
rect 71858 8571 72034 8605
rect 71858 8453 72034 8487
rect 70525 8379 70901 8413
rect 70525 8261 70901 8295
rect 70275 8115 70329 8187
rect 71858 8379 72234 8413
rect 71116 8319 71150 8353
rect 71500 8365 71555 8367
rect 71500 8307 71555 8365
rect 70525 8143 70901 8177
rect 71858 8261 72234 8295
rect 71215 8247 71270 8249
rect 71215 8189 71270 8247
rect 71858 8143 72234 8177
rect 70525 8025 70901 8059
rect 72335 8142 72369 8176
rect 71736 8084 71770 8118
rect 72487 8115 72501 8173
rect 72501 8115 72533 8173
rect 71858 8025 72234 8059
rect 71346 7965 71380 7999
rect 70525 7907 70901 7941
rect 71858 7907 72234 7941
rect 70525 7789 70901 7823
rect 71858 7829 72034 7863
rect 71858 7711 72034 7745
rect 70525 7670 70901 7704
rect 70525 7552 70901 7586
rect 70525 7434 70901 7468
rect 70525 7316 70901 7350
rect 70725 7197 70901 7231
rect 70725 7079 70901 7113
rect 70725 6961 70901 6995
rect 71075 7009 71109 7043
rect 70725 6843 70901 6877
rect 70725 6261 70901 6295
rect 70725 6143 70901 6177
rect 70725 6025 70901 6059
rect 71216 6132 71271 6190
rect 71216 6130 71271 6132
rect 70725 5907 70901 5941
rect 70525 5820 70901 5854
rect 70525 5702 70901 5736
rect 70525 5584 70901 5618
rect 70525 5466 70901 5500
rect 70525 5353 70901 5387
rect 71858 5427 72034 5461
rect 71858 5309 72034 5343
rect 70525 5235 70901 5269
rect 70525 5117 70901 5151
rect 70275 4971 70329 5043
rect 71858 5235 72234 5269
rect 71116 5175 71150 5209
rect 71500 5221 71555 5223
rect 71500 5163 71555 5221
rect 70525 4999 70901 5033
rect 71858 5117 72234 5151
rect 71215 5103 71270 5105
rect 71215 5045 71270 5103
rect 71858 4999 72234 5033
rect 70525 4881 70901 4915
rect 72335 4998 72369 5032
rect 71736 4940 71770 4974
rect 72487 4971 72501 5029
rect 72501 4971 72533 5029
rect 71858 4881 72234 4915
rect 71346 4821 71380 4855
rect 70525 4763 70901 4797
rect 71858 4763 72234 4797
rect 70525 4645 70901 4679
rect 71858 4685 72034 4719
rect 71858 4567 72034 4601
rect 70525 4526 70901 4560
rect 70525 4408 70901 4442
rect 70525 4290 70901 4324
rect 70525 4172 70901 4206
rect 70725 4053 70901 4087
rect 70725 3935 70901 3969
rect 70725 3817 70901 3851
rect 71075 3865 71109 3899
rect 70725 3699 70901 3733
rect 68420 3331 68486 3399
rect 68192 3216 68287 3288
rect 71495 3253 71555 3302
rect 67325 3099 67359 3133
rect 67443 3099 67477 3133
rect 70721 3129 70897 3163
rect 65693 2908 65727 2942
rect 65508 2841 65542 2875
rect 67598 2976 67650 3022
rect 66341 2908 66375 2942
rect 70721 3011 70897 3045
rect 70721 2893 70897 2927
rect 65959 2824 65993 2858
rect 66077 2825 66111 2859
rect 66631 2840 66665 2874
rect 71212 3000 71267 3058
rect 71212 2998 71267 3000
rect 51008 2363 51042 2539
rect 51126 2363 51160 2539
rect 51244 2363 51278 2539
rect 51362 2363 51396 2539
rect 51480 2363 51514 2539
rect 51598 2363 51632 2539
rect 51716 2363 51750 2539
rect 51834 2363 51868 2539
rect 51952 2363 51986 2539
rect 52070 2363 52104 2539
rect 55196 2610 55263 2612
rect 55196 2463 55260 2610
rect 55260 2463 55263 2610
rect 57630 2364 57664 2540
rect 57748 2364 57782 2540
rect 57866 2364 57900 2540
rect 57984 2364 58018 2540
rect 58102 2364 58136 2540
rect 58220 2364 58254 2540
rect 58338 2364 58372 2540
rect 58456 2364 58490 2540
rect 58574 2364 58608 2540
rect 58692 2364 58726 2540
rect 61817 2462 61882 2610
rect 61882 2462 61884 2610
rect 61817 2461 61884 2462
rect 65361 2598 65395 2774
rect 65479 2598 65513 2774
rect 65781 2398 65815 2774
rect 65899 2398 65933 2774
rect 66017 2398 66051 2774
rect 66135 2398 66169 2774
rect 66253 2398 66287 2774
rect 66659 2598 66693 2774
rect 70721 2775 70897 2809
rect 66777 2598 66811 2774
rect 70521 2688 70897 2722
rect 70521 2570 70897 2604
rect 70521 2452 70897 2486
rect 70521 2334 70897 2368
rect 51775 2269 51809 2303
rect 58397 2270 58431 2304
rect 51657 2152 51691 2186
rect 51245 1726 51279 2102
rect 51363 1726 51397 2102
rect 51481 1726 51515 2102
rect 51598 1926 51632 2102
rect 51716 1926 51750 2102
rect 51824 1694 51973 1761
rect 52472 1746 52506 1922
rect 52590 1746 52624 1922
rect 52708 1746 52742 1922
rect 52826 1746 52860 1922
rect 52956 1746 52990 2122
rect 53074 1746 53108 2122
rect 53192 1746 53226 2122
rect 53310 1746 53344 2122
rect 53428 1746 53462 2122
rect 53546 1746 53580 2122
rect 53664 1746 53698 2122
rect 53793 1746 53827 1922
rect 53911 1746 53945 1922
rect 54029 1746 54063 1922
rect 54147 1746 54181 1922
rect 54370 1746 54404 1922
rect 54488 1746 54522 1922
rect 54606 1746 54640 1922
rect 54724 1746 54758 1922
rect 54854 1746 54888 2122
rect 54972 1746 55006 2122
rect 55090 1746 55124 2122
rect 55208 1746 55242 2122
rect 55326 1746 55360 2122
rect 58279 2153 58313 2187
rect 55444 1746 55478 2122
rect 55562 1746 55596 2122
rect 55691 1746 55725 1922
rect 55809 1746 55843 1922
rect 55927 1746 55961 1922
rect 56045 1746 56079 1922
rect 57867 1727 57901 2103
rect 57985 1727 58019 2103
rect 58103 1727 58137 2103
rect 58220 1927 58254 2103
rect 58338 1927 58372 2103
rect 51304 1642 51338 1676
rect 51422 1642 51456 1676
rect 58447 1701 58596 1768
rect 59094 1747 59128 1923
rect 59212 1747 59246 1923
rect 59330 1747 59364 1923
rect 59448 1747 59482 1923
rect 59578 1747 59612 2123
rect 59696 1747 59730 2123
rect 59814 1747 59848 2123
rect 59932 1747 59966 2123
rect 60050 1747 60084 2123
rect 60168 1747 60202 2123
rect 60286 1747 60320 2123
rect 60415 1747 60449 1923
rect 60533 1747 60567 1923
rect 60651 1747 60685 1923
rect 60769 1747 60803 1923
rect 60992 1747 61026 1923
rect 61110 1747 61144 1923
rect 61228 1747 61262 1923
rect 61346 1747 61380 1923
rect 61476 1747 61510 2123
rect 61594 1747 61628 2123
rect 61712 1747 61746 2123
rect 61830 1747 61864 2123
rect 61948 1747 61982 2123
rect 62066 1747 62100 2123
rect 62184 1747 62218 2123
rect 65975 2125 66110 2227
rect 70521 2221 70897 2255
rect 71854 2295 72030 2329
rect 71854 2177 72030 2211
rect 70521 2103 70897 2137
rect 70521 1985 70897 2019
rect 62313 1747 62347 1923
rect 62431 1747 62465 1923
rect 62549 1747 62583 1923
rect 62667 1747 62701 1923
rect 70271 1839 70325 1911
rect 71854 2103 72230 2137
rect 71112 2043 71146 2077
rect 71496 2089 71551 2091
rect 71496 2031 71551 2089
rect 70521 1867 70897 1901
rect 71854 1985 72230 2019
rect 71211 1971 71266 1973
rect 71211 1913 71266 1971
rect 71854 1867 72230 1901
rect 70521 1749 70897 1783
rect 57926 1643 57960 1677
rect 58044 1643 58078 1677
rect 63830 1572 63890 1634
rect 72331 1866 72365 1900
rect 71732 1808 71766 1842
rect 72483 1839 72497 1897
rect 72497 1839 72529 1897
rect 71854 1749 72230 1783
rect 71342 1689 71376 1723
rect 70521 1631 70897 1665
rect 71854 1631 72230 1665
rect 53936 1474 53970 1508
rect 70521 1513 70897 1547
rect 56043 1453 56077 1487
rect 60558 1475 60592 1509
rect 51480 1200 51544 1346
rect 51544 1200 51547 1346
rect 51480 1197 51547 1200
rect 52899 1053 52933 1429
rect 53017 1053 53051 1429
rect 51003 759 51037 935
rect 51121 759 51155 935
rect 51239 759 51273 935
rect 51357 759 51391 935
rect 51475 759 51509 935
rect 51593 759 51627 935
rect 51711 759 51745 935
rect 51829 759 51863 935
rect 51947 759 51981 935
rect 53135 1053 53169 1429
rect 53253 1053 53287 1429
rect 53371 1053 53405 1429
rect 53489 1053 53523 1429
rect 53607 1053 53641 1429
rect 54797 1053 54831 1429
rect 54915 1053 54949 1429
rect 55033 1053 55067 1429
rect 55151 1053 55185 1429
rect 55269 1053 55303 1429
rect 55387 1053 55421 1429
rect 62665 1454 62699 1488
rect 55505 1053 55539 1429
rect 58101 1201 58166 1346
rect 58166 1201 58168 1346
rect 58101 1197 58168 1201
rect 59521 1054 59555 1430
rect 59639 1054 59673 1430
rect 52065 759 52099 935
rect 52929 831 52963 865
rect 52744 764 52778 798
rect 53577 831 53611 865
rect 54827 831 54861 865
rect 53195 747 53229 781
rect 53313 748 53347 782
rect 53867 763 53901 797
rect 54642 764 54676 798
rect 56166 926 56298 1024
rect 55473 832 55507 866
rect 55093 747 55127 781
rect 55211 748 55245 782
rect 55765 763 55799 797
rect 57625 760 57659 936
rect 57743 760 57777 936
rect 57861 760 57895 936
rect 57979 760 58013 936
rect 58097 760 58131 936
rect 58215 760 58249 936
rect 58333 760 58367 936
rect 58451 760 58485 936
rect 58569 760 58603 936
rect 59757 1054 59791 1430
rect 59875 1054 59909 1430
rect 59993 1054 60027 1430
rect 60111 1054 60145 1430
rect 60229 1054 60263 1430
rect 61419 1054 61453 1430
rect 61537 1054 61571 1430
rect 61655 1054 61689 1430
rect 61773 1054 61807 1430
rect 61891 1054 61925 1430
rect 62009 1054 62043 1430
rect 62127 1054 62161 1430
rect 63489 1220 63523 1396
rect 63607 1220 63641 1396
rect 63725 1220 63759 1396
rect 63843 1220 63877 1396
rect 63961 1220 63995 1396
rect 64079 1220 64113 1396
rect 64197 1220 64231 1396
rect 64315 1220 64349 1396
rect 64433 1220 64467 1396
rect 71854 1553 72030 1587
rect 71854 1435 72030 1469
rect 64551 1220 64585 1396
rect 70521 1394 70897 1428
rect 70521 1276 70897 1310
rect 64256 1126 64290 1160
rect 70521 1158 70897 1192
rect 58687 760 58721 936
rect 59551 832 59585 866
rect 59366 765 59400 799
rect 60199 832 60233 866
rect 61449 832 61483 866
rect 59817 748 59851 782
rect 59935 749 59969 783
rect 60489 764 60523 798
rect 61264 765 61298 799
rect 62788 927 62920 1025
rect 64138 1009 64172 1043
rect 70521 1040 70897 1074
rect 62095 833 62129 867
rect 61715 748 61749 782
rect 61833 749 61867 783
rect 62387 764 62421 798
rect 51770 665 51804 699
rect 51652 548 51686 582
rect 52597 521 52631 697
rect 51240 122 51274 498
rect 51358 122 51392 498
rect 51476 122 51510 498
rect 51593 322 51627 498
rect 52715 521 52749 697
rect 51711 322 51745 498
rect 53017 321 53051 697
rect 53135 321 53169 697
rect 53253 321 53287 697
rect 53371 321 53405 697
rect 53489 321 53523 697
rect 53895 521 53929 697
rect 54013 521 54047 697
rect 54495 521 54529 697
rect 54613 521 54647 697
rect 54915 321 54949 697
rect 55033 321 55067 697
rect 55151 321 55185 697
rect 55269 321 55303 697
rect 55387 321 55421 697
rect 55793 521 55827 697
rect 55911 521 55945 697
rect 58392 666 58426 700
rect 58274 549 58308 583
rect 59219 522 59253 698
rect 51827 85 51973 152
rect 51973 85 51976 152
rect 57862 123 57896 499
rect 57980 123 58014 499
rect 58098 123 58132 499
rect 58215 323 58249 499
rect 59337 522 59371 698
rect 58333 323 58367 499
rect 59639 322 59673 698
rect 59757 322 59791 698
rect 59875 322 59909 698
rect 59993 322 60027 698
rect 60111 322 60145 698
rect 60517 522 60551 698
rect 60635 522 60669 698
rect 61117 522 61151 698
rect 61235 522 61269 698
rect 61537 322 61571 698
rect 61655 322 61689 698
rect 61773 322 61807 698
rect 61891 322 61925 698
rect 62009 322 62043 698
rect 62415 522 62449 698
rect 62533 522 62567 698
rect 63726 583 63760 959
rect 63844 583 63878 959
rect 63962 583 63996 959
rect 64079 783 64113 959
rect 64197 783 64231 959
rect 70721 921 70897 955
rect 70721 803 70897 837
rect 70721 685 70897 719
rect 71071 733 71105 767
rect 70721 567 70897 601
rect 63785 499 63819 533
rect 63903 499 63937 533
rect 64058 376 64110 422
rect 65870 355 66291 389
rect 65870 210 65933 355
rect 65933 210 66242 355
rect 66242 210 66291 355
rect 65870 189 66291 210
rect 68555 188 68648 254
rect 51299 38 51333 72
rect 51417 38 51451 72
rect 58438 84 58587 151
rect 50188 -165 50258 -97
rect 57921 39 57955 73
rect 58039 39 58073 73
rect 71495 109 71555 158
rect 53229 -150 53296 -1
rect 59857 -144 59924 5
rect 70721 -15 70897 19
rect 65236 -525 65270 -349
rect 65354 -525 65388 -349
rect 65472 -525 65506 -349
rect 65590 -525 65624 -349
rect 65720 -525 65754 -149
rect 65838 -525 65872 -149
rect 65956 -525 65990 -149
rect 66074 -525 66108 -149
rect 66192 -525 66226 -149
rect 66310 -525 66344 -149
rect 66428 -525 66462 -149
rect 67370 -176 67430 -114
rect 70721 -133 70897 -99
rect 70721 -251 70897 -217
rect 66557 -525 66591 -349
rect 66675 -525 66709 -349
rect 66793 -525 66827 -349
rect 66911 -525 66945 -349
rect 67029 -528 67063 -352
rect 67147 -528 67181 -352
rect 67265 -528 67299 -352
rect 67383 -528 67417 -352
rect 67501 -528 67535 -352
rect 67619 -528 67653 -352
rect 67737 -528 67771 -352
rect 67855 -528 67889 -352
rect 67973 -528 68007 -352
rect 71212 -144 71267 -86
rect 71212 -146 71267 -144
rect 68091 -528 68125 -352
rect 70721 -369 70897 -335
rect 70521 -456 70897 -422
rect 67796 -622 67830 -588
rect 70521 -574 70897 -540
rect 42174 -769 42226 -723
rect 48728 -764 48780 -718
rect 55377 -776 55429 -730
rect 65216 -758 65289 -687
rect 70521 -692 70897 -658
rect 66888 -741 66922 -707
rect 67678 -739 67712 -705
rect 41901 -880 41935 -846
rect 42019 -880 42053 -846
rect 48455 -875 48489 -841
rect 48573 -875 48607 -841
rect 55104 -887 55138 -853
rect 55222 -887 55256 -853
rect 65488 -860 65522 -826
rect 41842 -1306 41876 -930
rect 41960 -1306 41994 -930
rect 42078 -1306 42112 -930
rect 42195 -1306 42229 -1130
rect 42313 -1306 42347 -1130
rect 48396 -1301 48430 -925
rect 48514 -1301 48548 -925
rect 48632 -1301 48666 -925
rect 48749 -1301 48783 -1125
rect 48867 -1301 48901 -1125
rect 55045 -1313 55079 -937
rect 55163 -1313 55197 -937
rect 55281 -1313 55315 -937
rect 55398 -1313 55432 -1137
rect 55516 -1313 55550 -1137
rect 63837 -1273 63897 -1211
rect 65663 -1218 65697 -842
rect 65781 -1218 65815 -842
rect 65899 -1218 65933 -842
rect 66017 -1218 66051 -842
rect 66135 -1218 66169 -842
rect 66253 -1218 66287 -842
rect 66371 -1218 66405 -842
rect 66537 -1138 66599 -1047
rect 67266 -1165 67300 -789
rect 67384 -1165 67418 -789
rect 67502 -1165 67536 -789
rect 67619 -965 67653 -789
rect 67737 -965 67771 -789
rect 70521 -810 70897 -776
rect 70521 -923 70897 -889
rect 71854 -849 72030 -815
rect 71854 -967 72030 -933
rect 70521 -1041 70897 -1007
rect 70521 -1159 70897 -1125
rect 67325 -1249 67359 -1215
rect 67443 -1249 67477 -1215
rect 42254 -1390 42288 -1356
rect 48808 -1385 48842 -1351
rect 55457 -1397 55491 -1363
rect 42372 -1507 42406 -1473
rect 48926 -1502 48960 -1468
rect 55575 -1514 55609 -1480
rect 41605 -1743 41639 -1567
rect 41723 -1743 41757 -1567
rect 41841 -1743 41875 -1567
rect 41959 -1743 41993 -1567
rect 42077 -1743 42111 -1567
rect 42195 -1743 42229 -1567
rect 42313 -1743 42347 -1567
rect 42431 -1743 42465 -1567
rect 42549 -1743 42583 -1567
rect 42667 -1743 42701 -1567
rect 48159 -1738 48193 -1562
rect 48277 -1738 48311 -1562
rect 48395 -1738 48429 -1562
rect 48513 -1738 48547 -1562
rect 48631 -1738 48665 -1562
rect 48749 -1738 48783 -1562
rect 48867 -1738 48901 -1562
rect 48985 -1738 49019 -1562
rect 49103 -1738 49137 -1562
rect 49221 -1738 49255 -1562
rect 54808 -1750 54842 -1574
rect 54926 -1750 54960 -1574
rect 55044 -1750 55078 -1574
rect 55162 -1750 55196 -1574
rect 55280 -1750 55314 -1574
rect 55398 -1750 55432 -1574
rect 55516 -1750 55550 -1574
rect 55634 -1750 55668 -1574
rect 55752 -1750 55786 -1574
rect 55870 -1750 55904 -1574
rect 63496 -1625 63530 -1449
rect 63614 -1625 63648 -1449
rect 63732 -1625 63766 -1449
rect 63850 -1625 63884 -1449
rect 63968 -1625 64002 -1449
rect 64086 -1625 64120 -1449
rect 64204 -1625 64238 -1449
rect 64322 -1625 64356 -1449
rect 64440 -1625 64474 -1449
rect 64558 -1625 64592 -1449
rect 65693 -1440 65727 -1406
rect 65508 -1507 65542 -1473
rect 67598 -1372 67650 -1326
rect 70271 -1305 70325 -1233
rect 71854 -1041 72230 -1007
rect 71112 -1101 71146 -1067
rect 71496 -1055 71551 -1053
rect 71496 -1113 71551 -1055
rect 70521 -1277 70897 -1243
rect 71854 -1159 72230 -1125
rect 71211 -1173 71266 -1171
rect 71211 -1231 71266 -1173
rect 71854 -1277 72230 -1243
rect 66341 -1440 66375 -1406
rect 70521 -1395 70897 -1361
rect 65959 -1524 65993 -1490
rect 66077 -1523 66111 -1489
rect 66631 -1508 66665 -1474
rect 64263 -1719 64297 -1685
rect 65361 -1750 65395 -1574
rect 65479 -1750 65513 -1574
rect 64145 -1836 64179 -1802
rect 41946 -1981 42006 -1919
rect 48500 -1976 48560 -1914
rect 55149 -1988 55209 -1926
rect 63733 -2262 63767 -1886
rect 63851 -2262 63885 -1886
rect 63969 -2262 64003 -1886
rect 64086 -2062 64120 -1886
rect 64204 -2062 64238 -1886
rect 65781 -1950 65815 -1574
rect 65899 -1950 65933 -1574
rect 66017 -1950 66051 -1574
rect 66135 -1950 66169 -1574
rect 66253 -1950 66287 -1574
rect 66659 -1750 66693 -1574
rect 66777 -1750 66811 -1574
rect 72331 -1278 72365 -1244
rect 71732 -1336 71766 -1302
rect 72483 -1305 72497 -1247
rect 72497 -1305 72529 -1247
rect 71854 -1395 72230 -1361
rect 71342 -1455 71376 -1421
rect 70521 -1513 70897 -1479
rect 71854 -1513 72230 -1479
rect 70521 -1631 70897 -1597
rect 71854 -1591 72030 -1557
rect 71854 -1709 72030 -1675
rect 70521 -1750 70897 -1716
rect 70521 -1868 70897 -1834
rect 70521 -1986 70897 -1952
rect 70521 -2104 70897 -2070
rect 65975 -2223 66110 -2121
rect 70721 -2223 70897 -2189
rect 63792 -2346 63826 -2312
rect 63910 -2346 63944 -2312
rect 70721 -2341 70897 -2307
rect 64065 -2469 64117 -2423
rect 70721 -2459 70897 -2425
rect 71071 -2411 71105 -2377
rect 70721 -2577 70897 -2543
rect 31387 -2768 31563 -2734
rect 33773 -2809 33880 -2726
rect 36506 -2798 36650 -2732
rect 31387 -2886 31563 -2852
rect 1613 -3009 1647 -2975
rect 4757 -3009 4791 -2975
rect 7889 -3005 7923 -2971
rect 11033 -3005 11067 -2971
rect 14235 -3009 14269 -2975
rect 17379 -3009 17413 -2975
rect 20511 -3005 20545 -2971
rect 23655 -3005 23689 -2971
rect 30162 -3020 30338 -2986
rect 31059 -3052 31161 -2950
rect 1126 -3273 1160 -3097
rect 1244 -3273 1278 -3097
rect 1318 -3473 1352 -3097
rect 1436 -3473 1470 -3097
rect 1554 -3473 1588 -3097
rect 1672 -3473 1706 -3097
rect 1790 -3473 1824 -3097
rect 1868 -3273 1902 -3097
rect 1986 -3273 2020 -3097
rect 4270 -3273 4304 -3097
rect 4388 -3273 4422 -3097
rect 4462 -3473 4496 -3097
rect 4580 -3473 4614 -3097
rect 4698 -3473 4732 -3097
rect 4816 -3473 4850 -3097
rect 4934 -3473 4968 -3097
rect 5012 -3273 5046 -3097
rect 5130 -3273 5164 -3097
rect 7402 -3269 7436 -3093
rect 7520 -3269 7554 -3093
rect 7594 -3469 7628 -3093
rect 7712 -3469 7746 -3093
rect 7830 -3469 7864 -3093
rect 7948 -3469 7982 -3093
rect 8066 -3469 8100 -3093
rect 8144 -3269 8178 -3093
rect 8262 -3269 8296 -3093
rect 10546 -3269 10580 -3093
rect 10664 -3269 10698 -3093
rect 10738 -3469 10772 -3093
rect 10856 -3469 10890 -3093
rect 10974 -3469 11008 -3093
rect 11092 -3469 11126 -3093
rect 11210 -3469 11244 -3093
rect 11288 -3269 11322 -3093
rect 11406 -3269 11440 -3093
rect 13748 -3273 13782 -3097
rect 13866 -3273 13900 -3097
rect 13940 -3473 13974 -3097
rect 14058 -3473 14092 -3097
rect 14176 -3473 14210 -3097
rect 14294 -3473 14328 -3097
rect 14412 -3473 14446 -3097
rect 14490 -3273 14524 -3097
rect 14608 -3273 14642 -3097
rect 16892 -3273 16926 -3097
rect 17010 -3273 17044 -3097
rect 17084 -3473 17118 -3097
rect 17202 -3473 17236 -3097
rect 17320 -3473 17354 -3097
rect 17438 -3473 17472 -3097
rect 17556 -3473 17590 -3097
rect 17634 -3273 17668 -3097
rect 17752 -3273 17786 -3097
rect 20024 -3269 20058 -3093
rect 20142 -3269 20176 -3093
rect 20216 -3469 20250 -3093
rect 20334 -3469 20368 -3093
rect 20452 -3469 20486 -3093
rect 20570 -3469 20604 -3093
rect 20688 -3469 20722 -3093
rect 20766 -3269 20800 -3093
rect 20884 -3269 20918 -3093
rect 23168 -3269 23202 -3093
rect 23286 -3269 23320 -3093
rect 23360 -3469 23394 -3093
rect 23478 -3469 23512 -3093
rect 23596 -3469 23630 -3093
rect 23714 -3469 23748 -3093
rect 23832 -3469 23866 -3093
rect 23910 -3269 23944 -3093
rect 24028 -3269 24062 -3093
rect 1555 -3608 1589 -3574
rect 4699 -3608 4733 -3574
rect 7831 -3604 7865 -3570
rect 10975 -3604 11009 -3570
rect 14177 -3608 14211 -3574
rect 17321 -3608 17355 -3574
rect 20453 -3604 20487 -3570
rect 23597 -3604 23631 -3570
rect 1558 -3740 1616 -3726
rect 1558 -3772 1616 -3740
rect 4702 -3740 4760 -3726
rect 4702 -3772 4760 -3740
rect 7834 -3736 7892 -3722
rect 7834 -3768 7892 -3736
rect 10978 -3736 11036 -3722
rect 10978 -3768 11036 -3736
rect 14180 -3740 14238 -3726
rect 14180 -3772 14238 -3740
rect 17324 -3740 17382 -3726
rect 17324 -3772 17382 -3740
rect 20456 -3736 20514 -3722
rect 20456 -3768 20514 -3736
rect 23600 -3736 23658 -3722
rect 23600 -3768 23658 -3736
<< metal1 >>
rect 38134 25229 38296 25488
rect 38133 25215 38296 25229
rect 38133 25093 38149 25215
rect 38280 25093 38296 25215
rect 38133 25043 38296 25093
rect 39997 24819 40217 24839
rect 39997 24711 40041 24819
rect 40173 24711 40217 24819
rect 41794 24777 41850 24785
rect 39997 24669 40217 24711
rect 40868 24769 41850 24777
rect 40868 24735 41810 24769
rect 41844 24735 41850 24769
rect 42513 24765 42523 24873
rect 42655 24810 42665 24873
rect 42655 24799 42667 24810
rect 42655 24765 42668 24799
rect 42924 24789 42980 24791
rect 40868 24719 41850 24735
rect 42523 24727 42668 24765
rect 40868 24718 41847 24719
rect 39601 24639 40578 24669
rect 39601 24533 39633 24639
rect 39837 24533 39869 24639
rect 40073 24533 40105 24639
rect 40309 24533 40341 24639
rect 40544 24533 40578 24639
rect 39594 24521 39640 24533
rect 39594 24345 39600 24521
rect 39634 24345 39640 24521
rect 39594 24333 39640 24345
rect 39712 24521 39758 24533
rect 39712 24345 39718 24521
rect 39752 24345 39758 24521
rect 39712 24333 39758 24345
rect 39830 24521 39876 24533
rect 39830 24345 39836 24521
rect 39870 24345 39876 24521
rect 39830 24333 39876 24345
rect 39948 24521 39994 24533
rect 39948 24345 39954 24521
rect 39988 24345 39994 24521
rect 39948 24333 39994 24345
rect 40066 24521 40112 24533
rect 40066 24345 40072 24521
rect 40106 24345 40112 24521
rect 40066 24333 40112 24345
rect 40184 24521 40230 24533
rect 40184 24345 40190 24521
rect 40224 24345 40230 24521
rect 40184 24333 40230 24345
rect 40302 24521 40348 24533
rect 40302 24345 40308 24521
rect 40342 24345 40348 24521
rect 40302 24333 40348 24345
rect 40420 24521 40466 24533
rect 40420 24345 40426 24521
rect 40460 24345 40466 24521
rect 40420 24333 40466 24345
rect 40538 24521 40584 24533
rect 40538 24345 40544 24521
rect 40578 24345 40584 24521
rect 40538 24333 40584 24345
rect 40656 24521 40702 24533
rect 40656 24345 40662 24521
rect 40696 24345 40702 24521
rect 40656 24333 40702 24345
rect 39717 24239 39753 24333
rect 39953 24239 39989 24333
rect 40189 24240 40225 24333
rect 40351 24285 40417 24292
rect 40351 24251 40367 24285
rect 40401 24251 40417 24285
rect 40351 24240 40417 24251
rect 40189 24239 40417 24240
rect 39717 24210 40417 24239
rect 39717 24209 40299 24210
rect 28279 24172 28348 24175
rect -1698 24170 -439 24172
rect 843 24171 29859 24172
rect 180 24170 29859 24171
rect -1698 24169 29859 24170
rect 34099 24169 34498 24170
rect -1698 24163 34498 24169
rect -1698 24096 28285 24163
rect 28342 24096 34498 24163
rect 39837 24096 39871 24209
rect 40233 24168 40299 24209
rect 40233 24134 40249 24168
rect 40283 24134 40299 24168
rect 40233 24127 40299 24134
rect 40661 24128 40696 24333
rect 40868 24128 40935 24718
rect 42627 24695 42668 24727
rect 42914 24723 42924 24789
rect 42980 24723 42990 24789
rect 43660 24765 43670 24873
rect 43802 24810 43812 24873
rect 46510 24816 46730 24836
rect 43802 24799 43814 24810
rect 43802 24765 43815 24799
rect 43670 24727 43815 24765
rect 43774 24699 43815 24727
rect 42043 24667 42313 24695
rect 41784 24601 41794 24667
rect 41860 24601 41870 24667
rect 42043 24605 42077 24667
rect 42279 24605 42313 24667
rect 42397 24667 42668 24695
rect 43185 24671 43455 24699
rect 42397 24605 42431 24667
rect 42633 24605 42668 24667
rect 42809 24655 42980 24671
rect 42809 24621 42940 24655
rect 42974 24621 42980 24655
rect 42809 24605 42980 24621
rect 43185 24609 43219 24671
rect 43421 24609 43455 24671
rect 43539 24671 43815 24699
rect 43539 24609 43573 24671
rect 43775 24609 43815 24671
rect 46510 24708 46554 24816
rect 46686 24708 46730 24816
rect 48307 24774 48363 24782
rect 46510 24666 46730 24708
rect 47381 24766 48363 24774
rect 47381 24732 48323 24766
rect 48357 24732 48363 24766
rect 49026 24762 49036 24870
rect 49168 24807 49178 24870
rect 49168 24796 49180 24807
rect 49168 24762 49181 24796
rect 49437 24786 49493 24788
rect 47381 24716 48363 24732
rect 49036 24724 49181 24762
rect 47381 24715 48360 24716
rect 41919 24593 41965 24605
rect 41919 24217 41925 24593
rect 41959 24217 41965 24593
rect 41919 24205 41965 24217
rect 42037 24593 42083 24605
rect 42037 24217 42043 24593
rect 42077 24217 42083 24593
rect 42037 24205 42083 24217
rect 42155 24593 42201 24605
rect 42155 24217 42161 24593
rect 42195 24217 42201 24593
rect 42155 24205 42201 24217
rect 42273 24593 42319 24605
rect 42273 24217 42279 24593
rect 42313 24217 42319 24593
rect 42273 24205 42319 24217
rect 42391 24593 42437 24605
rect 42391 24217 42397 24593
rect 42431 24217 42437 24593
rect 42391 24205 42437 24217
rect 42509 24593 42555 24605
rect 42509 24217 42515 24593
rect 42549 24217 42555 24593
rect 42509 24205 42555 24217
rect 42627 24593 42673 24605
rect 42627 24217 42633 24593
rect 42667 24217 42673 24593
rect 42627 24205 42673 24217
rect 40661 24100 40935 24128
rect 40307 24096 40935 24100
rect -1698 24089 34498 24096
rect -557 24088 1173 24089
rect -557 24087 272 24088
rect 28279 24084 28348 24089
rect 28465 24088 28654 24089
rect 28406 24053 28475 24054
rect 27903 24052 29530 24053
rect -1699 24050 -439 24052
rect 843 24051 29530 24052
rect 180 24050 29530 24051
rect -1699 24042 29530 24050
rect -1699 23975 28412 24042
rect 28469 23975 29530 24042
rect 29572 23991 34498 24089
rect -1699 23969 29530 23975
rect -557 23968 1173 23969
rect 27903 23968 29530 23969
rect -557 23967 272 23968
rect 28406 23967 28654 23968
rect 28406 23963 28475 23967
rect 28528 23934 28597 23936
rect 27918 23933 29327 23934
rect -1699 23931 -439 23933
rect 843 23932 29327 23933
rect 180 23931 29327 23932
rect -1699 23924 29327 23931
rect -1699 23857 28534 23924
rect 28591 23857 29327 23924
rect -1699 23850 29327 23857
rect -557 23849 1173 23850
rect 27918 23849 29327 23850
rect -557 23848 272 23849
rect 28465 23848 28654 23849
rect 28528 23845 28597 23848
rect 28652 23813 28721 23814
rect 27991 23812 28600 23813
rect 28644 23812 29144 23813
rect 27991 23811 29144 23812
rect -1698 23809 -439 23811
rect 843 23810 29144 23811
rect 180 23809 29144 23810
rect -1698 23802 29144 23809
rect -1698 23735 28658 23802
rect 28715 23735 29144 23802
rect -1698 23728 29144 23735
rect -557 23727 1173 23728
rect -557 23726 272 23727
rect 27991 23725 29144 23728
rect 28465 23724 28721 23725
rect 28652 23723 28721 23724
rect 28774 23694 28843 23695
rect 27770 23693 28600 23694
rect 28644 23693 28918 23694
rect 27770 23692 28918 23693
rect -1699 23690 -439 23692
rect 843 23691 28918 23692
rect 180 23690 28918 23691
rect -1699 23683 28918 23690
rect -1699 23616 28780 23683
rect 28837 23616 28918 23683
rect -1699 23609 28918 23616
rect -557 23608 1173 23609
rect 28465 23608 28654 23609
rect -557 23607 272 23608
rect 28774 23604 28918 23609
rect 27972 23571 28600 23572
rect 28644 23571 28756 23572
rect -1698 23570 -439 23571
rect 101 23570 467 23571
rect 843 23570 28756 23571
rect -1698 23522 28756 23570
rect -1698 23488 28757 23522
rect -562 23487 1173 23488
rect -1699 23451 -439 23452
rect 101 23451 467 23452
rect 843 23451 28585 23452
rect -1699 23369 28585 23451
rect -562 23368 1173 23369
rect 28491 23368 28585 23369
rect -1698 23328 -439 23329
rect 101 23328 467 23329
rect 843 23328 28456 23329
rect -1698 23246 28456 23328
rect -562 23245 1173 23246
rect -1698 22909 -1159 23000
rect -1698 22908 -439 22909
rect 101 22908 467 22909
rect 843 22908 28349 22909
rect -1698 22826 28349 22908
rect -562 22825 1173 22826
rect -1698 22785 -439 22786
rect 101 22785 467 22786
rect 843 22785 28242 22786
rect -1698 22703 28242 22785
rect -1698 22601 -1157 22703
rect -562 22702 1173 22703
rect 4270 22180 4280 22240
rect 4360 22180 4370 22240
rect 4270 22140 4370 22180
rect 7414 22180 7424 22240
rect 7504 22180 7514 22240
rect 7414 22140 7514 22180
rect 10546 22176 10556 22236
rect 10636 22176 10646 22236
rect 3364 22083 5167 22140
rect 3364 21796 3401 22083
rect 3958 21996 3992 22083
rect 5133 21996 5167 22083
rect 6508 22083 8311 22140
rect 10546 22136 10646 22176
rect 13690 22176 13700 22236
rect 13780 22176 13790 22236
rect 13690 22136 13790 22176
rect 16892 22180 16902 22240
rect 16982 22180 16992 22240
rect 16892 22140 16992 22180
rect 20036 22180 20046 22240
rect 20126 22180 20136 22240
rect 20036 22140 20136 22180
rect 23168 22176 23178 22236
rect 23258 22176 23268 22236
rect 3479 21984 3525 21996
rect 3006 21784 3052 21796
rect 3006 21608 3012 21784
rect 3046 21608 3052 21784
rect 3006 21596 3052 21608
rect 3124 21784 3170 21796
rect 3124 21608 3130 21784
rect 3164 21608 3170 21784
rect 3124 21596 3170 21608
rect 3242 21784 3288 21796
rect 3242 21608 3248 21784
rect 3282 21608 3288 21784
rect 3242 21596 3288 21608
rect 3360 21784 3406 21796
rect 3360 21608 3366 21784
rect 3400 21608 3406 21784
rect 3360 21596 3406 21608
rect 3479 21608 3485 21984
rect 3519 21608 3525 21984
rect 3479 21596 3525 21608
rect 3597 21984 3643 21996
rect 3597 21608 3603 21984
rect 3637 21608 3643 21984
rect 3597 21596 3643 21608
rect 3715 21984 3761 21996
rect 3715 21608 3721 21984
rect 3755 21608 3761 21984
rect 3715 21596 3761 21608
rect 3833 21984 3879 21996
rect 3833 21608 3839 21984
rect 3873 21608 3879 21984
rect 3833 21596 3879 21608
rect 3952 21984 3998 21996
rect 3952 21608 3958 21984
rect 3992 21608 3998 21984
rect 3952 21596 3998 21608
rect 4070 21984 4116 21996
rect 4070 21608 4076 21984
rect 4110 21608 4116 21984
rect 4070 21596 4116 21608
rect 4188 21984 4234 21996
rect 4188 21608 4194 21984
rect 4228 21608 4234 21984
rect 4188 21596 4234 21608
rect 4306 21984 4352 21996
rect 4306 21608 4312 21984
rect 4346 21608 4352 21984
rect 4306 21596 4352 21608
rect 4424 21984 4470 21996
rect 4424 21608 4430 21984
rect 4464 21608 4470 21984
rect 4424 21596 4470 21608
rect 4542 21984 4588 21996
rect 4542 21608 4548 21984
rect 4582 21608 4588 21984
rect 4542 21596 4588 21608
rect 4660 21984 4706 21996
rect 4660 21608 4666 21984
rect 4700 21608 4706 21984
rect 4660 21596 4706 21608
rect 4773 21984 4819 21996
rect 4773 21608 4779 21984
rect 4813 21608 4819 21984
rect 4773 21596 4819 21608
rect 4891 21984 4937 21996
rect 4891 21608 4897 21984
rect 4931 21608 4937 21984
rect 4891 21596 4937 21608
rect 5009 21984 5055 21996
rect 5009 21608 5015 21984
rect 5049 21608 5055 21984
rect 5009 21596 5055 21608
rect 5127 21984 5173 21996
rect 5127 21608 5133 21984
rect 5167 21796 5173 21984
rect 6508 21796 6545 22083
rect 7102 21996 7136 22083
rect 8277 21996 8311 22083
rect 9640 22079 11443 22136
rect 6623 21984 6669 21996
rect 5167 21784 5260 21796
rect 5167 21608 5220 21784
rect 5254 21608 5260 21784
rect 5127 21596 5260 21608
rect 5332 21784 5378 21796
rect 5332 21608 5338 21784
rect 5372 21608 5378 21784
rect 5332 21596 5378 21608
rect 5450 21784 5496 21796
rect 5450 21608 5456 21784
rect 5490 21608 5496 21784
rect 5450 21596 5496 21608
rect 5568 21784 5614 21796
rect 5568 21608 5574 21784
rect 5608 21608 5614 21784
rect 5568 21596 5614 21608
rect 6150 21784 6196 21796
rect 6150 21608 6156 21784
rect 6190 21608 6196 21784
rect 6150 21596 6196 21608
rect 6268 21784 6314 21796
rect 6268 21608 6274 21784
rect 6308 21608 6314 21784
rect 6268 21596 6314 21608
rect 6386 21784 6432 21796
rect 6386 21608 6392 21784
rect 6426 21608 6432 21784
rect 6386 21596 6432 21608
rect 6504 21784 6550 21796
rect 6504 21608 6510 21784
rect 6544 21608 6550 21784
rect 6504 21596 6550 21608
rect 6623 21608 6629 21984
rect 6663 21608 6669 21984
rect 6623 21596 6669 21608
rect 6741 21984 6787 21996
rect 6741 21608 6747 21984
rect 6781 21608 6787 21984
rect 6741 21596 6787 21608
rect 6859 21984 6905 21996
rect 6859 21608 6865 21984
rect 6899 21608 6905 21984
rect 6859 21596 6905 21608
rect 6977 21984 7023 21996
rect 6977 21608 6983 21984
rect 7017 21608 7023 21984
rect 6977 21596 7023 21608
rect 7096 21984 7142 21996
rect 7096 21608 7102 21984
rect 7136 21608 7142 21984
rect 7096 21596 7142 21608
rect 7214 21984 7260 21996
rect 7214 21608 7220 21984
rect 7254 21608 7260 21984
rect 7214 21596 7260 21608
rect 7332 21984 7378 21996
rect 7332 21608 7338 21984
rect 7372 21608 7378 21984
rect 7332 21596 7378 21608
rect 7450 21984 7496 21996
rect 7450 21608 7456 21984
rect 7490 21608 7496 21984
rect 7450 21596 7496 21608
rect 7568 21984 7614 21996
rect 7568 21608 7574 21984
rect 7608 21608 7614 21984
rect 7568 21596 7614 21608
rect 7686 21984 7732 21996
rect 7686 21608 7692 21984
rect 7726 21608 7732 21984
rect 7686 21596 7732 21608
rect 7804 21984 7850 21996
rect 7804 21608 7810 21984
rect 7844 21608 7850 21984
rect 7804 21596 7850 21608
rect 7917 21984 7963 21996
rect 7917 21608 7923 21984
rect 7957 21608 7963 21984
rect 7917 21596 7963 21608
rect 8035 21984 8081 21996
rect 8035 21608 8041 21984
rect 8075 21608 8081 21984
rect 8035 21596 8081 21608
rect 8153 21984 8199 21996
rect 8153 21608 8159 21984
rect 8193 21608 8199 21984
rect 8153 21596 8199 21608
rect 8271 21984 8317 21996
rect 8271 21608 8277 21984
rect 8311 21796 8317 21984
rect 8311 21784 8404 21796
rect 8311 21608 8364 21784
rect 8398 21608 8404 21784
rect 8271 21596 8404 21608
rect 8476 21784 8522 21796
rect 8476 21608 8482 21784
rect 8516 21608 8522 21784
rect 8476 21596 8522 21608
rect 8594 21784 8640 21796
rect 8594 21608 8600 21784
rect 8634 21608 8640 21784
rect 8594 21596 8640 21608
rect 8712 21784 8758 21796
rect 9640 21792 9677 22079
rect 10234 21992 10268 22079
rect 11409 21992 11443 22079
rect 12784 22079 14587 22136
rect 9755 21980 9801 21992
rect 8712 21608 8718 21784
rect 8752 21608 8758 21784
rect 8712 21596 8758 21608
rect 9282 21780 9328 21792
rect 9282 21604 9288 21780
rect 9322 21604 9328 21780
rect 3011 21242 3046 21596
rect 3485 21512 3519 21596
rect 4666 21512 4700 21596
rect 3485 21470 4700 21512
rect 3485 21450 3519 21470
rect 3162 21434 3519 21450
rect 3162 21400 3178 21434
rect 3212 21400 3519 21434
rect 5574 21410 5609 21596
rect 3162 21384 3519 21400
rect 4472 21393 5609 21410
rect 4472 21359 4488 21393
rect 4522 21359 5609 21393
rect 4472 21343 5609 21359
rect 2734 21234 3046 21242
rect 2734 21167 2748 21234
rect 2827 21167 3046 21234
rect 4342 21297 4434 21307
rect 4342 21235 4352 21297
rect 4422 21235 4434 21297
rect 4342 21222 4434 21235
rect 5427 21297 5519 21310
rect 5427 21234 5436 21297
rect 5507 21234 5519 21297
rect 5427 21225 5519 21234
rect 4122 21180 4187 21183
rect 4118 21177 4187 21180
rect 2734 21154 3046 21167
rect 3011 20834 3046 21154
rect 4112 21117 4122 21177
rect 4181 21117 4187 21177
rect 4118 21113 4187 21117
rect 4122 21111 4187 21113
rect 4460 21014 4552 21022
rect 4460 20949 4472 21014
rect 4540 20949 4552 21014
rect 4460 20937 4552 20949
rect 3011 20787 3915 20834
rect 5574 20833 5609 21343
rect 6155 21242 6190 21596
rect 6629 21512 6663 21596
rect 7810 21512 7844 21596
rect 6629 21470 7844 21512
rect 6629 21450 6663 21470
rect 6306 21434 6663 21450
rect 6306 21400 6322 21434
rect 6356 21400 6663 21434
rect 8718 21410 8753 21596
rect 9282 21592 9328 21604
rect 9400 21780 9446 21792
rect 9400 21604 9406 21780
rect 9440 21604 9446 21780
rect 9400 21592 9446 21604
rect 9518 21780 9564 21792
rect 9518 21604 9524 21780
rect 9558 21604 9564 21780
rect 9518 21592 9564 21604
rect 9636 21780 9682 21792
rect 9636 21604 9642 21780
rect 9676 21604 9682 21780
rect 9636 21592 9682 21604
rect 9755 21604 9761 21980
rect 9795 21604 9801 21980
rect 9755 21592 9801 21604
rect 9873 21980 9919 21992
rect 9873 21604 9879 21980
rect 9913 21604 9919 21980
rect 9873 21592 9919 21604
rect 9991 21980 10037 21992
rect 9991 21604 9997 21980
rect 10031 21604 10037 21980
rect 9991 21592 10037 21604
rect 10109 21980 10155 21992
rect 10109 21604 10115 21980
rect 10149 21604 10155 21980
rect 10109 21592 10155 21604
rect 10228 21980 10274 21992
rect 10228 21604 10234 21980
rect 10268 21604 10274 21980
rect 10228 21592 10274 21604
rect 10346 21980 10392 21992
rect 10346 21604 10352 21980
rect 10386 21604 10392 21980
rect 10346 21592 10392 21604
rect 10464 21980 10510 21992
rect 10464 21604 10470 21980
rect 10504 21604 10510 21980
rect 10464 21592 10510 21604
rect 10582 21980 10628 21992
rect 10582 21604 10588 21980
rect 10622 21604 10628 21980
rect 10582 21592 10628 21604
rect 10700 21980 10746 21992
rect 10700 21604 10706 21980
rect 10740 21604 10746 21980
rect 10700 21592 10746 21604
rect 10818 21980 10864 21992
rect 10818 21604 10824 21980
rect 10858 21604 10864 21980
rect 10818 21592 10864 21604
rect 10936 21980 10982 21992
rect 10936 21604 10942 21980
rect 10976 21604 10982 21980
rect 10936 21592 10982 21604
rect 11049 21980 11095 21992
rect 11049 21604 11055 21980
rect 11089 21604 11095 21980
rect 11049 21592 11095 21604
rect 11167 21980 11213 21992
rect 11167 21604 11173 21980
rect 11207 21604 11213 21980
rect 11167 21592 11213 21604
rect 11285 21980 11331 21992
rect 11285 21604 11291 21980
rect 11325 21604 11331 21980
rect 11285 21592 11331 21604
rect 11403 21980 11449 21992
rect 11403 21604 11409 21980
rect 11443 21792 11449 21980
rect 12784 21792 12821 22079
rect 13378 21992 13412 22079
rect 14553 21992 14587 22079
rect 15986 22083 17789 22140
rect 12899 21980 12945 21992
rect 11443 21780 11536 21792
rect 11443 21604 11496 21780
rect 11530 21604 11536 21780
rect 11403 21592 11536 21604
rect 11608 21780 11654 21792
rect 11608 21604 11614 21780
rect 11648 21604 11654 21780
rect 11608 21592 11654 21604
rect 11726 21780 11772 21792
rect 11726 21604 11732 21780
rect 11766 21604 11772 21780
rect 11726 21592 11772 21604
rect 11844 21780 11890 21792
rect 11844 21604 11850 21780
rect 11884 21604 11890 21780
rect 11844 21592 11890 21604
rect 12426 21780 12472 21792
rect 12426 21604 12432 21780
rect 12466 21604 12472 21780
rect 12426 21592 12472 21604
rect 12544 21780 12590 21792
rect 12544 21604 12550 21780
rect 12584 21604 12590 21780
rect 12544 21592 12590 21604
rect 12662 21780 12708 21792
rect 12662 21604 12668 21780
rect 12702 21604 12708 21780
rect 12662 21592 12708 21604
rect 12780 21780 12826 21792
rect 12780 21604 12786 21780
rect 12820 21604 12826 21780
rect 12780 21592 12826 21604
rect 12899 21604 12905 21980
rect 12939 21604 12945 21980
rect 12899 21592 12945 21604
rect 13017 21980 13063 21992
rect 13017 21604 13023 21980
rect 13057 21604 13063 21980
rect 13017 21592 13063 21604
rect 13135 21980 13181 21992
rect 13135 21604 13141 21980
rect 13175 21604 13181 21980
rect 13135 21592 13181 21604
rect 13253 21980 13299 21992
rect 13253 21604 13259 21980
rect 13293 21604 13299 21980
rect 13253 21592 13299 21604
rect 13372 21980 13418 21992
rect 13372 21604 13378 21980
rect 13412 21604 13418 21980
rect 13372 21592 13418 21604
rect 13490 21980 13536 21992
rect 13490 21604 13496 21980
rect 13530 21604 13536 21980
rect 13490 21592 13536 21604
rect 13608 21980 13654 21992
rect 13608 21604 13614 21980
rect 13648 21604 13654 21980
rect 13608 21592 13654 21604
rect 13726 21980 13772 21992
rect 13726 21604 13732 21980
rect 13766 21604 13772 21980
rect 13726 21592 13772 21604
rect 13844 21980 13890 21992
rect 13844 21604 13850 21980
rect 13884 21604 13890 21980
rect 13844 21592 13890 21604
rect 13962 21980 14008 21992
rect 13962 21604 13968 21980
rect 14002 21604 14008 21980
rect 13962 21592 14008 21604
rect 14080 21980 14126 21992
rect 14080 21604 14086 21980
rect 14120 21604 14126 21980
rect 14080 21592 14126 21604
rect 14193 21980 14239 21992
rect 14193 21604 14199 21980
rect 14233 21604 14239 21980
rect 14193 21592 14239 21604
rect 14311 21980 14357 21992
rect 14311 21604 14317 21980
rect 14351 21604 14357 21980
rect 14311 21592 14357 21604
rect 14429 21980 14475 21992
rect 14429 21604 14435 21980
rect 14469 21604 14475 21980
rect 14429 21592 14475 21604
rect 14547 21980 14593 21992
rect 14547 21604 14553 21980
rect 14587 21792 14593 21980
rect 15986 21796 16023 22083
rect 16580 21996 16614 22083
rect 17755 21996 17789 22083
rect 19130 22083 20933 22140
rect 23168 22136 23268 22176
rect 26312 22176 26322 22236
rect 26402 22176 26412 22236
rect 26312 22136 26412 22176
rect 16101 21984 16147 21996
rect 14587 21780 14680 21792
rect 14587 21604 14640 21780
rect 14674 21604 14680 21780
rect 14547 21592 14680 21604
rect 14752 21780 14798 21792
rect 14752 21604 14758 21780
rect 14792 21604 14798 21780
rect 14752 21592 14798 21604
rect 14870 21780 14916 21792
rect 14870 21604 14876 21780
rect 14910 21604 14916 21780
rect 14870 21592 14916 21604
rect 14988 21780 15034 21792
rect 14988 21604 14994 21780
rect 15028 21604 15034 21780
rect 14988 21592 15034 21604
rect 15628 21784 15674 21796
rect 15628 21608 15634 21784
rect 15668 21608 15674 21784
rect 15628 21596 15674 21608
rect 15746 21784 15792 21796
rect 15746 21608 15752 21784
rect 15786 21608 15792 21784
rect 15746 21596 15792 21608
rect 15864 21784 15910 21796
rect 15864 21608 15870 21784
rect 15904 21608 15910 21784
rect 15864 21596 15910 21608
rect 15982 21784 16028 21796
rect 15982 21608 15988 21784
rect 16022 21608 16028 21784
rect 15982 21596 16028 21608
rect 16101 21608 16107 21984
rect 16141 21608 16147 21984
rect 16101 21596 16147 21608
rect 16219 21984 16265 21996
rect 16219 21608 16225 21984
rect 16259 21608 16265 21984
rect 16219 21596 16265 21608
rect 16337 21984 16383 21996
rect 16337 21608 16343 21984
rect 16377 21608 16383 21984
rect 16337 21596 16383 21608
rect 16455 21984 16501 21996
rect 16455 21608 16461 21984
rect 16495 21608 16501 21984
rect 16455 21596 16501 21608
rect 16574 21984 16620 21996
rect 16574 21608 16580 21984
rect 16614 21608 16620 21984
rect 16574 21596 16620 21608
rect 16692 21984 16738 21996
rect 16692 21608 16698 21984
rect 16732 21608 16738 21984
rect 16692 21596 16738 21608
rect 16810 21984 16856 21996
rect 16810 21608 16816 21984
rect 16850 21608 16856 21984
rect 16810 21596 16856 21608
rect 16928 21984 16974 21996
rect 16928 21608 16934 21984
rect 16968 21608 16974 21984
rect 16928 21596 16974 21608
rect 17046 21984 17092 21996
rect 17046 21608 17052 21984
rect 17086 21608 17092 21984
rect 17046 21596 17092 21608
rect 17164 21984 17210 21996
rect 17164 21608 17170 21984
rect 17204 21608 17210 21984
rect 17164 21596 17210 21608
rect 17282 21984 17328 21996
rect 17282 21608 17288 21984
rect 17322 21608 17328 21984
rect 17282 21596 17328 21608
rect 17395 21984 17441 21996
rect 17395 21608 17401 21984
rect 17435 21608 17441 21984
rect 17395 21596 17441 21608
rect 17513 21984 17559 21996
rect 17513 21608 17519 21984
rect 17553 21608 17559 21984
rect 17513 21596 17559 21608
rect 17631 21984 17677 21996
rect 17631 21608 17637 21984
rect 17671 21608 17677 21984
rect 17631 21596 17677 21608
rect 17749 21984 17795 21996
rect 17749 21608 17755 21984
rect 17789 21796 17795 21984
rect 19130 21796 19167 22083
rect 19724 21996 19758 22083
rect 20899 21996 20933 22083
rect 22262 22079 24065 22136
rect 19245 21984 19291 21996
rect 17789 21784 17882 21796
rect 17789 21608 17842 21784
rect 17876 21608 17882 21784
rect 17749 21596 17882 21608
rect 17954 21784 18000 21796
rect 17954 21608 17960 21784
rect 17994 21608 18000 21784
rect 17954 21596 18000 21608
rect 18072 21784 18118 21796
rect 18072 21608 18078 21784
rect 18112 21608 18118 21784
rect 18072 21596 18118 21608
rect 18190 21784 18236 21796
rect 18190 21608 18196 21784
rect 18230 21608 18236 21784
rect 18190 21596 18236 21608
rect 18772 21784 18818 21796
rect 18772 21608 18778 21784
rect 18812 21608 18818 21784
rect 18772 21596 18818 21608
rect 18890 21784 18936 21796
rect 18890 21608 18896 21784
rect 18930 21608 18936 21784
rect 18890 21596 18936 21608
rect 19008 21784 19054 21796
rect 19008 21608 19014 21784
rect 19048 21608 19054 21784
rect 19008 21596 19054 21608
rect 19126 21784 19172 21796
rect 19126 21608 19132 21784
rect 19166 21608 19172 21784
rect 19126 21596 19172 21608
rect 19245 21608 19251 21984
rect 19285 21608 19291 21984
rect 19245 21596 19291 21608
rect 19363 21984 19409 21996
rect 19363 21608 19369 21984
rect 19403 21608 19409 21984
rect 19363 21596 19409 21608
rect 19481 21984 19527 21996
rect 19481 21608 19487 21984
rect 19521 21608 19527 21984
rect 19481 21596 19527 21608
rect 19599 21984 19645 21996
rect 19599 21608 19605 21984
rect 19639 21608 19645 21984
rect 19599 21596 19645 21608
rect 19718 21984 19764 21996
rect 19718 21608 19724 21984
rect 19758 21608 19764 21984
rect 19718 21596 19764 21608
rect 19836 21984 19882 21996
rect 19836 21608 19842 21984
rect 19876 21608 19882 21984
rect 19836 21596 19882 21608
rect 19954 21984 20000 21996
rect 19954 21608 19960 21984
rect 19994 21608 20000 21984
rect 19954 21596 20000 21608
rect 20072 21984 20118 21996
rect 20072 21608 20078 21984
rect 20112 21608 20118 21984
rect 20072 21596 20118 21608
rect 20190 21984 20236 21996
rect 20190 21608 20196 21984
rect 20230 21608 20236 21984
rect 20190 21596 20236 21608
rect 20308 21984 20354 21996
rect 20308 21608 20314 21984
rect 20348 21608 20354 21984
rect 20308 21596 20354 21608
rect 20426 21984 20472 21996
rect 20426 21608 20432 21984
rect 20466 21608 20472 21984
rect 20426 21596 20472 21608
rect 20539 21984 20585 21996
rect 20539 21608 20545 21984
rect 20579 21608 20585 21984
rect 20539 21596 20585 21608
rect 20657 21984 20703 21996
rect 20657 21608 20663 21984
rect 20697 21608 20703 21984
rect 20657 21596 20703 21608
rect 20775 21984 20821 21996
rect 20775 21608 20781 21984
rect 20815 21608 20821 21984
rect 20775 21596 20821 21608
rect 20893 21984 20939 21996
rect 20893 21608 20899 21984
rect 20933 21796 20939 21984
rect 20933 21784 21026 21796
rect 20933 21608 20986 21784
rect 21020 21608 21026 21784
rect 20893 21596 21026 21608
rect 21098 21784 21144 21796
rect 21098 21608 21104 21784
rect 21138 21608 21144 21784
rect 21098 21596 21144 21608
rect 21216 21784 21262 21796
rect 21216 21608 21222 21784
rect 21256 21608 21262 21784
rect 21216 21596 21262 21608
rect 21334 21784 21380 21796
rect 22262 21792 22299 22079
rect 22856 21992 22890 22079
rect 24031 21992 24065 22079
rect 25406 22079 27209 22136
rect 22377 21980 22423 21992
rect 21334 21608 21340 21784
rect 21374 21608 21380 21784
rect 21334 21596 21380 21608
rect 21904 21780 21950 21792
rect 21904 21604 21910 21780
rect 21944 21604 21950 21780
rect 6306 21384 6663 21400
rect 7616 21393 8753 21410
rect 7616 21359 7632 21393
rect 7666 21359 8753 21393
rect 7616 21343 8753 21359
rect 5692 21182 5762 21187
rect 5684 21114 5694 21182
rect 5751 21114 5762 21182
rect 6009 21147 6190 21242
rect 7486 21297 7578 21307
rect 7486 21235 7496 21297
rect 7566 21235 7578 21297
rect 7486 21222 7578 21235
rect 8571 21297 8663 21310
rect 8571 21234 8580 21297
rect 8651 21234 8663 21297
rect 8571 21225 8663 21234
rect 7266 21180 7331 21183
rect 7262 21177 7331 21180
rect 5692 21108 5762 21114
rect 6008 21096 6190 21147
rect 7256 21117 7266 21177
rect 7325 21117 7331 21177
rect 7262 21113 7331 21117
rect 7266 21111 7331 21113
rect 6008 20858 6103 21096
rect 3880 20663 3914 20787
rect 4237 20786 5609 20833
rect 6002 20801 6012 20858
rect 6065 20801 6103 20858
rect 6008 20793 6103 20801
rect 6155 20834 6190 21096
rect 7604 21014 7696 21022
rect 7604 20949 7616 21014
rect 7684 20949 7696 21014
rect 7604 20937 7696 20949
rect 6155 20787 7059 20834
rect 8718 20833 8753 21343
rect 9287 21238 9322 21592
rect 9761 21508 9795 21592
rect 10942 21508 10976 21592
rect 9761 21466 10976 21508
rect 9761 21446 9795 21466
rect 9438 21430 9795 21446
rect 9438 21396 9454 21430
rect 9488 21396 9795 21430
rect 11850 21406 11885 21592
rect 9438 21380 9795 21396
rect 10748 21389 11885 21406
rect 10748 21355 10764 21389
rect 10798 21355 11885 21389
rect 10748 21339 11885 21355
rect 8836 21182 8906 21187
rect 8828 21114 8838 21182
rect 8895 21114 8906 21182
rect 8836 21108 8906 21114
rect 9141 21092 9322 21238
rect 10618 21293 10710 21303
rect 10618 21231 10628 21293
rect 10698 21231 10710 21293
rect 10618 21218 10710 21231
rect 11703 21293 11795 21306
rect 11703 21230 11712 21293
rect 11783 21230 11795 21293
rect 11703 21221 11795 21230
rect 10398 21176 10463 21179
rect 10394 21173 10463 21176
rect 10388 21113 10398 21173
rect 10457 21113 10463 21173
rect 10394 21109 10463 21113
rect 10398 21107 10463 21109
rect 8836 21014 9012 21022
rect 8828 20946 8838 21014
rect 8895 20946 9012 21014
rect 8836 20938 9012 20946
rect 4237 20773 4303 20786
rect 4237 20739 4253 20773
rect 4287 20739 4303 20773
rect 4237 20723 4303 20739
rect 4741 20663 4775 20786
rect 7024 20663 7058 20787
rect 7381 20786 8753 20833
rect 7381 20773 7447 20786
rect 7381 20739 7397 20773
rect 7431 20739 7447 20773
rect 7381 20723 7447 20739
rect 7885 20663 7919 20786
rect 3874 20651 3920 20663
rect 3874 20475 3880 20651
rect 3914 20475 3920 20651
rect 3874 20463 3920 20475
rect 3992 20651 4116 20663
rect 3992 20475 3998 20651
rect 4032 20475 4076 20651
rect 3992 20463 4076 20475
rect 3998 20096 4032 20463
rect 4070 20275 4076 20463
rect 4110 20275 4116 20651
rect 4070 20263 4116 20275
rect 4188 20651 4234 20663
rect 4188 20275 4194 20651
rect 4228 20275 4234 20651
rect 4188 20263 4234 20275
rect 4306 20651 4352 20663
rect 4306 20275 4312 20651
rect 4346 20275 4352 20651
rect 4306 20263 4352 20275
rect 4424 20651 4470 20663
rect 4424 20275 4430 20651
rect 4464 20275 4470 20651
rect 4424 20263 4470 20275
rect 4542 20651 4662 20663
rect 4542 20275 4548 20651
rect 4582 20475 4622 20651
rect 4656 20475 4662 20651
rect 4582 20463 4662 20475
rect 4734 20651 4780 20663
rect 4734 20475 4740 20651
rect 4774 20475 4780 20651
rect 4734 20463 4780 20475
rect 7018 20651 7064 20663
rect 7018 20475 7024 20651
rect 7058 20475 7064 20651
rect 7018 20463 7064 20475
rect 7136 20651 7260 20663
rect 7136 20475 7142 20651
rect 7176 20475 7220 20651
rect 7136 20463 7220 20475
rect 4582 20275 4588 20463
rect 4542 20263 4588 20275
rect 4312 20190 4346 20263
rect 4295 20174 4361 20190
rect 4295 20140 4311 20174
rect 4345 20140 4361 20174
rect 4295 20124 4361 20140
rect 4622 20096 4656 20463
rect 3998 20044 4656 20096
rect 7142 20096 7176 20463
rect 7214 20275 7220 20463
rect 7254 20275 7260 20651
rect 7214 20263 7260 20275
rect 7332 20651 7378 20663
rect 7332 20275 7338 20651
rect 7372 20275 7378 20651
rect 7332 20263 7378 20275
rect 7450 20651 7496 20663
rect 7450 20275 7456 20651
rect 7490 20275 7496 20651
rect 7450 20263 7496 20275
rect 7568 20651 7614 20663
rect 7568 20275 7574 20651
rect 7608 20275 7614 20651
rect 7568 20263 7614 20275
rect 7686 20651 7806 20663
rect 7686 20275 7692 20651
rect 7726 20475 7766 20651
rect 7800 20475 7806 20651
rect 7726 20463 7806 20475
rect 7878 20651 7924 20663
rect 7878 20475 7884 20651
rect 7918 20475 7924 20651
rect 7878 20463 7924 20475
rect 7726 20275 7732 20463
rect 7686 20263 7732 20275
rect 7456 20190 7490 20263
rect 7439 20174 7505 20190
rect 7439 20140 7455 20174
rect 7489 20140 7505 20174
rect 7439 20124 7505 20140
rect 7766 20096 7800 20463
rect 7142 20044 7800 20096
rect 4266 20022 4358 20044
rect 4266 19970 4280 20022
rect 4346 19970 4358 20022
rect 4266 19966 4358 19970
rect 7410 20022 7502 20044
rect 7410 19970 7424 20022
rect 7490 19970 7502 20022
rect 7410 19966 7502 19970
rect 8939 19951 9012 20938
rect 9141 20731 9213 21092
rect 9287 20830 9322 21092
rect 10736 21010 10828 21018
rect 10736 20945 10748 21010
rect 10816 20945 10828 21010
rect 10736 20933 10828 20945
rect 9287 20783 10191 20830
rect 11850 20829 11885 21339
rect 12431 21238 12466 21592
rect 12905 21508 12939 21592
rect 14086 21508 14120 21592
rect 12905 21466 14120 21508
rect 12905 21446 12939 21466
rect 12582 21430 12939 21446
rect 12582 21396 12598 21430
rect 12632 21396 12939 21430
rect 14994 21406 15029 21592
rect 12582 21380 12939 21396
rect 13892 21389 15029 21406
rect 13892 21355 13908 21389
rect 13942 21355 15029 21389
rect 13892 21339 15029 21355
rect 11968 21178 12039 21183
rect 11960 21110 11970 21178
rect 12027 21110 12039 21178
rect 11968 21104 12039 21110
rect 12285 21092 12466 21238
rect 13762 21293 13854 21303
rect 13762 21231 13772 21293
rect 13842 21231 13854 21293
rect 13762 21218 13854 21231
rect 14847 21293 14939 21306
rect 14847 21230 14856 21293
rect 14927 21230 14939 21293
rect 14847 21221 14939 21230
rect 13542 21176 13607 21179
rect 13538 21173 13607 21176
rect 13532 21113 13542 21173
rect 13601 21113 13607 21173
rect 13538 21109 13607 21113
rect 13542 21107 13607 21109
rect 11968 21010 12144 21018
rect 11960 20942 11970 21010
rect 12027 20942 12144 21010
rect 11968 20934 12144 20942
rect 9136 20672 9146 20731
rect 9210 20672 9220 20731
rect 10156 20659 10190 20783
rect 10513 20782 11885 20829
rect 10513 20769 10579 20782
rect 10513 20735 10529 20769
rect 10563 20735 10579 20769
rect 10513 20719 10579 20735
rect 11017 20659 11051 20782
rect 10150 20647 10196 20659
rect 10150 20471 10156 20647
rect 10190 20471 10196 20647
rect 10150 20459 10196 20471
rect 10268 20647 10392 20659
rect 10268 20471 10274 20647
rect 10308 20471 10352 20647
rect 10268 20459 10352 20471
rect 10274 20092 10308 20459
rect 10346 20271 10352 20459
rect 10386 20271 10392 20647
rect 10346 20259 10392 20271
rect 10464 20647 10510 20659
rect 10464 20271 10470 20647
rect 10504 20271 10510 20647
rect 10464 20259 10510 20271
rect 10582 20647 10628 20659
rect 10582 20271 10588 20647
rect 10622 20271 10628 20647
rect 10582 20259 10628 20271
rect 10700 20647 10746 20659
rect 10700 20271 10706 20647
rect 10740 20271 10746 20647
rect 10700 20259 10746 20271
rect 10818 20647 10938 20659
rect 10818 20271 10824 20647
rect 10858 20471 10898 20647
rect 10932 20471 10938 20647
rect 10858 20459 10938 20471
rect 11010 20647 11056 20659
rect 11010 20471 11016 20647
rect 11050 20471 11056 20647
rect 11010 20459 11056 20471
rect 10858 20271 10864 20459
rect 10818 20259 10864 20271
rect 10588 20186 10622 20259
rect 10571 20170 10637 20186
rect 10571 20136 10587 20170
rect 10621 20136 10637 20170
rect 10571 20120 10637 20136
rect 10898 20092 10932 20459
rect 12061 20167 12144 20934
rect 12285 20578 12355 21092
rect 12431 20830 12466 21092
rect 13880 21010 13972 21018
rect 13880 20945 13892 21010
rect 13960 20945 13972 21010
rect 13880 20933 13972 20945
rect 12431 20783 13335 20830
rect 14994 20829 15029 21339
rect 15633 21242 15668 21596
rect 16107 21512 16141 21596
rect 17288 21512 17322 21596
rect 16107 21470 17322 21512
rect 16107 21450 16141 21470
rect 15784 21434 16141 21450
rect 15784 21400 15800 21434
rect 15834 21400 16141 21434
rect 18196 21410 18231 21596
rect 15784 21384 16141 21400
rect 17094 21393 18231 21410
rect 17094 21359 17110 21393
rect 17144 21359 18231 21393
rect 17094 21343 18231 21359
rect 15487 21096 15668 21242
rect 16964 21297 17056 21307
rect 16964 21235 16974 21297
rect 17044 21235 17056 21297
rect 16964 21222 17056 21235
rect 18049 21297 18141 21310
rect 18049 21234 18058 21297
rect 18129 21234 18141 21297
rect 18049 21225 18141 21234
rect 16744 21180 16809 21183
rect 16740 21177 16809 21180
rect 16734 21117 16744 21177
rect 16803 21117 16809 21177
rect 16740 21113 16809 21117
rect 16744 21111 16809 21113
rect 15112 21010 15288 21018
rect 15104 20942 15114 21010
rect 15171 20942 15288 21010
rect 15112 20934 15288 20942
rect 13300 20659 13334 20783
rect 13657 20782 15029 20829
rect 13657 20769 13723 20782
rect 13657 20735 13673 20769
rect 13707 20735 13723 20769
rect 13657 20719 13723 20735
rect 14161 20659 14195 20782
rect 13294 20647 13340 20659
rect 12280 20509 12290 20578
rect 12346 20509 12356 20578
rect 12285 20503 12355 20509
rect 13294 20471 13300 20647
rect 13334 20471 13340 20647
rect 13294 20459 13340 20471
rect 13412 20647 13536 20659
rect 13412 20471 13418 20647
rect 13452 20471 13496 20647
rect 13412 20459 13496 20471
rect 12061 20103 12084 20167
rect 12074 20100 12084 20103
rect 12141 20100 12151 20167
rect 10274 20040 10932 20092
rect 13418 20092 13452 20459
rect 13490 20271 13496 20459
rect 13530 20271 13536 20647
rect 13490 20259 13536 20271
rect 13608 20647 13654 20659
rect 13608 20271 13614 20647
rect 13648 20271 13654 20647
rect 13608 20259 13654 20271
rect 13726 20647 13772 20659
rect 13726 20271 13732 20647
rect 13766 20271 13772 20647
rect 13726 20259 13772 20271
rect 13844 20647 13890 20659
rect 13844 20271 13850 20647
rect 13884 20271 13890 20647
rect 13844 20259 13890 20271
rect 13962 20647 14082 20659
rect 13962 20271 13968 20647
rect 14002 20471 14042 20647
rect 14076 20471 14082 20647
rect 14002 20459 14082 20471
rect 14154 20647 14200 20659
rect 14154 20471 14160 20647
rect 14194 20471 14200 20647
rect 14154 20459 14200 20471
rect 14002 20271 14008 20459
rect 13962 20259 14008 20271
rect 13732 20186 13766 20259
rect 13715 20170 13781 20186
rect 13715 20136 13731 20170
rect 13765 20136 13781 20170
rect 13715 20120 13781 20136
rect 14042 20092 14076 20459
rect 15222 20302 15288 20934
rect 15488 20427 15581 21096
rect 15633 20834 15668 21096
rect 17082 21014 17174 21022
rect 17082 20949 17094 21014
rect 17162 20949 17174 21014
rect 17082 20937 17174 20949
rect 15633 20787 16537 20834
rect 18196 20833 18231 21343
rect 18777 21242 18812 21596
rect 19251 21512 19285 21596
rect 20432 21512 20466 21596
rect 19251 21470 20466 21512
rect 19251 21450 19285 21470
rect 18928 21434 19285 21450
rect 18928 21400 18944 21434
rect 18978 21400 19285 21434
rect 21340 21410 21375 21596
rect 21904 21592 21950 21604
rect 22022 21780 22068 21792
rect 22022 21604 22028 21780
rect 22062 21604 22068 21780
rect 22022 21592 22068 21604
rect 22140 21780 22186 21792
rect 22140 21604 22146 21780
rect 22180 21604 22186 21780
rect 22140 21592 22186 21604
rect 22258 21780 22304 21792
rect 22258 21604 22264 21780
rect 22298 21604 22304 21780
rect 22258 21592 22304 21604
rect 22377 21604 22383 21980
rect 22417 21604 22423 21980
rect 22377 21592 22423 21604
rect 22495 21980 22541 21992
rect 22495 21604 22501 21980
rect 22535 21604 22541 21980
rect 22495 21592 22541 21604
rect 22613 21980 22659 21992
rect 22613 21604 22619 21980
rect 22653 21604 22659 21980
rect 22613 21592 22659 21604
rect 22731 21980 22777 21992
rect 22731 21604 22737 21980
rect 22771 21604 22777 21980
rect 22731 21592 22777 21604
rect 22850 21980 22896 21992
rect 22850 21604 22856 21980
rect 22890 21604 22896 21980
rect 22850 21592 22896 21604
rect 22968 21980 23014 21992
rect 22968 21604 22974 21980
rect 23008 21604 23014 21980
rect 22968 21592 23014 21604
rect 23086 21980 23132 21992
rect 23086 21604 23092 21980
rect 23126 21604 23132 21980
rect 23086 21592 23132 21604
rect 23204 21980 23250 21992
rect 23204 21604 23210 21980
rect 23244 21604 23250 21980
rect 23204 21592 23250 21604
rect 23322 21980 23368 21992
rect 23322 21604 23328 21980
rect 23362 21604 23368 21980
rect 23322 21592 23368 21604
rect 23440 21980 23486 21992
rect 23440 21604 23446 21980
rect 23480 21604 23486 21980
rect 23440 21592 23486 21604
rect 23558 21980 23604 21992
rect 23558 21604 23564 21980
rect 23598 21604 23604 21980
rect 23558 21592 23604 21604
rect 23671 21980 23717 21992
rect 23671 21604 23677 21980
rect 23711 21604 23717 21980
rect 23671 21592 23717 21604
rect 23789 21980 23835 21992
rect 23789 21604 23795 21980
rect 23829 21604 23835 21980
rect 23789 21592 23835 21604
rect 23907 21980 23953 21992
rect 23907 21604 23913 21980
rect 23947 21604 23953 21980
rect 23907 21592 23953 21604
rect 24025 21980 24071 21992
rect 24025 21604 24031 21980
rect 24065 21792 24071 21980
rect 25406 21792 25443 22079
rect 26000 21992 26034 22079
rect 27175 21992 27209 22079
rect 25521 21980 25567 21992
rect 24065 21780 24158 21792
rect 24065 21604 24118 21780
rect 24152 21604 24158 21780
rect 24025 21592 24158 21604
rect 24230 21780 24276 21792
rect 24230 21604 24236 21780
rect 24270 21604 24276 21780
rect 24230 21592 24276 21604
rect 24348 21780 24394 21792
rect 24348 21604 24354 21780
rect 24388 21604 24394 21780
rect 24348 21592 24394 21604
rect 24466 21780 24512 21792
rect 24466 21604 24472 21780
rect 24506 21604 24512 21780
rect 24466 21592 24512 21604
rect 25048 21780 25094 21792
rect 25048 21604 25054 21780
rect 25088 21604 25094 21780
rect 25048 21592 25094 21604
rect 25166 21780 25212 21792
rect 25166 21604 25172 21780
rect 25206 21604 25212 21780
rect 25166 21592 25212 21604
rect 25284 21780 25330 21792
rect 25284 21604 25290 21780
rect 25324 21604 25330 21780
rect 25284 21592 25330 21604
rect 25402 21780 25448 21792
rect 25402 21604 25408 21780
rect 25442 21604 25448 21780
rect 25402 21592 25448 21604
rect 25521 21604 25527 21980
rect 25561 21604 25567 21980
rect 25521 21592 25567 21604
rect 25639 21980 25685 21992
rect 25639 21604 25645 21980
rect 25679 21604 25685 21980
rect 25639 21592 25685 21604
rect 25757 21980 25803 21992
rect 25757 21604 25763 21980
rect 25797 21604 25803 21980
rect 25757 21592 25803 21604
rect 25875 21980 25921 21992
rect 25875 21604 25881 21980
rect 25915 21604 25921 21980
rect 25875 21592 25921 21604
rect 25994 21980 26040 21992
rect 25994 21604 26000 21980
rect 26034 21604 26040 21980
rect 25994 21592 26040 21604
rect 26112 21980 26158 21992
rect 26112 21604 26118 21980
rect 26152 21604 26158 21980
rect 26112 21592 26158 21604
rect 26230 21980 26276 21992
rect 26230 21604 26236 21980
rect 26270 21604 26276 21980
rect 26230 21592 26276 21604
rect 26348 21980 26394 21992
rect 26348 21604 26354 21980
rect 26388 21604 26394 21980
rect 26348 21592 26394 21604
rect 26466 21980 26512 21992
rect 26466 21604 26472 21980
rect 26506 21604 26512 21980
rect 26466 21592 26512 21604
rect 26584 21980 26630 21992
rect 26584 21604 26590 21980
rect 26624 21604 26630 21980
rect 26584 21592 26630 21604
rect 26702 21980 26748 21992
rect 26702 21604 26708 21980
rect 26742 21604 26748 21980
rect 26702 21592 26748 21604
rect 26815 21980 26861 21992
rect 26815 21604 26821 21980
rect 26855 21604 26861 21980
rect 26815 21592 26861 21604
rect 26933 21980 26979 21992
rect 26933 21604 26939 21980
rect 26973 21604 26979 21980
rect 26933 21592 26979 21604
rect 27051 21980 27097 21992
rect 27051 21604 27057 21980
rect 27091 21604 27097 21980
rect 27051 21592 27097 21604
rect 27169 21980 27215 21992
rect 27169 21604 27175 21980
rect 27209 21792 27215 21980
rect 27209 21780 27302 21792
rect 27209 21604 27262 21780
rect 27296 21604 27302 21780
rect 27169 21592 27302 21604
rect 27374 21780 27420 21792
rect 27374 21604 27380 21780
rect 27414 21604 27420 21780
rect 27374 21592 27420 21604
rect 27492 21780 27538 21792
rect 27492 21604 27498 21780
rect 27532 21604 27538 21780
rect 27492 21592 27538 21604
rect 27610 21780 27656 21792
rect 27610 21604 27616 21780
rect 27650 21604 27656 21780
rect 27610 21592 27656 21604
rect 18928 21384 19285 21400
rect 20238 21393 21375 21410
rect 20238 21359 20254 21393
rect 20288 21359 21375 21393
rect 20238 21343 21375 21359
rect 18314 21182 18385 21190
rect 18306 21114 18316 21182
rect 18373 21114 18385 21182
rect 18314 21106 18385 21114
rect 18631 21096 18812 21242
rect 20108 21297 20200 21307
rect 20108 21235 20118 21297
rect 20188 21235 20200 21297
rect 20108 21222 20200 21235
rect 21193 21297 21285 21310
rect 21193 21234 21202 21297
rect 21273 21234 21285 21297
rect 21193 21225 21285 21234
rect 19888 21180 19953 21183
rect 19884 21177 19953 21180
rect 19878 21117 19888 21177
rect 19947 21117 19953 21177
rect 19884 21113 19953 21117
rect 19888 21111 19953 21113
rect 18314 21014 18490 21022
rect 18306 20946 18316 21014
rect 18373 20946 18490 21014
rect 18314 20938 18490 20946
rect 16502 20663 16536 20787
rect 16859 20786 18231 20833
rect 16859 20773 16925 20786
rect 16859 20739 16875 20773
rect 16909 20739 16925 20773
rect 16859 20723 16925 20739
rect 17363 20663 17397 20786
rect 16496 20651 16542 20663
rect 16496 20475 16502 20651
rect 16536 20475 16542 20651
rect 16496 20463 16542 20475
rect 16614 20651 16738 20663
rect 16614 20475 16620 20651
rect 16654 20475 16698 20651
rect 16614 20463 16698 20475
rect 15488 20359 15509 20427
rect 15571 20359 15581 20427
rect 15488 20354 15581 20359
rect 15213 20241 15223 20302
rect 15292 20241 15302 20302
rect 15213 20233 15302 20241
rect 13418 20040 14076 20092
rect 16620 20096 16654 20463
rect 16692 20275 16698 20463
rect 16732 20275 16738 20651
rect 16692 20263 16738 20275
rect 16810 20651 16856 20663
rect 16810 20275 16816 20651
rect 16850 20275 16856 20651
rect 16810 20263 16856 20275
rect 16928 20651 16974 20663
rect 16928 20275 16934 20651
rect 16968 20275 16974 20651
rect 16928 20263 16974 20275
rect 17046 20651 17092 20663
rect 17046 20275 17052 20651
rect 17086 20275 17092 20651
rect 17046 20263 17092 20275
rect 17164 20651 17284 20663
rect 17164 20275 17170 20651
rect 17204 20475 17244 20651
rect 17278 20475 17284 20651
rect 17204 20463 17284 20475
rect 17356 20651 17402 20663
rect 17356 20475 17362 20651
rect 17396 20475 17402 20651
rect 17356 20463 17402 20475
rect 18397 20526 18485 20938
rect 18397 20468 18408 20526
rect 18462 20468 18485 20526
rect 17204 20275 17210 20463
rect 17164 20263 17210 20275
rect 16934 20190 16968 20263
rect 16917 20174 16983 20190
rect 16917 20140 16933 20174
rect 16967 20140 16983 20174
rect 16917 20124 16983 20140
rect 17244 20096 17278 20463
rect 18397 20458 18485 20468
rect 18631 20279 18728 21096
rect 18777 20834 18812 21096
rect 20226 21014 20318 21022
rect 20226 20949 20238 21014
rect 20306 20949 20318 21014
rect 20226 20937 20318 20949
rect 18777 20787 19681 20834
rect 21340 20833 21375 21343
rect 21909 21238 21944 21592
rect 22383 21508 22417 21592
rect 23564 21508 23598 21592
rect 22383 21466 23598 21508
rect 22383 21446 22417 21466
rect 22060 21430 22417 21446
rect 22060 21396 22076 21430
rect 22110 21396 22417 21430
rect 24472 21406 24507 21592
rect 22060 21380 22417 21396
rect 23370 21389 24507 21406
rect 23370 21355 23386 21389
rect 23420 21355 24507 21389
rect 23370 21339 24507 21355
rect 24694 21343 24704 21396
rect 24764 21343 24774 21396
rect 21763 21092 21944 21238
rect 23240 21293 23332 21303
rect 23240 21231 23250 21293
rect 23320 21231 23332 21293
rect 23240 21218 23332 21231
rect 24325 21293 24417 21306
rect 24325 21230 24334 21293
rect 24405 21230 24417 21293
rect 24325 21221 24417 21230
rect 23020 21176 23085 21179
rect 23016 21173 23085 21176
rect 23010 21113 23020 21173
rect 23079 21113 23085 21173
rect 23016 21109 23085 21113
rect 23020 21107 23085 21109
rect 21458 21014 21634 21022
rect 21450 20946 21460 21014
rect 21517 20946 21634 21014
rect 21458 20938 21634 20946
rect 19646 20663 19680 20787
rect 20003 20786 21375 20833
rect 20003 20773 20069 20786
rect 20003 20739 20019 20773
rect 20053 20739 20069 20773
rect 20003 20723 20069 20739
rect 20507 20663 20541 20786
rect 19640 20651 19686 20663
rect 19640 20475 19646 20651
rect 19680 20475 19686 20651
rect 19640 20463 19686 20475
rect 19758 20651 19882 20663
rect 19758 20475 19764 20651
rect 19798 20475 19842 20651
rect 19758 20463 19842 20475
rect 18631 20222 18687 20279
rect 18746 20222 18756 20279
rect 18631 20221 18756 20222
rect 16620 20044 17278 20096
rect 19764 20096 19798 20463
rect 19836 20275 19842 20463
rect 19876 20275 19882 20651
rect 19836 20263 19882 20275
rect 19954 20651 20000 20663
rect 19954 20275 19960 20651
rect 19994 20275 20000 20651
rect 19954 20263 20000 20275
rect 20072 20651 20118 20663
rect 20072 20275 20078 20651
rect 20112 20275 20118 20651
rect 20072 20263 20118 20275
rect 20190 20651 20236 20663
rect 20190 20275 20196 20651
rect 20230 20275 20236 20651
rect 20190 20263 20236 20275
rect 20308 20651 20428 20663
rect 20308 20275 20314 20651
rect 20348 20475 20388 20651
rect 20422 20475 20428 20651
rect 20348 20463 20428 20475
rect 20500 20651 20546 20663
rect 20500 20475 20506 20651
rect 20540 20475 20546 20651
rect 21537 20631 21614 20938
rect 21530 20574 21540 20631
rect 21604 20574 21614 20631
rect 21537 20570 21614 20574
rect 20500 20463 20546 20475
rect 20348 20275 20354 20463
rect 20308 20263 20354 20275
rect 20078 20190 20112 20263
rect 20061 20174 20127 20190
rect 20061 20140 20077 20174
rect 20111 20140 20127 20174
rect 20061 20124 20127 20140
rect 20388 20096 20422 20463
rect 21763 20162 21851 21092
rect 21909 20830 21944 21092
rect 23358 21010 23450 21018
rect 23358 20945 23370 21010
rect 23438 20945 23450 21010
rect 23358 20933 23450 20945
rect 21909 20783 22813 20830
rect 24472 20829 24507 21339
rect 24703 21186 24766 21343
rect 25053 21238 25088 21592
rect 25527 21508 25561 21592
rect 26708 21508 26742 21592
rect 25527 21466 26742 21508
rect 25527 21446 25561 21466
rect 25204 21430 25561 21446
rect 25204 21396 25220 21430
rect 25254 21396 25561 21430
rect 27616 21406 27651 21592
rect 25204 21380 25561 21396
rect 26514 21389 27651 21406
rect 26514 21355 26530 21389
rect 26564 21355 27651 21389
rect 27728 21443 28055 21444
rect 27728 21381 27738 21443
rect 27792 21436 27952 21443
rect 28039 21436 28055 21443
rect 27792 21392 27950 21436
rect 28042 21392 28055 21436
rect 27792 21386 27952 21392
rect 28039 21386 28055 21392
rect 27792 21381 28055 21386
rect 26514 21339 27651 21355
rect 24590 21178 24766 21186
rect 24582 21110 24592 21178
rect 24649 21110 24766 21178
rect 24907 21120 25088 21238
rect 26384 21293 26476 21303
rect 26384 21231 26394 21293
rect 26464 21231 26476 21293
rect 26384 21218 26476 21231
rect 27469 21293 27561 21306
rect 27469 21230 27478 21293
rect 27549 21230 27561 21293
rect 27469 21221 27561 21230
rect 26164 21176 26229 21179
rect 26160 21173 26229 21176
rect 24590 21102 24766 21110
rect 24906 21092 25088 21120
rect 26154 21113 26164 21173
rect 26223 21113 26229 21173
rect 26160 21109 26229 21113
rect 26164 21107 26229 21109
rect 24590 21010 24766 21018
rect 24582 20942 24592 21010
rect 24649 20942 24766 21010
rect 24590 20934 24766 20942
rect 22778 20659 22812 20783
rect 23135 20782 24507 20829
rect 23135 20769 23201 20782
rect 23135 20735 23151 20769
rect 23185 20735 23201 20769
rect 23135 20719 23201 20735
rect 23639 20659 23673 20782
rect 24677 20772 24766 20934
rect 24674 20712 24684 20772
rect 24754 20712 24766 20772
rect 24677 20705 24766 20712
rect 22772 20647 22818 20659
rect 22772 20471 22778 20647
rect 22812 20471 22818 20647
rect 22772 20459 22818 20471
rect 22890 20647 23014 20659
rect 22890 20471 22896 20647
rect 22930 20471 22974 20647
rect 22890 20459 22974 20471
rect 21763 20096 21813 20162
rect 21872 20096 21882 20162
rect 19764 20044 20422 20096
rect 22896 20092 22930 20459
rect 22968 20271 22974 20459
rect 23008 20271 23014 20647
rect 22968 20259 23014 20271
rect 23086 20647 23132 20659
rect 23086 20271 23092 20647
rect 23126 20271 23132 20647
rect 23086 20259 23132 20271
rect 23204 20647 23250 20659
rect 23204 20271 23210 20647
rect 23244 20271 23250 20647
rect 23204 20259 23250 20271
rect 23322 20647 23368 20659
rect 23322 20271 23328 20647
rect 23362 20271 23368 20647
rect 23322 20259 23368 20271
rect 23440 20647 23560 20659
rect 23440 20271 23446 20647
rect 23480 20471 23520 20647
rect 23554 20471 23560 20647
rect 23480 20459 23560 20471
rect 23632 20647 23678 20659
rect 23632 20471 23638 20647
rect 23672 20471 23678 20647
rect 23632 20459 23678 20471
rect 23480 20271 23486 20459
rect 23440 20259 23486 20271
rect 23210 20186 23244 20259
rect 23193 20170 23259 20186
rect 23193 20136 23209 20170
rect 23243 20136 23259 20170
rect 23193 20120 23259 20136
rect 23520 20092 23554 20459
rect 10542 20018 10634 20040
rect 10542 19966 10556 20018
rect 10622 19966 10634 20018
rect 10542 19962 10634 19966
rect 13686 20018 13778 20040
rect 13686 19966 13700 20018
rect 13766 19966 13778 20018
rect 16888 20022 16980 20044
rect 16888 19970 16902 20022
rect 16968 19970 16980 20022
rect 16888 19966 16980 19970
rect 20032 20022 20124 20044
rect 22896 20040 23554 20092
rect 20032 19970 20046 20022
rect 20112 19970 20124 20022
rect 20032 19966 20124 19970
rect 23164 20018 23256 20040
rect 23164 19966 23178 20018
rect 23244 19966 23256 20018
rect 13686 19962 13778 19966
rect 23164 19962 23256 19966
rect 8932 19875 8942 19951
rect 9012 19875 9022 19951
rect 24906 19882 24967 21092
rect 25053 20830 25088 21092
rect 26502 21010 26594 21018
rect 26502 20945 26514 21010
rect 26582 20945 26594 21010
rect 26502 20933 26594 20945
rect 25053 20783 25957 20830
rect 27616 20829 27651 21339
rect 28158 21302 28242 22703
rect 27734 21294 28242 21302
rect 27726 21226 27736 21294
rect 27793 21226 28242 21294
rect 27734 21218 28242 21226
rect 27891 21018 28056 21019
rect 27734 21010 28056 21018
rect 27726 20942 27736 21010
rect 27793 21009 28056 21010
rect 27793 20998 27957 21009
rect 28037 20998 28056 21009
rect 27793 20954 27950 20998
rect 28042 20954 28056 20998
rect 27793 20947 27957 20954
rect 28037 20947 28056 20954
rect 27793 20942 28056 20947
rect 27734 20934 28056 20942
rect 27891 20933 28056 20934
rect 25922 20659 25956 20783
rect 26279 20782 27651 20829
rect 26279 20769 26345 20782
rect 26279 20735 26295 20769
rect 26329 20735 26345 20769
rect 26279 20719 26345 20735
rect 26783 20659 26817 20782
rect 27729 20768 28056 20769
rect 27729 20706 27739 20768
rect 27793 20758 28056 20768
rect 27793 20714 27950 20758
rect 28042 20714 28056 20758
rect 27793 20706 28056 20714
rect 27936 20663 28057 20671
rect 25916 20647 25962 20659
rect 25916 20471 25922 20647
rect 25956 20471 25962 20647
rect 25916 20459 25962 20471
rect 26034 20647 26158 20659
rect 26034 20471 26040 20647
rect 26074 20471 26118 20647
rect 26034 20459 26118 20471
rect 26040 20092 26074 20459
rect 26112 20271 26118 20459
rect 26152 20271 26158 20647
rect 26112 20259 26158 20271
rect 26230 20647 26276 20659
rect 26230 20271 26236 20647
rect 26270 20271 26276 20647
rect 26230 20259 26276 20271
rect 26348 20647 26394 20659
rect 26348 20271 26354 20647
rect 26388 20271 26394 20647
rect 26348 20259 26394 20271
rect 26466 20647 26512 20659
rect 26466 20271 26472 20647
rect 26506 20271 26512 20647
rect 26466 20259 26512 20271
rect 26584 20647 26704 20659
rect 26584 20271 26590 20647
rect 26624 20471 26664 20647
rect 26698 20471 26704 20647
rect 26624 20459 26704 20471
rect 26776 20647 26822 20659
rect 26776 20471 26782 20647
rect 26816 20471 26822 20647
rect 27936 20634 27956 20663
rect 27729 20633 27956 20634
rect 27729 20571 27739 20633
rect 27793 20622 27956 20633
rect 28038 20622 28057 20663
rect 27793 20578 27951 20622
rect 28043 20589 28057 20622
rect 28043 20578 28056 20589
rect 27793 20571 28056 20578
rect 26776 20459 26822 20471
rect 27727 20521 28054 20522
rect 27727 20459 27737 20521
rect 27791 20464 27949 20521
rect 28039 20512 28054 20521
rect 28042 20468 28054 20512
rect 28039 20464 28054 20468
rect 27791 20459 28054 20464
rect 26624 20271 26630 20459
rect 26584 20259 26630 20271
rect 26354 20186 26388 20259
rect 26337 20170 26403 20186
rect 26337 20136 26353 20170
rect 26387 20136 26403 20170
rect 26337 20120 26403 20136
rect 26664 20092 26698 20459
rect 27727 20396 28054 20397
rect 27727 20334 27737 20396
rect 27791 20392 28054 20396
rect 27791 20339 27945 20392
rect 28046 20339 28056 20392
rect 27791 20334 28054 20339
rect 28158 20239 28242 21218
rect 28273 20650 28349 22826
rect 28377 21177 28456 23246
rect 28494 21603 28585 23368
rect 28645 22050 28757 23488
rect 28803 22475 28918 23604
rect 29033 22909 29144 23725
rect 29221 23332 29327 23849
rect 29429 23745 29530 23968
rect 29429 23744 29729 23745
rect 29429 23656 34330 23744
rect 29429 23655 29531 23656
rect 29569 23561 34330 23656
rect 34404 23729 34498 23991
rect 39831 24084 39877 24096
rect 34404 23691 38948 23729
rect 39831 23708 39837 24084
rect 39871 23708 39877 24084
rect 39831 23696 39877 23708
rect 39949 24084 39995 24096
rect 39949 23708 39955 24084
rect 39989 23708 39995 24084
rect 39949 23696 39995 23708
rect 40067 24084 40113 24096
rect 40067 23708 40073 24084
rect 40107 23732 40113 24084
rect 40184 24084 40230 24096
rect 40184 23908 40190 24084
rect 40224 23908 40230 24084
rect 40184 23896 40230 23908
rect 40302 24084 40935 24096
rect 40302 23908 40308 24084
rect 40342 24071 40935 24084
rect 41925 24163 41959 24205
rect 42161 24163 42195 24205
rect 41925 24135 42195 24163
rect 42279 24164 42313 24205
rect 42515 24164 42549 24205
rect 42279 24135 42549 24164
rect 41925 24087 41959 24135
rect 40342 23908 40348 24071
rect 41925 24057 41988 24087
rect 40302 23896 40348 23908
rect 41953 23965 41988 24057
rect 41953 23929 42180 23965
rect 42450 23954 42460 24051
rect 42559 23954 42569 24051
rect 42633 24022 42667 24205
rect 42633 23968 42742 24022
rect 40190 23780 40225 23896
rect 41953 23822 41988 23929
rect 42114 23895 42180 23929
rect 42114 23861 42130 23895
rect 42164 23861 42180 23895
rect 42461 23953 42558 23954
rect 42461 23886 42518 23953
rect 42114 23855 42180 23861
rect 42355 23850 42624 23886
rect 42355 23822 42388 23850
rect 42591 23822 42624 23850
rect 42708 23822 42742 23968
rect 41829 23810 41875 23822
rect 40321 23780 40429 23790
rect 40190 23732 40321 23780
rect 40107 23708 40321 23732
rect 40067 23696 40321 23708
rect 40073 23692 40321 23696
rect 34404 23664 39709 23691
rect 34404 23658 39946 23664
rect 34404 23624 39896 23658
rect 39930 23624 39946 23658
rect 34404 23608 39946 23624
rect 39998 23658 40064 23664
rect 39998 23624 40014 23658
rect 40048 23624 40064 23658
rect 40247 23648 40321 23692
rect 40321 23638 40429 23648
rect 34404 23592 39709 23608
rect 34404 23591 39646 23592
rect 34404 23587 39181 23591
rect 38659 23586 38948 23587
rect 29221 23331 29710 23332
rect 29221 23198 34190 23331
rect 29221 23197 29327 23198
rect 29566 23140 34190 23198
rect 29033 22907 29635 22909
rect 33563 22907 34046 22908
rect 29033 22852 34046 22907
rect 29033 22803 33822 22852
rect 33876 22803 34046 22852
rect 29033 22802 34046 22803
rect 29033 22801 29144 22802
rect 29572 22721 34046 22802
rect 29572 22719 33627 22721
rect 28803 22431 33883 22475
rect 28803 22370 33666 22431
rect 28804 22369 33666 22370
rect 29569 22360 33666 22369
rect 33735 22360 33883 22431
rect 29569 22289 33883 22360
rect 28904 22050 28976 22051
rect 28645 22039 33744 22050
rect 28645 21963 28910 22039
rect 28970 22007 33744 22039
rect 28970 21963 33519 22007
rect 28645 21953 33519 21963
rect 28904 21951 28976 21953
rect 29566 21936 33519 21953
rect 33590 21936 33744 22007
rect 29566 21868 33744 21936
rect 28494 21602 29655 21603
rect 28494 21584 33615 21602
rect 28494 21508 29049 21584
rect 29109 21547 33615 21584
rect 29109 21508 33376 21547
rect 28494 21497 33376 21508
rect 29043 21496 29115 21497
rect 29572 21486 33376 21497
rect 33447 21486 33615 21547
rect 29572 21416 33615 21486
rect 33541 21216 33615 21416
rect 32597 21177 33482 21178
rect 28377 21165 33482 21177
rect 28377 21089 29192 21165
rect 29252 21089 33482 21165
rect 28377 21079 33482 21089
rect 29186 21077 29258 21079
rect 29569 20986 33482 21079
rect 28529 20865 28603 20867
rect 28525 20813 28535 20865
rect 28595 20813 28605 20865
rect 32575 20741 33329 20742
rect 29566 20650 33329 20741
rect 28273 20640 33329 20650
rect 28273 20586 28883 20640
rect 28274 20572 28883 20586
rect 28958 20572 33329 20640
rect 28274 20565 33329 20572
rect 32575 20563 33329 20565
rect 32590 20328 33170 20331
rect 29568 20306 33170 20328
rect 29568 20239 32926 20306
rect 28158 20222 32926 20239
rect 27722 20155 28049 20156
rect 27722 20093 27732 20155
rect 27786 20153 28049 20155
rect 28158 20154 29020 20222
rect 29090 20169 32926 20222
rect 33084 20169 33170 20306
rect 29090 20154 33170 20169
rect 27786 20150 28054 20153
rect 27786 20098 27945 20150
rect 28045 20098 28055 20150
rect 28158 20145 33170 20154
rect 28158 20144 29640 20145
rect 27786 20097 28054 20098
rect 27786 20093 28049 20097
rect 26040 20040 26698 20092
rect 26308 20018 26400 20040
rect 26308 19966 26322 20018
rect 26388 19966 26400 20018
rect 26308 19962 26400 19966
rect 27725 19933 28052 19934
rect 24906 19801 24932 19882
rect 25005 19801 25015 19882
rect 27725 19871 27735 19933
rect 27789 19929 28052 19933
rect 27789 19875 27945 19929
rect 28043 19875 28053 19929
rect 27789 19873 28053 19875
rect 29565 19907 32650 19908
rect 27789 19871 28052 19873
rect 24906 19800 24967 19801
rect 29565 19800 33035 19907
rect 28351 19793 33035 19800
rect 28351 19724 28779 19793
rect 28832 19724 33035 19793
rect 28351 19715 33035 19724
rect -1695 19562 -1391 19571
rect -1695 19498 -1493 19562
rect -1401 19498 -1391 19562
rect -1695 19488 -1391 19498
rect -1695 19447 -1391 19456
rect -1695 19383 -1493 19447
rect -1401 19383 -1391 19447
rect -1695 19373 -1391 19383
rect -1695 19326 -1391 19335
rect -1695 19262 -1493 19326
rect -1401 19262 -1391 19326
rect -1695 19252 -1391 19262
rect -1695 19207 -1391 19216
rect -1695 19143 -1493 19207
rect -1401 19143 -1391 19207
rect -1695 19133 -1391 19143
rect -1695 19093 -1391 19102
rect -1695 19029 -1493 19093
rect -1401 19029 -1391 19093
rect -1695 19019 -1391 19029
rect -1695 18979 -1391 18988
rect -1695 18915 -1493 18979
rect -1401 18915 -1391 18979
rect -1695 18905 -1391 18915
rect -1694 18864 -1390 18873
rect -1694 18800 -1492 18864
rect -1400 18800 -1390 18864
rect -1694 18790 -1390 18800
rect -1695 18750 -1390 18759
rect -1695 18686 -1492 18750
rect -1400 18686 -1390 18750
rect -1695 18676 -1390 18686
rect 28351 18646 28420 19715
rect 29562 19373 32900 19468
rect 28448 19365 32900 19373
rect 28448 19327 28671 19365
rect 27816 18636 28420 18646
rect 5302 18615 15114 18621
rect 5302 18561 15050 18615
rect 15104 18561 15114 18615
rect 27816 18577 27826 18636
rect 27886 18577 28420 18636
rect 27816 18565 28420 18577
rect 28449 19300 28671 19327
rect 28724 19300 32900 19365
rect 28449 19294 32900 19300
rect 28449 19292 29641 19294
rect 5302 18557 15114 18561
rect 4612 17046 4716 17052
rect 4612 16974 4624 17046
rect 4704 16974 4716 17046
rect 4612 16968 4716 16974
rect 5302 16970 5402 18557
rect 14929 18527 27395 18528
rect 4646 16912 4681 16968
rect 5302 16936 5318 16970
rect 5352 16936 5402 16970
rect 4520 16871 4790 16912
rect 5302 16911 5402 16936
rect 5440 18522 27395 18527
rect 5440 18468 14956 18522
rect 15010 18468 27395 18522
rect 5440 18464 27395 18468
rect 5440 18463 15020 18464
rect 4520 16808 4554 16871
rect 4756 16808 4790 16871
rect 4874 16871 5144 16899
rect 5440 16883 5504 18463
rect 6470 18430 16649 18435
rect 6470 18376 16588 18430
rect 16642 18376 16649 18430
rect 6470 18371 16649 18376
rect 5780 17046 5884 17052
rect 5780 16974 5792 17046
rect 5872 16974 5884 17046
rect 5780 16968 5884 16974
rect 6470 16970 6570 18371
rect 27000 18342 27119 18343
rect 25767 18341 27119 18342
rect 5814 16912 5849 16968
rect 6470 16936 6486 16970
rect 6520 16936 6570 16970
rect 4874 16808 4908 16871
rect 5110 16808 5144 16871
rect 5302 16862 5504 16883
rect 5302 16828 5318 16862
rect 5352 16828 5504 16862
rect 5302 16811 5504 16828
rect 5688 16871 5958 16912
rect 6470 16910 6570 16936
rect 6603 18335 27142 18341
rect 6603 18281 16413 18335
rect 16467 18281 27142 18335
rect 6603 18278 27142 18281
rect 6603 18277 16777 18278
rect 5688 16810 5722 16871
rect 5924 16810 5958 16871
rect 6042 16871 6312 16899
rect 6603 16882 6667 18277
rect 7638 18245 18113 18249
rect 7638 18191 18049 18245
rect 18103 18191 18113 18245
rect 7638 18185 18113 18191
rect 6948 17046 7052 17052
rect 6948 16974 6960 17046
rect 7040 16974 7052 17046
rect 6948 16968 7052 16974
rect 7638 16970 7738 18185
rect 17892 18155 26913 18157
rect 6982 16912 7017 16968
rect 7638 16936 7654 16970
rect 7688 16936 7738 16970
rect 6042 16810 6076 16871
rect 6278 16810 6312 16871
rect 6470 16862 6667 16882
rect 6470 16828 6486 16862
rect 6520 16828 6667 16862
rect 6470 16818 6667 16828
rect 6856 16871 7126 16912
rect 7638 16910 7738 16936
rect 7766 18151 26913 18155
rect 7766 18097 17911 18151
rect 17965 18097 26913 18151
rect 7766 18093 26913 18097
rect 7766 18091 17975 18093
rect 4514 16796 4560 16808
rect 4514 16420 4520 16796
rect 4554 16420 4560 16796
rect 4514 16408 4560 16420
rect 4632 16796 4678 16808
rect 4632 16420 4638 16796
rect 4672 16420 4678 16796
rect 4632 16408 4678 16420
rect 4750 16796 4796 16808
rect 4750 16420 4756 16796
rect 4790 16420 4796 16796
rect 4750 16408 4796 16420
rect 4868 16796 4914 16808
rect 4868 16420 4874 16796
rect 4908 16420 4914 16796
rect 4868 16408 4914 16420
rect 4986 16796 5032 16808
rect 4986 16420 4992 16796
rect 5026 16420 5032 16796
rect 4986 16408 5032 16420
rect 5104 16796 5150 16808
rect 5104 16420 5110 16796
rect 5144 16420 5150 16796
rect 5104 16408 5150 16420
rect 5222 16796 5268 16808
rect 5222 16420 5228 16796
rect 5262 16420 5268 16796
rect 5222 16408 5268 16420
rect 5682 16798 5728 16810
rect 5682 16422 5688 16798
rect 5722 16422 5728 16798
rect 5682 16410 5728 16422
rect 5800 16798 5846 16810
rect 5800 16422 5806 16798
rect 5840 16422 5846 16798
rect 5800 16410 5846 16422
rect 5918 16798 5964 16810
rect 5918 16422 5924 16798
rect 5958 16422 5964 16798
rect 5918 16410 5964 16422
rect 6036 16798 6082 16810
rect 6036 16422 6042 16798
rect 6076 16422 6082 16798
rect 6036 16410 6082 16422
rect 6154 16798 6200 16810
rect 6154 16422 6160 16798
rect 6194 16422 6200 16798
rect 6154 16410 6200 16422
rect 6272 16798 6318 16810
rect 6272 16422 6278 16798
rect 6312 16422 6318 16798
rect 6272 16410 6318 16422
rect 6390 16798 6436 16810
rect 6390 16422 6396 16798
rect 6430 16422 6436 16798
rect 6470 16730 6570 16818
rect 6856 16808 6890 16871
rect 7092 16808 7126 16871
rect 7210 16871 7480 16899
rect 7766 16882 7830 18091
rect 8806 18057 19615 18063
rect 8806 18003 19551 18057
rect 19605 18003 19615 18057
rect 8806 17999 19615 18003
rect 8806 17072 8870 17999
rect 8956 17967 19439 17969
rect 8956 17963 26741 17967
rect 8956 17909 19372 17963
rect 19426 17909 26741 17963
rect 8956 17905 19439 17909
rect 8116 17046 8220 17052
rect 8116 16974 8128 17046
rect 8208 16974 8220 17046
rect 8116 16968 8220 16974
rect 8806 16970 8906 17072
rect 8150 16912 8185 16968
rect 8806 16936 8822 16970
rect 8856 16936 8906 16970
rect 7210 16808 7244 16871
rect 7446 16808 7480 16871
rect 7638 16862 7830 16882
rect 7638 16828 7654 16862
rect 7688 16828 7830 16862
rect 7638 16818 7830 16828
rect 8024 16871 8294 16912
rect 8806 16910 8906 16936
rect 6850 16796 6896 16808
rect 6390 16410 6436 16422
rect 6850 16420 6856 16796
rect 6890 16420 6896 16796
rect 4520 16226 4554 16408
rect 4638 16368 4672 16408
rect 4874 16368 4908 16408
rect 4638 16339 4908 16368
rect 4992 16367 5026 16408
rect 5228 16367 5262 16408
rect 4992 16339 5262 16367
rect 5228 16291 5262 16339
rect 4445 16215 4554 16226
rect 5199 16261 5262 16291
rect 4445 16172 4553 16215
rect 4445 16020 4479 16172
rect 5199 16169 5234 16261
rect 5688 16226 5722 16410
rect 5806 16368 5840 16410
rect 6042 16368 6076 16410
rect 5806 16339 6076 16368
rect 6160 16367 6194 16410
rect 6396 16367 6430 16410
rect 6850 16408 6896 16420
rect 6968 16796 7014 16808
rect 6968 16420 6974 16796
rect 7008 16420 7014 16796
rect 6968 16408 7014 16420
rect 7086 16796 7132 16808
rect 7086 16420 7092 16796
rect 7126 16420 7132 16796
rect 7086 16408 7132 16420
rect 7204 16796 7250 16808
rect 7204 16420 7210 16796
rect 7244 16420 7250 16796
rect 7204 16408 7250 16420
rect 7322 16796 7368 16808
rect 7322 16420 7328 16796
rect 7362 16420 7368 16796
rect 7322 16408 7368 16420
rect 7440 16796 7486 16808
rect 7440 16420 7446 16796
rect 7480 16420 7486 16796
rect 7440 16408 7486 16420
rect 7558 16796 7604 16808
rect 7558 16420 7564 16796
rect 7598 16420 7604 16796
rect 7638 16730 7738 16818
rect 8024 16810 8058 16871
rect 8260 16810 8294 16871
rect 8378 16871 8648 16899
rect 8956 16882 9020 17905
rect 9980 17873 21071 17877
rect 9980 17819 21007 17873
rect 21061 17819 21071 17873
rect 9980 17814 21071 17819
rect 9980 17813 15025 17814
rect 9980 17070 10044 17813
rect 26464 17784 26538 17785
rect 15391 17783 26538 17784
rect 10154 17778 26538 17783
rect 10154 17724 20879 17778
rect 20933 17724 26538 17778
rect 10154 17720 26538 17724
rect 10154 17719 15118 17720
rect 9290 17044 9394 17050
rect 9290 16972 9302 17044
rect 9382 16972 9394 17044
rect 9290 16966 9394 16972
rect 9980 16968 10080 17070
rect 9324 16910 9359 16966
rect 9980 16934 9996 16968
rect 10030 16934 10080 16968
rect 8378 16810 8412 16871
rect 8614 16810 8648 16871
rect 8806 16862 9020 16882
rect 8806 16828 8822 16862
rect 8856 16828 9020 16862
rect 8806 16818 9020 16828
rect 9198 16869 9468 16910
rect 9980 16908 10080 16934
rect 8018 16798 8064 16810
rect 7558 16408 7604 16420
rect 8018 16422 8024 16798
rect 8058 16422 8064 16798
rect 8018 16410 8064 16422
rect 8136 16798 8182 16810
rect 8136 16422 8142 16798
rect 8176 16422 8182 16798
rect 8136 16410 8182 16422
rect 8254 16798 8300 16810
rect 8254 16422 8260 16798
rect 8294 16422 8300 16798
rect 8254 16410 8300 16422
rect 8372 16798 8418 16810
rect 8372 16422 8378 16798
rect 8412 16422 8418 16798
rect 8372 16410 8418 16422
rect 8490 16798 8536 16810
rect 8490 16422 8496 16798
rect 8530 16422 8536 16798
rect 8490 16410 8536 16422
rect 8608 16798 8654 16810
rect 8608 16422 8614 16798
rect 8648 16422 8654 16798
rect 8608 16410 8654 16422
rect 8726 16798 8772 16810
rect 8726 16422 8732 16798
rect 8766 16422 8772 16798
rect 8806 16730 8906 16818
rect 9198 16808 9232 16869
rect 9434 16808 9468 16869
rect 9552 16869 9822 16897
rect 10154 16880 10218 17719
rect 15388 17691 22521 17692
rect 11148 17687 22521 17691
rect 11148 17633 22460 17687
rect 22514 17633 22521 17687
rect 11148 17628 22521 17633
rect 11148 17627 14942 17628
rect 11148 17070 11212 17627
rect 15388 17597 26341 17598
rect 11325 17592 26341 17597
rect 11325 17538 22329 17592
rect 22383 17543 26341 17592
rect 22383 17538 22392 17543
rect 11325 17534 22392 17538
rect 11325 17533 14942 17534
rect 10458 17044 10562 17050
rect 10458 16972 10470 17044
rect 10550 16972 10562 17044
rect 10458 16966 10562 16972
rect 11148 16968 11248 17070
rect 10492 16910 10527 16966
rect 11148 16934 11164 16968
rect 11198 16934 11248 16968
rect 9552 16808 9586 16869
rect 9788 16808 9822 16869
rect 9980 16860 10218 16880
rect 9980 16826 9996 16860
rect 10030 16826 10218 16860
rect 9980 16816 10218 16826
rect 10366 16869 10636 16910
rect 11148 16908 11248 16934
rect 9192 16796 9238 16808
rect 8726 16410 8772 16422
rect 9192 16420 9198 16796
rect 9232 16420 9238 16796
rect 6160 16339 6430 16367
rect 6396 16291 6430 16339
rect 5007 16133 5234 16169
rect 5007 16099 5073 16133
rect 5007 16065 5023 16099
rect 5057 16065 5073 16099
rect 5007 16059 5073 16065
rect 5199 16026 5234 16133
rect 5613 16172 5722 16226
rect 6367 16261 6430 16291
rect 4563 16020 4596 16025
rect 4799 16020 4832 16024
rect 4439 16008 4485 16020
rect 4439 15832 4445 16008
rect 4479 15832 4485 16008
rect 4439 15820 4485 15832
rect 4557 16008 4603 16020
rect 4557 15832 4563 16008
rect 4597 15832 4603 16008
rect 4557 15820 4603 15832
rect 4675 16008 4721 16020
rect 4675 15832 4681 16008
rect 4715 15832 4721 16008
rect 4675 15820 4721 15832
rect 4793 16008 4839 16020
rect 4793 15832 4799 16008
rect 4833 15959 4839 16008
rect 4958 16014 5004 16026
rect 4958 15959 4964 16014
rect 4833 15871 4964 15959
rect 4833 15832 4839 15871
rect 4793 15820 4839 15832
rect 4958 15838 4964 15871
rect 4998 15838 5004 16014
rect 4958 15826 5004 15838
rect 5076 16014 5122 16026
rect 5076 15838 5082 16014
rect 5116 15838 5122 16014
rect 5076 15826 5122 15838
rect 5194 16014 5240 16026
rect 5194 15838 5200 16014
rect 5234 15838 5240 16014
rect 5194 15826 5240 15838
rect 5312 16014 5358 16026
rect 5613 16019 5647 16172
rect 6367 16169 6402 16261
rect 6856 16226 6890 16408
rect 6974 16368 7008 16408
rect 7210 16368 7244 16408
rect 6974 16339 7244 16368
rect 7328 16367 7362 16408
rect 7564 16367 7598 16408
rect 7328 16339 7598 16367
rect 7564 16291 7598 16339
rect 6175 16133 6402 16169
rect 6175 16099 6241 16133
rect 6175 16065 6191 16099
rect 6225 16065 6241 16099
rect 6175 16059 6241 16065
rect 6367 16026 6402 16133
rect 6781 16172 6890 16226
rect 7535 16261 7598 16291
rect 5731 16019 5764 16023
rect 5967 16019 6000 16023
rect 5312 15838 5318 16014
rect 5352 15838 5358 16014
rect 5312 15826 5358 15838
rect 5607 16007 5653 16019
rect 5607 15831 5613 16007
rect 5647 15831 5653 16007
rect 4446 15788 4479 15820
rect 4682 15788 4715 15820
rect 4446 15752 4715 15788
rect 5082 15787 5116 15826
rect 5318 15787 5352 15826
rect 5607 15819 5653 15831
rect 5725 16007 5771 16019
rect 5725 15831 5731 16007
rect 5765 15831 5771 16007
rect 5725 15819 5771 15831
rect 5843 16007 5889 16019
rect 5843 15831 5849 16007
rect 5883 15831 5889 16007
rect 5843 15819 5889 15831
rect 5961 16007 6007 16019
rect 5961 15831 5967 16007
rect 6001 15959 6007 16007
rect 6126 16014 6172 16026
rect 6126 15959 6132 16014
rect 6001 15871 6132 15959
rect 6001 15831 6007 15871
rect 5961 15819 6007 15831
rect 6126 15838 6132 15871
rect 6166 15838 6172 16014
rect 6126 15826 6172 15838
rect 6244 16014 6290 16026
rect 6244 15838 6250 16014
rect 6284 15838 6290 16014
rect 6244 15826 6290 15838
rect 6362 16014 6408 16026
rect 6362 15838 6368 16014
rect 6402 15838 6408 16014
rect 6362 15826 6408 15838
rect 6480 16014 6526 16026
rect 6781 16019 6815 16172
rect 7535 16169 7570 16261
rect 8024 16226 8058 16410
rect 8142 16368 8176 16410
rect 8378 16368 8412 16410
rect 8142 16339 8412 16368
rect 8496 16367 8530 16410
rect 8732 16367 8766 16410
rect 9192 16408 9238 16420
rect 9310 16796 9356 16808
rect 9310 16420 9316 16796
rect 9350 16420 9356 16796
rect 9310 16408 9356 16420
rect 9428 16796 9474 16808
rect 9428 16420 9434 16796
rect 9468 16420 9474 16796
rect 9428 16408 9474 16420
rect 9546 16796 9592 16808
rect 9546 16420 9552 16796
rect 9586 16420 9592 16796
rect 9546 16408 9592 16420
rect 9664 16796 9710 16808
rect 9664 16420 9670 16796
rect 9704 16420 9710 16796
rect 9664 16408 9710 16420
rect 9782 16796 9828 16808
rect 9782 16420 9788 16796
rect 9822 16420 9828 16796
rect 9782 16408 9828 16420
rect 9900 16796 9946 16808
rect 9900 16420 9906 16796
rect 9940 16420 9946 16796
rect 9980 16728 10080 16816
rect 10366 16806 10400 16869
rect 10602 16806 10636 16869
rect 10720 16869 10990 16897
rect 11325 16880 11389 17533
rect 16520 17505 23959 17506
rect 12316 17501 23959 17505
rect 12316 17447 23905 17501
rect 23959 17447 23969 17501
rect 12316 17442 23959 17447
rect 12316 17441 14944 17442
rect 12316 17070 12380 17441
rect 25576 17412 26102 17413
rect 16520 17411 26111 17412
rect 12472 17408 26111 17411
rect 12472 17354 23795 17408
rect 23849 17354 26111 17408
rect 12472 17348 26111 17354
rect 12472 17347 14944 17348
rect 11626 17044 11730 17050
rect 11626 16972 11638 17044
rect 11718 16972 11730 17044
rect 11626 16966 11730 16972
rect 12316 16968 12416 17070
rect 11660 16910 11695 16966
rect 12316 16934 12332 16968
rect 12366 16934 12416 16968
rect 10720 16806 10754 16869
rect 10956 16806 10990 16869
rect 11148 16860 11389 16880
rect 11148 16826 11164 16860
rect 11198 16826 11389 16860
rect 11148 16816 11389 16826
rect 11534 16869 11804 16910
rect 12316 16908 12416 16934
rect 10360 16794 10406 16806
rect 9900 16408 9946 16420
rect 10360 16418 10366 16794
rect 10400 16418 10406 16794
rect 8496 16339 8766 16367
rect 8732 16291 8766 16339
rect 7343 16133 7570 16169
rect 7343 16099 7409 16133
rect 7343 16065 7359 16099
rect 7393 16065 7409 16099
rect 7343 16059 7409 16065
rect 7535 16024 7570 16133
rect 7949 16172 8058 16226
rect 8703 16261 8766 16291
rect 6899 16019 6932 16024
rect 7135 16019 7168 16023
rect 6480 15838 6486 16014
rect 6520 15838 6526 16014
rect 6480 15826 6526 15838
rect 6775 16007 6821 16019
rect 6775 15831 6781 16007
rect 6815 15831 6821 16007
rect 5082 15748 5352 15787
rect 5614 15788 5647 15819
rect 5850 15788 5883 15819
rect 5614 15752 5883 15788
rect 6250 15787 6284 15826
rect 6486 15787 6520 15826
rect 6775 15819 6821 15831
rect 6893 16007 6939 16019
rect 6893 15831 6899 16007
rect 6933 15831 6939 16007
rect 6893 15819 6939 15831
rect 7011 16007 7057 16019
rect 7011 15831 7017 16007
rect 7051 15831 7057 16007
rect 7011 15819 7057 15831
rect 7129 16007 7175 16019
rect 7129 15831 7135 16007
rect 7169 15959 7175 16007
rect 7294 16012 7340 16024
rect 7294 15959 7300 16012
rect 7169 15871 7300 15959
rect 7169 15831 7175 15871
rect 7129 15819 7175 15831
rect 7294 15836 7300 15871
rect 7334 15836 7340 16012
rect 7294 15824 7340 15836
rect 7412 16012 7458 16024
rect 7412 15836 7418 16012
rect 7452 15836 7458 16012
rect 7412 15824 7458 15836
rect 7530 16012 7576 16024
rect 7530 15836 7536 16012
rect 7570 15836 7576 16012
rect 7530 15824 7576 15836
rect 7648 16012 7694 16024
rect 7949 16020 7983 16172
rect 8703 16169 8738 16261
rect 9198 16224 9232 16408
rect 9316 16366 9350 16408
rect 9552 16366 9586 16408
rect 9316 16337 9586 16366
rect 9670 16365 9704 16408
rect 9906 16365 9940 16408
rect 10360 16406 10406 16418
rect 10478 16794 10524 16806
rect 10478 16418 10484 16794
rect 10518 16418 10524 16794
rect 10478 16406 10524 16418
rect 10596 16794 10642 16806
rect 10596 16418 10602 16794
rect 10636 16418 10642 16794
rect 10596 16406 10642 16418
rect 10714 16794 10760 16806
rect 10714 16418 10720 16794
rect 10754 16418 10760 16794
rect 10714 16406 10760 16418
rect 10832 16794 10878 16806
rect 10832 16418 10838 16794
rect 10872 16418 10878 16794
rect 10832 16406 10878 16418
rect 10950 16794 10996 16806
rect 10950 16418 10956 16794
rect 10990 16418 10996 16794
rect 10950 16406 10996 16418
rect 11068 16794 11114 16806
rect 11068 16418 11074 16794
rect 11108 16418 11114 16794
rect 11148 16728 11248 16816
rect 11534 16808 11568 16869
rect 11770 16808 11804 16869
rect 11888 16869 12158 16897
rect 12472 16880 12536 17347
rect 13484 17255 25569 17319
rect 13484 17070 13548 17255
rect 13629 17161 25330 17225
rect 12794 17044 12898 17050
rect 12794 16972 12806 17044
rect 12886 16972 12898 17044
rect 12794 16966 12898 16972
rect 13484 16968 13584 17070
rect 12828 16910 12863 16966
rect 13484 16934 13500 16968
rect 13534 16934 13584 16968
rect 11888 16808 11922 16869
rect 12124 16808 12158 16869
rect 12316 16860 12536 16880
rect 12316 16826 12332 16860
rect 12366 16826 12536 16860
rect 12316 16816 12536 16826
rect 12702 16869 12972 16910
rect 13484 16908 13584 16934
rect 11528 16796 11574 16808
rect 11068 16406 11114 16418
rect 11528 16420 11534 16796
rect 11568 16420 11574 16796
rect 11528 16408 11574 16420
rect 11646 16796 11692 16808
rect 11646 16420 11652 16796
rect 11686 16420 11692 16796
rect 11646 16408 11692 16420
rect 11764 16796 11810 16808
rect 11764 16420 11770 16796
rect 11804 16420 11810 16796
rect 11764 16408 11810 16420
rect 11882 16796 11928 16808
rect 11882 16420 11888 16796
rect 11922 16420 11928 16796
rect 11882 16408 11928 16420
rect 12000 16796 12046 16808
rect 12000 16420 12006 16796
rect 12040 16420 12046 16796
rect 12000 16408 12046 16420
rect 12118 16796 12164 16808
rect 12118 16420 12124 16796
rect 12158 16420 12164 16796
rect 12118 16408 12164 16420
rect 12236 16796 12282 16808
rect 12236 16420 12242 16796
rect 12276 16420 12282 16796
rect 12316 16728 12416 16816
rect 12702 16808 12736 16869
rect 12938 16808 12972 16869
rect 13056 16869 13326 16897
rect 13056 16808 13090 16869
rect 13292 16808 13326 16869
rect 13484 16860 13584 16880
rect 13484 16826 13500 16860
rect 13534 16826 13584 16860
rect 12696 16796 12742 16808
rect 12236 16408 12282 16420
rect 12696 16420 12702 16796
rect 12736 16420 12742 16796
rect 12696 16408 12742 16420
rect 12814 16796 12860 16808
rect 12814 16420 12820 16796
rect 12854 16420 12860 16796
rect 12814 16408 12860 16420
rect 12932 16796 12978 16808
rect 12932 16420 12938 16796
rect 12972 16420 12978 16796
rect 12932 16408 12978 16420
rect 13050 16796 13096 16808
rect 13050 16420 13056 16796
rect 13090 16420 13096 16796
rect 13050 16408 13096 16420
rect 13168 16796 13214 16808
rect 13168 16420 13174 16796
rect 13208 16420 13214 16796
rect 13168 16408 13214 16420
rect 13286 16796 13332 16808
rect 13286 16420 13292 16796
rect 13326 16420 13332 16796
rect 13286 16408 13332 16420
rect 13404 16796 13450 16808
rect 13404 16420 13410 16796
rect 13444 16420 13450 16796
rect 13484 16797 13584 16826
rect 13629 16797 13684 17161
rect 25267 16962 25330 17161
rect 13484 16728 13684 16797
rect 14458 16839 14594 16859
rect 14458 16777 14498 16839
rect 14558 16777 14594 16839
rect 14458 16749 14594 16777
rect 15906 16839 16042 16859
rect 15906 16777 15946 16839
rect 16006 16777 16042 16839
rect 15906 16749 16042 16777
rect 17404 16837 17540 16857
rect 17404 16775 17444 16837
rect 17504 16775 17540 16837
rect 13921 16719 14898 16749
rect 13921 16613 13955 16719
rect 14158 16613 14190 16719
rect 14394 16613 14426 16719
rect 14630 16613 14662 16719
rect 14866 16613 14898 16719
rect 15369 16719 16346 16749
rect 17404 16747 17540 16775
rect 18852 16837 18988 16857
rect 18852 16775 18892 16837
rect 18952 16775 18988 16837
rect 18852 16747 18988 16775
rect 20372 16839 20508 16859
rect 20372 16777 20412 16839
rect 20472 16777 20508 16839
rect 20372 16749 20508 16777
rect 21820 16839 21956 16859
rect 21820 16777 21860 16839
rect 21920 16777 21956 16839
rect 21820 16749 21956 16777
rect 23318 16837 23454 16857
rect 23318 16775 23358 16837
rect 23418 16775 23454 16837
rect 15369 16613 15403 16719
rect 15606 16613 15638 16719
rect 15842 16613 15874 16719
rect 16078 16613 16110 16719
rect 16314 16613 16346 16719
rect 16867 16717 17844 16747
rect 13404 16408 13450 16420
rect 13797 16601 13843 16613
rect 13797 16425 13803 16601
rect 13837 16425 13843 16601
rect 13797 16413 13843 16425
rect 13915 16601 13961 16613
rect 13915 16425 13921 16601
rect 13955 16425 13961 16601
rect 13915 16413 13961 16425
rect 14033 16601 14079 16613
rect 14033 16425 14039 16601
rect 14073 16425 14079 16601
rect 14033 16413 14079 16425
rect 14151 16601 14197 16613
rect 14151 16425 14157 16601
rect 14191 16425 14197 16601
rect 14151 16413 14197 16425
rect 14269 16601 14315 16613
rect 14269 16425 14275 16601
rect 14309 16425 14315 16601
rect 14269 16413 14315 16425
rect 14387 16601 14433 16613
rect 14387 16425 14393 16601
rect 14427 16425 14433 16601
rect 14387 16413 14433 16425
rect 14505 16601 14551 16613
rect 14505 16425 14511 16601
rect 14545 16425 14551 16601
rect 14505 16413 14551 16425
rect 14623 16601 14669 16613
rect 14623 16425 14629 16601
rect 14663 16425 14669 16601
rect 14623 16413 14669 16425
rect 14741 16601 14787 16613
rect 14741 16425 14747 16601
rect 14781 16425 14787 16601
rect 14741 16413 14787 16425
rect 14859 16601 14905 16613
rect 14859 16425 14865 16601
rect 14899 16425 14905 16601
rect 14859 16413 14905 16425
rect 15245 16601 15291 16613
rect 15245 16425 15251 16601
rect 15285 16425 15291 16601
rect 15245 16413 15291 16425
rect 15363 16601 15409 16613
rect 15363 16425 15369 16601
rect 15403 16425 15409 16601
rect 15363 16413 15409 16425
rect 15481 16601 15527 16613
rect 15481 16425 15487 16601
rect 15521 16425 15527 16601
rect 15481 16413 15527 16425
rect 15599 16601 15645 16613
rect 15599 16425 15605 16601
rect 15639 16425 15645 16601
rect 15599 16413 15645 16425
rect 15717 16601 15763 16613
rect 15717 16425 15723 16601
rect 15757 16425 15763 16601
rect 15717 16413 15763 16425
rect 15835 16601 15881 16613
rect 15835 16425 15841 16601
rect 15875 16425 15881 16601
rect 15835 16413 15881 16425
rect 15953 16601 15999 16613
rect 15953 16425 15959 16601
rect 15993 16425 15999 16601
rect 15953 16413 15999 16425
rect 16071 16601 16117 16613
rect 16071 16425 16077 16601
rect 16111 16425 16117 16601
rect 16071 16413 16117 16425
rect 16189 16601 16235 16613
rect 16189 16425 16195 16601
rect 16229 16425 16235 16601
rect 16189 16413 16235 16425
rect 16307 16601 16353 16613
rect 16867 16611 16901 16717
rect 17104 16611 17136 16717
rect 17340 16611 17372 16717
rect 17576 16611 17608 16717
rect 17812 16611 17844 16717
rect 18315 16717 19292 16747
rect 18315 16611 18349 16717
rect 18552 16611 18584 16717
rect 18788 16611 18820 16717
rect 19024 16611 19056 16717
rect 19260 16611 19292 16717
rect 19835 16719 20812 16749
rect 19835 16613 19869 16719
rect 20072 16613 20104 16719
rect 20308 16613 20340 16719
rect 20544 16613 20576 16719
rect 20780 16613 20812 16719
rect 21283 16719 22260 16749
rect 23318 16747 23454 16775
rect 24766 16837 24902 16857
rect 24766 16775 24806 16837
rect 24866 16775 24902 16837
rect 24766 16747 24902 16775
rect 21283 16613 21317 16719
rect 21520 16613 21552 16719
rect 21756 16613 21788 16719
rect 21992 16613 22024 16719
rect 22228 16613 22260 16719
rect 22781 16717 23758 16747
rect 16307 16425 16313 16601
rect 16347 16425 16353 16601
rect 16307 16413 16353 16425
rect 16743 16599 16789 16611
rect 16743 16423 16749 16599
rect 16783 16423 16789 16599
rect 9670 16337 9940 16365
rect 9906 16289 9940 16337
rect 8511 16133 8738 16169
rect 8511 16099 8577 16133
rect 8511 16065 8527 16099
rect 8561 16065 8577 16099
rect 8511 16059 8577 16065
rect 8703 16024 8738 16133
rect 9123 16170 9232 16224
rect 9877 16259 9940 16289
rect 9123 16024 9157 16170
rect 9877 16167 9912 16259
rect 10366 16224 10400 16406
rect 10484 16366 10518 16406
rect 10720 16366 10754 16406
rect 10484 16337 10754 16366
rect 10838 16365 10872 16406
rect 11074 16365 11108 16406
rect 10838 16337 11108 16365
rect 11074 16289 11108 16337
rect 9685 16131 9912 16167
rect 9685 16097 9751 16131
rect 9685 16063 9701 16097
rect 9735 16063 9751 16097
rect 9685 16057 9751 16063
rect 9241 16024 9274 16028
rect 9477 16024 9510 16028
rect 9877 16024 9912 16131
rect 10291 16170 10400 16224
rect 11045 16259 11108 16289
rect 10291 16024 10325 16170
rect 11045 16167 11080 16259
rect 11534 16224 11568 16408
rect 11652 16366 11686 16408
rect 11888 16366 11922 16408
rect 11652 16337 11922 16366
rect 12006 16365 12040 16408
rect 12242 16365 12276 16408
rect 12006 16337 12276 16365
rect 12242 16289 12276 16337
rect 10853 16131 11080 16167
rect 10853 16097 10919 16131
rect 10853 16063 10869 16097
rect 10903 16063 10919 16097
rect 10853 16057 10919 16063
rect 10409 16024 10442 16028
rect 10645 16024 10678 16028
rect 11045 16024 11080 16131
rect 11459 16170 11568 16224
rect 12213 16259 12276 16289
rect 11459 16024 11493 16170
rect 12213 16167 12248 16259
rect 12702 16224 12736 16408
rect 12820 16366 12854 16408
rect 13056 16366 13090 16408
rect 12820 16337 13090 16366
rect 13174 16365 13208 16408
rect 13410 16365 13444 16408
rect 13174 16337 13444 16365
rect 13410 16289 13444 16337
rect 12021 16131 12248 16167
rect 12021 16097 12087 16131
rect 12021 16063 12037 16097
rect 12071 16063 12087 16097
rect 12021 16057 12087 16063
rect 11577 16024 11610 16028
rect 11813 16024 11846 16028
rect 12213 16024 12248 16131
rect 12627 16170 12736 16224
rect 13381 16259 13444 16289
rect 8067 16020 8100 16024
rect 8303 16020 8336 16024
rect 7648 15836 7654 16012
rect 7688 15836 7694 16012
rect 7648 15824 7694 15836
rect 7944 16008 7990 16020
rect 7944 15832 7950 16008
rect 7984 15832 7990 16008
rect 6250 15748 6520 15787
rect 6782 15788 6815 15819
rect 7018 15788 7051 15819
rect 6782 15752 7051 15788
rect 7418 15787 7452 15824
rect 7654 15787 7688 15824
rect 7944 15820 7990 15832
rect 8062 16008 8108 16020
rect 8062 15832 8068 16008
rect 8102 15832 8108 16008
rect 8062 15820 8108 15832
rect 8180 16008 8226 16020
rect 8180 15832 8186 16008
rect 8220 15832 8226 16008
rect 8180 15820 8226 15832
rect 8298 16008 8344 16020
rect 8298 15832 8304 16008
rect 8338 15959 8344 16008
rect 8462 16012 8508 16024
rect 8462 15959 8468 16012
rect 8338 15871 8468 15959
rect 8338 15832 8344 15871
rect 8298 15820 8344 15832
rect 8462 15836 8468 15871
rect 8502 15836 8508 16012
rect 8462 15824 8508 15836
rect 8580 16012 8626 16024
rect 8580 15836 8586 16012
rect 8620 15836 8626 16012
rect 8580 15824 8626 15836
rect 8698 16012 8744 16024
rect 8698 15836 8704 16012
rect 8738 15836 8744 16012
rect 8698 15824 8744 15836
rect 8816 16012 8862 16024
rect 8816 15836 8822 16012
rect 8856 15836 8862 16012
rect 8816 15824 8862 15836
rect 9116 16012 9162 16024
rect 9116 15836 9122 16012
rect 9156 15836 9162 16012
rect 9116 15824 9162 15836
rect 9234 16012 9280 16024
rect 9234 15836 9240 16012
rect 9274 15836 9280 16012
rect 9234 15824 9280 15836
rect 9352 16012 9398 16024
rect 9352 15836 9358 16012
rect 9392 15836 9398 16012
rect 9352 15824 9398 15836
rect 9470 16012 9516 16024
rect 9470 15836 9476 16012
rect 9510 15957 9516 16012
rect 9636 16012 9682 16024
rect 9636 15957 9642 16012
rect 9510 15869 9642 15957
rect 9510 15836 9516 15869
rect 9470 15824 9516 15836
rect 9636 15836 9642 15869
rect 9676 15836 9682 16012
rect 9636 15824 9682 15836
rect 9754 16012 9800 16024
rect 9754 15836 9760 16012
rect 9794 15836 9800 16012
rect 9754 15824 9800 15836
rect 9872 16012 9918 16024
rect 9872 15836 9878 16012
rect 9912 15836 9918 16012
rect 9872 15824 9918 15836
rect 9990 16012 10036 16024
rect 9990 15836 9996 16012
rect 10030 15836 10036 16012
rect 9990 15824 10036 15836
rect 10285 16012 10331 16024
rect 10285 15836 10291 16012
rect 10325 15836 10331 16012
rect 10285 15824 10331 15836
rect 10403 16012 10449 16024
rect 10403 15836 10409 16012
rect 10443 15836 10449 16012
rect 10403 15824 10449 15836
rect 10521 16012 10567 16024
rect 10521 15836 10527 16012
rect 10561 15836 10567 16012
rect 10521 15824 10567 15836
rect 10639 16012 10685 16024
rect 10639 15836 10645 16012
rect 10679 15957 10685 16012
rect 10804 16012 10850 16024
rect 10804 15957 10810 16012
rect 10679 15869 10810 15957
rect 10679 15836 10685 15869
rect 10639 15824 10685 15836
rect 10804 15836 10810 15869
rect 10844 15836 10850 16012
rect 10804 15824 10850 15836
rect 10922 16012 10968 16024
rect 10922 15836 10928 16012
rect 10962 15836 10968 16012
rect 10922 15824 10968 15836
rect 11040 16012 11086 16024
rect 11040 15836 11046 16012
rect 11080 15836 11086 16012
rect 11040 15824 11086 15836
rect 11158 16012 11204 16024
rect 11158 15836 11164 16012
rect 11198 15836 11204 16012
rect 11158 15824 11204 15836
rect 11453 16012 11499 16024
rect 11453 15836 11459 16012
rect 11493 15836 11499 16012
rect 11453 15824 11499 15836
rect 11571 16012 11617 16024
rect 11571 15836 11577 16012
rect 11611 15836 11617 16012
rect 11571 15824 11617 15836
rect 11689 16012 11735 16024
rect 11689 15836 11695 16012
rect 11729 15836 11735 16012
rect 11689 15824 11735 15836
rect 11807 16012 11853 16024
rect 11807 15836 11813 16012
rect 11847 15957 11853 16012
rect 11972 16012 12018 16024
rect 11972 15957 11978 16012
rect 11847 15869 11978 15957
rect 11847 15836 11853 15869
rect 11807 15824 11853 15836
rect 11972 15836 11978 15869
rect 12012 15836 12018 16012
rect 11972 15824 12018 15836
rect 12090 16012 12136 16024
rect 12090 15836 12096 16012
rect 12130 15836 12136 16012
rect 12090 15824 12136 15836
rect 12208 16012 12254 16024
rect 12208 15836 12214 16012
rect 12248 15836 12254 16012
rect 12208 15824 12254 15836
rect 12326 16012 12372 16024
rect 12627 16018 12661 16170
rect 13381 16167 13416 16259
rect 13189 16131 13416 16167
rect 13189 16097 13255 16131
rect 13189 16063 13205 16097
rect 13239 16063 13255 16097
rect 13189 16057 13255 16063
rect 12745 16018 12778 16049
rect 13381 16022 13416 16131
rect 13803 16180 13838 16413
rect 14082 16365 14148 16372
rect 14082 16331 14098 16365
rect 14132 16331 14148 16365
rect 14082 16320 14148 16331
rect 14274 16320 14310 16413
rect 14082 16319 14310 16320
rect 14510 16319 14546 16413
rect 14746 16319 14782 16413
rect 14082 16290 14782 16319
rect 14200 16289 14782 16290
rect 14200 16248 14266 16289
rect 14200 16214 14216 16248
rect 14250 16214 14266 16248
rect 14200 16207 14266 16214
rect 13803 16176 14192 16180
rect 14628 16176 14662 16289
rect 15251 16180 15286 16413
rect 15530 16365 15596 16372
rect 15530 16331 15546 16365
rect 15580 16331 15596 16365
rect 15530 16320 15596 16331
rect 15722 16320 15758 16413
rect 15530 16319 15758 16320
rect 15958 16319 15994 16413
rect 16194 16319 16230 16413
rect 16743 16411 16789 16423
rect 16861 16599 16907 16611
rect 16861 16423 16867 16599
rect 16901 16423 16907 16599
rect 16861 16411 16907 16423
rect 16979 16599 17025 16611
rect 16979 16423 16985 16599
rect 17019 16423 17025 16599
rect 16979 16411 17025 16423
rect 17097 16599 17143 16611
rect 17097 16423 17103 16599
rect 17137 16423 17143 16599
rect 17097 16411 17143 16423
rect 17215 16599 17261 16611
rect 17215 16423 17221 16599
rect 17255 16423 17261 16599
rect 17215 16411 17261 16423
rect 17333 16599 17379 16611
rect 17333 16423 17339 16599
rect 17373 16423 17379 16599
rect 17333 16411 17379 16423
rect 17451 16599 17497 16611
rect 17451 16423 17457 16599
rect 17491 16423 17497 16599
rect 17451 16411 17497 16423
rect 17569 16599 17615 16611
rect 17569 16423 17575 16599
rect 17609 16423 17615 16599
rect 17569 16411 17615 16423
rect 17687 16599 17733 16611
rect 17687 16423 17693 16599
rect 17727 16423 17733 16599
rect 17687 16411 17733 16423
rect 17805 16599 17851 16611
rect 17805 16423 17811 16599
rect 17845 16423 17851 16599
rect 17805 16411 17851 16423
rect 18191 16599 18237 16611
rect 18191 16423 18197 16599
rect 18231 16423 18237 16599
rect 18191 16411 18237 16423
rect 18309 16599 18355 16611
rect 18309 16423 18315 16599
rect 18349 16423 18355 16599
rect 18309 16411 18355 16423
rect 18427 16599 18473 16611
rect 18427 16423 18433 16599
rect 18467 16423 18473 16599
rect 18427 16411 18473 16423
rect 18545 16599 18591 16611
rect 18545 16423 18551 16599
rect 18585 16423 18591 16599
rect 18545 16411 18591 16423
rect 18663 16599 18709 16611
rect 18663 16423 18669 16599
rect 18703 16423 18709 16599
rect 18663 16411 18709 16423
rect 18781 16599 18827 16611
rect 18781 16423 18787 16599
rect 18821 16423 18827 16599
rect 18781 16411 18827 16423
rect 18899 16599 18945 16611
rect 18899 16423 18905 16599
rect 18939 16423 18945 16599
rect 18899 16411 18945 16423
rect 19017 16599 19063 16611
rect 19017 16423 19023 16599
rect 19057 16423 19063 16599
rect 19017 16411 19063 16423
rect 19135 16599 19181 16611
rect 19135 16423 19141 16599
rect 19175 16423 19181 16599
rect 19135 16411 19181 16423
rect 19253 16599 19299 16611
rect 19253 16423 19259 16599
rect 19293 16423 19299 16599
rect 19253 16411 19299 16423
rect 19711 16601 19757 16613
rect 19711 16425 19717 16601
rect 19751 16425 19757 16601
rect 19711 16413 19757 16425
rect 19829 16601 19875 16613
rect 19829 16425 19835 16601
rect 19869 16425 19875 16601
rect 19829 16413 19875 16425
rect 19947 16601 19993 16613
rect 19947 16425 19953 16601
rect 19987 16425 19993 16601
rect 19947 16413 19993 16425
rect 20065 16601 20111 16613
rect 20065 16425 20071 16601
rect 20105 16425 20111 16601
rect 20065 16413 20111 16425
rect 20183 16601 20229 16613
rect 20183 16425 20189 16601
rect 20223 16425 20229 16601
rect 20183 16413 20229 16425
rect 20301 16601 20347 16613
rect 20301 16425 20307 16601
rect 20341 16425 20347 16601
rect 20301 16413 20347 16425
rect 20419 16601 20465 16613
rect 20419 16425 20425 16601
rect 20459 16425 20465 16601
rect 20419 16413 20465 16425
rect 20537 16601 20583 16613
rect 20537 16425 20543 16601
rect 20577 16425 20583 16601
rect 20537 16413 20583 16425
rect 20655 16601 20701 16613
rect 20655 16425 20661 16601
rect 20695 16425 20701 16601
rect 20655 16413 20701 16425
rect 20773 16601 20819 16613
rect 20773 16425 20779 16601
rect 20813 16425 20819 16601
rect 20773 16413 20819 16425
rect 21159 16601 21205 16613
rect 21159 16425 21165 16601
rect 21199 16425 21205 16601
rect 21159 16413 21205 16425
rect 21277 16601 21323 16613
rect 21277 16425 21283 16601
rect 21317 16425 21323 16601
rect 21277 16413 21323 16425
rect 21395 16601 21441 16613
rect 21395 16425 21401 16601
rect 21435 16425 21441 16601
rect 21395 16413 21441 16425
rect 21513 16601 21559 16613
rect 21513 16425 21519 16601
rect 21553 16425 21559 16601
rect 21513 16413 21559 16425
rect 21631 16601 21677 16613
rect 21631 16425 21637 16601
rect 21671 16425 21677 16601
rect 21631 16413 21677 16425
rect 21749 16601 21795 16613
rect 21749 16425 21755 16601
rect 21789 16425 21795 16601
rect 21749 16413 21795 16425
rect 21867 16601 21913 16613
rect 21867 16425 21873 16601
rect 21907 16425 21913 16601
rect 21867 16413 21913 16425
rect 21985 16601 22031 16613
rect 21985 16425 21991 16601
rect 22025 16425 22031 16601
rect 21985 16413 22031 16425
rect 22103 16601 22149 16613
rect 22103 16425 22109 16601
rect 22143 16425 22149 16601
rect 22103 16413 22149 16425
rect 22221 16601 22267 16613
rect 22781 16611 22815 16717
rect 23018 16611 23050 16717
rect 23254 16611 23286 16717
rect 23490 16611 23522 16717
rect 23726 16611 23758 16717
rect 24229 16717 25206 16747
rect 24229 16611 24263 16717
rect 24466 16611 24498 16717
rect 24702 16611 24734 16717
rect 24938 16611 24970 16717
rect 25174 16611 25206 16717
rect 22221 16425 22227 16601
rect 22261 16425 22267 16601
rect 22221 16413 22267 16425
rect 22657 16599 22703 16611
rect 22657 16423 22663 16599
rect 22697 16423 22703 16599
rect 15530 16290 16230 16319
rect 15648 16289 16230 16290
rect 15648 16248 15714 16289
rect 15648 16214 15664 16248
rect 15698 16214 15714 16248
rect 15648 16207 15714 16214
rect 15251 16176 15640 16180
rect 16076 16176 16110 16289
rect 16749 16178 16784 16411
rect 17028 16363 17094 16370
rect 17028 16329 17044 16363
rect 17078 16329 17094 16363
rect 17028 16318 17094 16329
rect 17220 16318 17256 16411
rect 17028 16317 17256 16318
rect 17456 16317 17492 16411
rect 17692 16317 17728 16411
rect 17028 16288 17728 16317
rect 17146 16287 17728 16288
rect 17146 16246 17212 16287
rect 17146 16212 17162 16246
rect 17196 16212 17212 16246
rect 17146 16205 17212 16212
rect 13803 16164 14197 16176
rect 13803 16151 14157 16164
rect 12326 15836 12332 16012
rect 12366 15836 12372 16012
rect 12326 15824 12372 15836
rect 12620 16006 12666 16018
rect 12620 15830 12626 16006
rect 12660 15830 12666 16006
rect 7418 15748 7688 15787
rect 7950 15788 7983 15820
rect 8186 15788 8219 15820
rect 7950 15752 8219 15788
rect 8586 15787 8620 15824
rect 8822 15787 8856 15824
rect 8586 15748 8856 15787
rect 9124 15786 9157 15824
rect 9360 15786 9393 15824
rect 9124 15750 9393 15786
rect 9760 15785 9794 15824
rect 9996 15785 10030 15824
rect 5118 15720 5152 15748
rect 6286 15720 6320 15748
rect 7454 15720 7488 15748
rect 8622 15720 8656 15748
rect 9760 15746 10030 15785
rect 10292 15786 10325 15824
rect 10528 15786 10561 15824
rect 10292 15750 10561 15786
rect 10928 15785 10962 15824
rect 11164 15785 11198 15824
rect 10928 15746 11198 15785
rect 11460 15786 11493 15824
rect 11696 15786 11729 15824
rect 11460 15750 11729 15786
rect 12096 15785 12130 15824
rect 12332 15785 12366 15824
rect 12620 15818 12666 15830
rect 12738 16006 12784 16018
rect 12738 15830 12744 16006
rect 12778 15830 12784 16006
rect 12738 15818 12784 15830
rect 12856 16006 12902 16018
rect 12856 15830 12862 16006
rect 12896 15830 12902 16006
rect 12856 15818 12902 15830
rect 12974 16006 13020 16018
rect 12974 15830 12980 16006
rect 13014 15957 13020 16006
rect 13140 16010 13186 16022
rect 13140 15957 13146 16010
rect 13014 15869 13146 15957
rect 13014 15830 13020 15869
rect 12974 15818 13020 15830
rect 13140 15834 13146 15869
rect 13180 15834 13186 16010
rect 13140 15822 13186 15834
rect 13258 16010 13304 16022
rect 13258 15834 13264 16010
rect 13298 15834 13304 16010
rect 13258 15822 13304 15834
rect 13376 16010 13422 16022
rect 13376 15834 13382 16010
rect 13416 15834 13422 16010
rect 13376 15822 13422 15834
rect 13494 16010 13540 16022
rect 13494 15834 13500 16010
rect 13534 15834 13540 16010
rect 13494 15822 13540 15834
rect 12096 15746 12366 15785
rect 12628 15786 12661 15818
rect 12864 15786 12897 15818
rect 12628 15750 12897 15786
rect 13264 15785 13298 15822
rect 13500 15785 13534 15822
rect 13264 15746 13534 15785
rect 5096 15708 5174 15720
rect 5096 15638 5102 15708
rect 5168 15638 5174 15708
rect 5096 15626 5174 15638
rect 6264 15708 6342 15720
rect 6264 15638 6270 15708
rect 6336 15638 6342 15708
rect 6264 15626 6342 15638
rect 7432 15708 7510 15720
rect 7432 15638 7438 15708
rect 7504 15638 7510 15708
rect 7432 15626 7510 15638
rect 8600 15708 8678 15720
rect 9796 15718 9830 15746
rect 10964 15718 10998 15746
rect 12132 15718 12166 15746
rect 13300 15718 13334 15746
rect 8600 15638 8606 15708
rect 8672 15638 8678 15708
rect 8600 15626 8678 15638
rect 9774 15706 9852 15718
rect 9774 15636 9780 15706
rect 9846 15636 9852 15706
rect 9774 15624 9852 15636
rect 10942 15706 11020 15718
rect 10942 15636 10948 15706
rect 11014 15636 11020 15706
rect 10942 15624 11020 15636
rect 12110 15706 12188 15718
rect 12110 15636 12116 15706
rect 12182 15636 12188 15706
rect 12110 15624 12188 15636
rect 13278 15706 13356 15718
rect 13278 15636 13284 15706
rect 13350 15636 13356 15706
rect 13278 15624 13356 15636
rect 13803 15562 13907 16151
rect 14151 15988 14157 16151
rect 14191 15988 14197 16164
rect 14151 15976 14197 15988
rect 14269 16164 14315 16176
rect 14269 15988 14275 16164
rect 14309 15988 14315 16164
rect 14269 15981 14315 15988
rect 14266 15976 14315 15981
rect 14386 16164 14432 16176
rect 14266 15815 14309 15976
rect 14386 15815 14392 16164
rect 14266 15788 14392 15815
rect 14426 15788 14432 16164
rect 14266 15776 14432 15788
rect 14504 16164 14550 16176
rect 14504 15788 14510 16164
rect 14544 15788 14550 16164
rect 14504 15776 14550 15788
rect 14622 16164 14668 16176
rect 14622 15788 14628 16164
rect 14662 15788 14668 16164
rect 15251 16164 15645 16176
rect 15251 16151 15605 16164
rect 14708 16030 14808 16036
rect 14706 15942 14716 16030
rect 14802 15942 14812 16030
rect 14708 15936 14808 15942
rect 14622 15776 14668 15788
rect 14266 15772 14426 15776
rect 14266 15635 14342 15772
rect 14730 15744 14784 15936
rect 14820 15901 14920 15908
rect 14820 15813 14830 15901
rect 14916 15813 14926 15901
rect 14820 15808 14920 15813
rect 14435 15738 14501 15744
rect 14435 15704 14451 15738
rect 14485 15704 14501 15738
rect 14435 15659 14501 15704
rect 14553 15738 14784 15744
rect 14553 15704 14569 15738
rect 14603 15704 14784 15738
rect 14553 15688 14784 15704
rect 14844 15659 14898 15808
rect 14435 15651 14898 15659
rect 14264 15575 14274 15635
rect 14336 15575 14346 15635
rect 14434 15619 14898 15651
rect 12407 15514 13907 15562
rect 12407 15509 12445 15514
rect 9287 15437 12445 15509
rect 15251 15486 15355 16151
rect 15599 15988 15605 16151
rect 15639 15988 15645 16164
rect 15599 15976 15645 15988
rect 15717 16164 15763 16176
rect 15717 15988 15723 16164
rect 15757 15988 15763 16164
rect 15717 15981 15763 15988
rect 15714 15976 15763 15981
rect 15834 16164 15880 16176
rect 15714 15815 15757 15976
rect 15834 15815 15840 16164
rect 15714 15788 15840 15815
rect 15874 15788 15880 16164
rect 15714 15776 15880 15788
rect 15952 16164 15998 16176
rect 15952 15788 15958 16164
rect 15992 15788 15998 16164
rect 15952 15776 15998 15788
rect 16070 16164 16116 16176
rect 16070 15788 16076 16164
rect 16110 15788 16116 16164
rect 16749 16174 17138 16178
rect 17574 16174 17608 16287
rect 18197 16178 18232 16411
rect 18476 16363 18542 16370
rect 18476 16329 18492 16363
rect 18526 16329 18542 16363
rect 18476 16318 18542 16329
rect 18668 16318 18704 16411
rect 18476 16317 18704 16318
rect 18904 16317 18940 16411
rect 19140 16317 19176 16411
rect 18476 16288 19176 16317
rect 18594 16287 19176 16288
rect 18594 16246 18660 16287
rect 18594 16212 18610 16246
rect 18644 16212 18660 16246
rect 18594 16205 18660 16212
rect 18197 16174 18586 16178
rect 19022 16174 19056 16287
rect 19717 16180 19752 16413
rect 19996 16365 20062 16372
rect 19996 16331 20012 16365
rect 20046 16331 20062 16365
rect 19996 16320 20062 16331
rect 20188 16320 20224 16413
rect 19996 16319 20224 16320
rect 20424 16319 20460 16413
rect 20660 16319 20696 16413
rect 19996 16290 20696 16319
rect 20114 16289 20696 16290
rect 20114 16248 20180 16289
rect 20114 16214 20130 16248
rect 20164 16214 20180 16248
rect 20114 16207 20180 16214
rect 19717 16176 20106 16180
rect 20542 16176 20576 16289
rect 21165 16180 21200 16413
rect 21444 16365 21510 16372
rect 21444 16331 21460 16365
rect 21494 16331 21510 16365
rect 21444 16320 21510 16331
rect 21636 16320 21672 16413
rect 21444 16319 21672 16320
rect 21872 16319 21908 16413
rect 22108 16319 22144 16413
rect 22657 16411 22703 16423
rect 22775 16599 22821 16611
rect 22775 16423 22781 16599
rect 22815 16423 22821 16599
rect 22775 16411 22821 16423
rect 22893 16599 22939 16611
rect 22893 16423 22899 16599
rect 22933 16423 22939 16599
rect 22893 16411 22939 16423
rect 23011 16599 23057 16611
rect 23011 16423 23017 16599
rect 23051 16423 23057 16599
rect 23011 16411 23057 16423
rect 23129 16599 23175 16611
rect 23129 16423 23135 16599
rect 23169 16423 23175 16599
rect 23129 16411 23175 16423
rect 23247 16599 23293 16611
rect 23247 16423 23253 16599
rect 23287 16423 23293 16599
rect 23247 16411 23293 16423
rect 23365 16599 23411 16611
rect 23365 16423 23371 16599
rect 23405 16423 23411 16599
rect 23365 16411 23411 16423
rect 23483 16599 23529 16611
rect 23483 16423 23489 16599
rect 23523 16423 23529 16599
rect 23483 16411 23529 16423
rect 23601 16599 23647 16611
rect 23601 16423 23607 16599
rect 23641 16423 23647 16599
rect 23601 16411 23647 16423
rect 23719 16599 23765 16611
rect 23719 16423 23725 16599
rect 23759 16423 23765 16599
rect 23719 16411 23765 16423
rect 24105 16599 24151 16611
rect 24105 16423 24111 16599
rect 24145 16423 24151 16599
rect 24105 16411 24151 16423
rect 24223 16599 24269 16611
rect 24223 16423 24229 16599
rect 24263 16423 24269 16599
rect 24223 16411 24269 16423
rect 24341 16599 24387 16611
rect 24341 16423 24347 16599
rect 24381 16423 24387 16599
rect 24341 16411 24387 16423
rect 24459 16599 24505 16611
rect 24459 16423 24465 16599
rect 24499 16423 24505 16599
rect 24459 16411 24505 16423
rect 24577 16599 24623 16611
rect 24577 16423 24583 16599
rect 24617 16423 24623 16599
rect 24577 16411 24623 16423
rect 24695 16599 24741 16611
rect 24695 16423 24701 16599
rect 24735 16423 24741 16599
rect 24695 16411 24741 16423
rect 24813 16599 24859 16611
rect 24813 16423 24819 16599
rect 24853 16423 24859 16599
rect 24813 16411 24859 16423
rect 24931 16599 24977 16611
rect 24931 16423 24937 16599
rect 24971 16423 24977 16599
rect 24931 16411 24977 16423
rect 25049 16599 25095 16611
rect 25049 16423 25055 16599
rect 25089 16423 25095 16599
rect 25049 16411 25095 16423
rect 25167 16599 25213 16611
rect 25167 16423 25173 16599
rect 25207 16423 25213 16599
rect 25167 16411 25213 16423
rect 21444 16290 22144 16319
rect 21562 16289 22144 16290
rect 21562 16248 21628 16289
rect 21562 16214 21578 16248
rect 21612 16214 21628 16248
rect 21562 16207 21628 16214
rect 21165 16176 21554 16180
rect 21990 16176 22024 16289
rect 22663 16178 22698 16411
rect 22942 16363 23008 16370
rect 22942 16329 22958 16363
rect 22992 16329 23008 16363
rect 22942 16318 23008 16329
rect 23134 16318 23170 16411
rect 22942 16317 23170 16318
rect 23370 16317 23406 16411
rect 23606 16317 23642 16411
rect 22942 16288 23642 16317
rect 23060 16287 23642 16288
rect 23060 16246 23126 16287
rect 23060 16212 23076 16246
rect 23110 16212 23126 16246
rect 23060 16205 23126 16212
rect 16749 16162 17143 16174
rect 16749 16149 17103 16162
rect 16156 16014 16256 16036
rect 16156 15960 16180 16014
rect 16234 15960 16256 16014
rect 16156 15936 16256 15960
rect 16070 15776 16116 15788
rect 15714 15772 15874 15776
rect 15714 15635 15790 15772
rect 16178 15744 16232 15936
rect 16268 15884 16368 15908
rect 16268 15830 16292 15884
rect 16346 15830 16368 15884
rect 16268 15808 16368 15830
rect 15883 15738 15949 15744
rect 15883 15704 15899 15738
rect 15933 15704 15949 15738
rect 15883 15659 15949 15704
rect 16001 15738 16232 15744
rect 16001 15704 16017 15738
rect 16051 15704 16232 15738
rect 16001 15688 16232 15704
rect 16292 15659 16346 15808
rect 15883 15651 16346 15659
rect 15712 15575 15722 15635
rect 15784 15575 15794 15635
rect 15882 15619 16346 15651
rect 16749 15496 16853 16149
rect 17097 15986 17103 16149
rect 17137 15986 17143 16162
rect 17097 15974 17143 15986
rect 17215 16162 17261 16174
rect 17215 15986 17221 16162
rect 17255 15986 17261 16162
rect 17215 15979 17261 15986
rect 17212 15974 17261 15979
rect 17332 16162 17378 16174
rect 17212 15813 17255 15974
rect 17332 15813 17338 16162
rect 17212 15786 17338 15813
rect 17372 15786 17378 16162
rect 17212 15774 17378 15786
rect 17450 16162 17496 16174
rect 17450 15786 17456 16162
rect 17490 15786 17496 16162
rect 17450 15774 17496 15786
rect 17568 16162 17614 16174
rect 17568 15786 17574 16162
rect 17608 15786 17614 16162
rect 18197 16162 18591 16174
rect 18197 16149 18551 16162
rect 17654 16016 17754 16034
rect 17654 15962 17677 16016
rect 17731 15962 17754 16016
rect 17654 15934 17754 15962
rect 17568 15774 17614 15786
rect 17212 15770 17372 15774
rect 17212 15633 17288 15770
rect 17676 15742 17730 15934
rect 17766 15878 17866 15906
rect 17766 15824 17789 15878
rect 17843 15824 17866 15878
rect 17766 15806 17866 15824
rect 17381 15736 17447 15742
rect 17381 15702 17397 15736
rect 17431 15702 17447 15736
rect 17381 15657 17447 15702
rect 17499 15736 17730 15742
rect 17499 15702 17515 15736
rect 17549 15702 17730 15736
rect 17499 15686 17730 15702
rect 17790 15657 17844 15806
rect 17381 15649 17844 15657
rect 17210 15573 17220 15633
rect 17282 15573 17292 15633
rect 17380 15617 17844 15649
rect 12477 15438 15355 15486
rect 9287 15407 9359 15437
rect 12477 15409 12524 15438
rect 15686 15436 16853 15496
rect 15686 15409 15745 15436
rect 6306 15335 9359 15407
rect 9397 15336 12524 15409
rect 12552 15336 15745 15409
rect 18197 15407 18301 16149
rect 18545 15986 18551 16149
rect 18585 15986 18591 16162
rect 18545 15974 18591 15986
rect 18663 16162 18709 16174
rect 18663 15986 18669 16162
rect 18703 15986 18709 16162
rect 18663 15979 18709 15986
rect 18660 15974 18709 15979
rect 18780 16162 18826 16174
rect 18660 15813 18703 15974
rect 18780 15813 18786 16162
rect 18660 15786 18786 15813
rect 18820 15786 18826 16162
rect 18660 15774 18826 15786
rect 18898 16162 18944 16174
rect 18898 15786 18904 16162
rect 18938 15786 18944 16162
rect 18898 15774 18944 15786
rect 19016 16162 19062 16174
rect 19016 15786 19022 16162
rect 19056 15786 19062 16162
rect 19717 16164 20111 16176
rect 19717 16151 20071 16164
rect 19102 16009 19202 16034
rect 19102 15955 19125 16009
rect 19179 15955 19202 16009
rect 19102 15934 19202 15955
rect 19016 15774 19062 15786
rect 18660 15770 18820 15774
rect 18660 15633 18736 15770
rect 19124 15742 19178 15934
rect 19214 15884 19314 15906
rect 19214 15830 19241 15884
rect 19295 15830 19314 15884
rect 19214 15806 19314 15830
rect 18829 15736 18895 15742
rect 18829 15702 18845 15736
rect 18879 15702 18895 15736
rect 18829 15657 18895 15702
rect 18947 15736 19178 15742
rect 18947 15702 18963 15736
rect 18997 15702 19178 15736
rect 18947 15686 19178 15702
rect 19238 15657 19292 15806
rect 18829 15649 19292 15657
rect 18658 15573 18668 15633
rect 18730 15573 18740 15633
rect 18828 15617 19292 15649
rect 6306 15307 6378 15335
rect 9397 15307 9476 15336
rect 12552 15307 12638 15336
rect 15777 15334 18301 15407
rect 19717 15402 19821 16151
rect 20065 15988 20071 16151
rect 20105 15988 20111 16164
rect 20065 15976 20111 15988
rect 20183 16164 20229 16176
rect 20183 15988 20189 16164
rect 20223 15988 20229 16164
rect 20183 15981 20229 15988
rect 20180 15976 20229 15981
rect 20300 16164 20346 16176
rect 20180 15815 20223 15976
rect 20300 15815 20306 16164
rect 20180 15788 20306 15815
rect 20340 15788 20346 16164
rect 20180 15776 20346 15788
rect 20418 16164 20464 16176
rect 20418 15788 20424 16164
rect 20458 15788 20464 16164
rect 20418 15776 20464 15788
rect 20536 16164 20582 16176
rect 20536 15788 20542 16164
rect 20576 15788 20582 16164
rect 21165 16164 21559 16176
rect 21165 16151 21519 16164
rect 20622 16014 20722 16036
rect 20622 15960 20644 16014
rect 20698 15960 20722 16014
rect 20622 15936 20722 15960
rect 20536 15776 20582 15788
rect 20180 15772 20340 15776
rect 20180 15635 20256 15772
rect 20644 15744 20698 15936
rect 20734 15884 20834 15908
rect 20734 15830 20757 15884
rect 20811 15830 20834 15884
rect 20734 15808 20834 15830
rect 20349 15738 20415 15744
rect 20349 15704 20365 15738
rect 20399 15704 20415 15738
rect 20349 15659 20415 15704
rect 20467 15738 20698 15744
rect 20467 15704 20483 15738
rect 20517 15704 20698 15738
rect 20467 15688 20698 15704
rect 20758 15659 20812 15808
rect 20349 15651 20812 15659
rect 20178 15575 20188 15635
rect 20250 15575 20260 15635
rect 20348 15619 20812 15651
rect 15777 15307 15851 15334
rect 3263 15235 6378 15307
rect 6407 15235 9476 15307
rect 1768 15042 1778 15102
rect 1858 15042 1868 15102
rect 1768 15002 1868 15042
rect 862 14945 2665 15002
rect 862 14658 899 14945
rect 1456 14858 1490 14945
rect 2631 14858 2665 14945
rect 977 14846 1023 14858
rect 504 14646 550 14658
rect 504 14470 510 14646
rect 544 14470 550 14646
rect 504 14458 550 14470
rect 622 14646 668 14658
rect 622 14470 628 14646
rect 662 14470 668 14646
rect 622 14458 668 14470
rect 740 14646 786 14658
rect 740 14470 746 14646
rect 780 14470 786 14646
rect 740 14458 786 14470
rect 858 14646 904 14658
rect 858 14470 864 14646
rect 898 14470 904 14646
rect 858 14458 904 14470
rect 977 14470 983 14846
rect 1017 14470 1023 14846
rect 977 14458 1023 14470
rect 1095 14846 1141 14858
rect 1095 14470 1101 14846
rect 1135 14470 1141 14846
rect 1095 14458 1141 14470
rect 1213 14846 1259 14858
rect 1213 14470 1219 14846
rect 1253 14470 1259 14846
rect 1213 14458 1259 14470
rect 1331 14846 1377 14858
rect 1331 14470 1337 14846
rect 1371 14470 1377 14846
rect 1331 14458 1377 14470
rect 1450 14846 1496 14858
rect 1450 14470 1456 14846
rect 1490 14470 1496 14846
rect 1450 14458 1496 14470
rect 1568 14846 1614 14858
rect 1568 14470 1574 14846
rect 1608 14470 1614 14846
rect 1568 14458 1614 14470
rect 1686 14846 1732 14858
rect 1686 14470 1692 14846
rect 1726 14470 1732 14846
rect 1686 14458 1732 14470
rect 1804 14846 1850 14858
rect 1804 14470 1810 14846
rect 1844 14470 1850 14846
rect 1804 14458 1850 14470
rect 1922 14846 1968 14858
rect 1922 14470 1928 14846
rect 1962 14470 1968 14846
rect 1922 14458 1968 14470
rect 2040 14846 2086 14858
rect 2040 14470 2046 14846
rect 2080 14470 2086 14846
rect 2040 14458 2086 14470
rect 2158 14846 2204 14858
rect 2158 14470 2164 14846
rect 2198 14470 2204 14846
rect 2158 14458 2204 14470
rect 2271 14846 2317 14858
rect 2271 14470 2277 14846
rect 2311 14470 2317 14846
rect 2271 14458 2317 14470
rect 2389 14846 2435 14858
rect 2389 14470 2395 14846
rect 2429 14470 2435 14846
rect 2389 14458 2435 14470
rect 2507 14846 2553 14858
rect 2507 14470 2513 14846
rect 2547 14470 2553 14846
rect 2507 14458 2553 14470
rect 2625 14846 2671 14858
rect 2625 14470 2631 14846
rect 2665 14658 2671 14846
rect 2665 14646 2758 14658
rect 2665 14470 2718 14646
rect 2752 14470 2758 14646
rect 2625 14458 2758 14470
rect 2830 14646 2876 14658
rect 2830 14470 2836 14646
rect 2870 14470 2876 14646
rect 2830 14458 2876 14470
rect 2948 14646 2994 14658
rect 2948 14470 2954 14646
rect 2988 14470 2994 14646
rect 2948 14458 2994 14470
rect 3066 14646 3112 14658
rect 3066 14470 3072 14646
rect 3106 14470 3112 14646
rect 3066 14458 3112 14470
rect 509 14104 544 14458
rect 983 14374 1017 14458
rect 2164 14374 2198 14458
rect 983 14332 2198 14374
rect 983 14312 1017 14332
rect 660 14296 1017 14312
rect 660 14262 676 14296
rect 710 14262 1017 14296
rect 3072 14272 3107 14458
rect 660 14246 1017 14262
rect 1970 14255 3107 14272
rect 1970 14221 1986 14255
rect 2020 14221 3107 14255
rect 1970 14205 3107 14221
rect 363 13958 544 14104
rect 1840 14159 1932 14169
rect 1840 14097 1850 14159
rect 1920 14097 1932 14159
rect 1840 14084 1932 14097
rect 2925 14159 3017 14172
rect 2925 14096 2934 14159
rect 3005 14096 3017 14159
rect 2925 14087 3017 14096
rect 1620 14042 1685 14045
rect 1616 14039 1685 14042
rect 1610 13979 1620 14039
rect 1679 13979 1685 14039
rect 1616 13975 1685 13979
rect 1620 13973 1685 13975
rect 363 12705 443 13958
rect 509 13696 544 13958
rect 1958 13876 2050 13884
rect 1958 13811 1970 13876
rect 2038 13811 2050 13876
rect 1958 13799 2050 13811
rect 509 13649 1413 13696
rect 3072 13695 3107 14205
rect 3263 14052 3350 15235
rect 4912 15042 4922 15102
rect 5002 15042 5012 15102
rect 4912 15002 5012 15042
rect 4006 14945 5809 15002
rect 4006 14658 4043 14945
rect 4600 14858 4634 14945
rect 5775 14858 5809 14945
rect 4121 14846 4167 14858
rect 3648 14646 3694 14658
rect 3648 14470 3654 14646
rect 3688 14470 3694 14646
rect 3648 14458 3694 14470
rect 3766 14646 3812 14658
rect 3766 14470 3772 14646
rect 3806 14470 3812 14646
rect 3766 14458 3812 14470
rect 3884 14646 3930 14658
rect 3884 14470 3890 14646
rect 3924 14470 3930 14646
rect 3884 14458 3930 14470
rect 4002 14646 4048 14658
rect 4002 14470 4008 14646
rect 4042 14470 4048 14646
rect 4002 14458 4048 14470
rect 4121 14470 4127 14846
rect 4161 14470 4167 14846
rect 4121 14458 4167 14470
rect 4239 14846 4285 14858
rect 4239 14470 4245 14846
rect 4279 14470 4285 14846
rect 4239 14458 4285 14470
rect 4357 14846 4403 14858
rect 4357 14470 4363 14846
rect 4397 14470 4403 14846
rect 4357 14458 4403 14470
rect 4475 14846 4521 14858
rect 4475 14470 4481 14846
rect 4515 14470 4521 14846
rect 4475 14458 4521 14470
rect 4594 14846 4640 14858
rect 4594 14470 4600 14846
rect 4634 14470 4640 14846
rect 4594 14458 4640 14470
rect 4712 14846 4758 14858
rect 4712 14470 4718 14846
rect 4752 14470 4758 14846
rect 4712 14458 4758 14470
rect 4830 14846 4876 14858
rect 4830 14470 4836 14846
rect 4870 14470 4876 14846
rect 4830 14458 4876 14470
rect 4948 14846 4994 14858
rect 4948 14470 4954 14846
rect 4988 14470 4994 14846
rect 4948 14458 4994 14470
rect 5066 14846 5112 14858
rect 5066 14470 5072 14846
rect 5106 14470 5112 14846
rect 5066 14458 5112 14470
rect 5184 14846 5230 14858
rect 5184 14470 5190 14846
rect 5224 14470 5230 14846
rect 5184 14458 5230 14470
rect 5302 14846 5348 14858
rect 5302 14470 5308 14846
rect 5342 14470 5348 14846
rect 5302 14458 5348 14470
rect 5415 14846 5461 14858
rect 5415 14470 5421 14846
rect 5455 14470 5461 14846
rect 5415 14458 5461 14470
rect 5533 14846 5579 14858
rect 5533 14470 5539 14846
rect 5573 14470 5579 14846
rect 5533 14458 5579 14470
rect 5651 14846 5697 14858
rect 5651 14470 5657 14846
rect 5691 14470 5697 14846
rect 5651 14458 5697 14470
rect 5769 14846 5815 14858
rect 5769 14470 5775 14846
rect 5809 14658 5815 14846
rect 5809 14646 5902 14658
rect 5809 14470 5862 14646
rect 5896 14470 5902 14646
rect 5769 14458 5902 14470
rect 5974 14646 6020 14658
rect 5974 14470 5980 14646
rect 6014 14470 6020 14646
rect 5974 14458 6020 14470
rect 6092 14646 6138 14658
rect 6092 14470 6098 14646
rect 6132 14470 6138 14646
rect 6092 14458 6138 14470
rect 6210 14646 6256 14658
rect 6210 14470 6216 14646
rect 6250 14470 6256 14646
rect 6210 14458 6256 14470
rect 3653 14104 3688 14458
rect 4127 14374 4161 14458
rect 5308 14374 5342 14458
rect 4127 14332 5342 14374
rect 4127 14312 4161 14332
rect 3804 14296 4161 14312
rect 3804 14262 3820 14296
rect 3854 14262 4161 14296
rect 6216 14272 6251 14458
rect 3804 14246 4161 14262
rect 5114 14255 6251 14272
rect 5114 14221 5130 14255
rect 5164 14221 6251 14255
rect 5114 14205 6251 14221
rect 3190 14044 3350 14052
rect 3182 13976 3192 14044
rect 3249 13976 3350 14044
rect 3190 13968 3350 13976
rect 3509 13958 3688 14104
rect 4984 14159 5076 14169
rect 4984 14097 4994 14159
rect 5064 14097 5076 14159
rect 4984 14084 5076 14097
rect 6069 14159 6161 14172
rect 6069 14096 6078 14159
rect 6149 14096 6161 14159
rect 6069 14087 6161 14096
rect 4764 14042 4829 14045
rect 4760 14039 4829 14042
rect 4754 13979 4764 14039
rect 4823 13979 4829 14039
rect 4760 13975 4829 13979
rect 4764 13973 4829 13975
rect 3190 13876 3260 13884
rect 3182 13808 3192 13876
rect 3249 13808 3260 13876
rect 3190 13800 3260 13808
rect 1378 13525 1412 13649
rect 1735 13648 3107 13695
rect 1735 13635 1801 13648
rect 1735 13601 1751 13635
rect 1785 13601 1801 13635
rect 1735 13585 1801 13601
rect 2239 13525 2273 13648
rect 1372 13513 1418 13525
rect 1372 13337 1378 13513
rect 1412 13337 1418 13513
rect 1372 13325 1418 13337
rect 1490 13513 1614 13525
rect 1490 13337 1496 13513
rect 1530 13337 1574 13513
rect 1490 13325 1574 13337
rect 1496 12958 1530 13325
rect 1568 13137 1574 13325
rect 1608 13137 1614 13513
rect 1568 13125 1614 13137
rect 1686 13513 1732 13525
rect 1686 13137 1692 13513
rect 1726 13137 1732 13513
rect 1686 13125 1732 13137
rect 1804 13513 1850 13525
rect 1804 13137 1810 13513
rect 1844 13137 1850 13513
rect 1804 13125 1850 13137
rect 1922 13513 1968 13525
rect 1922 13137 1928 13513
rect 1962 13137 1968 13513
rect 1922 13125 1968 13137
rect 2040 13513 2160 13525
rect 2040 13137 2046 13513
rect 2080 13337 2120 13513
rect 2154 13337 2160 13513
rect 2080 13325 2160 13337
rect 2232 13513 2278 13525
rect 2232 13337 2238 13513
rect 2272 13337 2278 13513
rect 2232 13325 2278 13337
rect 2080 13137 2086 13325
rect 2040 13125 2086 13137
rect 1810 13052 1844 13125
rect 1793 13036 1859 13052
rect 1793 13002 1809 13036
rect 1843 13002 1859 13036
rect 1793 12986 1859 13002
rect 2120 12958 2154 13325
rect 1496 12906 2154 12958
rect 1764 12884 1856 12906
rect 1764 12832 1778 12884
rect 1844 12832 1856 12884
rect 1764 12828 1856 12832
rect 363 12637 3366 12705
rect 1768 12308 1778 12368
rect 1858 12308 1868 12368
rect 1768 12268 1868 12308
rect 862 12211 2665 12268
rect 862 11924 899 12211
rect 1456 12124 1490 12211
rect 2631 12124 2665 12211
rect 977 12112 1023 12124
rect 504 11912 550 11924
rect 504 11736 510 11912
rect 544 11736 550 11912
rect 504 11724 550 11736
rect 622 11912 668 11924
rect 622 11736 628 11912
rect 662 11736 668 11912
rect 622 11724 668 11736
rect 740 11912 786 11924
rect 740 11736 746 11912
rect 780 11736 786 11912
rect 740 11724 786 11736
rect 858 11912 904 11924
rect 858 11736 864 11912
rect 898 11736 904 11912
rect 858 11724 904 11736
rect 977 11736 983 12112
rect 1017 11736 1023 12112
rect 977 11724 1023 11736
rect 1095 12112 1141 12124
rect 1095 11736 1101 12112
rect 1135 11736 1141 12112
rect 1095 11724 1141 11736
rect 1213 12112 1259 12124
rect 1213 11736 1219 12112
rect 1253 11736 1259 12112
rect 1213 11724 1259 11736
rect 1331 12112 1377 12124
rect 1331 11736 1337 12112
rect 1371 11736 1377 12112
rect 1331 11724 1377 11736
rect 1450 12112 1496 12124
rect 1450 11736 1456 12112
rect 1490 11736 1496 12112
rect 1450 11724 1496 11736
rect 1568 12112 1614 12124
rect 1568 11736 1574 12112
rect 1608 11736 1614 12112
rect 1568 11724 1614 11736
rect 1686 12112 1732 12124
rect 1686 11736 1692 12112
rect 1726 11736 1732 12112
rect 1686 11724 1732 11736
rect 1804 12112 1850 12124
rect 1804 11736 1810 12112
rect 1844 11736 1850 12112
rect 1804 11724 1850 11736
rect 1922 12112 1968 12124
rect 1922 11736 1928 12112
rect 1962 11736 1968 12112
rect 1922 11724 1968 11736
rect 2040 12112 2086 12124
rect 2040 11736 2046 12112
rect 2080 11736 2086 12112
rect 2040 11724 2086 11736
rect 2158 12112 2204 12124
rect 2158 11736 2164 12112
rect 2198 11736 2204 12112
rect 2158 11724 2204 11736
rect 2271 12112 2317 12124
rect 2271 11736 2277 12112
rect 2311 11736 2317 12112
rect 2271 11724 2317 11736
rect 2389 12112 2435 12124
rect 2389 11736 2395 12112
rect 2429 11736 2435 12112
rect 2389 11724 2435 11736
rect 2507 12112 2553 12124
rect 2507 11736 2513 12112
rect 2547 11736 2553 12112
rect 2507 11724 2553 11736
rect 2625 12112 2671 12124
rect 2625 11736 2631 12112
rect 2665 11924 2671 12112
rect 2665 11912 2758 11924
rect 2665 11736 2718 11912
rect 2752 11736 2758 11912
rect 2625 11724 2758 11736
rect 2830 11912 2876 11924
rect 2830 11736 2836 11912
rect 2870 11736 2876 11912
rect 2830 11724 2876 11736
rect 2948 11912 2994 11924
rect 2948 11736 2954 11912
rect 2988 11736 2994 11912
rect 2948 11724 2994 11736
rect 3066 11912 3112 11924
rect 3066 11736 3072 11912
rect 3106 11736 3112 11912
rect 3066 11724 3112 11736
rect 509 11370 544 11724
rect 983 11640 1017 11724
rect 2164 11640 2198 11724
rect 983 11598 2198 11640
rect 983 11578 1017 11598
rect 660 11562 1017 11578
rect 660 11528 676 11562
rect 710 11528 1017 11562
rect 3072 11538 3107 11724
rect 660 11512 1017 11528
rect 1970 11521 3107 11538
rect 1970 11487 1986 11521
rect 2020 11487 3107 11521
rect 1970 11471 3107 11487
rect 64 11361 544 11370
rect 64 11232 80 11361
rect 191 11232 544 11361
rect 1840 11425 1932 11435
rect 1840 11363 1850 11425
rect 1920 11363 1932 11425
rect 1840 11350 1932 11363
rect 2925 11425 3017 11438
rect 2925 11362 2934 11425
rect 3005 11362 3017 11425
rect 2925 11353 3017 11362
rect 1620 11308 1685 11311
rect 1616 11305 1685 11308
rect 1610 11245 1620 11305
rect 1679 11245 1685 11305
rect 1616 11241 1685 11245
rect 1620 11239 1685 11241
rect 64 11224 544 11232
rect 509 10962 544 11224
rect 1958 11142 2050 11150
rect 1958 11077 1970 11142
rect 2038 11077 2050 11142
rect 1958 11065 2050 11077
rect -570 10937 173 10950
rect -570 10936 142 10937
rect -570 10879 -547 10936
rect -425 10879 142 10936
rect -570 10867 142 10879
rect 201 10867 211 10937
rect 509 10915 1413 10962
rect 3072 10961 3107 11471
rect 3295 11318 3366 12637
rect 3509 12704 3600 13958
rect 3653 13696 3688 13958
rect 5102 13876 5194 13884
rect 5102 13811 5114 13876
rect 5182 13811 5194 13876
rect 5102 13799 5194 13811
rect 3653 13649 4557 13696
rect 6216 13695 6251 14205
rect 6407 14052 6494 15235
rect 9538 15234 12638 15307
rect 12684 15234 15851 15307
rect 18876 15330 19821 15402
rect 18876 15306 18955 15330
rect 15884 15234 18955 15306
rect 21165 15302 21269 16151
rect 21513 15988 21519 16151
rect 21553 15988 21559 16164
rect 21513 15976 21559 15988
rect 21631 16164 21677 16176
rect 21631 15988 21637 16164
rect 21671 15988 21677 16164
rect 21631 15981 21677 15988
rect 21628 15976 21677 15981
rect 21748 16164 21794 16176
rect 21628 15815 21671 15976
rect 21748 15815 21754 16164
rect 21628 15788 21754 15815
rect 21788 15788 21794 16164
rect 21628 15776 21794 15788
rect 21866 16164 21912 16176
rect 21866 15788 21872 16164
rect 21906 15788 21912 16164
rect 21866 15776 21912 15788
rect 21984 16164 22030 16176
rect 21984 15788 21990 16164
rect 22024 15788 22030 16164
rect 22663 16174 23052 16178
rect 23488 16174 23522 16287
rect 24111 16178 24146 16411
rect 24390 16363 24456 16370
rect 24390 16329 24406 16363
rect 24440 16329 24456 16363
rect 24390 16318 24456 16329
rect 24582 16318 24618 16411
rect 24390 16317 24618 16318
rect 24818 16317 24854 16411
rect 25054 16317 25090 16411
rect 24390 16288 25090 16317
rect 24508 16287 25090 16288
rect 24508 16246 24574 16287
rect 24508 16212 24524 16246
rect 24558 16212 24574 16246
rect 24508 16205 24574 16212
rect 24111 16174 24500 16178
rect 24936 16174 24970 16287
rect 22663 16162 23057 16174
rect 22663 16149 23017 16162
rect 22070 16011 22170 16036
rect 22070 15957 22094 16011
rect 22148 15957 22170 16011
rect 22070 15936 22170 15957
rect 21984 15776 22030 15788
rect 21628 15772 21788 15776
rect 21628 15635 21704 15772
rect 22092 15744 22146 15936
rect 22182 15879 22282 15908
rect 22182 15825 22205 15879
rect 22259 15825 22282 15879
rect 22182 15808 22282 15825
rect 21797 15738 21863 15744
rect 21797 15704 21813 15738
rect 21847 15704 21863 15738
rect 21797 15659 21863 15704
rect 21915 15738 22146 15744
rect 21915 15704 21931 15738
rect 21965 15704 22146 15738
rect 21915 15688 22146 15704
rect 22206 15659 22260 15808
rect 21797 15651 22260 15659
rect 21626 15575 21636 15635
rect 21698 15575 21708 15635
rect 21796 15619 22260 15651
rect 22663 15338 22767 16149
rect 23011 15986 23017 16149
rect 23051 15986 23057 16162
rect 23011 15974 23057 15986
rect 23129 16162 23175 16174
rect 23129 15986 23135 16162
rect 23169 15986 23175 16162
rect 23129 15979 23175 15986
rect 23126 15974 23175 15979
rect 23246 16162 23292 16174
rect 23126 15813 23169 15974
rect 23246 15813 23252 16162
rect 23126 15786 23252 15813
rect 23286 15786 23292 16162
rect 23126 15774 23292 15786
rect 23364 16162 23410 16174
rect 23364 15786 23370 16162
rect 23404 15786 23410 16162
rect 23364 15774 23410 15786
rect 23482 16162 23528 16174
rect 23482 15786 23488 16162
rect 23522 15786 23528 16162
rect 24111 16162 24505 16174
rect 24111 16156 24465 16162
rect 24110 16149 24465 16156
rect 23568 16012 23668 16034
rect 24110 16016 24218 16149
rect 23568 15958 23588 16012
rect 23642 15958 23668 16012
rect 23568 15934 23668 15958
rect 24109 15994 24218 16016
rect 23482 15774 23528 15786
rect 23126 15770 23286 15774
rect 23126 15633 23202 15770
rect 23590 15742 23644 15934
rect 23680 15881 23780 15906
rect 23680 15826 23703 15881
rect 23757 15826 23780 15881
rect 23680 15806 23780 15826
rect 23295 15736 23361 15742
rect 23295 15702 23311 15736
rect 23345 15702 23361 15736
rect 23295 15657 23361 15702
rect 23413 15736 23644 15742
rect 23413 15702 23429 15736
rect 23463 15702 23644 15736
rect 23413 15686 23644 15702
rect 23704 15657 23758 15806
rect 23295 15649 23758 15657
rect 23124 15573 23134 15633
rect 23196 15573 23206 15633
rect 23294 15617 23758 15649
rect 24109 15467 24217 15994
rect 24459 15986 24465 16149
rect 24499 15986 24505 16162
rect 24459 15974 24505 15986
rect 24577 16162 24623 16174
rect 24577 15986 24583 16162
rect 24617 15986 24623 16162
rect 24577 15979 24623 15986
rect 24574 15974 24623 15979
rect 24694 16162 24740 16174
rect 24574 15813 24617 15974
rect 24694 15813 24700 16162
rect 24574 15786 24700 15813
rect 24734 15786 24740 16162
rect 24574 15774 24740 15786
rect 24812 16162 24858 16174
rect 24812 15786 24818 16162
rect 24852 15786 24858 16162
rect 24812 15774 24858 15786
rect 24930 16162 24976 16174
rect 24930 15786 24936 16162
rect 24970 15786 24976 16162
rect 25266 16107 25330 16962
rect 25506 16182 25569 17255
rect 25506 16181 25711 16182
rect 25506 16122 25630 16181
rect 25701 16122 25711 16181
rect 25266 16085 25425 16107
rect 25266 16034 25346 16085
rect 25016 16021 25346 16034
rect 25415 16021 25425 16085
rect 25016 16010 25425 16021
rect 25016 15934 25330 16010
rect 24930 15774 24976 15786
rect 24574 15770 24734 15774
rect 24574 15633 24650 15770
rect 25038 15742 25092 15934
rect 25506 15906 25569 16122
rect 25128 15806 25569 15906
rect 24743 15736 24809 15742
rect 24743 15702 24759 15736
rect 24793 15702 24809 15736
rect 24743 15657 24809 15702
rect 24861 15736 25092 15742
rect 24861 15702 24877 15736
rect 24911 15702 25092 15736
rect 24861 15686 25092 15702
rect 25152 15657 25206 15806
rect 24743 15649 25206 15657
rect 24572 15573 24582 15633
rect 24644 15573 24654 15633
rect 24742 15617 25206 15649
rect 19028 15234 21269 15302
rect 22177 15245 22767 15338
rect 24111 15338 24217 15467
rect 24111 15292 25409 15338
rect 24112 15245 25409 15292
rect 8044 15038 8054 15098
rect 8134 15038 8144 15098
rect 8044 14998 8144 15038
rect 7138 14941 8941 14998
rect 7138 14654 7175 14941
rect 7732 14854 7766 14941
rect 8907 14854 8941 14941
rect 7253 14842 7299 14854
rect 6780 14642 6826 14654
rect 6780 14466 6786 14642
rect 6820 14466 6826 14642
rect 6780 14454 6826 14466
rect 6898 14642 6944 14654
rect 6898 14466 6904 14642
rect 6938 14466 6944 14642
rect 6898 14454 6944 14466
rect 7016 14642 7062 14654
rect 7016 14466 7022 14642
rect 7056 14466 7062 14642
rect 7016 14454 7062 14466
rect 7134 14642 7180 14654
rect 7134 14466 7140 14642
rect 7174 14466 7180 14642
rect 7134 14454 7180 14466
rect 7253 14466 7259 14842
rect 7293 14466 7299 14842
rect 7253 14454 7299 14466
rect 7371 14842 7417 14854
rect 7371 14466 7377 14842
rect 7411 14466 7417 14842
rect 7371 14454 7417 14466
rect 7489 14842 7535 14854
rect 7489 14466 7495 14842
rect 7529 14466 7535 14842
rect 7489 14454 7535 14466
rect 7607 14842 7653 14854
rect 7607 14466 7613 14842
rect 7647 14466 7653 14842
rect 7607 14454 7653 14466
rect 7726 14842 7772 14854
rect 7726 14466 7732 14842
rect 7766 14466 7772 14842
rect 7726 14454 7772 14466
rect 7844 14842 7890 14854
rect 7844 14466 7850 14842
rect 7884 14466 7890 14842
rect 7844 14454 7890 14466
rect 7962 14842 8008 14854
rect 7962 14466 7968 14842
rect 8002 14466 8008 14842
rect 7962 14454 8008 14466
rect 8080 14842 8126 14854
rect 8080 14466 8086 14842
rect 8120 14466 8126 14842
rect 8080 14454 8126 14466
rect 8198 14842 8244 14854
rect 8198 14466 8204 14842
rect 8238 14466 8244 14842
rect 8198 14454 8244 14466
rect 8316 14842 8362 14854
rect 8316 14466 8322 14842
rect 8356 14466 8362 14842
rect 8316 14454 8362 14466
rect 8434 14842 8480 14854
rect 8434 14466 8440 14842
rect 8474 14466 8480 14842
rect 8434 14454 8480 14466
rect 8547 14842 8593 14854
rect 8547 14466 8553 14842
rect 8587 14466 8593 14842
rect 8547 14454 8593 14466
rect 8665 14842 8711 14854
rect 8665 14466 8671 14842
rect 8705 14466 8711 14842
rect 8665 14454 8711 14466
rect 8783 14842 8829 14854
rect 8783 14466 8789 14842
rect 8823 14466 8829 14842
rect 8783 14454 8829 14466
rect 8901 14842 8947 14854
rect 8901 14466 8907 14842
rect 8941 14654 8947 14842
rect 8941 14642 9034 14654
rect 8941 14466 8994 14642
rect 9028 14466 9034 14642
rect 8901 14454 9034 14466
rect 9106 14642 9152 14654
rect 9106 14466 9112 14642
rect 9146 14466 9152 14642
rect 9106 14454 9152 14466
rect 9224 14642 9270 14654
rect 9224 14466 9230 14642
rect 9264 14466 9270 14642
rect 9224 14454 9270 14466
rect 9342 14642 9388 14654
rect 9342 14466 9348 14642
rect 9382 14466 9388 14642
rect 9342 14454 9388 14466
rect 6785 14100 6820 14454
rect 7259 14370 7293 14454
rect 8440 14370 8474 14454
rect 7259 14328 8474 14370
rect 7259 14308 7293 14328
rect 6936 14292 7293 14308
rect 6936 14258 6952 14292
rect 6986 14258 7293 14292
rect 9348 14268 9383 14454
rect 6936 14242 7293 14258
rect 8246 14251 9383 14268
rect 8246 14217 8262 14251
rect 8296 14217 9383 14251
rect 8246 14201 9383 14217
rect 6334 14044 6494 14052
rect 6326 13976 6336 14044
rect 6393 13976 6494 14044
rect 6334 13968 6494 13976
rect 6639 13967 6820 14100
rect 8116 14155 8208 14165
rect 8116 14093 8126 14155
rect 8196 14093 8208 14155
rect 8116 14080 8208 14093
rect 9201 14155 9293 14168
rect 9201 14092 9210 14155
rect 9281 14092 9293 14155
rect 9201 14083 9293 14092
rect 7896 14038 7961 14041
rect 7892 14035 7961 14038
rect 7886 13975 7896 14035
rect 7955 13975 7961 14035
rect 7892 13971 7961 13975
rect 7896 13969 7961 13971
rect 6638 13954 6820 13967
rect 6334 13876 6405 13884
rect 6326 13808 6336 13876
rect 6393 13808 6405 13876
rect 6334 13800 6405 13808
rect 4522 13525 4556 13649
rect 4879 13648 6251 13695
rect 4879 13635 4945 13648
rect 4879 13601 4895 13635
rect 4929 13601 4945 13635
rect 4879 13585 4945 13601
rect 5383 13525 5417 13648
rect 4516 13513 4562 13525
rect 4516 13337 4522 13513
rect 4556 13337 4562 13513
rect 4516 13325 4562 13337
rect 4634 13513 4758 13525
rect 4634 13337 4640 13513
rect 4674 13337 4718 13513
rect 4634 13325 4718 13337
rect 4640 12958 4674 13325
rect 4712 13137 4718 13325
rect 4752 13137 4758 13513
rect 4712 13125 4758 13137
rect 4830 13513 4876 13525
rect 4830 13137 4836 13513
rect 4870 13137 4876 13513
rect 4830 13125 4876 13137
rect 4948 13513 4994 13525
rect 4948 13137 4954 13513
rect 4988 13137 4994 13513
rect 4948 13125 4994 13137
rect 5066 13513 5112 13525
rect 5066 13137 5072 13513
rect 5106 13137 5112 13513
rect 5066 13125 5112 13137
rect 5184 13513 5304 13525
rect 5184 13137 5190 13513
rect 5224 13337 5264 13513
rect 5298 13337 5304 13513
rect 5224 13325 5304 13337
rect 5376 13513 5422 13525
rect 5376 13337 5382 13513
rect 5416 13337 5422 13513
rect 5376 13325 5422 13337
rect 5224 13137 5230 13325
rect 5184 13125 5230 13137
rect 4954 13052 4988 13125
rect 4937 13036 5003 13052
rect 4937 13002 4953 13036
rect 4987 13002 5003 13036
rect 4937 12986 5003 13002
rect 5264 12958 5298 13325
rect 4640 12906 5298 12958
rect 4908 12884 5000 12906
rect 4908 12832 4922 12884
rect 4988 12832 5000 12884
rect 4908 12828 5000 12832
rect 6638 12704 6741 13954
rect 6785 13692 6820 13954
rect 8234 13872 8326 13880
rect 8234 13807 8246 13872
rect 8314 13807 8326 13872
rect 8234 13795 8326 13807
rect 6785 13645 7689 13692
rect 9348 13691 9383 14201
rect 9538 14048 9625 15234
rect 11188 15038 11198 15098
rect 11278 15038 11288 15098
rect 11188 14998 11288 15038
rect 10282 14941 12085 14998
rect 10282 14654 10319 14941
rect 10876 14854 10910 14941
rect 12051 14854 12085 14941
rect 10397 14842 10443 14854
rect 9924 14642 9970 14654
rect 9924 14466 9930 14642
rect 9964 14466 9970 14642
rect 9924 14454 9970 14466
rect 10042 14642 10088 14654
rect 10042 14466 10048 14642
rect 10082 14466 10088 14642
rect 10042 14454 10088 14466
rect 10160 14642 10206 14654
rect 10160 14466 10166 14642
rect 10200 14466 10206 14642
rect 10160 14454 10206 14466
rect 10278 14642 10324 14654
rect 10278 14466 10284 14642
rect 10318 14466 10324 14642
rect 10278 14454 10324 14466
rect 10397 14466 10403 14842
rect 10437 14466 10443 14842
rect 10397 14454 10443 14466
rect 10515 14842 10561 14854
rect 10515 14466 10521 14842
rect 10555 14466 10561 14842
rect 10515 14454 10561 14466
rect 10633 14842 10679 14854
rect 10633 14466 10639 14842
rect 10673 14466 10679 14842
rect 10633 14454 10679 14466
rect 10751 14842 10797 14854
rect 10751 14466 10757 14842
rect 10791 14466 10797 14842
rect 10751 14454 10797 14466
rect 10870 14842 10916 14854
rect 10870 14466 10876 14842
rect 10910 14466 10916 14842
rect 10870 14454 10916 14466
rect 10988 14842 11034 14854
rect 10988 14466 10994 14842
rect 11028 14466 11034 14842
rect 10988 14454 11034 14466
rect 11106 14842 11152 14854
rect 11106 14466 11112 14842
rect 11146 14466 11152 14842
rect 11106 14454 11152 14466
rect 11224 14842 11270 14854
rect 11224 14466 11230 14842
rect 11264 14466 11270 14842
rect 11224 14454 11270 14466
rect 11342 14842 11388 14854
rect 11342 14466 11348 14842
rect 11382 14466 11388 14842
rect 11342 14454 11388 14466
rect 11460 14842 11506 14854
rect 11460 14466 11466 14842
rect 11500 14466 11506 14842
rect 11460 14454 11506 14466
rect 11578 14842 11624 14854
rect 11578 14466 11584 14842
rect 11618 14466 11624 14842
rect 11578 14454 11624 14466
rect 11691 14842 11737 14854
rect 11691 14466 11697 14842
rect 11731 14466 11737 14842
rect 11691 14454 11737 14466
rect 11809 14842 11855 14854
rect 11809 14466 11815 14842
rect 11849 14466 11855 14842
rect 11809 14454 11855 14466
rect 11927 14842 11973 14854
rect 11927 14466 11933 14842
rect 11967 14466 11973 14842
rect 11927 14454 11973 14466
rect 12045 14842 12091 14854
rect 12045 14466 12051 14842
rect 12085 14654 12091 14842
rect 12085 14642 12178 14654
rect 12085 14466 12138 14642
rect 12172 14466 12178 14642
rect 12045 14454 12178 14466
rect 12250 14642 12296 14654
rect 12250 14466 12256 14642
rect 12290 14466 12296 14642
rect 12250 14454 12296 14466
rect 12368 14642 12414 14654
rect 12368 14466 12374 14642
rect 12408 14466 12414 14642
rect 12368 14454 12414 14466
rect 12486 14642 12532 14654
rect 12486 14466 12492 14642
rect 12526 14466 12532 14642
rect 12486 14454 12532 14466
rect 9929 14100 9964 14454
rect 10403 14370 10437 14454
rect 11584 14370 11618 14454
rect 10403 14328 11618 14370
rect 10403 14308 10437 14328
rect 10080 14292 10437 14308
rect 10080 14258 10096 14292
rect 10130 14258 10437 14292
rect 12492 14268 12527 14454
rect 10080 14242 10437 14258
rect 11390 14251 12527 14268
rect 11390 14217 11406 14251
rect 11440 14217 12527 14251
rect 11390 14201 12527 14217
rect 9466 14040 9625 14048
rect 9458 13972 9468 14040
rect 9525 13972 9625 14040
rect 9466 13964 9625 13972
rect 9783 13954 9964 14100
rect 11260 14155 11352 14165
rect 11260 14093 11270 14155
rect 11340 14093 11352 14155
rect 11260 14080 11352 14093
rect 12345 14155 12437 14168
rect 12345 14092 12354 14155
rect 12425 14092 12437 14155
rect 12345 14083 12437 14092
rect 11040 14038 11105 14041
rect 11036 14035 11105 14038
rect 11030 13975 11040 14035
rect 11099 13975 11105 14035
rect 11036 13971 11105 13975
rect 11040 13969 11105 13971
rect 9466 13872 9536 13880
rect 9458 13804 9468 13872
rect 9525 13804 9536 13872
rect 9466 13796 9536 13804
rect 7654 13521 7688 13645
rect 8011 13644 9383 13691
rect 8011 13631 8077 13644
rect 8011 13597 8027 13631
rect 8061 13597 8077 13631
rect 8011 13581 8077 13597
rect 8515 13521 8549 13644
rect 7648 13509 7694 13521
rect 7648 13333 7654 13509
rect 7688 13333 7694 13509
rect 7648 13321 7694 13333
rect 7766 13509 7890 13521
rect 7766 13333 7772 13509
rect 7806 13333 7850 13509
rect 7766 13321 7850 13333
rect 7772 12954 7806 13321
rect 7844 13133 7850 13321
rect 7884 13133 7890 13509
rect 7844 13121 7890 13133
rect 7962 13509 8008 13521
rect 7962 13133 7968 13509
rect 8002 13133 8008 13509
rect 7962 13121 8008 13133
rect 8080 13509 8126 13521
rect 8080 13133 8086 13509
rect 8120 13133 8126 13509
rect 8080 13121 8126 13133
rect 8198 13509 8244 13521
rect 8198 13133 8204 13509
rect 8238 13133 8244 13509
rect 8198 13121 8244 13133
rect 8316 13509 8436 13521
rect 8316 13133 8322 13509
rect 8356 13333 8396 13509
rect 8430 13333 8436 13509
rect 8356 13321 8436 13333
rect 8508 13509 8554 13521
rect 8508 13333 8514 13509
rect 8548 13333 8554 13509
rect 8508 13321 8554 13333
rect 8356 13133 8362 13321
rect 8316 13121 8362 13133
rect 8086 13048 8120 13121
rect 8069 13032 8135 13048
rect 8069 12998 8085 13032
rect 8119 12998 8135 13032
rect 8069 12982 8135 12998
rect 8396 12954 8430 13321
rect 7772 12902 8430 12954
rect 8040 12880 8132 12902
rect 8040 12828 8054 12880
rect 8120 12828 8132 12880
rect 8040 12824 8132 12828
rect 9783 12704 9870 13954
rect 9929 13692 9964 13954
rect 9929 13645 10833 13692
rect 12492 13691 12527 14201
rect 12684 14048 12771 15234
rect 14390 15042 14400 15102
rect 14480 15042 14490 15102
rect 14390 15002 14490 15042
rect 13484 14945 15287 15002
rect 13484 14658 13521 14945
rect 14078 14858 14112 14945
rect 15253 14858 15287 14945
rect 13599 14846 13645 14858
rect 13126 14646 13172 14658
rect 13126 14470 13132 14646
rect 13166 14470 13172 14646
rect 13126 14458 13172 14470
rect 13244 14646 13290 14658
rect 13244 14470 13250 14646
rect 13284 14470 13290 14646
rect 13244 14458 13290 14470
rect 13362 14646 13408 14658
rect 13362 14470 13368 14646
rect 13402 14470 13408 14646
rect 13362 14458 13408 14470
rect 13480 14646 13526 14658
rect 13480 14470 13486 14646
rect 13520 14470 13526 14646
rect 13480 14458 13526 14470
rect 13599 14470 13605 14846
rect 13639 14470 13645 14846
rect 13599 14458 13645 14470
rect 13717 14846 13763 14858
rect 13717 14470 13723 14846
rect 13757 14470 13763 14846
rect 13717 14458 13763 14470
rect 13835 14846 13881 14858
rect 13835 14470 13841 14846
rect 13875 14470 13881 14846
rect 13835 14458 13881 14470
rect 13953 14846 13999 14858
rect 13953 14470 13959 14846
rect 13993 14470 13999 14846
rect 13953 14458 13999 14470
rect 14072 14846 14118 14858
rect 14072 14470 14078 14846
rect 14112 14470 14118 14846
rect 14072 14458 14118 14470
rect 14190 14846 14236 14858
rect 14190 14470 14196 14846
rect 14230 14470 14236 14846
rect 14190 14458 14236 14470
rect 14308 14846 14354 14858
rect 14308 14470 14314 14846
rect 14348 14470 14354 14846
rect 14308 14458 14354 14470
rect 14426 14846 14472 14858
rect 14426 14470 14432 14846
rect 14466 14470 14472 14846
rect 14426 14458 14472 14470
rect 14544 14846 14590 14858
rect 14544 14470 14550 14846
rect 14584 14470 14590 14846
rect 14544 14458 14590 14470
rect 14662 14846 14708 14858
rect 14662 14470 14668 14846
rect 14702 14470 14708 14846
rect 14662 14458 14708 14470
rect 14780 14846 14826 14858
rect 14780 14470 14786 14846
rect 14820 14470 14826 14846
rect 14780 14458 14826 14470
rect 14893 14846 14939 14858
rect 14893 14470 14899 14846
rect 14933 14470 14939 14846
rect 14893 14458 14939 14470
rect 15011 14846 15057 14858
rect 15011 14470 15017 14846
rect 15051 14470 15057 14846
rect 15011 14458 15057 14470
rect 15129 14846 15175 14858
rect 15129 14470 15135 14846
rect 15169 14470 15175 14846
rect 15129 14458 15175 14470
rect 15247 14846 15293 14858
rect 15247 14470 15253 14846
rect 15287 14658 15293 14846
rect 15287 14646 15380 14658
rect 15287 14470 15340 14646
rect 15374 14470 15380 14646
rect 15247 14458 15380 14470
rect 15452 14646 15498 14658
rect 15452 14470 15458 14646
rect 15492 14470 15498 14646
rect 15452 14458 15498 14470
rect 15570 14646 15616 14658
rect 15570 14470 15576 14646
rect 15610 14470 15616 14646
rect 15570 14458 15616 14470
rect 15688 14646 15734 14658
rect 15688 14470 15694 14646
rect 15728 14470 15734 14646
rect 15688 14458 15734 14470
rect 13131 14104 13166 14458
rect 13605 14374 13639 14458
rect 14786 14374 14820 14458
rect 13605 14332 14820 14374
rect 13605 14312 13639 14332
rect 13282 14296 13639 14312
rect 13282 14262 13298 14296
rect 13332 14262 13639 14296
rect 15694 14272 15729 14458
rect 13282 14246 13639 14262
rect 14592 14255 15729 14272
rect 14592 14221 14608 14255
rect 14642 14221 15729 14255
rect 14592 14205 15729 14221
rect 12610 14040 12771 14048
rect 12602 13972 12612 14040
rect 12669 13972 12771 14040
rect 12610 13964 12771 13972
rect 10798 13521 10832 13645
rect 11155 13644 12527 13691
rect 12990 13958 13166 14104
rect 14462 14159 14554 14169
rect 14462 14097 14472 14159
rect 14542 14097 14554 14159
rect 14462 14084 14554 14097
rect 15547 14159 15639 14172
rect 15547 14096 15556 14159
rect 15627 14096 15639 14159
rect 15547 14087 15639 14096
rect 14242 14042 14307 14045
rect 14238 14039 14307 14042
rect 14232 13979 14242 14039
rect 14301 13979 14307 14039
rect 14238 13975 14307 13979
rect 14242 13973 14307 13975
rect 11155 13631 11221 13644
rect 11155 13597 11171 13631
rect 11205 13597 11221 13631
rect 11155 13581 11221 13597
rect 11659 13521 11693 13644
rect 10792 13509 10838 13521
rect 10792 13333 10798 13509
rect 10832 13333 10838 13509
rect 10792 13321 10838 13333
rect 10910 13509 11034 13521
rect 10910 13333 10916 13509
rect 10950 13333 10994 13509
rect 10910 13321 10994 13333
rect 10916 12954 10950 13321
rect 10988 13133 10994 13321
rect 11028 13133 11034 13509
rect 10988 13121 11034 13133
rect 11106 13509 11152 13521
rect 11106 13133 11112 13509
rect 11146 13133 11152 13509
rect 11106 13121 11152 13133
rect 11224 13509 11270 13521
rect 11224 13133 11230 13509
rect 11264 13133 11270 13509
rect 11224 13121 11270 13133
rect 11342 13509 11388 13521
rect 11342 13133 11348 13509
rect 11382 13133 11388 13509
rect 11342 13121 11388 13133
rect 11460 13509 11580 13521
rect 11460 13133 11466 13509
rect 11500 13333 11540 13509
rect 11574 13333 11580 13509
rect 11500 13321 11580 13333
rect 11652 13509 11698 13521
rect 11652 13333 11658 13509
rect 11692 13333 11698 13509
rect 11652 13321 11698 13333
rect 11500 13133 11506 13321
rect 11460 13121 11506 13133
rect 11230 13048 11264 13121
rect 11213 13032 11279 13048
rect 11213 12998 11229 13032
rect 11263 12998 11279 13032
rect 11213 12982 11279 12998
rect 11540 12954 11574 13321
rect 10916 12902 11574 12954
rect 11184 12880 11276 12902
rect 11184 12828 11198 12880
rect 11264 12828 11276 12880
rect 11184 12824 11276 12828
rect 12990 12704 13062 13958
rect 13131 13696 13166 13958
rect 13131 13649 14035 13696
rect 15694 13695 15729 14205
rect 15884 14052 15971 15234
rect 17534 15042 17544 15102
rect 17624 15042 17634 15102
rect 17534 15002 17634 15042
rect 16628 14945 18431 15002
rect 16628 14658 16665 14945
rect 17222 14858 17256 14945
rect 18397 14858 18431 14945
rect 16743 14846 16789 14858
rect 16270 14646 16316 14658
rect 16270 14470 16276 14646
rect 16310 14470 16316 14646
rect 16270 14458 16316 14470
rect 16388 14646 16434 14658
rect 16388 14470 16394 14646
rect 16428 14470 16434 14646
rect 16388 14458 16434 14470
rect 16506 14646 16552 14658
rect 16506 14470 16512 14646
rect 16546 14470 16552 14646
rect 16506 14458 16552 14470
rect 16624 14646 16670 14658
rect 16624 14470 16630 14646
rect 16664 14470 16670 14646
rect 16624 14458 16670 14470
rect 16743 14470 16749 14846
rect 16783 14470 16789 14846
rect 16743 14458 16789 14470
rect 16861 14846 16907 14858
rect 16861 14470 16867 14846
rect 16901 14470 16907 14846
rect 16861 14458 16907 14470
rect 16979 14846 17025 14858
rect 16979 14470 16985 14846
rect 17019 14470 17025 14846
rect 16979 14458 17025 14470
rect 17097 14846 17143 14858
rect 17097 14470 17103 14846
rect 17137 14470 17143 14846
rect 17097 14458 17143 14470
rect 17216 14846 17262 14858
rect 17216 14470 17222 14846
rect 17256 14470 17262 14846
rect 17216 14458 17262 14470
rect 17334 14846 17380 14858
rect 17334 14470 17340 14846
rect 17374 14470 17380 14846
rect 17334 14458 17380 14470
rect 17452 14846 17498 14858
rect 17452 14470 17458 14846
rect 17492 14470 17498 14846
rect 17452 14458 17498 14470
rect 17570 14846 17616 14858
rect 17570 14470 17576 14846
rect 17610 14470 17616 14846
rect 17570 14458 17616 14470
rect 17688 14846 17734 14858
rect 17688 14470 17694 14846
rect 17728 14470 17734 14846
rect 17688 14458 17734 14470
rect 17806 14846 17852 14858
rect 17806 14470 17812 14846
rect 17846 14470 17852 14846
rect 17806 14458 17852 14470
rect 17924 14846 17970 14858
rect 17924 14470 17930 14846
rect 17964 14470 17970 14846
rect 17924 14458 17970 14470
rect 18037 14846 18083 14858
rect 18037 14470 18043 14846
rect 18077 14470 18083 14846
rect 18037 14458 18083 14470
rect 18155 14846 18201 14858
rect 18155 14470 18161 14846
rect 18195 14470 18201 14846
rect 18155 14458 18201 14470
rect 18273 14846 18319 14858
rect 18273 14470 18279 14846
rect 18313 14470 18319 14846
rect 18273 14458 18319 14470
rect 18391 14846 18437 14858
rect 18391 14470 18397 14846
rect 18431 14658 18437 14846
rect 18431 14646 18524 14658
rect 18431 14470 18484 14646
rect 18518 14470 18524 14646
rect 18391 14458 18524 14470
rect 18596 14646 18642 14658
rect 18596 14470 18602 14646
rect 18636 14470 18642 14646
rect 18596 14458 18642 14470
rect 18714 14646 18760 14658
rect 18714 14470 18720 14646
rect 18754 14470 18760 14646
rect 18714 14458 18760 14470
rect 18832 14646 18878 14658
rect 18832 14470 18838 14646
rect 18872 14470 18878 14646
rect 18832 14458 18878 14470
rect 16275 14104 16310 14458
rect 16749 14374 16783 14458
rect 17930 14374 17964 14458
rect 16749 14332 17964 14374
rect 16749 14312 16783 14332
rect 16426 14296 16783 14312
rect 16426 14262 16442 14296
rect 16476 14262 16783 14296
rect 18838 14272 18873 14458
rect 16426 14246 16783 14262
rect 17736 14255 18873 14272
rect 17736 14221 17752 14255
rect 17786 14221 18873 14255
rect 17736 14205 18873 14221
rect 15812 14044 15971 14052
rect 15804 13976 15814 14044
rect 15871 13976 15971 14044
rect 15812 13968 15971 13976
rect 14000 13525 14034 13649
rect 14357 13648 15729 13695
rect 16130 13958 16310 14104
rect 17606 14159 17698 14169
rect 17606 14097 17616 14159
rect 17686 14097 17698 14159
rect 17606 14084 17698 14097
rect 18691 14159 18783 14172
rect 18691 14096 18700 14159
rect 18771 14096 18783 14159
rect 18691 14087 18783 14096
rect 17386 14042 17451 14045
rect 17382 14039 17451 14042
rect 17376 13979 17386 14039
rect 17445 13979 17451 14039
rect 17382 13975 17451 13979
rect 17386 13973 17451 13975
rect 14357 13635 14423 13648
rect 14357 13601 14373 13635
rect 14407 13601 14423 13635
rect 14357 13585 14423 13601
rect 14861 13525 14895 13648
rect 13994 13513 14040 13525
rect 13994 13337 14000 13513
rect 14034 13337 14040 13513
rect 13994 13325 14040 13337
rect 14112 13513 14236 13525
rect 14112 13337 14118 13513
rect 14152 13337 14196 13513
rect 14112 13325 14196 13337
rect 14118 12958 14152 13325
rect 14190 13137 14196 13325
rect 14230 13137 14236 13513
rect 14190 13125 14236 13137
rect 14308 13513 14354 13525
rect 14308 13137 14314 13513
rect 14348 13137 14354 13513
rect 14308 13125 14354 13137
rect 14426 13513 14472 13525
rect 14426 13137 14432 13513
rect 14466 13137 14472 13513
rect 14426 13125 14472 13137
rect 14544 13513 14590 13525
rect 14544 13137 14550 13513
rect 14584 13137 14590 13513
rect 14544 13125 14590 13137
rect 14662 13513 14782 13525
rect 14662 13137 14668 13513
rect 14702 13337 14742 13513
rect 14776 13337 14782 13513
rect 14702 13325 14782 13337
rect 14854 13513 14900 13525
rect 14854 13337 14860 13513
rect 14894 13337 14900 13513
rect 14854 13325 14900 13337
rect 14702 13137 14708 13325
rect 14662 13125 14708 13137
rect 14432 13052 14466 13125
rect 14415 13036 14481 13052
rect 14415 13002 14431 13036
rect 14465 13002 14481 13036
rect 14415 12986 14481 13002
rect 14742 12958 14776 13325
rect 14118 12906 14776 12958
rect 14386 12884 14478 12906
rect 14386 12832 14400 12884
rect 14466 12832 14478 12884
rect 14386 12828 14478 12832
rect 3509 12636 6510 12704
rect 6638 12636 9642 12704
rect 9783 12636 12786 12704
rect 12990 12636 15988 12704
rect 16130 12701 16202 13958
rect 16275 13696 16310 13958
rect 17724 13876 17816 13884
rect 17724 13811 17736 13876
rect 17804 13811 17816 13876
rect 17724 13799 17816 13811
rect 16275 13649 17179 13696
rect 18838 13695 18873 14205
rect 19028 14052 19115 15234
rect 20666 15038 20676 15098
rect 20756 15038 20766 15098
rect 20666 14998 20766 15038
rect 19760 14941 21563 14998
rect 19760 14654 19797 14941
rect 20354 14854 20388 14941
rect 21529 14854 21563 14941
rect 19875 14842 19921 14854
rect 19402 14642 19448 14654
rect 19402 14466 19408 14642
rect 19442 14466 19448 14642
rect 19402 14454 19448 14466
rect 19520 14642 19566 14654
rect 19520 14466 19526 14642
rect 19560 14466 19566 14642
rect 19520 14454 19566 14466
rect 19638 14642 19684 14654
rect 19638 14466 19644 14642
rect 19678 14466 19684 14642
rect 19638 14454 19684 14466
rect 19756 14642 19802 14654
rect 19756 14466 19762 14642
rect 19796 14466 19802 14642
rect 19756 14454 19802 14466
rect 19875 14466 19881 14842
rect 19915 14466 19921 14842
rect 19875 14454 19921 14466
rect 19993 14842 20039 14854
rect 19993 14466 19999 14842
rect 20033 14466 20039 14842
rect 19993 14454 20039 14466
rect 20111 14842 20157 14854
rect 20111 14466 20117 14842
rect 20151 14466 20157 14842
rect 20111 14454 20157 14466
rect 20229 14842 20275 14854
rect 20229 14466 20235 14842
rect 20269 14466 20275 14842
rect 20229 14454 20275 14466
rect 20348 14842 20394 14854
rect 20348 14466 20354 14842
rect 20388 14466 20394 14842
rect 20348 14454 20394 14466
rect 20466 14842 20512 14854
rect 20466 14466 20472 14842
rect 20506 14466 20512 14842
rect 20466 14454 20512 14466
rect 20584 14842 20630 14854
rect 20584 14466 20590 14842
rect 20624 14466 20630 14842
rect 20584 14454 20630 14466
rect 20702 14842 20748 14854
rect 20702 14466 20708 14842
rect 20742 14466 20748 14842
rect 20702 14454 20748 14466
rect 20820 14842 20866 14854
rect 20820 14466 20826 14842
rect 20860 14466 20866 14842
rect 20820 14454 20866 14466
rect 20938 14842 20984 14854
rect 20938 14466 20944 14842
rect 20978 14466 20984 14842
rect 20938 14454 20984 14466
rect 21056 14842 21102 14854
rect 21056 14466 21062 14842
rect 21096 14466 21102 14842
rect 21056 14454 21102 14466
rect 21169 14842 21215 14854
rect 21169 14466 21175 14842
rect 21209 14466 21215 14842
rect 21169 14454 21215 14466
rect 21287 14842 21333 14854
rect 21287 14466 21293 14842
rect 21327 14466 21333 14842
rect 21287 14454 21333 14466
rect 21405 14842 21451 14854
rect 21405 14466 21411 14842
rect 21445 14466 21451 14842
rect 21405 14454 21451 14466
rect 21523 14842 21569 14854
rect 21523 14466 21529 14842
rect 21563 14654 21569 14842
rect 21563 14642 21656 14654
rect 21563 14466 21616 14642
rect 21650 14466 21656 14642
rect 21523 14454 21656 14466
rect 21728 14642 21774 14654
rect 21728 14466 21734 14642
rect 21768 14466 21774 14642
rect 21728 14454 21774 14466
rect 21846 14642 21892 14654
rect 21846 14466 21852 14642
rect 21886 14466 21892 14642
rect 21846 14454 21892 14466
rect 21964 14642 22010 14654
rect 21964 14466 21970 14642
rect 22004 14466 22010 14642
rect 21964 14454 22010 14466
rect 19407 14100 19442 14454
rect 19881 14370 19915 14454
rect 21062 14370 21096 14454
rect 19881 14328 21096 14370
rect 19881 14308 19915 14328
rect 19558 14292 19915 14308
rect 19558 14258 19574 14292
rect 19608 14258 19915 14292
rect 21970 14268 22005 14454
rect 19558 14242 19915 14258
rect 20868 14251 22005 14268
rect 20868 14217 20884 14251
rect 20918 14217 22005 14251
rect 20868 14201 22005 14217
rect 18956 14044 19115 14052
rect 18948 13976 18958 14044
rect 19015 13976 19115 14044
rect 18956 13968 19115 13976
rect 19261 13954 19442 14100
rect 20738 14155 20830 14165
rect 20738 14093 20748 14155
rect 20818 14093 20830 14155
rect 20738 14080 20830 14093
rect 21823 14155 21915 14168
rect 21823 14092 21832 14155
rect 21903 14092 21915 14155
rect 21823 14083 21915 14092
rect 20518 14038 20583 14041
rect 20514 14035 20583 14038
rect 20508 13975 20518 14035
rect 20577 13975 20583 14035
rect 20514 13971 20583 13975
rect 20518 13969 20583 13971
rect 18956 13876 19028 13884
rect 18948 13808 18958 13876
rect 19015 13808 19028 13876
rect 18956 13800 19028 13808
rect 17144 13525 17178 13649
rect 17501 13648 18873 13695
rect 17501 13635 17567 13648
rect 17501 13601 17517 13635
rect 17551 13601 17567 13635
rect 17501 13585 17567 13601
rect 18005 13525 18039 13648
rect 17138 13513 17184 13525
rect 17138 13337 17144 13513
rect 17178 13337 17184 13513
rect 17138 13325 17184 13337
rect 17256 13513 17380 13525
rect 17256 13337 17262 13513
rect 17296 13337 17340 13513
rect 17256 13325 17340 13337
rect 17262 12958 17296 13325
rect 17334 13137 17340 13325
rect 17374 13137 17380 13513
rect 17334 13125 17380 13137
rect 17452 13513 17498 13525
rect 17452 13137 17458 13513
rect 17492 13137 17498 13513
rect 17452 13125 17498 13137
rect 17570 13513 17616 13525
rect 17570 13137 17576 13513
rect 17610 13137 17616 13513
rect 17570 13125 17616 13137
rect 17688 13513 17734 13525
rect 17688 13137 17694 13513
rect 17728 13137 17734 13513
rect 17688 13125 17734 13137
rect 17806 13513 17926 13525
rect 17806 13137 17812 13513
rect 17846 13337 17886 13513
rect 17920 13337 17926 13513
rect 17846 13325 17926 13337
rect 17998 13513 18044 13525
rect 17998 13337 18004 13513
rect 18038 13337 18044 13513
rect 17998 13325 18044 13337
rect 17846 13137 17852 13325
rect 17806 13125 17852 13137
rect 17576 13052 17610 13125
rect 17559 13036 17625 13052
rect 17559 13002 17575 13036
rect 17609 13002 17625 13036
rect 17559 12986 17625 13002
rect 17886 12958 17920 13325
rect 17262 12906 17920 12958
rect 17530 12884 17622 12906
rect 17530 12832 17544 12884
rect 17610 12832 17622 12884
rect 17530 12828 17622 12832
rect 19263 12701 19335 13954
rect 19407 13692 19442 13954
rect 20856 13872 20948 13880
rect 20856 13807 20868 13872
rect 20936 13807 20948 13872
rect 20856 13795 20948 13807
rect 19407 13645 20311 13692
rect 21970 13691 22005 14201
rect 22177 14048 22264 15245
rect 24112 15244 24248 15245
rect 23810 15038 23820 15098
rect 23900 15038 23910 15098
rect 23810 14998 23910 15038
rect 22904 14941 24707 14998
rect 22904 14654 22941 14941
rect 23498 14854 23532 14941
rect 24673 14854 24707 14941
rect 23019 14842 23065 14854
rect 22546 14642 22592 14654
rect 22546 14466 22552 14642
rect 22586 14466 22592 14642
rect 22546 14454 22592 14466
rect 22664 14642 22710 14654
rect 22664 14466 22670 14642
rect 22704 14466 22710 14642
rect 22664 14454 22710 14466
rect 22782 14642 22828 14654
rect 22782 14466 22788 14642
rect 22822 14466 22828 14642
rect 22782 14454 22828 14466
rect 22900 14642 22946 14654
rect 22900 14466 22906 14642
rect 22940 14466 22946 14642
rect 22900 14454 22946 14466
rect 23019 14466 23025 14842
rect 23059 14466 23065 14842
rect 23019 14454 23065 14466
rect 23137 14842 23183 14854
rect 23137 14466 23143 14842
rect 23177 14466 23183 14842
rect 23137 14454 23183 14466
rect 23255 14842 23301 14854
rect 23255 14466 23261 14842
rect 23295 14466 23301 14842
rect 23255 14454 23301 14466
rect 23373 14842 23419 14854
rect 23373 14466 23379 14842
rect 23413 14466 23419 14842
rect 23373 14454 23419 14466
rect 23492 14842 23538 14854
rect 23492 14466 23498 14842
rect 23532 14466 23538 14842
rect 23492 14454 23538 14466
rect 23610 14842 23656 14854
rect 23610 14466 23616 14842
rect 23650 14466 23656 14842
rect 23610 14454 23656 14466
rect 23728 14842 23774 14854
rect 23728 14466 23734 14842
rect 23768 14466 23774 14842
rect 23728 14454 23774 14466
rect 23846 14842 23892 14854
rect 23846 14466 23852 14842
rect 23886 14466 23892 14842
rect 23846 14454 23892 14466
rect 23964 14842 24010 14854
rect 23964 14466 23970 14842
rect 24004 14466 24010 14842
rect 23964 14454 24010 14466
rect 24082 14842 24128 14854
rect 24082 14466 24088 14842
rect 24122 14466 24128 14842
rect 24082 14454 24128 14466
rect 24200 14842 24246 14854
rect 24200 14466 24206 14842
rect 24240 14466 24246 14842
rect 24200 14454 24246 14466
rect 24313 14842 24359 14854
rect 24313 14466 24319 14842
rect 24353 14466 24359 14842
rect 24313 14454 24359 14466
rect 24431 14842 24477 14854
rect 24431 14466 24437 14842
rect 24471 14466 24477 14842
rect 24431 14454 24477 14466
rect 24549 14842 24595 14854
rect 24549 14466 24555 14842
rect 24589 14466 24595 14842
rect 24549 14454 24595 14466
rect 24667 14842 24713 14854
rect 24667 14466 24673 14842
rect 24707 14654 24713 14842
rect 24707 14642 24800 14654
rect 24707 14466 24760 14642
rect 24794 14466 24800 14642
rect 24667 14454 24800 14466
rect 24872 14642 24918 14654
rect 24872 14466 24878 14642
rect 24912 14466 24918 14642
rect 24872 14454 24918 14466
rect 24990 14642 25036 14654
rect 24990 14466 24996 14642
rect 25030 14466 25036 14642
rect 24990 14454 25036 14466
rect 25108 14642 25154 14654
rect 25108 14466 25114 14642
rect 25148 14466 25154 14642
rect 25108 14454 25154 14466
rect 22551 14100 22586 14454
rect 23025 14370 23059 14454
rect 24206 14370 24240 14454
rect 23025 14328 24240 14370
rect 23025 14308 23059 14328
rect 22702 14292 23059 14308
rect 22702 14258 22718 14292
rect 22752 14258 23059 14292
rect 25114 14268 25149 14454
rect 22702 14242 23059 14258
rect 24012 14251 25149 14268
rect 24012 14217 24028 14251
rect 24062 14217 25149 14251
rect 24012 14201 25149 14217
rect 22088 14040 22264 14048
rect 22080 13972 22090 14040
rect 22147 13972 22264 14040
rect 22088 13964 22264 13972
rect 22405 13954 22586 14100
rect 23882 14155 23974 14165
rect 23882 14093 23892 14155
rect 23962 14093 23974 14155
rect 23882 14080 23974 14093
rect 24967 14155 25059 14168
rect 24967 14092 24976 14155
rect 25047 14092 25059 14155
rect 24967 14083 25059 14092
rect 23662 14038 23727 14041
rect 23658 14035 23727 14038
rect 23652 13975 23662 14035
rect 23721 13975 23727 14035
rect 23658 13971 23727 13975
rect 23662 13969 23727 13971
rect 22088 13872 22158 13880
rect 22080 13804 22090 13872
rect 22147 13804 22158 13872
rect 22088 13796 22158 13804
rect 20276 13521 20310 13645
rect 20633 13644 22005 13691
rect 20633 13631 20699 13644
rect 20633 13597 20649 13631
rect 20683 13597 20699 13631
rect 20633 13581 20699 13597
rect 21137 13521 21171 13644
rect 20270 13509 20316 13521
rect 20270 13333 20276 13509
rect 20310 13333 20316 13509
rect 20270 13321 20316 13333
rect 20388 13509 20512 13521
rect 20388 13333 20394 13509
rect 20428 13333 20472 13509
rect 20388 13321 20472 13333
rect 20394 12954 20428 13321
rect 20466 13133 20472 13321
rect 20506 13133 20512 13509
rect 20466 13121 20512 13133
rect 20584 13509 20630 13521
rect 20584 13133 20590 13509
rect 20624 13133 20630 13509
rect 20584 13121 20630 13133
rect 20702 13509 20748 13521
rect 20702 13133 20708 13509
rect 20742 13133 20748 13509
rect 20702 13121 20748 13133
rect 20820 13509 20866 13521
rect 20820 13133 20826 13509
rect 20860 13133 20866 13509
rect 20820 13121 20866 13133
rect 20938 13509 21058 13521
rect 20938 13133 20944 13509
rect 20978 13333 21018 13509
rect 21052 13333 21058 13509
rect 20978 13321 21058 13333
rect 21130 13509 21176 13521
rect 21130 13333 21136 13509
rect 21170 13333 21176 13509
rect 21130 13321 21176 13333
rect 20978 13133 20984 13321
rect 20938 13121 20984 13133
rect 20708 13048 20742 13121
rect 20691 13032 20757 13048
rect 20691 12998 20707 13032
rect 20741 12998 20757 13032
rect 20691 12982 20757 12998
rect 21018 12954 21052 13321
rect 20394 12902 21052 12954
rect 20662 12880 20754 12902
rect 20662 12828 20676 12880
rect 20742 12828 20754 12880
rect 20662 12824 20754 12828
rect 16130 12636 19132 12701
rect 19263 12636 22264 12701
rect 22406 12700 22478 13954
rect 22551 13692 22586 13954
rect 24000 13872 24092 13880
rect 24000 13807 24012 13872
rect 24080 13807 24092 13872
rect 24000 13795 24092 13807
rect 22551 13645 23455 13692
rect 25114 13691 25149 14201
rect 25322 14048 25409 15245
rect 25817 14158 25927 14165
rect 25817 14080 25828 14158
rect 25232 14040 25409 14048
rect 25224 13972 25234 14040
rect 25291 13972 25409 14040
rect 25232 13964 25409 13972
rect 25818 14070 25828 14080
rect 25911 14070 25927 14158
rect 25232 13872 25305 13880
rect 25224 13804 25234 13872
rect 25291 13804 25305 13872
rect 25232 13796 25305 13804
rect 23420 13521 23454 13645
rect 23777 13644 25149 13691
rect 23777 13631 23843 13644
rect 23777 13597 23793 13631
rect 23827 13597 23843 13631
rect 23777 13581 23843 13597
rect 24281 13521 24315 13644
rect 23414 13509 23460 13521
rect 23414 13333 23420 13509
rect 23454 13333 23460 13509
rect 23414 13321 23460 13333
rect 23532 13509 23656 13521
rect 23532 13333 23538 13509
rect 23572 13333 23616 13509
rect 23532 13321 23616 13333
rect 23538 12954 23572 13321
rect 23610 13133 23616 13321
rect 23650 13133 23656 13509
rect 23610 13121 23656 13133
rect 23728 13509 23774 13521
rect 23728 13133 23734 13509
rect 23768 13133 23774 13509
rect 23728 13121 23774 13133
rect 23846 13509 23892 13521
rect 23846 13133 23852 13509
rect 23886 13133 23892 13509
rect 23846 13121 23892 13133
rect 23964 13509 24010 13521
rect 23964 13133 23970 13509
rect 24004 13133 24010 13509
rect 23964 13121 24010 13133
rect 24082 13509 24202 13521
rect 24082 13133 24088 13509
rect 24122 13333 24162 13509
rect 24196 13333 24202 13509
rect 24122 13321 24202 13333
rect 24274 13509 24320 13521
rect 24274 13333 24280 13509
rect 24314 13333 24320 13509
rect 24274 13321 24320 13333
rect 24122 13133 24128 13321
rect 24082 13121 24128 13133
rect 23852 13048 23886 13121
rect 23835 13032 23901 13048
rect 23835 12998 23851 13032
rect 23885 12998 23901 13032
rect 23835 12982 23901 12998
rect 24162 12954 24196 13321
rect 23538 12902 24196 12954
rect 23806 12880 23898 12902
rect 23806 12828 23820 12880
rect 23886 12828 23898 12880
rect 23806 12824 23898 12828
rect 22406 12636 25408 12700
rect 4912 12308 4922 12368
rect 5002 12308 5012 12368
rect 4912 12268 5012 12308
rect 4006 12211 5809 12268
rect 4006 11924 4043 12211
rect 4600 12124 4634 12211
rect 5775 12124 5809 12211
rect 4121 12112 4167 12124
rect 3648 11912 3694 11924
rect 3648 11736 3654 11912
rect 3688 11736 3694 11912
rect 3648 11724 3694 11736
rect 3766 11912 3812 11924
rect 3766 11736 3772 11912
rect 3806 11736 3812 11912
rect 3766 11724 3812 11736
rect 3884 11912 3930 11924
rect 3884 11736 3890 11912
rect 3924 11736 3930 11912
rect 3884 11724 3930 11736
rect 4002 11912 4048 11924
rect 4002 11736 4008 11912
rect 4042 11736 4048 11912
rect 4002 11724 4048 11736
rect 4121 11736 4127 12112
rect 4161 11736 4167 12112
rect 4121 11724 4167 11736
rect 4239 12112 4285 12124
rect 4239 11736 4245 12112
rect 4279 11736 4285 12112
rect 4239 11724 4285 11736
rect 4357 12112 4403 12124
rect 4357 11736 4363 12112
rect 4397 11736 4403 12112
rect 4357 11724 4403 11736
rect 4475 12112 4521 12124
rect 4475 11736 4481 12112
rect 4515 11736 4521 12112
rect 4475 11724 4521 11736
rect 4594 12112 4640 12124
rect 4594 11736 4600 12112
rect 4634 11736 4640 12112
rect 4594 11724 4640 11736
rect 4712 12112 4758 12124
rect 4712 11736 4718 12112
rect 4752 11736 4758 12112
rect 4712 11724 4758 11736
rect 4830 12112 4876 12124
rect 4830 11736 4836 12112
rect 4870 11736 4876 12112
rect 4830 11724 4876 11736
rect 4948 12112 4994 12124
rect 4948 11736 4954 12112
rect 4988 11736 4994 12112
rect 4948 11724 4994 11736
rect 5066 12112 5112 12124
rect 5066 11736 5072 12112
rect 5106 11736 5112 12112
rect 5066 11724 5112 11736
rect 5184 12112 5230 12124
rect 5184 11736 5190 12112
rect 5224 11736 5230 12112
rect 5184 11724 5230 11736
rect 5302 12112 5348 12124
rect 5302 11736 5308 12112
rect 5342 11736 5348 12112
rect 5302 11724 5348 11736
rect 5415 12112 5461 12124
rect 5415 11736 5421 12112
rect 5455 11736 5461 12112
rect 5415 11724 5461 11736
rect 5533 12112 5579 12124
rect 5533 11736 5539 12112
rect 5573 11736 5579 12112
rect 5533 11724 5579 11736
rect 5651 12112 5697 12124
rect 5651 11736 5657 12112
rect 5691 11736 5697 12112
rect 5651 11724 5697 11736
rect 5769 12112 5815 12124
rect 5769 11736 5775 12112
rect 5809 11924 5815 12112
rect 5809 11912 5902 11924
rect 5809 11736 5862 11912
rect 5896 11736 5902 11912
rect 5769 11724 5902 11736
rect 5974 11912 6020 11924
rect 5974 11736 5980 11912
rect 6014 11736 6020 11912
rect 5974 11724 6020 11736
rect 6092 11912 6138 11924
rect 6092 11736 6098 11912
rect 6132 11736 6138 11912
rect 6092 11724 6138 11736
rect 6210 11912 6256 11924
rect 6210 11736 6216 11912
rect 6250 11736 6256 11912
rect 6210 11724 6256 11736
rect 3653 11370 3688 11724
rect 4127 11640 4161 11724
rect 5308 11640 5342 11724
rect 4127 11598 5342 11640
rect 4127 11578 4161 11598
rect 3804 11562 4161 11578
rect 3804 11528 3820 11562
rect 3854 11528 4161 11562
rect 6216 11538 6251 11724
rect 3804 11512 4161 11528
rect 5114 11521 6251 11538
rect 5114 11487 5130 11521
rect 5164 11487 6251 11521
rect 5114 11471 6251 11487
rect 3190 11310 3366 11318
rect 3182 11242 3192 11310
rect 3249 11242 3366 11310
rect 3190 11234 3366 11242
rect 3507 11224 3688 11370
rect 4984 11425 5076 11435
rect 4984 11363 4994 11425
rect 5064 11363 5076 11425
rect 4984 11350 5076 11363
rect 6069 11425 6161 11438
rect 6069 11362 6078 11425
rect 6149 11362 6161 11425
rect 6069 11353 6161 11362
rect 4764 11308 4829 11311
rect 4760 11305 4829 11308
rect 4754 11245 4764 11305
rect 4823 11245 4829 11305
rect 4760 11241 4829 11245
rect 4764 11239 4829 11241
rect 3190 11142 3318 11150
rect 3182 11074 3192 11142
rect 3249 11074 3318 11142
rect 3190 11066 3318 11074
rect -570 10860 173 10867
rect 64 10859 168 10860
rect 1378 10791 1412 10915
rect 1735 10914 3107 10961
rect 1735 10901 1801 10914
rect 1735 10867 1751 10901
rect 1785 10867 1801 10901
rect 1735 10851 1801 10867
rect 2239 10791 2273 10914
rect 1372 10779 1418 10791
rect -808 10758 132 10760
rect -808 10745 213 10758
rect -808 10744 141 10745
rect -808 10687 -783 10744
rect -661 10687 141 10744
rect -808 10682 141 10687
rect 202 10682 213 10745
rect -808 10673 213 10682
rect 64 10672 213 10673
rect 1372 10603 1378 10779
rect 1412 10603 1418 10779
rect 1372 10591 1418 10603
rect 1490 10779 1614 10791
rect 1490 10603 1496 10779
rect 1530 10603 1574 10779
rect 1490 10591 1574 10603
rect -1068 10525 215 10542
rect -1068 10516 141 10525
rect -1068 10459 -1048 10516
rect -926 10459 141 10516
rect 203 10459 215 10525
rect -1068 10447 215 10459
rect -1068 10443 132 10447
rect -1275 10346 110 10347
rect -1275 10331 213 10346
rect -1275 10274 -1255 10331
rect -1133 10329 213 10331
rect -1133 10274 140 10329
rect -1275 10271 140 10274
rect 203 10271 213 10329
rect -1275 10260 213 10271
rect -1275 10255 110 10260
rect 1496 10224 1530 10591
rect 1568 10403 1574 10591
rect 1608 10403 1614 10779
rect 1568 10391 1614 10403
rect 1686 10779 1732 10791
rect 1686 10403 1692 10779
rect 1726 10403 1732 10779
rect 1686 10391 1732 10403
rect 1804 10779 1850 10791
rect 1804 10403 1810 10779
rect 1844 10403 1850 10779
rect 1804 10391 1850 10403
rect 1922 10779 1968 10791
rect 1922 10403 1928 10779
rect 1962 10403 1968 10779
rect 1922 10391 1968 10403
rect 2040 10779 2160 10791
rect 2040 10403 2046 10779
rect 2080 10603 2120 10779
rect 2154 10603 2160 10779
rect 2080 10591 2160 10603
rect 2232 10779 2278 10791
rect 2232 10603 2238 10779
rect 2272 10603 2278 10779
rect 2232 10591 2278 10603
rect 2080 10403 2086 10591
rect 2040 10391 2086 10403
rect 1810 10318 1844 10391
rect 1793 10302 1859 10318
rect 1793 10268 1809 10302
rect 1843 10268 1859 10302
rect 1793 10252 1859 10268
rect 2120 10224 2154 10591
rect 1496 10172 2154 10224
rect 1764 10150 1856 10172
rect 1764 10098 1778 10150
rect 1844 10098 1856 10150
rect 1764 10094 1856 10098
rect -1531 9986 215 10004
rect -1531 9984 140 9986
rect -1531 9927 -1515 9984
rect -1393 9927 140 9984
rect -1531 9925 140 9927
rect 204 9925 215 9986
rect -1531 9914 215 9925
rect -1531 9912 116 9914
rect 3267 9875 3318 11066
rect 3507 10930 3603 11224
rect 3507 10859 3520 10930
rect 3591 10859 3603 10930
rect 3653 10962 3688 11224
rect 5102 11142 5194 11150
rect 5102 11077 5114 11142
rect 5182 11077 5194 11142
rect 5102 11065 5194 11077
rect 3653 10915 4557 10962
rect 6216 10961 6251 11471
rect 6439 11318 6510 12636
rect 8044 12304 8054 12364
rect 8134 12304 8144 12364
rect 8044 12264 8144 12304
rect 7138 12207 8941 12264
rect 7138 11920 7175 12207
rect 7732 12120 7766 12207
rect 8907 12120 8941 12207
rect 7253 12108 7299 12120
rect 6780 11908 6826 11920
rect 6780 11732 6786 11908
rect 6820 11732 6826 11908
rect 6780 11720 6826 11732
rect 6898 11908 6944 11920
rect 6898 11732 6904 11908
rect 6938 11732 6944 11908
rect 6898 11720 6944 11732
rect 7016 11908 7062 11920
rect 7016 11732 7022 11908
rect 7056 11732 7062 11908
rect 7016 11720 7062 11732
rect 7134 11908 7180 11920
rect 7134 11732 7140 11908
rect 7174 11732 7180 11908
rect 7134 11720 7180 11732
rect 7253 11732 7259 12108
rect 7293 11732 7299 12108
rect 7253 11720 7299 11732
rect 7371 12108 7417 12120
rect 7371 11732 7377 12108
rect 7411 11732 7417 12108
rect 7371 11720 7417 11732
rect 7489 12108 7535 12120
rect 7489 11732 7495 12108
rect 7529 11732 7535 12108
rect 7489 11720 7535 11732
rect 7607 12108 7653 12120
rect 7607 11732 7613 12108
rect 7647 11732 7653 12108
rect 7607 11720 7653 11732
rect 7726 12108 7772 12120
rect 7726 11732 7732 12108
rect 7766 11732 7772 12108
rect 7726 11720 7772 11732
rect 7844 12108 7890 12120
rect 7844 11732 7850 12108
rect 7884 11732 7890 12108
rect 7844 11720 7890 11732
rect 7962 12108 8008 12120
rect 7962 11732 7968 12108
rect 8002 11732 8008 12108
rect 7962 11720 8008 11732
rect 8080 12108 8126 12120
rect 8080 11732 8086 12108
rect 8120 11732 8126 12108
rect 8080 11720 8126 11732
rect 8198 12108 8244 12120
rect 8198 11732 8204 12108
rect 8238 11732 8244 12108
rect 8198 11720 8244 11732
rect 8316 12108 8362 12120
rect 8316 11732 8322 12108
rect 8356 11732 8362 12108
rect 8316 11720 8362 11732
rect 8434 12108 8480 12120
rect 8434 11732 8440 12108
rect 8474 11732 8480 12108
rect 8434 11720 8480 11732
rect 8547 12108 8593 12120
rect 8547 11732 8553 12108
rect 8587 11732 8593 12108
rect 8547 11720 8593 11732
rect 8665 12108 8711 12120
rect 8665 11732 8671 12108
rect 8705 11732 8711 12108
rect 8665 11720 8711 11732
rect 8783 12108 8829 12120
rect 8783 11732 8789 12108
rect 8823 11732 8829 12108
rect 8783 11720 8829 11732
rect 8901 12108 8947 12120
rect 8901 11732 8907 12108
rect 8941 11920 8947 12108
rect 8941 11908 9034 11920
rect 8941 11732 8994 11908
rect 9028 11732 9034 11908
rect 8901 11720 9034 11732
rect 9106 11908 9152 11920
rect 9106 11732 9112 11908
rect 9146 11732 9152 11908
rect 9106 11720 9152 11732
rect 9224 11908 9270 11920
rect 9224 11732 9230 11908
rect 9264 11732 9270 11908
rect 9224 11720 9270 11732
rect 9342 11908 9388 11920
rect 9342 11732 9348 11908
rect 9382 11732 9388 11908
rect 9342 11720 9388 11732
rect 6785 11366 6820 11720
rect 7259 11636 7293 11720
rect 8440 11636 8474 11720
rect 7259 11594 8474 11636
rect 7259 11574 7293 11594
rect 6936 11558 7293 11574
rect 6936 11524 6952 11558
rect 6986 11524 7293 11558
rect 9348 11534 9383 11720
rect 6936 11508 7293 11524
rect 8246 11517 9383 11534
rect 8246 11483 8262 11517
rect 8296 11483 9383 11517
rect 8246 11467 9383 11483
rect 6334 11310 6510 11318
rect 6326 11242 6336 11310
rect 6393 11242 6510 11310
rect 6334 11234 6510 11242
rect 6639 11220 6820 11366
rect 8116 11421 8208 11431
rect 8116 11359 8126 11421
rect 8196 11359 8208 11421
rect 8116 11346 8208 11359
rect 9201 11421 9293 11434
rect 9201 11358 9210 11421
rect 9281 11358 9293 11421
rect 9201 11349 9293 11358
rect 7896 11304 7961 11307
rect 7892 11301 7961 11304
rect 7886 11241 7896 11301
rect 7955 11241 7961 11301
rect 7892 11237 7961 11241
rect 7896 11235 7961 11237
rect 6334 11142 6502 11150
rect 6326 11074 6336 11142
rect 6393 11074 6502 11142
rect 6334 11066 6502 11074
rect 3507 10849 3603 10859
rect 4522 10791 4556 10915
rect 4879 10914 6251 10961
rect 4879 10901 4945 10914
rect 4879 10867 4895 10901
rect 4929 10867 4945 10901
rect 4879 10851 4945 10867
rect 5383 10791 5417 10914
rect 4516 10779 4562 10791
rect 4516 10603 4522 10779
rect 4556 10603 4562 10779
rect 4516 10591 4562 10603
rect 4634 10779 4758 10791
rect 4634 10603 4640 10779
rect 4674 10603 4718 10779
rect 4634 10591 4718 10603
rect 4640 10224 4674 10591
rect 4712 10403 4718 10591
rect 4752 10403 4758 10779
rect 4712 10391 4758 10403
rect 4830 10779 4876 10791
rect 4830 10403 4836 10779
rect 4870 10403 4876 10779
rect 4830 10391 4876 10403
rect 4948 10779 4994 10791
rect 4948 10403 4954 10779
rect 4988 10403 4994 10779
rect 4948 10391 4994 10403
rect 5066 10779 5112 10791
rect 5066 10403 5072 10779
rect 5106 10403 5112 10779
rect 5066 10391 5112 10403
rect 5184 10779 5304 10791
rect 5184 10403 5190 10779
rect 5224 10603 5264 10779
rect 5298 10603 5304 10779
rect 5224 10591 5304 10603
rect 5376 10779 5422 10791
rect 5376 10603 5382 10779
rect 5416 10603 5422 10779
rect 5376 10591 5422 10603
rect 5224 10403 5230 10591
rect 5184 10391 5230 10403
rect 4954 10318 4988 10391
rect 4937 10302 5003 10318
rect 4937 10268 4953 10302
rect 4987 10268 5003 10302
rect 4937 10252 5003 10268
rect 5264 10224 5298 10591
rect 4640 10172 5298 10224
rect 4908 10150 5000 10172
rect 4908 10098 4922 10150
rect 4988 10098 5000 10150
rect 4908 10094 5000 10098
rect 6422 9875 6502 11066
rect 6639 10771 6729 11220
rect 6785 10958 6820 11220
rect 8234 11138 8326 11146
rect 8234 11073 8246 11138
rect 8314 11073 8326 11138
rect 8234 11061 8326 11073
rect 6785 10911 7689 10958
rect 9348 10957 9383 11467
rect 9466 11422 9532 11430
rect 9458 11354 9468 11422
rect 9525 11354 9532 11422
rect 9466 11346 9532 11354
rect 9571 11314 9642 12636
rect 11188 12304 11198 12364
rect 11278 12304 11288 12364
rect 11188 12264 11288 12304
rect 10282 12207 12085 12264
rect 10282 11920 10319 12207
rect 10876 12120 10910 12207
rect 12051 12120 12085 12207
rect 10397 12108 10443 12120
rect 9924 11908 9970 11920
rect 9924 11732 9930 11908
rect 9964 11732 9970 11908
rect 9924 11720 9970 11732
rect 10042 11908 10088 11920
rect 10042 11732 10048 11908
rect 10082 11732 10088 11908
rect 10042 11720 10088 11732
rect 10160 11908 10206 11920
rect 10160 11732 10166 11908
rect 10200 11732 10206 11908
rect 10160 11720 10206 11732
rect 10278 11908 10324 11920
rect 10278 11732 10284 11908
rect 10318 11732 10324 11908
rect 10278 11720 10324 11732
rect 10397 11732 10403 12108
rect 10437 11732 10443 12108
rect 10397 11720 10443 11732
rect 10515 12108 10561 12120
rect 10515 11732 10521 12108
rect 10555 11732 10561 12108
rect 10515 11720 10561 11732
rect 10633 12108 10679 12120
rect 10633 11732 10639 12108
rect 10673 11732 10679 12108
rect 10633 11720 10679 11732
rect 10751 12108 10797 12120
rect 10751 11732 10757 12108
rect 10791 11732 10797 12108
rect 10751 11720 10797 11732
rect 10870 12108 10916 12120
rect 10870 11732 10876 12108
rect 10910 11732 10916 12108
rect 10870 11720 10916 11732
rect 10988 12108 11034 12120
rect 10988 11732 10994 12108
rect 11028 11732 11034 12108
rect 10988 11720 11034 11732
rect 11106 12108 11152 12120
rect 11106 11732 11112 12108
rect 11146 11732 11152 12108
rect 11106 11720 11152 11732
rect 11224 12108 11270 12120
rect 11224 11732 11230 12108
rect 11264 11732 11270 12108
rect 11224 11720 11270 11732
rect 11342 12108 11388 12120
rect 11342 11732 11348 12108
rect 11382 11732 11388 12108
rect 11342 11720 11388 11732
rect 11460 12108 11506 12120
rect 11460 11732 11466 12108
rect 11500 11732 11506 12108
rect 11460 11720 11506 11732
rect 11578 12108 11624 12120
rect 11578 11732 11584 12108
rect 11618 11732 11624 12108
rect 11578 11720 11624 11732
rect 11691 12108 11737 12120
rect 11691 11732 11697 12108
rect 11731 11732 11737 12108
rect 11691 11720 11737 11732
rect 11809 12108 11855 12120
rect 11809 11732 11815 12108
rect 11849 11732 11855 12108
rect 11809 11720 11855 11732
rect 11927 12108 11973 12120
rect 11927 11732 11933 12108
rect 11967 11732 11973 12108
rect 11927 11720 11973 11732
rect 12045 12108 12091 12120
rect 12045 11732 12051 12108
rect 12085 11920 12091 12108
rect 12085 11908 12178 11920
rect 12085 11732 12138 11908
rect 12172 11732 12178 11908
rect 12045 11720 12178 11732
rect 12250 11908 12296 11920
rect 12250 11732 12256 11908
rect 12290 11732 12296 11908
rect 12250 11720 12296 11732
rect 12368 11908 12414 11920
rect 12368 11732 12374 11908
rect 12408 11732 12414 11908
rect 12368 11720 12414 11732
rect 12486 11908 12532 11920
rect 12486 11732 12492 11908
rect 12526 11732 12532 11908
rect 12486 11720 12532 11732
rect 9929 11366 9964 11720
rect 10403 11636 10437 11720
rect 11584 11636 11618 11720
rect 10403 11594 11618 11636
rect 10403 11574 10437 11594
rect 10080 11558 10437 11574
rect 10080 11524 10096 11558
rect 10130 11524 10437 11558
rect 12492 11534 12527 11720
rect 10080 11508 10437 11524
rect 11390 11517 12527 11534
rect 11390 11483 11406 11517
rect 11440 11483 12527 11517
rect 11390 11467 12527 11483
rect 9466 11306 9642 11314
rect 9458 11238 9468 11306
rect 9525 11238 9642 11306
rect 9783 11269 9964 11366
rect 11260 11421 11352 11431
rect 11260 11359 11270 11421
rect 11340 11359 11352 11421
rect 11260 11346 11352 11359
rect 12345 11421 12437 11434
rect 12345 11358 12354 11421
rect 12425 11358 12437 11421
rect 12345 11349 12437 11358
rect 11040 11304 11105 11307
rect 11036 11301 11105 11304
rect 9466 11230 9642 11238
rect 9781 11220 9964 11269
rect 11030 11241 11040 11301
rect 11099 11241 11105 11301
rect 11036 11237 11105 11241
rect 11040 11235 11105 11237
rect 9466 11138 9618 11146
rect 9458 11070 9468 11138
rect 9525 11070 9618 11138
rect 9466 11062 9618 11070
rect 7654 10787 7688 10911
rect 8011 10910 9383 10957
rect 8011 10897 8077 10910
rect 8011 10863 8027 10897
rect 8061 10863 8077 10897
rect 8011 10847 8077 10863
rect 8515 10787 8549 10910
rect 7648 10775 7694 10787
rect 6639 10678 6650 10771
rect 6720 10678 6730 10771
rect 6639 10670 6729 10678
rect 7648 10599 7654 10775
rect 7688 10599 7694 10775
rect 7648 10587 7694 10599
rect 7766 10775 7890 10787
rect 7766 10599 7772 10775
rect 7806 10599 7850 10775
rect 7766 10587 7850 10599
rect 7772 10220 7806 10587
rect 7844 10399 7850 10587
rect 7884 10399 7890 10775
rect 7844 10387 7890 10399
rect 7962 10775 8008 10787
rect 7962 10399 7968 10775
rect 8002 10399 8008 10775
rect 7962 10387 8008 10399
rect 8080 10775 8126 10787
rect 8080 10399 8086 10775
rect 8120 10399 8126 10775
rect 8080 10387 8126 10399
rect 8198 10775 8244 10787
rect 8198 10399 8204 10775
rect 8238 10399 8244 10775
rect 8198 10387 8244 10399
rect 8316 10775 8436 10787
rect 8316 10399 8322 10775
rect 8356 10599 8396 10775
rect 8430 10599 8436 10775
rect 8356 10587 8436 10599
rect 8508 10775 8554 10787
rect 8508 10599 8514 10775
rect 8548 10599 8554 10775
rect 8508 10587 8554 10599
rect 8356 10399 8362 10587
rect 8316 10387 8362 10399
rect 8086 10314 8120 10387
rect 8069 10298 8135 10314
rect 8069 10264 8085 10298
rect 8119 10264 8135 10298
rect 8069 10248 8135 10264
rect 8396 10220 8430 10587
rect 7772 10168 8430 10220
rect 8040 10146 8132 10168
rect 8040 10094 8054 10146
rect 8120 10094 8132 10146
rect 8040 10090 8132 10094
rect 9561 9876 9618 11062
rect 9781 10540 9879 11220
rect 9929 10958 9964 11220
rect 11378 11138 11470 11146
rect 11378 11073 11390 11138
rect 11458 11073 11470 11138
rect 11378 11061 11470 11073
rect 9929 10911 10833 10958
rect 12492 10957 12527 11467
rect 12715 11314 12786 12636
rect 14390 12308 14400 12368
rect 14480 12308 14490 12368
rect 14390 12268 14490 12308
rect 13484 12211 15287 12268
rect 13484 11924 13521 12211
rect 14078 12124 14112 12211
rect 15253 12124 15287 12211
rect 13599 12112 13645 12124
rect 13126 11912 13172 11924
rect 13126 11736 13132 11912
rect 13166 11736 13172 11912
rect 13126 11724 13172 11736
rect 13244 11912 13290 11924
rect 13244 11736 13250 11912
rect 13284 11736 13290 11912
rect 13244 11724 13290 11736
rect 13362 11912 13408 11924
rect 13362 11736 13368 11912
rect 13402 11736 13408 11912
rect 13362 11724 13408 11736
rect 13480 11912 13526 11924
rect 13480 11736 13486 11912
rect 13520 11736 13526 11912
rect 13480 11724 13526 11736
rect 13599 11736 13605 12112
rect 13639 11736 13645 12112
rect 13599 11724 13645 11736
rect 13717 12112 13763 12124
rect 13717 11736 13723 12112
rect 13757 11736 13763 12112
rect 13717 11724 13763 11736
rect 13835 12112 13881 12124
rect 13835 11736 13841 12112
rect 13875 11736 13881 12112
rect 13835 11724 13881 11736
rect 13953 12112 13999 12124
rect 13953 11736 13959 12112
rect 13993 11736 13999 12112
rect 13953 11724 13999 11736
rect 14072 12112 14118 12124
rect 14072 11736 14078 12112
rect 14112 11736 14118 12112
rect 14072 11724 14118 11736
rect 14190 12112 14236 12124
rect 14190 11736 14196 12112
rect 14230 11736 14236 12112
rect 14190 11724 14236 11736
rect 14308 12112 14354 12124
rect 14308 11736 14314 12112
rect 14348 11736 14354 12112
rect 14308 11724 14354 11736
rect 14426 12112 14472 12124
rect 14426 11736 14432 12112
rect 14466 11736 14472 12112
rect 14426 11724 14472 11736
rect 14544 12112 14590 12124
rect 14544 11736 14550 12112
rect 14584 11736 14590 12112
rect 14544 11724 14590 11736
rect 14662 12112 14708 12124
rect 14662 11736 14668 12112
rect 14702 11736 14708 12112
rect 14662 11724 14708 11736
rect 14780 12112 14826 12124
rect 14780 11736 14786 12112
rect 14820 11736 14826 12112
rect 14780 11724 14826 11736
rect 14893 12112 14939 12124
rect 14893 11736 14899 12112
rect 14933 11736 14939 12112
rect 14893 11724 14939 11736
rect 15011 12112 15057 12124
rect 15011 11736 15017 12112
rect 15051 11736 15057 12112
rect 15011 11724 15057 11736
rect 15129 12112 15175 12124
rect 15129 11736 15135 12112
rect 15169 11736 15175 12112
rect 15129 11724 15175 11736
rect 15247 12112 15293 12124
rect 15247 11736 15253 12112
rect 15287 11924 15293 12112
rect 15287 11912 15380 11924
rect 15287 11736 15340 11912
rect 15374 11736 15380 11912
rect 15247 11724 15380 11736
rect 15452 11912 15498 11924
rect 15452 11736 15458 11912
rect 15492 11736 15498 11912
rect 15452 11724 15498 11736
rect 15570 11912 15616 11924
rect 15570 11736 15576 11912
rect 15610 11736 15616 11912
rect 15570 11724 15616 11736
rect 15688 11912 15734 11924
rect 15688 11736 15694 11912
rect 15728 11736 15734 11912
rect 15688 11724 15734 11736
rect 13131 11370 13166 11724
rect 13605 11640 13639 11724
rect 14786 11640 14820 11724
rect 13605 11598 14820 11640
rect 13605 11578 13639 11598
rect 13282 11562 13639 11578
rect 13282 11528 13298 11562
rect 13332 11528 13639 11562
rect 15694 11538 15729 11724
rect 13282 11512 13639 11528
rect 14592 11521 15729 11538
rect 14592 11487 14608 11521
rect 14642 11487 15729 11521
rect 14592 11471 15729 11487
rect 12610 11306 12786 11314
rect 12602 11238 12612 11306
rect 12669 11238 12786 11306
rect 12610 11230 12786 11238
rect 12985 11224 13166 11370
rect 14462 11425 14554 11435
rect 14462 11363 14472 11425
rect 14542 11363 14554 11425
rect 14462 11350 14554 11363
rect 15547 11425 15639 11438
rect 15547 11362 15556 11425
rect 15627 11362 15639 11425
rect 15547 11353 15639 11362
rect 14242 11308 14307 11311
rect 14238 11305 14307 11308
rect 14232 11245 14242 11305
rect 14301 11245 14307 11305
rect 14238 11241 14307 11245
rect 14242 11239 14307 11241
rect 12610 11138 12786 11146
rect 12602 11070 12612 11138
rect 12669 11070 12786 11138
rect 12610 11062 12786 11070
rect 10798 10787 10832 10911
rect 11155 10910 12527 10957
rect 11155 10897 11221 10910
rect 11155 10863 11171 10897
rect 11205 10863 11221 10897
rect 11155 10847 11221 10863
rect 11659 10787 11693 10910
rect 10792 10775 10838 10787
rect 10792 10599 10798 10775
rect 10832 10599 10838 10775
rect 10792 10587 10838 10599
rect 10910 10775 11034 10787
rect 10910 10599 10916 10775
rect 10950 10599 10994 10775
rect 10910 10587 10994 10599
rect 9773 10445 9783 10540
rect 9879 10445 9889 10540
rect 10916 10220 10950 10587
rect 10988 10399 10994 10587
rect 11028 10399 11034 10775
rect 10988 10387 11034 10399
rect 11106 10775 11152 10787
rect 11106 10399 11112 10775
rect 11146 10399 11152 10775
rect 11106 10387 11152 10399
rect 11224 10775 11270 10787
rect 11224 10399 11230 10775
rect 11264 10399 11270 10775
rect 11224 10387 11270 10399
rect 11342 10775 11388 10787
rect 11342 10399 11348 10775
rect 11382 10399 11388 10775
rect 11342 10387 11388 10399
rect 11460 10775 11580 10787
rect 11460 10399 11466 10775
rect 11500 10599 11540 10775
rect 11574 10599 11580 10775
rect 11500 10587 11580 10599
rect 11652 10775 11698 10787
rect 11652 10599 11658 10775
rect 11692 10599 11698 10775
rect 11652 10587 11698 10599
rect 11500 10399 11506 10587
rect 11460 10387 11506 10399
rect 11230 10314 11264 10387
rect 11213 10298 11279 10314
rect 11213 10264 11229 10298
rect 11263 10264 11279 10298
rect 11213 10248 11279 10264
rect 11540 10220 11574 10587
rect 10916 10168 11574 10220
rect 11184 10146 11276 10168
rect 11184 10094 11198 10146
rect 11264 10094 11276 10146
rect 11184 10090 11276 10094
rect 12710 9876 12786 11062
rect 12986 10336 13079 11224
rect 13131 10962 13166 11224
rect 14580 11142 14672 11150
rect 14580 11077 14592 11142
rect 14660 11077 14672 11142
rect 14580 11065 14672 11077
rect 13131 10915 14035 10962
rect 15694 10961 15729 11471
rect 15917 11318 15988 12636
rect 17534 12308 17544 12368
rect 17624 12308 17634 12368
rect 17534 12268 17634 12308
rect 16628 12211 18431 12268
rect 16628 11924 16665 12211
rect 17222 12124 17256 12211
rect 18397 12124 18431 12211
rect 16743 12112 16789 12124
rect 16270 11912 16316 11924
rect 16270 11736 16276 11912
rect 16310 11736 16316 11912
rect 16270 11724 16316 11736
rect 16388 11912 16434 11924
rect 16388 11736 16394 11912
rect 16428 11736 16434 11912
rect 16388 11724 16434 11736
rect 16506 11912 16552 11924
rect 16506 11736 16512 11912
rect 16546 11736 16552 11912
rect 16506 11724 16552 11736
rect 16624 11912 16670 11924
rect 16624 11736 16630 11912
rect 16664 11736 16670 11912
rect 16624 11724 16670 11736
rect 16743 11736 16749 12112
rect 16783 11736 16789 12112
rect 16743 11724 16789 11736
rect 16861 12112 16907 12124
rect 16861 11736 16867 12112
rect 16901 11736 16907 12112
rect 16861 11724 16907 11736
rect 16979 12112 17025 12124
rect 16979 11736 16985 12112
rect 17019 11736 17025 12112
rect 16979 11724 17025 11736
rect 17097 12112 17143 12124
rect 17097 11736 17103 12112
rect 17137 11736 17143 12112
rect 17097 11724 17143 11736
rect 17216 12112 17262 12124
rect 17216 11736 17222 12112
rect 17256 11736 17262 12112
rect 17216 11724 17262 11736
rect 17334 12112 17380 12124
rect 17334 11736 17340 12112
rect 17374 11736 17380 12112
rect 17334 11724 17380 11736
rect 17452 12112 17498 12124
rect 17452 11736 17458 12112
rect 17492 11736 17498 12112
rect 17452 11724 17498 11736
rect 17570 12112 17616 12124
rect 17570 11736 17576 12112
rect 17610 11736 17616 12112
rect 17570 11724 17616 11736
rect 17688 12112 17734 12124
rect 17688 11736 17694 12112
rect 17728 11736 17734 12112
rect 17688 11724 17734 11736
rect 17806 12112 17852 12124
rect 17806 11736 17812 12112
rect 17846 11736 17852 12112
rect 17806 11724 17852 11736
rect 17924 12112 17970 12124
rect 17924 11736 17930 12112
rect 17964 11736 17970 12112
rect 17924 11724 17970 11736
rect 18037 12112 18083 12124
rect 18037 11736 18043 12112
rect 18077 11736 18083 12112
rect 18037 11724 18083 11736
rect 18155 12112 18201 12124
rect 18155 11736 18161 12112
rect 18195 11736 18201 12112
rect 18155 11724 18201 11736
rect 18273 12112 18319 12124
rect 18273 11736 18279 12112
rect 18313 11736 18319 12112
rect 18273 11724 18319 11736
rect 18391 12112 18437 12124
rect 18391 11736 18397 12112
rect 18431 11924 18437 12112
rect 18431 11912 18524 11924
rect 18431 11736 18484 11912
rect 18518 11736 18524 11912
rect 18391 11724 18524 11736
rect 18596 11912 18642 11924
rect 18596 11736 18602 11912
rect 18636 11736 18642 11912
rect 18596 11724 18642 11736
rect 18714 11912 18760 11924
rect 18714 11736 18720 11912
rect 18754 11736 18760 11912
rect 18714 11724 18760 11736
rect 18832 11912 18878 11924
rect 18832 11736 18838 11912
rect 18872 11736 18878 11912
rect 18832 11724 18878 11736
rect 16275 11370 16310 11724
rect 16749 11640 16783 11724
rect 17930 11640 17964 11724
rect 16749 11598 17964 11640
rect 16749 11578 16783 11598
rect 16426 11562 16783 11578
rect 16426 11528 16442 11562
rect 16476 11528 16783 11562
rect 18838 11538 18873 11724
rect 16426 11512 16783 11528
rect 17736 11521 18873 11538
rect 17736 11487 17752 11521
rect 17786 11487 18873 11521
rect 17736 11471 18873 11487
rect 15812 11310 15988 11318
rect 15804 11242 15814 11310
rect 15871 11242 15988 11310
rect 15812 11234 15988 11242
rect 16129 11224 16310 11370
rect 17606 11425 17698 11435
rect 17606 11363 17616 11425
rect 17686 11363 17698 11425
rect 17606 11350 17698 11363
rect 18691 11425 18783 11438
rect 18691 11362 18700 11425
rect 18771 11362 18783 11425
rect 18691 11353 18783 11362
rect 17386 11308 17451 11311
rect 17382 11305 17451 11308
rect 17376 11245 17386 11305
rect 17445 11245 17451 11305
rect 17382 11241 17451 11245
rect 17386 11239 17451 11241
rect 15812 11142 15964 11150
rect 15804 11074 15814 11142
rect 15871 11074 15964 11142
rect 15812 11066 15964 11074
rect 14000 10791 14034 10915
rect 14357 10914 15729 10961
rect 14357 10901 14423 10914
rect 14357 10867 14373 10901
rect 14407 10867 14423 10901
rect 14357 10851 14423 10867
rect 14861 10791 14895 10914
rect 13994 10779 14040 10791
rect 13994 10603 14000 10779
rect 14034 10603 14040 10779
rect 13994 10591 14040 10603
rect 14112 10779 14236 10791
rect 14112 10603 14118 10779
rect 14152 10603 14196 10779
rect 14112 10591 14196 10603
rect 12986 10267 13001 10336
rect 13079 10267 13089 10336
rect 14118 10224 14152 10591
rect 14190 10403 14196 10591
rect 14230 10403 14236 10779
rect 14190 10391 14236 10403
rect 14308 10779 14354 10791
rect 14308 10403 14314 10779
rect 14348 10403 14354 10779
rect 14308 10391 14354 10403
rect 14426 10779 14472 10791
rect 14426 10403 14432 10779
rect 14466 10403 14472 10779
rect 14426 10391 14472 10403
rect 14544 10779 14590 10791
rect 14544 10403 14550 10779
rect 14584 10403 14590 10779
rect 14544 10391 14590 10403
rect 14662 10779 14782 10791
rect 14662 10403 14668 10779
rect 14702 10603 14742 10779
rect 14776 10603 14782 10779
rect 14702 10591 14782 10603
rect 14854 10779 14900 10791
rect 14854 10603 14860 10779
rect 14894 10603 14900 10779
rect 14854 10591 14900 10603
rect 14702 10403 14708 10591
rect 14662 10391 14708 10403
rect 14432 10318 14466 10391
rect 14415 10302 14481 10318
rect 14415 10268 14431 10302
rect 14465 10268 14481 10302
rect 14415 10252 14481 10268
rect 14742 10224 14776 10591
rect 14118 10172 14776 10224
rect 14386 10150 14478 10172
rect 14386 10098 14400 10150
rect 14466 10098 14478 10150
rect 14386 10094 14478 10098
rect 1964 9874 3318 9875
rect -1752 9831 117 9833
rect -1752 9815 213 9831
rect -1752 9758 -1730 9815
rect -1608 9814 213 9815
rect -1608 9758 138 9814
rect -1752 9754 138 9758
rect 202 9754 213 9814
rect -1752 9744 213 9754
rect 62 9742 213 9744
rect 514 9813 3318 9874
rect 3517 9814 6502 9875
rect 6649 9815 9618 9876
rect 9934 9815 12786 9876
rect 15903 9875 15964 11066
rect 16129 9992 16220 11224
rect 16275 10962 16310 11224
rect 17724 11142 17816 11150
rect 17724 11077 17736 11142
rect 17804 11077 17816 11142
rect 17724 11065 17816 11077
rect 16275 10915 17179 10962
rect 18838 10961 18873 11471
rect 19061 11318 19132 12636
rect 20666 12304 20676 12364
rect 20756 12304 20766 12364
rect 20666 12264 20766 12304
rect 19760 12207 21563 12264
rect 19760 11920 19797 12207
rect 20354 12120 20388 12207
rect 21529 12120 21563 12207
rect 19875 12108 19921 12120
rect 19402 11908 19448 11920
rect 19402 11732 19408 11908
rect 19442 11732 19448 11908
rect 19402 11720 19448 11732
rect 19520 11908 19566 11920
rect 19520 11732 19526 11908
rect 19560 11732 19566 11908
rect 19520 11720 19566 11732
rect 19638 11908 19684 11920
rect 19638 11732 19644 11908
rect 19678 11732 19684 11908
rect 19638 11720 19684 11732
rect 19756 11908 19802 11920
rect 19756 11732 19762 11908
rect 19796 11732 19802 11908
rect 19756 11720 19802 11732
rect 19875 11732 19881 12108
rect 19915 11732 19921 12108
rect 19875 11720 19921 11732
rect 19993 12108 20039 12120
rect 19993 11732 19999 12108
rect 20033 11732 20039 12108
rect 19993 11720 20039 11732
rect 20111 12108 20157 12120
rect 20111 11732 20117 12108
rect 20151 11732 20157 12108
rect 20111 11720 20157 11732
rect 20229 12108 20275 12120
rect 20229 11732 20235 12108
rect 20269 11732 20275 12108
rect 20229 11720 20275 11732
rect 20348 12108 20394 12120
rect 20348 11732 20354 12108
rect 20388 11732 20394 12108
rect 20348 11720 20394 11732
rect 20466 12108 20512 12120
rect 20466 11732 20472 12108
rect 20506 11732 20512 12108
rect 20466 11720 20512 11732
rect 20584 12108 20630 12120
rect 20584 11732 20590 12108
rect 20624 11732 20630 12108
rect 20584 11720 20630 11732
rect 20702 12108 20748 12120
rect 20702 11732 20708 12108
rect 20742 11732 20748 12108
rect 20702 11720 20748 11732
rect 20820 12108 20866 12120
rect 20820 11732 20826 12108
rect 20860 11732 20866 12108
rect 20820 11720 20866 11732
rect 20938 12108 20984 12120
rect 20938 11732 20944 12108
rect 20978 11732 20984 12108
rect 20938 11720 20984 11732
rect 21056 12108 21102 12120
rect 21056 11732 21062 12108
rect 21096 11732 21102 12108
rect 21056 11720 21102 11732
rect 21169 12108 21215 12120
rect 21169 11732 21175 12108
rect 21209 11732 21215 12108
rect 21169 11720 21215 11732
rect 21287 12108 21333 12120
rect 21287 11732 21293 12108
rect 21327 11732 21333 12108
rect 21287 11720 21333 11732
rect 21405 12108 21451 12120
rect 21405 11732 21411 12108
rect 21445 11732 21451 12108
rect 21405 11720 21451 11732
rect 21523 12108 21569 12120
rect 21523 11732 21529 12108
rect 21563 11920 21569 12108
rect 21563 11908 21656 11920
rect 21563 11732 21616 11908
rect 21650 11732 21656 11908
rect 21523 11720 21656 11732
rect 21728 11908 21774 11920
rect 21728 11732 21734 11908
rect 21768 11732 21774 11908
rect 21728 11720 21774 11732
rect 21846 11908 21892 11920
rect 21846 11732 21852 11908
rect 21886 11732 21892 11908
rect 21846 11720 21892 11732
rect 21964 11908 22010 11920
rect 21964 11732 21970 11908
rect 22004 11732 22010 11908
rect 21964 11720 22010 11732
rect 19407 11366 19442 11720
rect 19881 11636 19915 11720
rect 21062 11636 21096 11720
rect 19881 11594 21096 11636
rect 19881 11574 19915 11594
rect 19558 11558 19915 11574
rect 19558 11524 19574 11558
rect 19608 11524 19915 11558
rect 21970 11534 22005 11720
rect 19558 11508 19915 11524
rect 20868 11517 22005 11534
rect 20868 11483 20884 11517
rect 20918 11483 22005 11517
rect 20868 11467 22005 11483
rect 18956 11310 19132 11318
rect 18948 11242 18958 11310
rect 19015 11242 19132 11310
rect 18956 11234 19132 11242
rect 19261 11238 19442 11366
rect 20738 11421 20830 11431
rect 20738 11359 20748 11421
rect 20818 11359 20830 11421
rect 20738 11346 20830 11359
rect 21823 11421 21915 11434
rect 21823 11358 21832 11421
rect 21903 11358 21915 11421
rect 21823 11349 21915 11358
rect 20518 11304 20583 11307
rect 20514 11301 20583 11304
rect 20508 11241 20518 11301
rect 20577 11241 20583 11301
rect 19260 11220 19442 11238
rect 20514 11237 20583 11241
rect 20518 11235 20583 11237
rect 18956 11142 19115 11150
rect 18948 11074 18958 11142
rect 19015 11074 19115 11142
rect 18956 11066 19115 11074
rect 17144 10791 17178 10915
rect 17501 10914 18873 10961
rect 17501 10901 17567 10914
rect 17501 10867 17517 10901
rect 17551 10867 17567 10901
rect 17501 10851 17567 10867
rect 18005 10791 18039 10914
rect 17138 10779 17184 10791
rect 17138 10603 17144 10779
rect 17178 10603 17184 10779
rect 17138 10591 17184 10603
rect 17256 10779 17380 10791
rect 17256 10603 17262 10779
rect 17296 10603 17340 10779
rect 17256 10591 17340 10603
rect 17262 10224 17296 10591
rect 17334 10403 17340 10591
rect 17374 10403 17380 10779
rect 17334 10391 17380 10403
rect 17452 10779 17498 10791
rect 17452 10403 17458 10779
rect 17492 10403 17498 10779
rect 17452 10391 17498 10403
rect 17570 10779 17616 10791
rect 17570 10403 17576 10779
rect 17610 10403 17616 10779
rect 17570 10391 17616 10403
rect 17688 10779 17734 10791
rect 17688 10403 17694 10779
rect 17728 10403 17734 10779
rect 17688 10391 17734 10403
rect 17806 10779 17926 10791
rect 17806 10403 17812 10779
rect 17846 10603 17886 10779
rect 17920 10603 17926 10779
rect 17846 10591 17926 10603
rect 17998 10779 18044 10791
rect 17998 10603 18004 10779
rect 18038 10603 18044 10779
rect 17998 10591 18044 10603
rect 17846 10403 17852 10591
rect 17806 10391 17852 10403
rect 17576 10318 17610 10391
rect 17559 10302 17625 10318
rect 17559 10268 17575 10302
rect 17609 10268 17625 10302
rect 17559 10252 17625 10268
rect 17886 10224 17920 10591
rect 17262 10172 17920 10224
rect 17530 10150 17622 10172
rect 17530 10098 17544 10150
rect 17610 10098 17622 10150
rect 17530 10094 17622 10098
rect 16129 9926 16159 9992
rect 16149 9924 16159 9926
rect 16226 9924 16236 9992
rect 19066 9875 19115 11066
rect 19260 10118 19358 11220
rect 19407 10958 19442 11220
rect 20856 11138 20948 11146
rect 20856 11073 20868 11138
rect 20936 11073 20948 11138
rect 20856 11061 20948 11073
rect 19407 10911 20311 10958
rect 21970 10957 22005 11467
rect 22193 11314 22264 12636
rect 23810 12304 23820 12364
rect 23900 12304 23910 12364
rect 23810 12264 23910 12304
rect 22904 12207 24707 12264
rect 22904 11920 22941 12207
rect 23498 12120 23532 12207
rect 24673 12120 24707 12207
rect 23019 12108 23065 12120
rect 22546 11908 22592 11920
rect 22546 11732 22552 11908
rect 22586 11732 22592 11908
rect 22546 11720 22592 11732
rect 22664 11908 22710 11920
rect 22664 11732 22670 11908
rect 22704 11732 22710 11908
rect 22664 11720 22710 11732
rect 22782 11908 22828 11920
rect 22782 11732 22788 11908
rect 22822 11732 22828 11908
rect 22782 11720 22828 11732
rect 22900 11908 22946 11920
rect 22900 11732 22906 11908
rect 22940 11732 22946 11908
rect 22900 11720 22946 11732
rect 23019 11732 23025 12108
rect 23059 11732 23065 12108
rect 23019 11720 23065 11732
rect 23137 12108 23183 12120
rect 23137 11732 23143 12108
rect 23177 11732 23183 12108
rect 23137 11720 23183 11732
rect 23255 12108 23301 12120
rect 23255 11732 23261 12108
rect 23295 11732 23301 12108
rect 23255 11720 23301 11732
rect 23373 12108 23419 12120
rect 23373 11732 23379 12108
rect 23413 11732 23419 12108
rect 23373 11720 23419 11732
rect 23492 12108 23538 12120
rect 23492 11732 23498 12108
rect 23532 11732 23538 12108
rect 23492 11720 23538 11732
rect 23610 12108 23656 12120
rect 23610 11732 23616 12108
rect 23650 11732 23656 12108
rect 23610 11720 23656 11732
rect 23728 12108 23774 12120
rect 23728 11732 23734 12108
rect 23768 11732 23774 12108
rect 23728 11720 23774 11732
rect 23846 12108 23892 12120
rect 23846 11732 23852 12108
rect 23886 11732 23892 12108
rect 23846 11720 23892 11732
rect 23964 12108 24010 12120
rect 23964 11732 23970 12108
rect 24004 11732 24010 12108
rect 23964 11720 24010 11732
rect 24082 12108 24128 12120
rect 24082 11732 24088 12108
rect 24122 11732 24128 12108
rect 24082 11720 24128 11732
rect 24200 12108 24246 12120
rect 24200 11732 24206 12108
rect 24240 11732 24246 12108
rect 24200 11720 24246 11732
rect 24313 12108 24359 12120
rect 24313 11732 24319 12108
rect 24353 11732 24359 12108
rect 24313 11720 24359 11732
rect 24431 12108 24477 12120
rect 24431 11732 24437 12108
rect 24471 11732 24477 12108
rect 24431 11720 24477 11732
rect 24549 12108 24595 12120
rect 24549 11732 24555 12108
rect 24589 11732 24595 12108
rect 24549 11720 24595 11732
rect 24667 12108 24713 12120
rect 24667 11732 24673 12108
rect 24707 11920 24713 12108
rect 24707 11908 24800 11920
rect 24707 11732 24760 11908
rect 24794 11732 24800 11908
rect 24667 11720 24800 11732
rect 24872 11908 24918 11920
rect 24872 11732 24878 11908
rect 24912 11732 24918 11908
rect 24872 11720 24918 11732
rect 24990 11908 25036 11920
rect 24990 11732 24996 11908
rect 25030 11732 25036 11908
rect 24990 11720 25036 11732
rect 25108 11908 25154 11920
rect 25108 11732 25114 11908
rect 25148 11732 25154 11908
rect 25108 11720 25154 11732
rect 22551 11366 22586 11720
rect 23025 11636 23059 11720
rect 24206 11636 24240 11720
rect 23025 11594 24240 11636
rect 23025 11574 23059 11594
rect 22702 11558 23059 11574
rect 22702 11524 22718 11558
rect 22752 11524 23059 11558
rect 25114 11534 25149 11720
rect 22702 11508 23059 11524
rect 24012 11517 25149 11534
rect 24012 11483 24028 11517
rect 24062 11483 25149 11517
rect 24012 11467 25149 11483
rect 22088 11306 22264 11314
rect 22080 11238 22090 11306
rect 22147 11238 22264 11306
rect 22088 11230 22264 11238
rect 22405 11220 22586 11366
rect 23882 11421 23974 11431
rect 23882 11359 23892 11421
rect 23962 11359 23974 11421
rect 23882 11346 23974 11359
rect 24967 11421 25059 11434
rect 24967 11358 24976 11421
rect 25047 11358 25059 11421
rect 24967 11349 25059 11358
rect 23662 11304 23727 11307
rect 23658 11301 23727 11304
rect 23652 11241 23662 11301
rect 23721 11241 23727 11301
rect 23658 11237 23727 11241
rect 23662 11235 23727 11237
rect 22088 11138 22264 11146
rect 22080 11070 22090 11138
rect 22147 11070 22264 11138
rect 22088 11065 22264 11070
rect 22088 11062 22265 11065
rect 20276 10787 20310 10911
rect 20633 10910 22005 10957
rect 20633 10897 20699 10910
rect 20633 10863 20649 10897
rect 20683 10863 20699 10897
rect 20633 10847 20699 10863
rect 21137 10787 21171 10910
rect 20270 10775 20316 10787
rect 20270 10599 20276 10775
rect 20310 10599 20316 10775
rect 20270 10587 20316 10599
rect 20388 10775 20512 10787
rect 20388 10599 20394 10775
rect 20428 10599 20472 10775
rect 20388 10587 20472 10599
rect 20394 10220 20428 10587
rect 20466 10399 20472 10587
rect 20506 10399 20512 10775
rect 20466 10387 20512 10399
rect 20584 10775 20630 10787
rect 20584 10399 20590 10775
rect 20624 10399 20630 10775
rect 20584 10387 20630 10399
rect 20702 10775 20748 10787
rect 20702 10399 20708 10775
rect 20742 10399 20748 10775
rect 20702 10387 20748 10399
rect 20820 10775 20866 10787
rect 20820 10399 20826 10775
rect 20860 10399 20866 10775
rect 20820 10387 20866 10399
rect 20938 10775 21058 10787
rect 20938 10399 20944 10775
rect 20978 10599 21018 10775
rect 21052 10599 21058 10775
rect 20978 10587 21058 10599
rect 21130 10775 21176 10787
rect 21130 10599 21136 10775
rect 21170 10599 21176 10775
rect 21130 10587 21176 10599
rect 20978 10399 20984 10587
rect 20938 10387 20984 10399
rect 20708 10314 20742 10387
rect 20691 10298 20757 10314
rect 20691 10264 20707 10298
rect 20741 10264 20757 10298
rect 20691 10248 20757 10264
rect 21018 10220 21052 10587
rect 20394 10168 21052 10220
rect 20662 10146 20754 10168
rect 19260 10068 19294 10118
rect 19284 10046 19294 10068
rect 19362 10046 19372 10118
rect 20662 10094 20676 10146
rect 20742 10094 20754 10146
rect 20662 10090 20754 10094
rect 22190 9875 22265 11062
rect 22405 10177 22478 11220
rect 22551 10958 22586 11220
rect 24000 11138 24092 11146
rect 24000 11073 24012 11138
rect 24080 11073 24092 11138
rect 24000 11061 24092 11073
rect 22551 10911 23455 10958
rect 25114 10957 25149 11467
rect 25336 11314 25408 12636
rect 25232 11306 25408 11314
rect 25224 11238 25234 11306
rect 25291 11238 25408 11306
rect 25818 11247 25927 14070
rect 25232 11230 25408 11238
rect 25232 11138 25408 11146
rect 25224 11070 25234 11138
rect 25291 11070 25408 11138
rect 25232 11062 25408 11070
rect 23420 10787 23454 10911
rect 23777 10910 25149 10957
rect 23777 10897 23843 10910
rect 23777 10863 23793 10897
rect 23827 10863 23843 10897
rect 23777 10847 23843 10863
rect 24281 10787 24315 10910
rect 23414 10775 23460 10787
rect 23414 10599 23420 10775
rect 23454 10599 23460 10775
rect 23414 10587 23460 10599
rect 23532 10775 23656 10787
rect 23532 10599 23538 10775
rect 23572 10599 23616 10775
rect 23532 10587 23616 10599
rect 23538 10220 23572 10587
rect 23610 10399 23616 10587
rect 23650 10399 23656 10775
rect 23610 10387 23656 10399
rect 23728 10775 23774 10787
rect 23728 10399 23734 10775
rect 23768 10399 23774 10775
rect 23728 10387 23774 10399
rect 23846 10775 23892 10787
rect 23846 10399 23852 10775
rect 23886 10399 23892 10775
rect 23846 10387 23892 10399
rect 23964 10775 24010 10787
rect 23964 10399 23970 10775
rect 24004 10399 24010 10775
rect 23964 10387 24010 10399
rect 24082 10775 24202 10787
rect 24082 10399 24088 10775
rect 24122 10599 24162 10775
rect 24196 10599 24202 10775
rect 24122 10587 24202 10599
rect 24274 10775 24320 10787
rect 24274 10599 24280 10775
rect 24314 10599 24320 10775
rect 24274 10587 24320 10599
rect 24122 10399 24128 10587
rect 24082 10387 24128 10399
rect 23852 10314 23886 10387
rect 23835 10298 23901 10314
rect 23835 10264 23851 10298
rect 23885 10264 23901 10298
rect 23835 10248 23901 10264
rect 24162 10220 24196 10587
rect 22398 10100 22408 10177
rect 22472 10100 22482 10177
rect 23538 10168 24196 10220
rect 23806 10146 23898 10168
rect 22405 10099 22478 10100
rect 23806 10094 23820 10146
rect 23886 10094 23898 10146
rect 23806 10090 23898 10094
rect -2012 9480 149 9482
rect -2012 9460 216 9480
rect -2012 9455 136 9460
rect -2012 9398 -1991 9455
rect -1869 9399 136 9455
rect 203 9399 216 9460
rect -1869 9398 216 9399
rect -2012 9386 216 9398
rect 514 9180 560 9813
rect 1778 9576 1788 9636
rect 1868 9576 1878 9636
rect 1778 9536 1878 9576
rect 872 9479 2675 9536
rect 872 9192 909 9479
rect 1466 9392 1500 9479
rect 2641 9392 2675 9479
rect 987 9380 1033 9392
rect 514 9004 520 9180
rect 554 9004 560 9180
rect 514 8992 560 9004
rect 632 9180 678 9192
rect 632 9004 638 9180
rect 672 9004 678 9180
rect 632 8992 678 9004
rect 750 9180 796 9192
rect 750 9004 756 9180
rect 790 9004 796 9180
rect 750 8992 796 9004
rect 868 9180 914 9192
rect 868 9004 874 9180
rect 908 9004 914 9180
rect 868 8992 914 9004
rect 987 9004 993 9380
rect 1027 9004 1033 9380
rect 987 8992 1033 9004
rect 1105 9380 1151 9392
rect 1105 9004 1111 9380
rect 1145 9004 1151 9380
rect 1105 8992 1151 9004
rect 1223 9380 1269 9392
rect 1223 9004 1229 9380
rect 1263 9004 1269 9380
rect 1223 8992 1269 9004
rect 1341 9380 1387 9392
rect 1341 9004 1347 9380
rect 1381 9004 1387 9380
rect 1341 8992 1387 9004
rect 1460 9380 1506 9392
rect 1460 9004 1466 9380
rect 1500 9004 1506 9380
rect 1460 8992 1506 9004
rect 1578 9380 1624 9392
rect 1578 9004 1584 9380
rect 1618 9004 1624 9380
rect 1578 8992 1624 9004
rect 1696 9380 1742 9392
rect 1696 9004 1702 9380
rect 1736 9004 1742 9380
rect 1696 8992 1742 9004
rect 1814 9380 1860 9392
rect 1814 9004 1820 9380
rect 1854 9004 1860 9380
rect 1814 8992 1860 9004
rect 1932 9380 1978 9392
rect 1932 9004 1938 9380
rect 1972 9004 1978 9380
rect 1932 8992 1978 9004
rect 2050 9380 2096 9392
rect 2050 9004 2056 9380
rect 2090 9004 2096 9380
rect 2050 8992 2096 9004
rect 2168 9380 2214 9392
rect 2168 9004 2174 9380
rect 2208 9004 2214 9380
rect 2168 8992 2214 9004
rect 2281 9380 2327 9392
rect 2281 9004 2287 9380
rect 2321 9004 2327 9380
rect 2281 8992 2327 9004
rect 2399 9380 2445 9392
rect 2399 9004 2405 9380
rect 2439 9004 2445 9380
rect 2399 8992 2445 9004
rect 2517 9380 2563 9392
rect 2517 9004 2523 9380
rect 2557 9004 2563 9380
rect 2517 8992 2563 9004
rect 2635 9380 2681 9392
rect 2635 9004 2641 9380
rect 2675 9192 2681 9380
rect 2675 9180 2768 9192
rect 2675 9004 2728 9180
rect 2762 9004 2768 9180
rect 2635 8992 2768 9004
rect 2840 9180 2886 9192
rect 2840 9004 2846 9180
rect 2880 9004 2886 9180
rect 2840 8992 2886 9004
rect 2958 9180 3004 9192
rect 2958 9004 2964 9180
rect 2998 9004 3004 9180
rect 2958 8992 3004 9004
rect 3076 9180 3122 9192
rect 3076 9004 3082 9180
rect 3116 9004 3122 9180
rect 3076 8992 3122 9004
rect 519 8638 554 8992
rect 993 8908 1027 8992
rect 2174 8908 2208 8992
rect 993 8866 2208 8908
rect 993 8846 1027 8866
rect 670 8830 1027 8846
rect 670 8796 686 8830
rect 720 8796 1027 8830
rect 3082 8806 3117 8992
rect 670 8780 1027 8796
rect 1980 8789 3117 8806
rect 1980 8755 1996 8789
rect 2030 8755 3117 8789
rect 1980 8739 3117 8755
rect 518 8492 554 8638
rect 1850 8693 1942 8703
rect 1850 8631 1860 8693
rect 1930 8631 1942 8693
rect 1850 8618 1942 8631
rect 2935 8693 3027 8706
rect 2935 8630 2944 8693
rect 3015 8630 3027 8693
rect 2935 8621 3027 8630
rect 1630 8576 1695 8579
rect 1626 8573 1695 8576
rect 1620 8513 1630 8573
rect 1689 8513 1695 8573
rect 1626 8509 1695 8513
rect 1630 8507 1695 8509
rect 519 8230 554 8492
rect 1968 8410 2060 8418
rect 1968 8345 1980 8410
rect 2048 8345 2060 8410
rect 1968 8333 2060 8345
rect 519 8183 1423 8230
rect 3082 8229 3117 8739
rect 3200 8694 3376 8702
rect 3192 8626 3202 8694
rect 3259 8626 3376 8694
rect 3200 8618 3376 8626
rect 3517 8638 3588 9814
rect 4922 9576 4932 9636
rect 5012 9576 5022 9636
rect 4922 9536 5022 9576
rect 4016 9479 5819 9536
rect 4016 9192 4053 9479
rect 4610 9392 4644 9479
rect 5785 9392 5819 9479
rect 4131 9380 4177 9392
rect 3658 9180 3704 9192
rect 3658 9004 3664 9180
rect 3698 9004 3704 9180
rect 3658 8992 3704 9004
rect 3776 9180 3822 9192
rect 3776 9004 3782 9180
rect 3816 9004 3822 9180
rect 3776 8992 3822 9004
rect 3894 9180 3940 9192
rect 3894 9004 3900 9180
rect 3934 9004 3940 9180
rect 3894 8992 3940 9004
rect 4012 9180 4058 9192
rect 4012 9004 4018 9180
rect 4052 9004 4058 9180
rect 4012 8992 4058 9004
rect 4131 9004 4137 9380
rect 4171 9004 4177 9380
rect 4131 8992 4177 9004
rect 4249 9380 4295 9392
rect 4249 9004 4255 9380
rect 4289 9004 4295 9380
rect 4249 8992 4295 9004
rect 4367 9380 4413 9392
rect 4367 9004 4373 9380
rect 4407 9004 4413 9380
rect 4367 8992 4413 9004
rect 4485 9380 4531 9392
rect 4485 9004 4491 9380
rect 4525 9004 4531 9380
rect 4485 8992 4531 9004
rect 4604 9380 4650 9392
rect 4604 9004 4610 9380
rect 4644 9004 4650 9380
rect 4604 8992 4650 9004
rect 4722 9380 4768 9392
rect 4722 9004 4728 9380
rect 4762 9004 4768 9380
rect 4722 8992 4768 9004
rect 4840 9380 4886 9392
rect 4840 9004 4846 9380
rect 4880 9004 4886 9380
rect 4840 8992 4886 9004
rect 4958 9380 5004 9392
rect 4958 9004 4964 9380
rect 4998 9004 5004 9380
rect 4958 8992 5004 9004
rect 5076 9380 5122 9392
rect 5076 9004 5082 9380
rect 5116 9004 5122 9380
rect 5076 8992 5122 9004
rect 5194 9380 5240 9392
rect 5194 9004 5200 9380
rect 5234 9004 5240 9380
rect 5194 8992 5240 9004
rect 5312 9380 5358 9392
rect 5312 9004 5318 9380
rect 5352 9004 5358 9380
rect 5312 8992 5358 9004
rect 5425 9380 5471 9392
rect 5425 9004 5431 9380
rect 5465 9004 5471 9380
rect 5425 8992 5471 9004
rect 5543 9380 5589 9392
rect 5543 9004 5549 9380
rect 5583 9004 5589 9380
rect 5543 8992 5589 9004
rect 5661 9380 5707 9392
rect 5661 9004 5667 9380
rect 5701 9004 5707 9380
rect 5661 8992 5707 9004
rect 5779 9380 5825 9392
rect 5779 9004 5785 9380
rect 5819 9192 5825 9380
rect 5819 9180 5912 9192
rect 5819 9004 5872 9180
rect 5906 9004 5912 9180
rect 5779 8992 5912 9004
rect 5984 9180 6030 9192
rect 5984 9004 5990 9180
rect 6024 9004 6030 9180
rect 5984 8992 6030 9004
rect 6102 9180 6148 9192
rect 6102 9004 6108 9180
rect 6142 9004 6148 9180
rect 6102 8992 6148 9004
rect 6220 9180 6266 9192
rect 6220 9004 6226 9180
rect 6260 9004 6266 9180
rect 6220 8992 6266 9004
rect 3663 8638 3698 8992
rect 4137 8908 4171 8992
rect 5318 8908 5352 8992
rect 4137 8866 5352 8908
rect 4137 8846 4171 8866
rect 3814 8830 4171 8846
rect 3814 8796 3830 8830
rect 3864 8796 4171 8830
rect 6226 8806 6261 8992
rect 3814 8780 4171 8796
rect 5124 8789 6261 8806
rect 5124 8755 5140 8789
rect 5174 8755 6261 8789
rect 5124 8739 6261 8755
rect 3200 8578 3270 8586
rect 3192 8510 3202 8578
rect 3259 8510 3270 8578
rect 3200 8502 3270 8510
rect 3517 8492 3698 8638
rect 4994 8693 5086 8703
rect 4994 8631 5004 8693
rect 5074 8631 5086 8693
rect 4994 8618 5086 8631
rect 6079 8693 6171 8706
rect 6079 8630 6088 8693
rect 6159 8630 6171 8693
rect 6079 8621 6171 8630
rect 4774 8576 4839 8579
rect 4770 8573 4839 8576
rect 4764 8513 4774 8573
rect 4833 8513 4839 8573
rect 4770 8509 4839 8513
rect 4774 8507 4839 8509
rect 3270 8418 3334 8419
rect 3200 8410 3334 8418
rect 3192 8342 3202 8410
rect 3259 8342 3334 8410
rect 3200 8334 3334 8342
rect 1388 8059 1422 8183
rect 1745 8182 3117 8229
rect 1745 8169 1811 8182
rect 1745 8135 1761 8169
rect 1795 8135 1811 8169
rect 1745 8119 1811 8135
rect 2249 8059 2283 8182
rect 1382 8047 1428 8059
rect 1382 7871 1388 8047
rect 1422 7871 1428 8047
rect 1382 7859 1428 7871
rect 1500 8047 1624 8059
rect 1500 7871 1506 8047
rect 1540 7871 1584 8047
rect 1500 7859 1584 7871
rect 1506 7492 1540 7859
rect 1578 7671 1584 7859
rect 1618 7671 1624 8047
rect 1578 7659 1624 7671
rect 1696 8047 1742 8059
rect 1696 7671 1702 8047
rect 1736 7671 1742 8047
rect 1696 7659 1742 7671
rect 1814 8047 1860 8059
rect 1814 7671 1820 8047
rect 1854 7671 1860 8047
rect 1814 7659 1860 7671
rect 1932 8047 1978 8059
rect 1932 7671 1938 8047
rect 1972 7671 1978 8047
rect 1932 7659 1978 7671
rect 2050 8047 2170 8059
rect 2050 7671 2056 8047
rect 2090 7871 2130 8047
rect 2164 7871 2170 8047
rect 2090 7859 2170 7871
rect 2242 8047 2288 8059
rect 2242 7871 2248 8047
rect 2282 7871 2288 8047
rect 2242 7859 2288 7871
rect 2090 7671 2096 7859
rect 2050 7659 2096 7671
rect 1820 7586 1854 7659
rect 1803 7570 1869 7586
rect 1803 7536 1819 7570
rect 1853 7536 1869 7570
rect 1803 7520 1869 7536
rect 2130 7492 2164 7859
rect 1506 7440 2164 7492
rect 1774 7418 1866 7440
rect 1774 7366 1788 7418
rect 1854 7366 1866 7418
rect 1774 7362 1866 7366
rect 3270 6954 3334 8334
rect 3663 8230 3698 8492
rect 5112 8410 5204 8418
rect 5112 8345 5124 8410
rect 5192 8345 5204 8410
rect 5112 8333 5204 8345
rect 3663 8183 4567 8230
rect 6226 8229 6261 8739
rect 6344 8694 6520 8702
rect 6336 8626 6346 8694
rect 6403 8626 6520 8694
rect 6344 8618 6520 8626
rect 6649 8634 6720 9815
rect 8054 9572 8064 9632
rect 8144 9572 8154 9632
rect 8054 9532 8154 9572
rect 7148 9475 8951 9532
rect 7148 9188 7185 9475
rect 7742 9388 7776 9475
rect 8917 9388 8951 9475
rect 7263 9376 7309 9388
rect 6790 9176 6836 9188
rect 6790 9000 6796 9176
rect 6830 9000 6836 9176
rect 6790 8988 6836 9000
rect 6908 9176 6954 9188
rect 6908 9000 6914 9176
rect 6948 9000 6954 9176
rect 6908 8988 6954 9000
rect 7026 9176 7072 9188
rect 7026 9000 7032 9176
rect 7066 9000 7072 9176
rect 7026 8988 7072 9000
rect 7144 9176 7190 9188
rect 7144 9000 7150 9176
rect 7184 9000 7190 9176
rect 7144 8988 7190 9000
rect 7263 9000 7269 9376
rect 7303 9000 7309 9376
rect 7263 8988 7309 9000
rect 7381 9376 7427 9388
rect 7381 9000 7387 9376
rect 7421 9000 7427 9376
rect 7381 8988 7427 9000
rect 7499 9376 7545 9388
rect 7499 9000 7505 9376
rect 7539 9000 7545 9376
rect 7499 8988 7545 9000
rect 7617 9376 7663 9388
rect 7617 9000 7623 9376
rect 7657 9000 7663 9376
rect 7617 8988 7663 9000
rect 7736 9376 7782 9388
rect 7736 9000 7742 9376
rect 7776 9000 7782 9376
rect 7736 8988 7782 9000
rect 7854 9376 7900 9388
rect 7854 9000 7860 9376
rect 7894 9000 7900 9376
rect 7854 8988 7900 9000
rect 7972 9376 8018 9388
rect 7972 9000 7978 9376
rect 8012 9000 8018 9376
rect 7972 8988 8018 9000
rect 8090 9376 8136 9388
rect 8090 9000 8096 9376
rect 8130 9000 8136 9376
rect 8090 8988 8136 9000
rect 8208 9376 8254 9388
rect 8208 9000 8214 9376
rect 8248 9000 8254 9376
rect 8208 8988 8254 9000
rect 8326 9376 8372 9388
rect 8326 9000 8332 9376
rect 8366 9000 8372 9376
rect 8326 8988 8372 9000
rect 8444 9376 8490 9388
rect 8444 9000 8450 9376
rect 8484 9000 8490 9376
rect 8444 8988 8490 9000
rect 8557 9376 8603 9388
rect 8557 9000 8563 9376
rect 8597 9000 8603 9376
rect 8557 8988 8603 9000
rect 8675 9376 8721 9388
rect 8675 9000 8681 9376
rect 8715 9000 8721 9376
rect 8675 8988 8721 9000
rect 8793 9376 8839 9388
rect 8793 9000 8799 9376
rect 8833 9000 8839 9376
rect 8793 8988 8839 9000
rect 8911 9376 8957 9388
rect 8911 9000 8917 9376
rect 8951 9188 8957 9376
rect 8951 9176 9044 9188
rect 8951 9000 9004 9176
rect 9038 9000 9044 9176
rect 8911 8988 9044 9000
rect 9116 9176 9162 9188
rect 9116 9000 9122 9176
rect 9156 9000 9162 9176
rect 9116 8988 9162 9000
rect 9234 9176 9280 9188
rect 9234 9000 9240 9176
rect 9274 9000 9280 9176
rect 9234 8988 9280 9000
rect 9352 9176 9398 9188
rect 9352 9000 9358 9176
rect 9392 9000 9398 9176
rect 9352 8988 9398 9000
rect 9934 9176 9980 9815
rect 12994 9814 15964 9875
rect 16139 9814 19115 9875
rect 11198 9572 11208 9632
rect 11288 9572 11298 9632
rect 11198 9532 11298 9572
rect 10292 9475 12095 9532
rect 10292 9188 10329 9475
rect 10886 9388 10920 9475
rect 12061 9388 12095 9475
rect 10407 9376 10453 9388
rect 9934 9000 9940 9176
rect 9974 9000 9980 9176
rect 9934 8988 9980 9000
rect 10052 9176 10098 9188
rect 10052 9000 10058 9176
rect 10092 9000 10098 9176
rect 10052 8988 10098 9000
rect 10170 9176 10216 9188
rect 10170 9000 10176 9176
rect 10210 9000 10216 9176
rect 10170 8988 10216 9000
rect 10288 9176 10334 9188
rect 10288 9000 10294 9176
rect 10328 9000 10334 9176
rect 10288 8988 10334 9000
rect 10407 9000 10413 9376
rect 10447 9000 10453 9376
rect 10407 8988 10453 9000
rect 10525 9376 10571 9388
rect 10525 9000 10531 9376
rect 10565 9000 10571 9376
rect 10525 8988 10571 9000
rect 10643 9376 10689 9388
rect 10643 9000 10649 9376
rect 10683 9000 10689 9376
rect 10643 8988 10689 9000
rect 10761 9376 10807 9388
rect 10761 9000 10767 9376
rect 10801 9000 10807 9376
rect 10761 8988 10807 9000
rect 10880 9376 10926 9388
rect 10880 9000 10886 9376
rect 10920 9000 10926 9376
rect 10880 8988 10926 9000
rect 10998 9376 11044 9388
rect 10998 9000 11004 9376
rect 11038 9000 11044 9376
rect 10998 8988 11044 9000
rect 11116 9376 11162 9388
rect 11116 9000 11122 9376
rect 11156 9000 11162 9376
rect 11116 8988 11162 9000
rect 11234 9376 11280 9388
rect 11234 9000 11240 9376
rect 11274 9000 11280 9376
rect 11234 8988 11280 9000
rect 11352 9376 11398 9388
rect 11352 9000 11358 9376
rect 11392 9000 11398 9376
rect 11352 8988 11398 9000
rect 11470 9376 11516 9388
rect 11470 9000 11476 9376
rect 11510 9000 11516 9376
rect 11470 8988 11516 9000
rect 11588 9376 11634 9388
rect 11588 9000 11594 9376
rect 11628 9000 11634 9376
rect 11588 8988 11634 9000
rect 11701 9376 11747 9388
rect 11701 9000 11707 9376
rect 11741 9000 11747 9376
rect 11701 8988 11747 9000
rect 11819 9376 11865 9388
rect 11819 9000 11825 9376
rect 11859 9000 11865 9376
rect 11819 8988 11865 9000
rect 11937 9376 11983 9388
rect 11937 9000 11943 9376
rect 11977 9000 11983 9376
rect 11937 8988 11983 9000
rect 12055 9376 12101 9388
rect 12055 9000 12061 9376
rect 12095 9188 12101 9376
rect 12095 9176 12188 9188
rect 12095 9000 12148 9176
rect 12182 9000 12188 9176
rect 12055 8988 12188 9000
rect 12260 9176 12306 9188
rect 12260 9000 12266 9176
rect 12300 9000 12306 9176
rect 12260 8988 12306 9000
rect 12378 9176 12424 9188
rect 12378 9000 12384 9176
rect 12418 9000 12424 9176
rect 12378 8988 12424 9000
rect 12496 9176 12542 9188
rect 12496 9000 12502 9176
rect 12536 9000 12542 9176
rect 12496 8988 12542 9000
rect 6795 8634 6830 8988
rect 7269 8904 7303 8988
rect 8450 8904 8484 8988
rect 7269 8862 8484 8904
rect 7269 8842 7303 8862
rect 6946 8826 7303 8842
rect 6946 8792 6962 8826
rect 6996 8792 7303 8826
rect 9358 8802 9393 8988
rect 6946 8776 7303 8792
rect 8256 8785 9393 8802
rect 8256 8751 8272 8785
rect 8306 8751 9393 8785
rect 8256 8735 9393 8751
rect 6344 8578 6414 8586
rect 6336 8510 6346 8578
rect 6403 8510 6414 8578
rect 6344 8502 6414 8510
rect 6649 8488 6830 8634
rect 8126 8689 8218 8699
rect 8126 8627 8136 8689
rect 8206 8627 8218 8689
rect 8126 8614 8218 8627
rect 9211 8689 9303 8702
rect 9211 8626 9220 8689
rect 9291 8626 9303 8689
rect 9211 8617 9303 8626
rect 7906 8572 7971 8575
rect 7902 8569 7971 8572
rect 7896 8509 7906 8569
rect 7965 8509 7971 8569
rect 7902 8505 7971 8509
rect 7906 8503 7971 8505
rect 6344 8410 6463 8418
rect 6336 8342 6346 8410
rect 6403 8342 6463 8410
rect 6344 8334 6463 8342
rect 4532 8059 4566 8183
rect 4889 8182 6261 8229
rect 4889 8169 4955 8182
rect 4889 8135 4905 8169
rect 4939 8135 4955 8169
rect 4889 8119 4955 8135
rect 5393 8059 5427 8182
rect 4526 8047 4572 8059
rect 4526 7871 4532 8047
rect 4566 7871 4572 8047
rect 4526 7859 4572 7871
rect 4644 8047 4768 8059
rect 4644 7871 4650 8047
rect 4684 7871 4728 8047
rect 4644 7859 4728 7871
rect 4650 7492 4684 7859
rect 4722 7671 4728 7859
rect 4762 7671 4768 8047
rect 4722 7659 4768 7671
rect 4840 8047 4886 8059
rect 4840 7671 4846 8047
rect 4880 7671 4886 8047
rect 4840 7659 4886 7671
rect 4958 8047 5004 8059
rect 4958 7671 4964 8047
rect 4998 7671 5004 8047
rect 4958 7659 5004 7671
rect 5076 8047 5122 8059
rect 5076 7671 5082 8047
rect 5116 7671 5122 8047
rect 5076 7659 5122 7671
rect 5194 8047 5314 8059
rect 5194 7671 5200 8047
rect 5234 7871 5274 8047
rect 5308 7871 5314 8047
rect 5234 7859 5314 7871
rect 5386 8047 5432 8059
rect 5386 7871 5392 8047
rect 5426 7871 5432 8047
rect 5386 7859 5432 7871
rect 5234 7671 5240 7859
rect 5194 7659 5240 7671
rect 4964 7586 4998 7659
rect 4947 7570 5013 7586
rect 4947 7536 4963 7570
rect 4997 7536 5013 7570
rect 4947 7520 5013 7536
rect 5274 7492 5308 7859
rect 4650 7440 5308 7492
rect 4918 7418 5010 7440
rect 4918 7366 4932 7418
rect 4998 7366 5010 7418
rect 4918 7362 5010 7366
rect 6415 7326 6463 8334
rect 6795 8226 6830 8488
rect 8244 8406 8336 8414
rect 8244 8341 8256 8406
rect 8324 8341 8336 8406
rect 8244 8329 8336 8341
rect 6795 8179 7699 8226
rect 9358 8225 9393 8735
rect 9476 8690 9652 8698
rect 9468 8622 9478 8690
rect 9535 8622 9652 8690
rect 9476 8614 9652 8622
rect 9476 8574 9547 8582
rect 9468 8506 9478 8574
rect 9535 8506 9547 8574
rect 9476 8498 9547 8506
rect 9546 8414 9594 8415
rect 9476 8406 9595 8414
rect 9468 8338 9478 8406
rect 9535 8338 9595 8406
rect 9476 8330 9595 8338
rect 7664 8055 7698 8179
rect 8021 8178 9393 8225
rect 8021 8165 8087 8178
rect 8021 8131 8037 8165
rect 8071 8131 8087 8165
rect 8021 8115 8087 8131
rect 8525 8055 8559 8178
rect 7658 8043 7704 8055
rect 7658 7867 7664 8043
rect 7698 7867 7704 8043
rect 7658 7855 7704 7867
rect 7776 8043 7900 8055
rect 7776 7867 7782 8043
rect 7816 7867 7860 8043
rect 7776 7855 7860 7867
rect 7782 7488 7816 7855
rect 7854 7667 7860 7855
rect 7894 7667 7900 8043
rect 7854 7655 7900 7667
rect 7972 8043 8018 8055
rect 7972 7667 7978 8043
rect 8012 7667 8018 8043
rect 7972 7655 8018 7667
rect 8090 8043 8136 8055
rect 8090 7667 8096 8043
rect 8130 7667 8136 8043
rect 8090 7655 8136 7667
rect 8208 8043 8254 8055
rect 8208 7667 8214 8043
rect 8248 7667 8254 8043
rect 8208 7655 8254 7667
rect 8326 8043 8446 8055
rect 8326 7667 8332 8043
rect 8366 7867 8406 8043
rect 8440 7867 8446 8043
rect 8366 7855 8446 7867
rect 8518 8043 8564 8055
rect 8518 7867 8524 8043
rect 8558 7867 8564 8043
rect 8518 7855 8564 7867
rect 8366 7667 8372 7855
rect 8326 7655 8372 7667
rect 8096 7582 8130 7655
rect 8079 7566 8145 7582
rect 8079 7532 8095 7566
rect 8129 7532 8145 7566
rect 8079 7516 8145 7532
rect 8406 7488 8440 7855
rect 7782 7436 8440 7488
rect 8050 7414 8142 7436
rect 8050 7362 8064 7414
rect 8130 7362 8142 7414
rect 8050 7358 8142 7362
rect 3003 6890 3334 6954
rect 3743 7278 6463 7326
rect 9546 7323 9594 8330
rect 9939 8226 9974 8988
rect 10413 8904 10447 8988
rect 11594 8904 11628 8988
rect 10413 8862 11628 8904
rect 10413 8842 10447 8862
rect 10090 8826 10447 8842
rect 10090 8792 10106 8826
rect 10140 8792 10447 8826
rect 12502 8802 12537 8988
rect 10090 8776 10447 8792
rect 11400 8785 12537 8802
rect 11400 8751 11416 8785
rect 11450 8751 12537 8785
rect 11400 8735 12537 8751
rect 11270 8689 11362 8699
rect 11270 8627 11280 8689
rect 11350 8627 11362 8689
rect 11270 8614 11362 8627
rect 12355 8689 12447 8702
rect 12355 8626 12364 8689
rect 12435 8626 12447 8689
rect 12355 8617 12447 8626
rect 11050 8572 11115 8575
rect 11046 8569 11115 8572
rect 11040 8509 11050 8569
rect 11109 8509 11115 8569
rect 11046 8505 11115 8509
rect 11050 8503 11115 8505
rect 11388 8406 11480 8414
rect 11388 8341 11400 8406
rect 11468 8341 11480 8406
rect 11388 8329 11480 8341
rect 9939 8179 10843 8226
rect 12502 8225 12537 8735
rect 12620 8690 12796 8698
rect 12612 8622 12622 8690
rect 12679 8622 12796 8690
rect 12994 8638 13065 9814
rect 14400 9576 14410 9636
rect 14490 9576 14500 9636
rect 14400 9536 14500 9576
rect 13494 9479 15297 9536
rect 13494 9192 13531 9479
rect 14088 9392 14122 9479
rect 15263 9392 15297 9479
rect 13609 9380 13655 9392
rect 13136 9180 13182 9192
rect 13136 9004 13142 9180
rect 13176 9004 13182 9180
rect 13136 8992 13182 9004
rect 13254 9180 13300 9192
rect 13254 9004 13260 9180
rect 13294 9004 13300 9180
rect 13254 8992 13300 9004
rect 13372 9180 13418 9192
rect 13372 9004 13378 9180
rect 13412 9004 13418 9180
rect 13372 8992 13418 9004
rect 13490 9180 13536 9192
rect 13490 9004 13496 9180
rect 13530 9004 13536 9180
rect 13490 8992 13536 9004
rect 13609 9004 13615 9380
rect 13649 9004 13655 9380
rect 13609 8992 13655 9004
rect 13727 9380 13773 9392
rect 13727 9004 13733 9380
rect 13767 9004 13773 9380
rect 13727 8992 13773 9004
rect 13845 9380 13891 9392
rect 13845 9004 13851 9380
rect 13885 9004 13891 9380
rect 13845 8992 13891 9004
rect 13963 9380 14009 9392
rect 13963 9004 13969 9380
rect 14003 9004 14009 9380
rect 13963 8992 14009 9004
rect 14082 9380 14128 9392
rect 14082 9004 14088 9380
rect 14122 9004 14128 9380
rect 14082 8992 14128 9004
rect 14200 9380 14246 9392
rect 14200 9004 14206 9380
rect 14240 9004 14246 9380
rect 14200 8992 14246 9004
rect 14318 9380 14364 9392
rect 14318 9004 14324 9380
rect 14358 9004 14364 9380
rect 14318 8992 14364 9004
rect 14436 9380 14482 9392
rect 14436 9004 14442 9380
rect 14476 9004 14482 9380
rect 14436 8992 14482 9004
rect 14554 9380 14600 9392
rect 14554 9004 14560 9380
rect 14594 9004 14600 9380
rect 14554 8992 14600 9004
rect 14672 9380 14718 9392
rect 14672 9004 14678 9380
rect 14712 9004 14718 9380
rect 14672 8992 14718 9004
rect 14790 9380 14836 9392
rect 14790 9004 14796 9380
rect 14830 9004 14836 9380
rect 14790 8992 14836 9004
rect 14903 9380 14949 9392
rect 14903 9004 14909 9380
rect 14943 9004 14949 9380
rect 14903 8992 14949 9004
rect 15021 9380 15067 9392
rect 15021 9004 15027 9380
rect 15061 9004 15067 9380
rect 15021 8992 15067 9004
rect 15139 9380 15185 9392
rect 15139 9004 15145 9380
rect 15179 9004 15185 9380
rect 15139 8992 15185 9004
rect 15257 9380 15303 9392
rect 15257 9004 15263 9380
rect 15297 9192 15303 9380
rect 15297 9180 15390 9192
rect 15297 9004 15350 9180
rect 15384 9004 15390 9180
rect 15257 8992 15390 9004
rect 15462 9180 15508 9192
rect 15462 9004 15468 9180
rect 15502 9004 15508 9180
rect 15462 8992 15508 9004
rect 15580 9180 15626 9192
rect 15580 9004 15586 9180
rect 15620 9004 15626 9180
rect 15580 8992 15626 9004
rect 15698 9180 15744 9192
rect 15698 9004 15704 9180
rect 15738 9004 15744 9180
rect 15698 8992 15744 9004
rect 13141 8638 13176 8992
rect 13615 8908 13649 8992
rect 14796 8908 14830 8992
rect 13615 8866 14830 8908
rect 13615 8846 13649 8866
rect 13292 8830 13649 8846
rect 13292 8796 13308 8830
rect 13342 8796 13649 8830
rect 15704 8806 15739 8992
rect 13292 8780 13649 8796
rect 14602 8789 15739 8806
rect 14602 8755 14618 8789
rect 14652 8755 15739 8789
rect 14602 8739 15739 8755
rect 12620 8614 12796 8622
rect 12620 8574 12690 8582
rect 12612 8506 12622 8574
rect 12679 8506 12690 8574
rect 12620 8498 12690 8506
rect 12995 8492 13176 8638
rect 14472 8693 14564 8703
rect 14472 8631 14482 8693
rect 14552 8631 14564 8693
rect 14472 8618 14564 8631
rect 15557 8693 15649 8706
rect 15557 8630 15566 8693
rect 15637 8630 15649 8693
rect 15557 8621 15649 8630
rect 14252 8576 14317 8579
rect 14248 8573 14317 8576
rect 14242 8513 14252 8573
rect 14311 8513 14317 8573
rect 14248 8509 14317 8513
rect 14252 8507 14317 8509
rect 12620 8406 12736 8414
rect 12612 8338 12622 8406
rect 12679 8338 12736 8406
rect 12620 8330 12736 8338
rect 10808 8055 10842 8179
rect 11165 8178 12537 8225
rect 11165 8165 11231 8178
rect 11165 8131 11181 8165
rect 11215 8131 11231 8165
rect 11165 8115 11231 8131
rect 11669 8055 11703 8178
rect 10802 8043 10848 8055
rect 10802 7867 10808 8043
rect 10842 7867 10848 8043
rect 10802 7855 10848 7867
rect 10920 8043 11044 8055
rect 10920 7867 10926 8043
rect 10960 7867 11004 8043
rect 10920 7855 11004 7867
rect 10926 7488 10960 7855
rect 10998 7667 11004 7855
rect 11038 7667 11044 8043
rect 10998 7655 11044 7667
rect 11116 8043 11162 8055
rect 11116 7667 11122 8043
rect 11156 7667 11162 8043
rect 11116 7655 11162 7667
rect 11234 8043 11280 8055
rect 11234 7667 11240 8043
rect 11274 7667 11280 8043
rect 11234 7655 11280 7667
rect 11352 8043 11398 8055
rect 11352 7667 11358 8043
rect 11392 7667 11398 8043
rect 11352 7655 11398 7667
rect 11470 8043 11590 8055
rect 11470 7667 11476 8043
rect 11510 7867 11550 8043
rect 11584 7867 11590 8043
rect 11510 7855 11590 7867
rect 11662 8043 11708 8055
rect 11662 7867 11668 8043
rect 11702 7867 11708 8043
rect 11662 7855 11708 7867
rect 11510 7667 11516 7855
rect 11470 7655 11516 7667
rect 11240 7582 11274 7655
rect 11223 7566 11289 7582
rect 11223 7532 11239 7566
rect 11273 7532 11289 7566
rect 11223 7516 11289 7532
rect 11550 7488 11584 7855
rect 10926 7436 11584 7488
rect 11194 7414 11286 7436
rect 11194 7362 11208 7414
rect 11274 7362 11286 7414
rect 11194 7358 11286 7362
rect 12688 7323 12736 8330
rect 13141 8230 13176 8492
rect 14590 8410 14682 8418
rect 14590 8345 14602 8410
rect 14670 8345 14682 8410
rect 14590 8333 14682 8345
rect 13141 8183 14045 8230
rect 15704 8229 15739 8739
rect 15822 8694 15998 8702
rect 15814 8626 15824 8694
rect 15881 8626 15998 8694
rect 15822 8618 15998 8626
rect 16139 8638 16210 9814
rect 19066 9812 19115 9814
rect 19271 9814 22265 9875
rect 25324 9874 25408 11062
rect 22414 9814 25408 9874
rect 25817 11099 25927 11247
rect 25817 11029 25837 11099
rect 25904 11029 25927 11099
rect 17544 9576 17554 9636
rect 17634 9576 17644 9636
rect 17544 9536 17644 9576
rect 16638 9479 18441 9536
rect 16638 9192 16675 9479
rect 17232 9392 17266 9479
rect 18407 9392 18441 9479
rect 16753 9380 16799 9392
rect 16280 9180 16326 9192
rect 16280 9004 16286 9180
rect 16320 9004 16326 9180
rect 16280 8992 16326 9004
rect 16398 9180 16444 9192
rect 16398 9004 16404 9180
rect 16438 9004 16444 9180
rect 16398 8992 16444 9004
rect 16516 9180 16562 9192
rect 16516 9004 16522 9180
rect 16556 9004 16562 9180
rect 16516 8992 16562 9004
rect 16634 9180 16680 9192
rect 16634 9004 16640 9180
rect 16674 9004 16680 9180
rect 16634 8992 16680 9004
rect 16753 9004 16759 9380
rect 16793 9004 16799 9380
rect 16753 8992 16799 9004
rect 16871 9380 16917 9392
rect 16871 9004 16877 9380
rect 16911 9004 16917 9380
rect 16871 8992 16917 9004
rect 16989 9380 17035 9392
rect 16989 9004 16995 9380
rect 17029 9004 17035 9380
rect 16989 8992 17035 9004
rect 17107 9380 17153 9392
rect 17107 9004 17113 9380
rect 17147 9004 17153 9380
rect 17107 8992 17153 9004
rect 17226 9380 17272 9392
rect 17226 9004 17232 9380
rect 17266 9004 17272 9380
rect 17226 8992 17272 9004
rect 17344 9380 17390 9392
rect 17344 9004 17350 9380
rect 17384 9004 17390 9380
rect 17344 8992 17390 9004
rect 17462 9380 17508 9392
rect 17462 9004 17468 9380
rect 17502 9004 17508 9380
rect 17462 8992 17508 9004
rect 17580 9380 17626 9392
rect 17580 9004 17586 9380
rect 17620 9004 17626 9380
rect 17580 8992 17626 9004
rect 17698 9380 17744 9392
rect 17698 9004 17704 9380
rect 17738 9004 17744 9380
rect 17698 8992 17744 9004
rect 17816 9380 17862 9392
rect 17816 9004 17822 9380
rect 17856 9004 17862 9380
rect 17816 8992 17862 9004
rect 17934 9380 17980 9392
rect 17934 9004 17940 9380
rect 17974 9004 17980 9380
rect 17934 8992 17980 9004
rect 18047 9380 18093 9392
rect 18047 9004 18053 9380
rect 18087 9004 18093 9380
rect 18047 8992 18093 9004
rect 18165 9380 18211 9392
rect 18165 9004 18171 9380
rect 18205 9004 18211 9380
rect 18165 8992 18211 9004
rect 18283 9380 18329 9392
rect 18283 9004 18289 9380
rect 18323 9004 18329 9380
rect 18283 8992 18329 9004
rect 18401 9380 18447 9392
rect 18401 9004 18407 9380
rect 18441 9192 18447 9380
rect 18441 9180 18534 9192
rect 18441 9004 18494 9180
rect 18528 9004 18534 9180
rect 18401 8992 18534 9004
rect 18606 9180 18652 9192
rect 18606 9004 18612 9180
rect 18646 9004 18652 9180
rect 18606 8992 18652 9004
rect 18724 9180 18770 9192
rect 18724 9004 18730 9180
rect 18764 9004 18770 9180
rect 18724 8992 18770 9004
rect 18842 9180 18888 9192
rect 18842 9004 18848 9180
rect 18882 9004 18888 9180
rect 18842 8992 18888 9004
rect 16285 8638 16320 8992
rect 16759 8908 16793 8992
rect 17940 8908 17974 8992
rect 16759 8866 17974 8908
rect 16759 8846 16793 8866
rect 16436 8830 16793 8846
rect 16436 8796 16452 8830
rect 16486 8796 16793 8830
rect 18848 8806 18883 8992
rect 16436 8780 16793 8796
rect 17746 8789 18883 8806
rect 17746 8755 17762 8789
rect 17796 8755 18883 8789
rect 17746 8739 18883 8755
rect 15822 8578 15892 8586
rect 15814 8510 15824 8578
rect 15881 8510 15892 8578
rect 15822 8502 15892 8510
rect 16139 8500 16320 8638
rect 17616 8693 17708 8703
rect 17616 8631 17626 8693
rect 17696 8631 17708 8693
rect 17616 8618 17708 8631
rect 18701 8693 18793 8706
rect 18701 8630 18710 8693
rect 18781 8630 18793 8693
rect 18701 8621 18793 8630
rect 17396 8576 17461 8579
rect 17392 8573 17461 8576
rect 17386 8513 17396 8573
rect 17455 8513 17461 8573
rect 17392 8509 17461 8513
rect 17396 8507 17461 8509
rect 15822 8410 15940 8418
rect 15814 8342 15824 8410
rect 15881 8342 15940 8410
rect 15822 8334 15940 8342
rect 14010 8059 14044 8183
rect 14367 8182 15739 8229
rect 14367 8169 14433 8182
rect 14367 8135 14383 8169
rect 14417 8135 14433 8169
rect 14367 8119 14433 8135
rect 14871 8059 14905 8182
rect 14004 8047 14050 8059
rect 14004 7871 14010 8047
rect 14044 7871 14050 8047
rect 14004 7859 14050 7871
rect 14122 8047 14246 8059
rect 14122 7871 14128 8047
rect 14162 7871 14206 8047
rect 14122 7859 14206 7871
rect 14128 7492 14162 7859
rect 14200 7671 14206 7859
rect 14240 7671 14246 8047
rect 14200 7659 14246 7671
rect 14318 8047 14364 8059
rect 14318 7671 14324 8047
rect 14358 7671 14364 8047
rect 14318 7659 14364 7671
rect 14436 8047 14482 8059
rect 14436 7671 14442 8047
rect 14476 7671 14482 8047
rect 14436 7659 14482 7671
rect 14554 8047 14600 8059
rect 14554 7671 14560 8047
rect 14594 7671 14600 8047
rect 14554 7659 14600 7671
rect 14672 8047 14792 8059
rect 14672 7671 14678 8047
rect 14712 7871 14752 8047
rect 14786 7871 14792 8047
rect 14712 7859 14792 7871
rect 14864 8047 14910 8059
rect 14864 7871 14870 8047
rect 14904 7871 14910 8047
rect 14864 7859 14910 7871
rect 14712 7671 14718 7859
rect 14672 7659 14718 7671
rect 14442 7586 14476 7659
rect 14425 7570 14491 7586
rect 14425 7536 14441 7570
rect 14475 7536 14491 7570
rect 14425 7520 14491 7536
rect 14752 7492 14786 7859
rect 14128 7440 14786 7492
rect 14396 7418 14488 7440
rect 14396 7366 14410 7418
rect 14476 7366 14488 7418
rect 14396 7362 14488 7366
rect 7987 7322 9594 7323
rect 3003 6285 3067 6890
rect 3273 6737 3283 6751
rect 3241 6731 3283 6737
rect 3359 6737 3369 6751
rect 3359 6731 3399 6737
rect 3241 6695 3277 6731
rect 3373 6695 3399 6731
rect 3241 6677 3283 6695
rect 3359 6677 3399 6695
rect 3241 6637 3399 6677
rect 3241 6591 3523 6637
rect 3123 6545 3169 6557
rect 3123 6369 3129 6545
rect 3163 6369 3169 6545
rect 3123 6367 3169 6369
rect 3121 6285 3169 6367
rect 3241 6545 3287 6591
rect 3241 6369 3247 6545
rect 3281 6369 3287 6545
rect 3241 6357 3287 6369
rect 3359 6545 3405 6557
rect 3359 6369 3365 6545
rect 3399 6369 3405 6545
rect 3359 6357 3405 6369
rect 3477 6545 3523 6591
rect 3477 6369 3483 6545
rect 3517 6369 3523 6545
rect 3477 6357 3523 6369
rect 3003 6221 3173 6285
rect 3743 6282 3807 7278
rect 6499 7274 9594 7322
rect 9622 7274 12736 7323
rect 15892 7320 15940 8334
rect 16285 8230 16320 8500
rect 17734 8410 17826 8418
rect 17734 8345 17746 8410
rect 17814 8345 17826 8410
rect 17734 8333 17826 8345
rect 16285 8183 17189 8230
rect 18848 8229 18883 8739
rect 18966 8694 19142 8702
rect 18958 8626 18968 8694
rect 19025 8626 19142 8694
rect 18966 8618 19142 8626
rect 19271 8634 19342 9814
rect 20676 9572 20686 9632
rect 20766 9572 20776 9632
rect 20676 9532 20776 9572
rect 19770 9475 21573 9532
rect 19770 9188 19807 9475
rect 20364 9388 20398 9475
rect 21539 9388 21573 9475
rect 19885 9376 19931 9388
rect 19412 9176 19458 9188
rect 19412 9000 19418 9176
rect 19452 9000 19458 9176
rect 19412 8988 19458 9000
rect 19530 9176 19576 9188
rect 19530 9000 19536 9176
rect 19570 9000 19576 9176
rect 19530 8988 19576 9000
rect 19648 9176 19694 9188
rect 19648 9000 19654 9176
rect 19688 9000 19694 9176
rect 19648 8988 19694 9000
rect 19766 9176 19812 9188
rect 19766 9000 19772 9176
rect 19806 9000 19812 9176
rect 19766 8988 19812 9000
rect 19885 9000 19891 9376
rect 19925 9000 19931 9376
rect 19885 8988 19931 9000
rect 20003 9376 20049 9388
rect 20003 9000 20009 9376
rect 20043 9000 20049 9376
rect 20003 8988 20049 9000
rect 20121 9376 20167 9388
rect 20121 9000 20127 9376
rect 20161 9000 20167 9376
rect 20121 8988 20167 9000
rect 20239 9376 20285 9388
rect 20239 9000 20245 9376
rect 20279 9000 20285 9376
rect 20239 8988 20285 9000
rect 20358 9376 20404 9388
rect 20358 9000 20364 9376
rect 20398 9000 20404 9376
rect 20358 8988 20404 9000
rect 20476 9376 20522 9388
rect 20476 9000 20482 9376
rect 20516 9000 20522 9376
rect 20476 8988 20522 9000
rect 20594 9376 20640 9388
rect 20594 9000 20600 9376
rect 20634 9000 20640 9376
rect 20594 8988 20640 9000
rect 20712 9376 20758 9388
rect 20712 9000 20718 9376
rect 20752 9000 20758 9376
rect 20712 8988 20758 9000
rect 20830 9376 20876 9388
rect 20830 9000 20836 9376
rect 20870 9000 20876 9376
rect 20830 8988 20876 9000
rect 20948 9376 20994 9388
rect 20948 9000 20954 9376
rect 20988 9000 20994 9376
rect 20948 8988 20994 9000
rect 21066 9376 21112 9388
rect 21066 9000 21072 9376
rect 21106 9000 21112 9376
rect 21066 8988 21112 9000
rect 21179 9376 21225 9388
rect 21179 9000 21185 9376
rect 21219 9000 21225 9376
rect 21179 8988 21225 9000
rect 21297 9376 21343 9388
rect 21297 9000 21303 9376
rect 21337 9000 21343 9376
rect 21297 8988 21343 9000
rect 21415 9376 21461 9388
rect 21415 9000 21421 9376
rect 21455 9000 21461 9376
rect 21415 8988 21461 9000
rect 21533 9376 21579 9388
rect 21533 9000 21539 9376
rect 21573 9188 21579 9376
rect 21573 9176 21666 9188
rect 21573 9000 21626 9176
rect 21660 9000 21666 9176
rect 21533 8988 21666 9000
rect 21738 9176 21784 9188
rect 21738 9000 21744 9176
rect 21778 9000 21784 9176
rect 21738 8988 21784 9000
rect 21856 9176 21902 9188
rect 21856 9000 21862 9176
rect 21896 9000 21902 9176
rect 21856 8988 21902 9000
rect 21974 9176 22020 9188
rect 21974 9000 21980 9176
rect 22014 9000 22020 9176
rect 21974 8988 22020 9000
rect 19417 8634 19452 8988
rect 19891 8904 19925 8988
rect 21072 8904 21106 8988
rect 19891 8862 21106 8904
rect 19891 8842 19925 8862
rect 19568 8826 19925 8842
rect 19568 8792 19584 8826
rect 19618 8792 19925 8826
rect 21980 8802 22015 8988
rect 19568 8776 19925 8792
rect 20878 8785 22015 8802
rect 20878 8751 20894 8785
rect 20928 8751 22015 8785
rect 20878 8735 22015 8751
rect 18966 8578 19037 8586
rect 18958 8510 18968 8578
rect 19025 8510 19037 8578
rect 18966 8502 19037 8510
rect 19271 8488 19452 8634
rect 20748 8689 20840 8699
rect 20748 8627 20758 8689
rect 20828 8627 20840 8689
rect 20748 8614 20840 8627
rect 21833 8689 21925 8702
rect 21833 8626 21842 8689
rect 21913 8626 21925 8689
rect 21833 8617 21925 8626
rect 20528 8572 20593 8575
rect 20524 8569 20593 8572
rect 20518 8509 20528 8569
rect 20587 8509 20593 8569
rect 20524 8505 20593 8509
rect 20528 8503 20593 8505
rect 18966 8410 19142 8418
rect 18958 8342 18968 8410
rect 19025 8342 19142 8410
rect 18966 8334 19142 8342
rect 17154 8059 17188 8183
rect 17511 8182 18883 8229
rect 17511 8169 17577 8182
rect 17511 8135 17527 8169
rect 17561 8135 17577 8169
rect 17511 8119 17577 8135
rect 18015 8059 18049 8182
rect 17148 8047 17194 8059
rect 17148 7871 17154 8047
rect 17188 7871 17194 8047
rect 17148 7859 17194 7871
rect 17266 8047 17390 8059
rect 17266 7871 17272 8047
rect 17306 7871 17350 8047
rect 17266 7859 17350 7871
rect 17272 7492 17306 7859
rect 17344 7671 17350 7859
rect 17384 7671 17390 8047
rect 17344 7659 17390 7671
rect 17462 8047 17508 8059
rect 17462 7671 17468 8047
rect 17502 7671 17508 8047
rect 17462 7659 17508 7671
rect 17580 8047 17626 8059
rect 17580 7671 17586 8047
rect 17620 7671 17626 8047
rect 17580 7659 17626 7671
rect 17698 8047 17744 8059
rect 17698 7671 17704 8047
rect 17738 7671 17744 8047
rect 17698 7659 17744 7671
rect 17816 8047 17936 8059
rect 17816 7671 17822 8047
rect 17856 7871 17896 8047
rect 17930 7871 17936 8047
rect 17856 7859 17936 7871
rect 18008 8047 18054 8059
rect 18008 7871 18014 8047
rect 18048 7871 18054 8047
rect 18008 7859 18054 7871
rect 17856 7671 17862 7859
rect 17816 7659 17862 7671
rect 17586 7586 17620 7659
rect 17569 7570 17635 7586
rect 17569 7536 17585 7570
rect 17619 7536 17635 7570
rect 17569 7520 17635 7536
rect 17896 7492 17930 7859
rect 17272 7440 17930 7492
rect 17540 7418 17632 7440
rect 17540 7366 17554 7418
rect 17620 7366 17632 7418
rect 17540 7362 17632 7366
rect 6499 7250 6547 7274
rect 4486 7202 6547 7250
rect 9622 7244 9670 7274
rect 12768 7272 15940 7320
rect 12768 7246 12816 7272
rect 4011 6737 4021 6751
rect 3979 6731 4021 6737
rect 4097 6737 4107 6751
rect 4097 6731 4137 6737
rect 3979 6695 4015 6731
rect 4111 6695 4137 6731
rect 3979 6677 4021 6695
rect 4097 6677 4137 6695
rect 3979 6637 4137 6677
rect 3979 6591 4261 6637
rect 3861 6545 3907 6557
rect 3861 6369 3867 6545
rect 3901 6369 3907 6545
rect 3861 6367 3907 6369
rect 3859 6282 3907 6367
rect 3979 6545 4025 6591
rect 3979 6369 3985 6545
rect 4019 6369 4025 6545
rect 3979 6357 4025 6369
rect 4097 6545 4143 6557
rect 4097 6369 4103 6545
rect 4137 6369 4143 6545
rect 4097 6357 4143 6369
rect 4215 6545 4261 6591
rect 4215 6369 4221 6545
rect 4255 6369 4261 6545
rect 4215 6357 4261 6369
rect 4486 6285 4550 7202
rect 6619 7196 9670 7244
rect 9698 7198 12816 7246
rect 19037 7244 19100 8334
rect 19417 8226 19452 8488
rect 20866 8406 20958 8414
rect 20866 8341 20878 8406
rect 20946 8341 20958 8406
rect 20866 8329 20958 8341
rect 19417 8179 20321 8226
rect 21980 8225 22015 8735
rect 22098 8690 22274 8698
rect 22090 8622 22100 8690
rect 22157 8622 22274 8690
rect 22414 8634 22486 9814
rect 23820 9572 23830 9632
rect 23910 9572 23920 9632
rect 23820 9532 23920 9572
rect 22914 9475 24717 9532
rect 22914 9188 22951 9475
rect 23508 9388 23542 9475
rect 24683 9388 24717 9475
rect 23029 9376 23075 9388
rect 22556 9176 22602 9188
rect 22556 9000 22562 9176
rect 22596 9000 22602 9176
rect 22556 8988 22602 9000
rect 22674 9176 22720 9188
rect 22674 9000 22680 9176
rect 22714 9000 22720 9176
rect 22674 8988 22720 9000
rect 22792 9176 22838 9188
rect 22792 9000 22798 9176
rect 22832 9000 22838 9176
rect 22792 8988 22838 9000
rect 22910 9176 22956 9188
rect 22910 9000 22916 9176
rect 22950 9000 22956 9176
rect 22910 8988 22956 9000
rect 23029 9000 23035 9376
rect 23069 9000 23075 9376
rect 23029 8988 23075 9000
rect 23147 9376 23193 9388
rect 23147 9000 23153 9376
rect 23187 9000 23193 9376
rect 23147 8988 23193 9000
rect 23265 9376 23311 9388
rect 23265 9000 23271 9376
rect 23305 9000 23311 9376
rect 23265 8988 23311 9000
rect 23383 9376 23429 9388
rect 23383 9000 23389 9376
rect 23423 9000 23429 9376
rect 23383 8988 23429 9000
rect 23502 9376 23548 9388
rect 23502 9000 23508 9376
rect 23542 9000 23548 9376
rect 23502 8988 23548 9000
rect 23620 9376 23666 9388
rect 23620 9000 23626 9376
rect 23660 9000 23666 9376
rect 23620 8988 23666 9000
rect 23738 9376 23784 9388
rect 23738 9000 23744 9376
rect 23778 9000 23784 9376
rect 23738 8988 23784 9000
rect 23856 9376 23902 9388
rect 23856 9000 23862 9376
rect 23896 9000 23902 9376
rect 23856 8988 23902 9000
rect 23974 9376 24020 9388
rect 23974 9000 23980 9376
rect 24014 9000 24020 9376
rect 23974 8988 24020 9000
rect 24092 9376 24138 9388
rect 24092 9000 24098 9376
rect 24132 9000 24138 9376
rect 24092 8988 24138 9000
rect 24210 9376 24256 9388
rect 24210 9000 24216 9376
rect 24250 9000 24256 9376
rect 24210 8988 24256 9000
rect 24323 9376 24369 9388
rect 24323 9000 24329 9376
rect 24363 9000 24369 9376
rect 24323 8988 24369 9000
rect 24441 9376 24487 9388
rect 24441 9000 24447 9376
rect 24481 9000 24487 9376
rect 24441 8988 24487 9000
rect 24559 9376 24605 9388
rect 24559 9000 24565 9376
rect 24599 9000 24605 9376
rect 24559 8988 24605 9000
rect 24677 9376 24723 9388
rect 24677 9000 24683 9376
rect 24717 9188 24723 9376
rect 24717 9176 24810 9188
rect 24717 9000 24770 9176
rect 24804 9000 24810 9176
rect 24677 8988 24810 9000
rect 24882 9176 24928 9188
rect 24882 9000 24888 9176
rect 24922 9000 24928 9176
rect 24882 8988 24928 9000
rect 25000 9176 25046 9188
rect 25000 9000 25006 9176
rect 25040 9000 25046 9176
rect 25000 8988 25046 9000
rect 25118 9176 25164 9188
rect 25118 9000 25124 9176
rect 25158 9000 25164 9176
rect 25118 8988 25164 9000
rect 22561 8634 22596 8988
rect 23035 8904 23069 8988
rect 24216 8904 24250 8988
rect 23035 8862 24250 8904
rect 23035 8842 23069 8862
rect 22712 8826 23069 8842
rect 22712 8792 22728 8826
rect 22762 8792 23069 8826
rect 25124 8802 25159 8988
rect 22712 8776 23069 8792
rect 24022 8785 25159 8802
rect 24022 8751 24038 8785
rect 24072 8751 25159 8785
rect 24022 8735 25159 8751
rect 22414 8626 22596 8634
rect 22098 8614 22274 8622
rect 22098 8574 22169 8582
rect 22090 8506 22100 8574
rect 22157 8506 22169 8574
rect 22098 8498 22169 8506
rect 22415 8488 22596 8626
rect 23892 8689 23984 8699
rect 23892 8627 23902 8689
rect 23972 8627 23984 8689
rect 23892 8614 23984 8627
rect 24977 8689 25069 8702
rect 24977 8626 24986 8689
rect 25057 8626 25069 8689
rect 24977 8617 25069 8626
rect 23672 8572 23737 8575
rect 23668 8569 23737 8572
rect 23662 8509 23672 8569
rect 23731 8509 23737 8569
rect 23668 8505 23737 8509
rect 23672 8503 23737 8505
rect 22098 8406 22232 8414
rect 22090 8338 22100 8406
rect 22157 8338 22232 8406
rect 22098 8330 22232 8338
rect 20286 8055 20320 8179
rect 20643 8178 22015 8225
rect 20643 8165 20709 8178
rect 20643 8131 20659 8165
rect 20693 8131 20709 8165
rect 20643 8115 20709 8131
rect 21147 8055 21181 8178
rect 20280 8043 20326 8055
rect 20280 7867 20286 8043
rect 20320 7867 20326 8043
rect 20280 7855 20326 7867
rect 20398 8043 20522 8055
rect 20398 7867 20404 8043
rect 20438 7867 20482 8043
rect 20398 7855 20482 7867
rect 20404 7488 20438 7855
rect 20476 7667 20482 7855
rect 20516 7667 20522 8043
rect 20476 7655 20522 7667
rect 20594 8043 20640 8055
rect 20594 7667 20600 8043
rect 20634 7667 20640 8043
rect 20594 7655 20640 7667
rect 20712 8043 20758 8055
rect 20712 7667 20718 8043
rect 20752 7667 20758 8043
rect 20712 7655 20758 7667
rect 20830 8043 20876 8055
rect 20830 7667 20836 8043
rect 20870 7667 20876 8043
rect 20830 7655 20876 7667
rect 20948 8043 21068 8055
rect 20948 7667 20954 8043
rect 20988 7867 21028 8043
rect 21062 7867 21068 8043
rect 20988 7855 21068 7867
rect 21140 8043 21186 8055
rect 21140 7867 21146 8043
rect 21180 7867 21186 8043
rect 21140 7855 21186 7867
rect 20988 7667 20994 7855
rect 20948 7655 20994 7667
rect 20718 7582 20752 7655
rect 20701 7566 20767 7582
rect 20701 7532 20717 7566
rect 20751 7532 20767 7566
rect 20701 7516 20767 7532
rect 21028 7488 21062 7855
rect 20404 7436 21062 7488
rect 20672 7414 20764 7436
rect 20672 7362 20686 7414
rect 20752 7362 20764 7414
rect 20672 7358 20764 7362
rect 6619 7172 6667 7196
rect 5219 7124 6667 7172
rect 9698 7168 9741 7198
rect 12844 7196 19100 7244
rect 12844 7170 12892 7196
rect 4749 6737 4759 6751
rect 4717 6731 4759 6737
rect 4835 6737 4845 6751
rect 4835 6731 4875 6737
rect 4717 6695 4753 6731
rect 4849 6695 4875 6731
rect 4717 6677 4759 6695
rect 4835 6677 4875 6695
rect 4717 6637 4875 6677
rect 4717 6591 4999 6637
rect 4599 6545 4645 6557
rect 4599 6369 4605 6545
rect 4639 6369 4645 6545
rect 4599 6367 4645 6369
rect 4597 6285 4645 6367
rect 4717 6545 4763 6591
rect 4717 6369 4723 6545
rect 4757 6369 4763 6545
rect 4717 6357 4763 6369
rect 4835 6545 4881 6557
rect 4835 6369 4841 6545
rect 4875 6369 4881 6545
rect 4835 6357 4881 6369
rect 4953 6545 4999 6591
rect 4953 6369 4959 6545
rect 4993 6369 4999 6545
rect 4953 6357 4999 6369
rect 5219 6285 5283 7124
rect 6695 7120 9741 7168
rect 9769 7122 12892 7170
rect 6695 7096 6743 7120
rect 5963 7048 6743 7096
rect 9769 7091 9817 7122
rect 5487 6737 5497 6751
rect 5455 6731 5497 6737
rect 5573 6737 5583 6751
rect 5573 6731 5613 6737
rect 5455 6695 5491 6731
rect 5587 6695 5613 6731
rect 5455 6677 5497 6695
rect 5573 6677 5613 6695
rect 5455 6637 5613 6677
rect 5455 6591 5737 6637
rect 5337 6545 5383 6557
rect 5337 6369 5343 6545
rect 5377 6369 5383 6545
rect 5337 6367 5383 6369
rect 5335 6285 5383 6367
rect 5455 6545 5501 6591
rect 5455 6369 5461 6545
rect 5495 6369 5501 6545
rect 5455 6357 5501 6369
rect 5573 6545 5619 6557
rect 5573 6369 5579 6545
rect 5613 6369 5619 6545
rect 5573 6357 5619 6369
rect 5691 6545 5737 6591
rect 5691 6369 5697 6545
rect 5731 6369 5737 6545
rect 5691 6357 5737 6369
rect 5963 6285 6027 7048
rect 6771 7043 9817 7091
rect 6771 6987 6819 7043
rect 22168 7008 22232 8330
rect 22561 8226 22596 8488
rect 24010 8406 24102 8414
rect 24010 8341 24022 8406
rect 24090 8341 24102 8406
rect 24010 8329 24102 8341
rect 22561 8179 23465 8226
rect 25124 8225 25159 8735
rect 25817 8698 25927 11029
rect 25242 8690 25927 8698
rect 25234 8622 25244 8690
rect 25301 8622 25927 8690
rect 25242 8614 25927 8622
rect 25242 8574 25317 8582
rect 25234 8506 25244 8574
rect 25301 8506 25317 8574
rect 25242 8498 25317 8506
rect 25242 8406 25376 8414
rect 25234 8338 25244 8406
rect 25301 8338 25376 8406
rect 25242 8330 25376 8338
rect 23430 8055 23464 8179
rect 23787 8178 25159 8225
rect 23787 8165 23853 8178
rect 23787 8131 23803 8165
rect 23837 8131 23853 8165
rect 23787 8115 23853 8131
rect 24291 8055 24325 8178
rect 23424 8043 23470 8055
rect 23424 7867 23430 8043
rect 23464 7867 23470 8043
rect 23424 7855 23470 7867
rect 23542 8043 23666 8055
rect 23542 7867 23548 8043
rect 23582 7867 23626 8043
rect 23542 7855 23626 7867
rect 23548 7488 23582 7855
rect 23620 7667 23626 7855
rect 23660 7667 23666 8043
rect 23620 7655 23666 7667
rect 23738 8043 23784 8055
rect 23738 7667 23744 8043
rect 23778 7667 23784 8043
rect 23738 7655 23784 7667
rect 23856 8043 23902 8055
rect 23856 7667 23862 8043
rect 23896 7667 23902 8043
rect 23856 7655 23902 7667
rect 23974 8043 24020 8055
rect 23974 7667 23980 8043
rect 24014 7667 24020 8043
rect 23974 7655 24020 7667
rect 24092 8043 24212 8055
rect 24092 7667 24098 8043
rect 24132 7867 24172 8043
rect 24206 7867 24212 8043
rect 24132 7855 24212 7867
rect 24284 8043 24330 8055
rect 24284 7867 24290 8043
rect 24324 7867 24330 8043
rect 24284 7855 24330 7867
rect 24132 7667 24138 7855
rect 24092 7655 24138 7667
rect 23862 7582 23896 7655
rect 23845 7566 23911 7582
rect 23845 7532 23861 7566
rect 23895 7532 23911 7566
rect 23845 7516 23911 7532
rect 24172 7488 24206 7855
rect 23548 7436 24206 7488
rect 23816 7414 23908 7436
rect 23816 7362 23830 7414
rect 23896 7362 23908 7414
rect 23816 7358 23908 7362
rect 6732 6959 6819 6987
rect 7457 6960 22232 7008
rect 6227 6737 6237 6751
rect 6195 6731 6237 6737
rect 6313 6737 6323 6751
rect 6313 6731 6353 6737
rect 6195 6695 6231 6731
rect 6327 6695 6353 6731
rect 6195 6677 6237 6695
rect 6313 6677 6353 6695
rect 6195 6637 6353 6677
rect 6195 6591 6477 6637
rect 6077 6545 6123 6557
rect 6077 6369 6083 6545
rect 6117 6369 6123 6545
rect 6077 6367 6123 6369
rect 6075 6285 6123 6367
rect 6195 6545 6241 6591
rect 6195 6369 6201 6545
rect 6235 6369 6241 6545
rect 6195 6357 6241 6369
rect 6313 6545 6359 6557
rect 6313 6369 6319 6545
rect 6353 6369 6359 6545
rect 6313 6357 6359 6369
rect 6431 6545 6477 6591
rect 6431 6369 6437 6545
rect 6471 6369 6477 6545
rect 6431 6357 6477 6369
rect 6732 6286 6780 6959
rect 6969 6737 6979 6751
rect 6937 6731 6979 6737
rect 7055 6737 7065 6751
rect 7055 6731 7095 6737
rect 6937 6695 6973 6731
rect 7069 6695 7095 6731
rect 6937 6677 6979 6695
rect 7055 6677 7095 6695
rect 6937 6637 7095 6677
rect 6937 6591 7219 6637
rect 6819 6547 6865 6559
rect 6819 6371 6825 6547
rect 6859 6371 6865 6547
rect 6819 6367 6865 6371
rect 6817 6286 6865 6367
rect 6937 6547 6983 6591
rect 6937 6371 6943 6547
rect 6977 6371 6983 6547
rect 6937 6359 6983 6371
rect 7055 6547 7101 6559
rect 7055 6371 7061 6547
rect 7095 6371 7101 6547
rect 7055 6359 7101 6371
rect 7173 6547 7219 6591
rect 7173 6371 7179 6547
rect 7213 6371 7219 6547
rect 7173 6359 7219 6371
rect 3481 6269 3531 6281
rect 3295 6263 3487 6269
rect 3295 6229 3307 6263
rect 3341 6229 3487 6263
rect 3295 6223 3487 6229
rect 3525 6223 3531 6269
rect 3121 6175 3169 6221
rect 3481 6211 3531 6223
rect 3743 6218 3914 6282
rect 4220 6269 4268 6281
rect 4033 6263 4226 6269
rect 4033 6229 4045 6263
rect 4079 6229 4226 6263
rect 4033 6223 4226 6229
rect 4262 6223 4268 6269
rect 3859 6175 3907 6218
rect 4220 6211 4268 6223
rect 4486 6221 4649 6285
rect 4771 6263 4853 6269
rect 4771 6229 4783 6263
rect 4817 6229 4853 6263
rect 4771 6223 4853 6229
rect 5219 6221 5387 6285
rect 5509 6263 5589 6269
rect 5509 6229 5521 6263
rect 5555 6229 5589 6263
rect 5509 6223 5589 6229
rect 5963 6221 6127 6285
rect 6249 6263 6329 6269
rect 6249 6229 6261 6263
rect 6295 6229 6329 6263
rect 6249 6223 6329 6229
rect 6732 6224 6869 6286
rect 7457 6284 7521 6960
rect 25312 6899 25376 8330
rect 8201 6851 25376 6899
rect 7707 6737 7717 6751
rect 7675 6731 7717 6737
rect 7793 6737 7803 6751
rect 7793 6731 7833 6737
rect 7675 6695 7711 6731
rect 7807 6695 7833 6731
rect 7675 6677 7717 6695
rect 7793 6677 7833 6695
rect 7675 6637 7833 6677
rect 7675 6591 7957 6637
rect 7557 6551 7603 6563
rect 7557 6375 7563 6551
rect 7597 6375 7603 6551
rect 7557 6367 7603 6375
rect 7555 6284 7603 6367
rect 7675 6551 7721 6591
rect 7675 6375 7681 6551
rect 7715 6375 7721 6551
rect 7675 6363 7721 6375
rect 7793 6551 7839 6563
rect 7793 6375 7799 6551
rect 7833 6375 7839 6551
rect 7793 6363 7839 6375
rect 7911 6551 7957 6591
rect 7911 6375 7917 6551
rect 7951 6375 7957 6551
rect 7911 6363 7957 6375
rect 6991 6263 7070 6269
rect 6991 6229 7003 6263
rect 7037 6229 7070 6263
rect 4597 6175 4645 6221
rect 5335 6175 5383 6221
rect 6075 6175 6123 6221
rect 6817 6175 6865 6224
rect 6991 6223 7070 6229
rect 7457 6220 7607 6284
rect 8201 6282 8265 6851
rect 8445 6739 8455 6753
rect 8413 6733 8455 6739
rect 8531 6739 8541 6753
rect 8531 6733 8571 6739
rect 8413 6697 8449 6733
rect 8545 6697 8571 6733
rect 8413 6679 8455 6697
rect 8531 6679 8571 6697
rect 8413 6639 8571 6679
rect 10051 6676 10061 6698
rect 10019 6644 10061 6676
rect 10115 6676 10125 6698
rect 10115 6644 10153 6676
rect 12119 6674 12129 6696
rect 8413 6593 8695 6639
rect 10019 6593 10153 6644
rect 12087 6642 12129 6674
rect 12183 6674 12193 6696
rect 14188 6676 14198 6698
rect 12183 6642 12221 6674
rect 8295 6547 8341 6559
rect 8295 6371 8301 6547
rect 8335 6371 8341 6547
rect 8295 6369 8341 6371
rect 8293 6282 8341 6369
rect 8413 6547 8459 6593
rect 8413 6371 8419 6547
rect 8453 6371 8459 6547
rect 8413 6359 8459 6371
rect 8531 6547 8577 6559
rect 8531 6371 8537 6547
rect 8571 6371 8577 6547
rect 8531 6359 8577 6371
rect 8649 6547 8695 6593
rect 8649 6371 8655 6547
rect 8689 6371 8695 6547
rect 8649 6359 8695 6371
rect 9351 6550 10824 6593
rect 12087 6591 12221 6642
rect 14156 6644 14198 6676
rect 14252 6676 14262 6698
rect 14252 6644 14290 6676
rect 16256 6674 16266 6696
rect 14156 6593 14290 6644
rect 16224 6642 16266 6674
rect 16320 6674 16330 6696
rect 18325 6674 18335 6696
rect 16320 6642 16358 6674
rect 7729 6263 7815 6269
rect 7729 6229 7741 6263
rect 7775 6229 7815 6263
rect 7729 6223 7815 6229
rect 8201 6221 8345 6282
rect 8467 6265 8544 6271
rect 8467 6231 8479 6265
rect 8513 6231 8544 6265
rect 9351 6247 9385 6550
rect 9716 6447 9750 6550
rect 9952 6447 9986 6550
rect 10188 6447 10222 6550
rect 10424 6447 10458 6550
rect 9710 6435 9756 6447
rect 8467 6225 8544 6231
rect 9227 6235 9273 6247
rect 7555 6175 7603 6220
rect 8293 6177 8341 6221
rect 3121 6163 3287 6175
rect 3121 6145 3247 6163
rect 3241 5987 3247 6145
rect 3281 5987 3287 6163
rect 3241 5975 3287 5987
rect 3359 6163 3405 6175
rect 3359 5987 3365 6163
rect 3399 5987 3405 6163
rect 3859 6163 4025 6175
rect 3859 6145 3985 6163
rect 3359 5869 3405 5987
rect 3979 5987 3985 6145
rect 4019 5987 4025 6163
rect 3979 5975 4025 5987
rect 4097 6163 4143 6175
rect 4097 5987 4103 6163
rect 4137 5987 4143 6163
rect 4597 6159 4763 6175
rect 4597 6145 4723 6159
rect 4097 5869 4143 5987
rect 4717 5983 4723 6145
rect 4757 5983 4763 6159
rect 4717 5971 4763 5983
rect 4835 6159 4881 6171
rect 4835 5983 4841 6159
rect 4875 5983 4881 6159
rect 5335 6159 5501 6175
rect 5335 6145 5461 6159
rect 4835 5869 4881 5983
rect 5455 5983 5461 6145
rect 5495 5983 5501 6159
rect 5455 5971 5501 5983
rect 5573 6159 5619 6171
rect 5573 5983 5579 6159
rect 5613 5983 5619 6159
rect 6075 6159 6241 6175
rect 6075 6145 6201 6159
rect 5573 5869 5619 5983
rect 6195 5983 6201 6145
rect 6235 5983 6241 6159
rect 6195 5971 6241 5983
rect 6313 6159 6359 6171
rect 6313 5983 6319 6159
rect 6353 5983 6359 6159
rect 6817 6159 6983 6175
rect 6817 6145 6943 6159
rect 6313 5869 6359 5983
rect 6937 5983 6943 6145
rect 6977 5983 6983 6159
rect 6937 5971 6983 5983
rect 7055 6159 7101 6171
rect 7055 5983 7061 6159
rect 7095 5983 7101 6159
rect 7555 6163 7721 6175
rect 7555 6145 7681 6163
rect 7055 5869 7101 5983
rect 7675 5987 7681 6145
rect 7715 5987 7721 6163
rect 7675 5975 7721 5987
rect 7793 6163 7839 6175
rect 7793 5987 7799 6163
rect 7833 5987 7839 6163
rect 8293 6161 8459 6177
rect 8293 6147 8419 6161
rect 7793 5869 7839 5987
rect 8413 5985 8419 6147
rect 8453 5985 8459 6161
rect 8413 5973 8459 5985
rect 8531 6161 8577 6173
rect 8531 5985 8537 6161
rect 8571 5985 8577 6161
rect 9227 6059 9233 6235
rect 9267 6059 9273 6235
rect 9227 6047 9273 6059
rect 9345 6235 9391 6247
rect 9345 6059 9351 6235
rect 9385 6059 9391 6235
rect 9345 6047 9391 6059
rect 9463 6235 9509 6247
rect 9463 6059 9469 6235
rect 9503 6059 9509 6235
rect 9463 6047 9509 6059
rect 9581 6235 9627 6247
rect 9710 6235 9716 6435
rect 9581 6059 9587 6235
rect 9621 6059 9716 6235
rect 9750 6059 9756 6435
rect 9581 6047 9627 6059
rect 9710 6047 9756 6059
rect 9828 6435 9874 6447
rect 9828 6059 9834 6435
rect 9868 6059 9874 6435
rect 9828 6047 9874 6059
rect 9946 6435 9992 6447
rect 9946 6059 9952 6435
rect 9986 6059 9992 6435
rect 9946 6047 9992 6059
rect 10064 6435 10110 6447
rect 10064 6059 10070 6435
rect 10104 6059 10110 6435
rect 10064 6047 10110 6059
rect 10182 6435 10228 6447
rect 10182 6059 10188 6435
rect 10222 6059 10228 6435
rect 10182 6047 10228 6059
rect 10300 6435 10346 6447
rect 10300 6059 10306 6435
rect 10340 6059 10346 6435
rect 10300 6047 10346 6059
rect 10418 6435 10464 6447
rect 10418 6059 10424 6435
rect 10458 6235 10464 6435
rect 10790 6247 10824 6550
rect 11419 6548 12892 6591
rect 10548 6235 10594 6247
rect 10458 6059 10554 6235
rect 10588 6059 10594 6235
rect 10418 6047 10464 6059
rect 10548 6047 10594 6059
rect 10666 6235 10712 6247
rect 10666 6059 10672 6235
rect 10706 6059 10712 6235
rect 10666 6047 10712 6059
rect 10784 6235 10830 6247
rect 10784 6059 10790 6235
rect 10824 6059 10830 6235
rect 10784 6047 10830 6059
rect 10902 6235 10948 6247
rect 11419 6245 11453 6548
rect 11784 6445 11818 6548
rect 12020 6445 12054 6548
rect 12256 6445 12290 6548
rect 12492 6445 12526 6548
rect 11778 6433 11824 6445
rect 10902 6059 10908 6235
rect 10942 6059 10948 6235
rect 10902 6047 10948 6059
rect 11295 6233 11341 6245
rect 11295 6057 11301 6233
rect 11335 6057 11341 6233
rect 8531 5871 8577 5985
rect 9233 6013 9267 6047
rect 9469 6013 9503 6047
rect 9233 5978 9503 6013
rect 10070 6013 10104 6047
rect 10306 6013 10340 6047
rect 10908 6013 10942 6047
rect 11295 6045 11341 6057
rect 11413 6233 11459 6245
rect 11413 6057 11419 6233
rect 11453 6057 11459 6233
rect 11413 6045 11459 6057
rect 11531 6233 11577 6245
rect 11531 6057 11537 6233
rect 11571 6057 11577 6233
rect 11531 6045 11577 6057
rect 11649 6233 11695 6245
rect 11778 6233 11784 6433
rect 11649 6057 11655 6233
rect 11689 6057 11784 6233
rect 11818 6057 11824 6433
rect 11649 6045 11695 6057
rect 11778 6045 11824 6057
rect 11896 6433 11942 6445
rect 11896 6057 11902 6433
rect 11936 6057 11942 6433
rect 11896 6045 11942 6057
rect 12014 6433 12060 6445
rect 12014 6057 12020 6433
rect 12054 6057 12060 6433
rect 12014 6045 12060 6057
rect 12132 6433 12178 6445
rect 12132 6057 12138 6433
rect 12172 6057 12178 6433
rect 12132 6045 12178 6057
rect 12250 6433 12296 6445
rect 12250 6057 12256 6433
rect 12290 6057 12296 6433
rect 12250 6045 12296 6057
rect 12368 6433 12414 6445
rect 12368 6057 12374 6433
rect 12408 6057 12414 6433
rect 12368 6045 12414 6057
rect 12486 6433 12532 6445
rect 12486 6057 12492 6433
rect 12526 6233 12532 6433
rect 12858 6245 12892 6548
rect 13488 6550 14961 6593
rect 16224 6591 16358 6642
rect 18293 6642 18335 6674
rect 18389 6674 18399 6696
rect 18389 6642 18427 6674
rect 20393 6672 20403 6694
rect 18293 6591 18427 6642
rect 20361 6640 20403 6672
rect 20457 6672 20467 6694
rect 22462 6674 22472 6696
rect 20457 6640 20495 6672
rect 13488 6247 13522 6550
rect 13853 6447 13887 6550
rect 14089 6447 14123 6550
rect 14325 6447 14359 6550
rect 14561 6447 14595 6550
rect 13847 6435 13893 6447
rect 12616 6233 12662 6245
rect 12526 6057 12622 6233
rect 12656 6057 12662 6233
rect 12486 6045 12532 6057
rect 12616 6045 12662 6057
rect 12734 6233 12780 6245
rect 12734 6057 12740 6233
rect 12774 6057 12780 6233
rect 12734 6045 12780 6057
rect 12852 6233 12898 6245
rect 12852 6057 12858 6233
rect 12892 6057 12898 6233
rect 12852 6045 12898 6057
rect 12970 6233 13016 6245
rect 12970 6057 12976 6233
rect 13010 6057 13016 6233
rect 12970 6045 13016 6057
rect 13364 6235 13410 6247
rect 13364 6059 13370 6235
rect 13404 6059 13410 6235
rect 13364 6047 13410 6059
rect 13482 6235 13528 6247
rect 13482 6059 13488 6235
rect 13522 6059 13528 6235
rect 13482 6047 13528 6059
rect 13600 6235 13646 6247
rect 13600 6059 13606 6235
rect 13640 6059 13646 6235
rect 13600 6047 13646 6059
rect 13718 6235 13764 6247
rect 13847 6235 13853 6435
rect 13718 6059 13724 6235
rect 13758 6059 13853 6235
rect 13887 6059 13893 6435
rect 13718 6047 13764 6059
rect 13847 6047 13893 6059
rect 13965 6435 14011 6447
rect 13965 6059 13971 6435
rect 14005 6059 14011 6435
rect 13965 6047 14011 6059
rect 14083 6435 14129 6447
rect 14083 6059 14089 6435
rect 14123 6059 14129 6435
rect 14083 6047 14129 6059
rect 14201 6435 14247 6447
rect 14201 6059 14207 6435
rect 14241 6059 14247 6435
rect 14201 6047 14247 6059
rect 14319 6435 14365 6447
rect 14319 6059 14325 6435
rect 14359 6059 14365 6435
rect 14319 6047 14365 6059
rect 14437 6435 14483 6447
rect 14437 6059 14443 6435
rect 14477 6059 14483 6435
rect 14437 6047 14483 6059
rect 14555 6435 14601 6447
rect 14555 6059 14561 6435
rect 14595 6235 14601 6435
rect 14927 6247 14961 6550
rect 15556 6548 17029 6591
rect 14685 6235 14731 6247
rect 14595 6059 14691 6235
rect 14725 6059 14731 6235
rect 14555 6047 14601 6059
rect 14685 6047 14731 6059
rect 14803 6235 14849 6247
rect 14803 6059 14809 6235
rect 14843 6059 14849 6235
rect 14803 6047 14849 6059
rect 14921 6235 14967 6247
rect 14921 6059 14927 6235
rect 14961 6059 14967 6235
rect 14921 6047 14967 6059
rect 15039 6235 15085 6247
rect 15556 6245 15590 6548
rect 15921 6445 15955 6548
rect 16157 6445 16191 6548
rect 16393 6445 16427 6548
rect 16629 6445 16663 6548
rect 15915 6433 15961 6445
rect 15039 6059 15045 6235
rect 15079 6059 15085 6235
rect 15039 6047 15085 6059
rect 15432 6233 15478 6245
rect 15432 6057 15438 6233
rect 15472 6057 15478 6233
rect 10070 5978 10340 6013
rect 10783 5978 10942 6013
rect 11301 6011 11335 6045
rect 11537 6011 11571 6045
rect 3323 5803 3333 5869
rect 3435 5803 3445 5869
rect 4061 5803 4071 5869
rect 4173 5803 4183 5869
rect 4799 5803 4809 5869
rect 4911 5803 4921 5869
rect 5537 5803 5547 5869
rect 5649 5803 5659 5869
rect 6277 5803 6287 5869
rect 6389 5803 6399 5869
rect 7019 5803 7029 5869
rect 7131 5803 7141 5869
rect 7757 5803 7767 5869
rect 7869 5803 7879 5869
rect 8495 5805 8505 5871
rect 8607 5805 8617 5871
rect 9189 5338 9315 5344
rect 9189 5236 9201 5338
rect 9303 5236 9315 5338
rect 9189 5230 9315 5236
rect 9367 5195 9401 5978
rect 10070 5916 10104 5978
rect 9469 5890 9547 5896
rect 9469 5836 9481 5890
rect 9535 5836 9547 5890
rect 9469 5830 9547 5836
rect 9773 5878 10515 5916
rect 9773 5754 9807 5878
rect 10009 5754 10043 5878
rect 10245 5754 10279 5878
rect 10481 5754 10515 5878
rect 9767 5742 9813 5754
rect 9767 5366 9773 5742
rect 9807 5366 9813 5742
rect 9767 5354 9813 5366
rect 9885 5742 9931 5754
rect 9885 5366 9891 5742
rect 9925 5366 9931 5742
rect 9885 5354 9931 5366
rect 10003 5742 10049 5754
rect 10003 5366 10009 5742
rect 10043 5366 10049 5742
rect 10003 5354 10049 5366
rect 10121 5742 10167 5754
rect 10121 5366 10127 5742
rect 10161 5366 10167 5742
rect 10121 5354 10167 5366
rect 10239 5742 10285 5754
rect 10239 5366 10245 5742
rect 10279 5366 10285 5742
rect 10239 5354 10285 5366
rect 10357 5742 10403 5754
rect 10357 5366 10363 5742
rect 10397 5366 10403 5742
rect 10357 5354 10403 5366
rect 10475 5742 10521 5754
rect 10475 5366 10481 5742
rect 10515 5366 10521 5742
rect 10475 5354 10521 5366
rect 9367 5194 9674 5195
rect 10783 5194 10817 5978
rect 11301 5976 11571 6011
rect 12138 6011 12172 6045
rect 12374 6011 12408 6045
rect 12976 6011 13010 6045
rect 12138 5976 12408 6011
rect 12851 5976 13010 6011
rect 13370 6013 13404 6047
rect 13606 6013 13640 6047
rect 13370 5978 13640 6013
rect 14207 6013 14241 6047
rect 14443 6013 14477 6047
rect 15045 6013 15079 6047
rect 15432 6045 15478 6057
rect 15550 6233 15596 6245
rect 15550 6057 15556 6233
rect 15590 6057 15596 6233
rect 15550 6045 15596 6057
rect 15668 6233 15714 6245
rect 15668 6057 15674 6233
rect 15708 6057 15714 6233
rect 15668 6045 15714 6057
rect 15786 6233 15832 6245
rect 15915 6233 15921 6433
rect 15786 6057 15792 6233
rect 15826 6057 15921 6233
rect 15955 6057 15961 6433
rect 15786 6045 15832 6057
rect 15915 6045 15961 6057
rect 16033 6433 16079 6445
rect 16033 6057 16039 6433
rect 16073 6057 16079 6433
rect 16033 6045 16079 6057
rect 16151 6433 16197 6445
rect 16151 6057 16157 6433
rect 16191 6057 16197 6433
rect 16151 6045 16197 6057
rect 16269 6433 16315 6445
rect 16269 6057 16275 6433
rect 16309 6057 16315 6433
rect 16269 6045 16315 6057
rect 16387 6433 16433 6445
rect 16387 6057 16393 6433
rect 16427 6057 16433 6433
rect 16387 6045 16433 6057
rect 16505 6433 16551 6445
rect 16505 6057 16511 6433
rect 16545 6057 16551 6433
rect 16505 6045 16551 6057
rect 16623 6433 16669 6445
rect 16623 6057 16629 6433
rect 16663 6233 16669 6433
rect 16995 6245 17029 6548
rect 17625 6548 19098 6591
rect 20361 6589 20495 6640
rect 22430 6642 22472 6674
rect 22526 6674 22536 6696
rect 22526 6642 22564 6674
rect 24530 6672 24540 6694
rect 22430 6591 22564 6642
rect 24498 6640 24540 6672
rect 24594 6672 24604 6694
rect 24594 6640 24632 6672
rect 17625 6245 17659 6548
rect 17990 6445 18024 6548
rect 18226 6445 18260 6548
rect 18462 6445 18496 6548
rect 18698 6445 18732 6548
rect 17984 6433 18030 6445
rect 16753 6233 16799 6245
rect 16663 6057 16759 6233
rect 16793 6057 16799 6233
rect 16623 6045 16669 6057
rect 16753 6045 16799 6057
rect 16871 6233 16917 6245
rect 16871 6057 16877 6233
rect 16911 6057 16917 6233
rect 16871 6045 16917 6057
rect 16989 6233 17035 6245
rect 16989 6057 16995 6233
rect 17029 6057 17035 6233
rect 16989 6045 17035 6057
rect 17107 6233 17153 6245
rect 17107 6057 17113 6233
rect 17147 6057 17153 6233
rect 17107 6045 17153 6057
rect 17501 6233 17547 6245
rect 17501 6057 17507 6233
rect 17541 6057 17547 6233
rect 17501 6045 17547 6057
rect 17619 6233 17665 6245
rect 17619 6057 17625 6233
rect 17659 6057 17665 6233
rect 17619 6045 17665 6057
rect 17737 6233 17783 6245
rect 17737 6057 17743 6233
rect 17777 6057 17783 6233
rect 17737 6045 17783 6057
rect 17855 6233 17901 6245
rect 17984 6233 17990 6433
rect 17855 6057 17861 6233
rect 17895 6057 17990 6233
rect 18024 6057 18030 6433
rect 17855 6045 17901 6057
rect 17984 6045 18030 6057
rect 18102 6433 18148 6445
rect 18102 6057 18108 6433
rect 18142 6057 18148 6433
rect 18102 6045 18148 6057
rect 18220 6433 18266 6445
rect 18220 6057 18226 6433
rect 18260 6057 18266 6433
rect 18220 6045 18266 6057
rect 18338 6433 18384 6445
rect 18338 6057 18344 6433
rect 18378 6057 18384 6433
rect 18338 6045 18384 6057
rect 18456 6433 18502 6445
rect 18456 6057 18462 6433
rect 18496 6057 18502 6433
rect 18456 6045 18502 6057
rect 18574 6433 18620 6445
rect 18574 6057 18580 6433
rect 18614 6057 18620 6433
rect 18574 6045 18620 6057
rect 18692 6433 18738 6445
rect 18692 6057 18698 6433
rect 18732 6233 18738 6433
rect 19064 6245 19098 6548
rect 19693 6546 21166 6589
rect 18822 6233 18868 6245
rect 18732 6057 18828 6233
rect 18862 6057 18868 6233
rect 18692 6045 18738 6057
rect 18822 6045 18868 6057
rect 18940 6233 18986 6245
rect 18940 6057 18946 6233
rect 18980 6057 18986 6233
rect 18940 6045 18986 6057
rect 19058 6233 19104 6245
rect 19058 6057 19064 6233
rect 19098 6057 19104 6233
rect 19058 6045 19104 6057
rect 19176 6233 19222 6245
rect 19693 6243 19727 6546
rect 20058 6443 20092 6546
rect 20294 6443 20328 6546
rect 20530 6443 20564 6546
rect 20766 6443 20800 6546
rect 20052 6431 20098 6443
rect 19176 6057 19182 6233
rect 19216 6057 19222 6233
rect 19176 6045 19222 6057
rect 19569 6231 19615 6243
rect 19569 6055 19575 6231
rect 19609 6055 19615 6231
rect 14207 5978 14477 6013
rect 14920 5978 15079 6013
rect 15438 6011 15472 6045
rect 15674 6011 15708 6045
rect 10847 5830 10857 5896
rect 10923 5830 10997 5896
rect 10930 5706 10994 5707
rect 10857 5700 10994 5706
rect 10857 5640 10869 5700
rect 10935 5640 10994 5700
rect 10857 5634 10994 5640
rect 9367 5189 9787 5194
rect 10501 5189 10817 5194
rect 9367 5178 9854 5189
rect 9367 5151 9803 5178
rect 9367 5150 9674 5151
rect 9367 5022 9401 5150
rect 9787 5144 9803 5151
rect 9837 5144 9854 5178
rect 9787 5138 9854 5144
rect 10434 5178 10817 5189
rect 10434 5144 10451 5178
rect 10485 5151 10817 5178
rect 10485 5144 10501 5151
rect 10434 5138 10501 5144
rect 9507 5110 9563 5122
rect 10620 5111 10676 5123
rect 10620 5110 10636 5111
rect 9507 5076 9513 5110
rect 9547 5095 10117 5110
rect 9547 5076 10067 5095
rect 9507 5061 10067 5076
rect 10101 5061 10117 5095
rect 9507 5060 9563 5061
rect 10050 5051 10117 5061
rect 10169 5094 10636 5110
rect 10169 5060 10185 5094
rect 10219 5077 10636 5094
rect 10670 5077 10676 5111
rect 10219 5061 10676 5077
rect 10219 5060 10235 5061
rect 10169 5053 10235 5060
rect 10783 5022 10817 5151
rect 9361 5010 9407 5022
rect 9361 4834 9367 5010
rect 9401 4834 9407 5010
rect 9361 4822 9407 4834
rect 9479 5010 9525 5022
rect 9479 4834 9485 5010
rect 9519 4834 9525 5010
rect 9479 4822 9525 4834
rect 9885 5010 9931 5022
rect 453 4635 590 4650
rect 453 4566 483 4635
rect 563 4566 590 4635
rect 233 4483 369 4496
rect 233 4405 257 4483
rect 352 4405 369 4483
rect -19 4287 108 4302
rect -19 4213 3 4287
rect 84 4213 108 4287
rect -19 4171 108 4213
rect -809 4079 108 4171
rect -809 4078 98 4079
rect -2003 3349 -1993 3408
rect -1872 3349 -1862 3408
rect -1530 3110 -1520 3173
rect -1404 3110 -1394 3173
rect -1268 2993 -1258 3060
rect -1137 2993 -1127 3060
rect -1059 2863 -1049 2945
rect -925 2863 -915 2945
rect -809 -604 -669 4078
rect -574 3954 -434 3955
rect 233 3954 369 4405
rect -574 3861 369 3954
rect -574 -317 -434 3861
rect 453 3773 590 4566
rect 9486 4528 9519 4822
rect 9885 4634 9891 5010
rect 9925 4634 9931 5010
rect 9885 4622 9931 4634
rect 10003 5010 10049 5022
rect 10003 4634 10009 5010
rect 10043 4634 10049 5010
rect 10003 4622 10049 4634
rect 10121 5010 10167 5022
rect 10121 4634 10127 5010
rect 10161 4634 10167 5010
rect 10121 4622 10167 4634
rect 10239 5010 10285 5022
rect 10239 4634 10245 5010
rect 10279 4634 10285 5010
rect 10239 4622 10285 4634
rect 10357 5010 10403 5022
rect 10357 4634 10363 5010
rect 10397 4634 10403 5010
rect 10659 5010 10705 5022
rect 10659 4834 10665 5010
rect 10699 4834 10705 5010
rect 10659 4822 10705 4834
rect 10777 5010 10823 5022
rect 10777 4834 10783 5010
rect 10817 4834 10823 5010
rect 10777 4822 10823 4834
rect 10357 4622 10403 4634
rect 10009 4528 10043 4622
rect 10666 4528 10700 4822
rect 9486 4496 10700 4528
rect 10075 4474 10207 4496
rect 10075 4416 10111 4474
rect 10173 4416 10207 4474
rect 10075 4411 10207 4416
rect -310 3666 590 3773
rect -310 3665 512 3666
rect -574 -479 -550 -317
rect -446 -479 -434 -317
rect -309 -155 -142 3665
rect 10930 3415 10994 5634
rect 11257 5336 11383 5342
rect 11257 5234 11269 5336
rect 11371 5234 11383 5336
rect 11257 5228 11383 5234
rect 11435 5193 11469 5976
rect 12138 5914 12172 5976
rect 11537 5888 11615 5894
rect 11537 5834 11549 5888
rect 11603 5834 11615 5888
rect 11537 5828 11615 5834
rect 11841 5876 12583 5914
rect 11841 5752 11875 5876
rect 12077 5752 12111 5876
rect 12313 5752 12347 5876
rect 12549 5752 12583 5876
rect 11835 5740 11881 5752
rect 11835 5364 11841 5740
rect 11875 5364 11881 5740
rect 11835 5352 11881 5364
rect 11953 5740 11999 5752
rect 11953 5364 11959 5740
rect 11993 5364 11999 5740
rect 11953 5352 11999 5364
rect 12071 5740 12117 5752
rect 12071 5364 12077 5740
rect 12111 5364 12117 5740
rect 12071 5352 12117 5364
rect 12189 5740 12235 5752
rect 12189 5364 12195 5740
rect 12229 5364 12235 5740
rect 12189 5352 12235 5364
rect 12307 5740 12353 5752
rect 12307 5364 12313 5740
rect 12347 5364 12353 5740
rect 12307 5352 12353 5364
rect 12425 5740 12471 5752
rect 12425 5364 12431 5740
rect 12465 5364 12471 5740
rect 12425 5352 12471 5364
rect 12543 5740 12589 5752
rect 12543 5364 12549 5740
rect 12583 5364 12589 5740
rect 12543 5352 12589 5364
rect 11435 5192 11742 5193
rect 12851 5192 12885 5976
rect 12915 5828 12925 5894
rect 12991 5828 13065 5894
rect 12925 5698 13065 5704
rect 12925 5638 12937 5698
rect 13003 5638 13065 5698
rect 12925 5632 13065 5638
rect 11435 5187 11855 5192
rect 12569 5187 12885 5192
rect 11435 5176 11922 5187
rect 11435 5149 11871 5176
rect 11435 5148 11742 5149
rect 11435 5020 11469 5148
rect 11855 5142 11871 5149
rect 11905 5142 11922 5176
rect 11855 5136 11922 5142
rect 12502 5176 12885 5187
rect 12502 5142 12519 5176
rect 12553 5149 12885 5176
rect 12553 5142 12569 5149
rect 12502 5136 12569 5142
rect 11575 5108 11631 5120
rect 12688 5109 12744 5121
rect 12688 5108 12704 5109
rect 11575 5074 11581 5108
rect 11615 5093 12185 5108
rect 11615 5074 12135 5093
rect 11575 5059 12135 5074
rect 12169 5059 12185 5093
rect 11575 5058 11631 5059
rect 12118 5049 12185 5059
rect 12237 5092 12704 5108
rect 12237 5058 12253 5092
rect 12287 5075 12704 5092
rect 12738 5075 12744 5109
rect 12287 5059 12744 5075
rect 12287 5058 12303 5059
rect 12237 5051 12303 5058
rect 12851 5020 12885 5149
rect 11429 5008 11475 5020
rect 11429 4832 11435 5008
rect 11469 4832 11475 5008
rect 11429 4820 11475 4832
rect 11547 5008 11593 5020
rect 11547 4832 11553 5008
rect 11587 4832 11593 5008
rect 11547 4820 11593 4832
rect 11953 5008 11999 5020
rect 11554 4526 11587 4820
rect 11953 4632 11959 5008
rect 11993 4632 11999 5008
rect 11953 4620 11999 4632
rect 12071 5008 12117 5020
rect 12071 4632 12077 5008
rect 12111 4632 12117 5008
rect 12071 4620 12117 4632
rect 12189 5008 12235 5020
rect 12189 4632 12195 5008
rect 12229 4632 12235 5008
rect 12189 4620 12235 4632
rect 12307 5008 12353 5020
rect 12307 4632 12313 5008
rect 12347 4632 12353 5008
rect 12307 4620 12353 4632
rect 12425 5008 12471 5020
rect 12425 4632 12431 5008
rect 12465 4632 12471 5008
rect 12727 5008 12773 5020
rect 12727 4832 12733 5008
rect 12767 4832 12773 5008
rect 12727 4820 12773 4832
rect 12845 5008 12891 5020
rect 12845 4832 12851 5008
rect 12885 4832 12891 5008
rect 12845 4820 12891 4832
rect 12425 4620 12471 4632
rect 12077 4526 12111 4620
rect 12734 4526 12768 4820
rect 11554 4494 12768 4526
rect 12143 4472 12275 4494
rect 12143 4414 12179 4472
rect 12241 4414 12275 4472
rect 12143 4409 12275 4414
rect 13001 3503 13065 5632
rect 13326 5338 13452 5344
rect 13326 5236 13338 5338
rect 13440 5236 13452 5338
rect 13326 5230 13452 5236
rect 13504 5195 13538 5978
rect 14207 5916 14241 5978
rect 13606 5890 13684 5896
rect 13606 5836 13618 5890
rect 13672 5836 13684 5890
rect 13606 5830 13684 5836
rect 13910 5878 14652 5916
rect 13910 5754 13944 5878
rect 14146 5754 14180 5878
rect 14382 5754 14416 5878
rect 14618 5754 14652 5878
rect 13904 5742 13950 5754
rect 13904 5366 13910 5742
rect 13944 5366 13950 5742
rect 13904 5354 13950 5366
rect 14022 5742 14068 5754
rect 14022 5366 14028 5742
rect 14062 5366 14068 5742
rect 14022 5354 14068 5366
rect 14140 5742 14186 5754
rect 14140 5366 14146 5742
rect 14180 5366 14186 5742
rect 14140 5354 14186 5366
rect 14258 5742 14304 5754
rect 14258 5366 14264 5742
rect 14298 5366 14304 5742
rect 14258 5354 14304 5366
rect 14376 5742 14422 5754
rect 14376 5366 14382 5742
rect 14416 5366 14422 5742
rect 14376 5354 14422 5366
rect 14494 5742 14540 5754
rect 14494 5366 14500 5742
rect 14534 5366 14540 5742
rect 14494 5354 14540 5366
rect 14612 5742 14658 5754
rect 14612 5366 14618 5742
rect 14652 5366 14658 5742
rect 14612 5354 14658 5366
rect 13504 5194 13811 5195
rect 14920 5194 14954 5978
rect 15438 5976 15708 6011
rect 16275 6011 16309 6045
rect 16511 6011 16545 6045
rect 17113 6011 17147 6045
rect 16275 5976 16545 6011
rect 16988 5976 17147 6011
rect 17507 6011 17541 6045
rect 17743 6011 17777 6045
rect 17507 5976 17777 6011
rect 18344 6011 18378 6045
rect 18580 6011 18614 6045
rect 19182 6011 19216 6045
rect 19569 6043 19615 6055
rect 19687 6231 19733 6243
rect 19687 6055 19693 6231
rect 19727 6055 19733 6231
rect 19687 6043 19733 6055
rect 19805 6231 19851 6243
rect 19805 6055 19811 6231
rect 19845 6055 19851 6231
rect 19805 6043 19851 6055
rect 19923 6231 19969 6243
rect 20052 6231 20058 6431
rect 19923 6055 19929 6231
rect 19963 6055 20058 6231
rect 20092 6055 20098 6431
rect 19923 6043 19969 6055
rect 20052 6043 20098 6055
rect 20170 6431 20216 6443
rect 20170 6055 20176 6431
rect 20210 6055 20216 6431
rect 20170 6043 20216 6055
rect 20288 6431 20334 6443
rect 20288 6055 20294 6431
rect 20328 6055 20334 6431
rect 20288 6043 20334 6055
rect 20406 6431 20452 6443
rect 20406 6055 20412 6431
rect 20446 6055 20452 6431
rect 20406 6043 20452 6055
rect 20524 6431 20570 6443
rect 20524 6055 20530 6431
rect 20564 6055 20570 6431
rect 20524 6043 20570 6055
rect 20642 6431 20688 6443
rect 20642 6055 20648 6431
rect 20682 6055 20688 6431
rect 20642 6043 20688 6055
rect 20760 6431 20806 6443
rect 20760 6055 20766 6431
rect 20800 6231 20806 6431
rect 21132 6243 21166 6546
rect 21762 6548 23235 6591
rect 24498 6589 24632 6640
rect 21762 6245 21796 6548
rect 22127 6445 22161 6548
rect 22363 6445 22397 6548
rect 22599 6445 22633 6548
rect 22835 6445 22869 6548
rect 22121 6433 22167 6445
rect 20890 6231 20936 6243
rect 20800 6055 20896 6231
rect 20930 6055 20936 6231
rect 20760 6043 20806 6055
rect 20890 6043 20936 6055
rect 21008 6231 21054 6243
rect 21008 6055 21014 6231
rect 21048 6055 21054 6231
rect 21008 6043 21054 6055
rect 21126 6231 21172 6243
rect 21126 6055 21132 6231
rect 21166 6055 21172 6231
rect 21126 6043 21172 6055
rect 21244 6231 21290 6243
rect 21244 6055 21250 6231
rect 21284 6055 21290 6231
rect 21244 6043 21290 6055
rect 21638 6233 21684 6245
rect 21638 6057 21644 6233
rect 21678 6057 21684 6233
rect 21638 6045 21684 6057
rect 21756 6233 21802 6245
rect 21756 6057 21762 6233
rect 21796 6057 21802 6233
rect 21756 6045 21802 6057
rect 21874 6233 21920 6245
rect 21874 6057 21880 6233
rect 21914 6057 21920 6233
rect 21874 6045 21920 6057
rect 21992 6233 22038 6245
rect 22121 6233 22127 6433
rect 21992 6057 21998 6233
rect 22032 6057 22127 6233
rect 22161 6057 22167 6433
rect 21992 6045 22038 6057
rect 22121 6045 22167 6057
rect 22239 6433 22285 6445
rect 22239 6057 22245 6433
rect 22279 6057 22285 6433
rect 22239 6045 22285 6057
rect 22357 6433 22403 6445
rect 22357 6057 22363 6433
rect 22397 6057 22403 6433
rect 22357 6045 22403 6057
rect 22475 6433 22521 6445
rect 22475 6057 22481 6433
rect 22515 6057 22521 6433
rect 22475 6045 22521 6057
rect 22593 6433 22639 6445
rect 22593 6057 22599 6433
rect 22633 6057 22639 6433
rect 22593 6045 22639 6057
rect 22711 6433 22757 6445
rect 22711 6057 22717 6433
rect 22751 6057 22757 6433
rect 22711 6045 22757 6057
rect 22829 6433 22875 6445
rect 22829 6057 22835 6433
rect 22869 6233 22875 6433
rect 23201 6245 23235 6548
rect 23830 6546 25303 6589
rect 22959 6233 23005 6245
rect 22869 6057 22965 6233
rect 22999 6057 23005 6233
rect 22829 6045 22875 6057
rect 22959 6045 23005 6057
rect 23077 6233 23123 6245
rect 23077 6057 23083 6233
rect 23117 6057 23123 6233
rect 23077 6045 23123 6057
rect 23195 6233 23241 6245
rect 23195 6057 23201 6233
rect 23235 6057 23241 6233
rect 23195 6045 23241 6057
rect 23313 6233 23359 6245
rect 23830 6243 23864 6546
rect 24195 6443 24229 6546
rect 24431 6443 24465 6546
rect 24667 6443 24701 6546
rect 24903 6443 24937 6546
rect 24189 6431 24235 6443
rect 23313 6057 23319 6233
rect 23353 6057 23359 6233
rect 23313 6045 23359 6057
rect 23706 6231 23752 6243
rect 23706 6055 23712 6231
rect 23746 6055 23752 6231
rect 18344 5976 18614 6011
rect 19057 5976 19216 6011
rect 19575 6009 19609 6043
rect 19811 6009 19845 6043
rect 14984 5830 14994 5896
rect 15060 5830 15134 5896
rect 14994 5700 15164 5706
rect 14994 5640 15006 5700
rect 15072 5640 15164 5700
rect 14994 5634 15164 5640
rect 13504 5189 13924 5194
rect 14638 5189 14954 5194
rect 13504 5178 13991 5189
rect 13504 5151 13940 5178
rect 13504 5150 13811 5151
rect 13504 5022 13538 5150
rect 13924 5144 13940 5151
rect 13974 5144 13991 5178
rect 13924 5138 13991 5144
rect 14571 5178 14954 5189
rect 14571 5144 14588 5178
rect 14622 5151 14954 5178
rect 14622 5144 14638 5151
rect 14571 5138 14638 5144
rect 13644 5110 13700 5122
rect 14757 5111 14813 5123
rect 14757 5110 14773 5111
rect 13644 5076 13650 5110
rect 13684 5095 14254 5110
rect 13684 5076 14204 5095
rect 13644 5061 14204 5076
rect 14238 5061 14254 5095
rect 13644 5060 13700 5061
rect 14187 5051 14254 5061
rect 14306 5094 14773 5110
rect 14306 5060 14322 5094
rect 14356 5077 14773 5094
rect 14807 5077 14813 5111
rect 14356 5061 14813 5077
rect 14356 5060 14372 5061
rect 14306 5053 14372 5060
rect 14920 5022 14954 5151
rect 13498 5010 13544 5022
rect 13498 4834 13504 5010
rect 13538 4834 13544 5010
rect 13498 4822 13544 4834
rect 13616 5010 13662 5022
rect 13616 4834 13622 5010
rect 13656 4834 13662 5010
rect 13616 4822 13662 4834
rect 14022 5010 14068 5022
rect 13623 4528 13656 4822
rect 14022 4634 14028 5010
rect 14062 4634 14068 5010
rect 14022 4622 14068 4634
rect 14140 5010 14186 5022
rect 14140 4634 14146 5010
rect 14180 4634 14186 5010
rect 14140 4622 14186 4634
rect 14258 5010 14304 5022
rect 14258 4634 14264 5010
rect 14298 4634 14304 5010
rect 14258 4622 14304 4634
rect 14376 5010 14422 5022
rect 14376 4634 14382 5010
rect 14416 4634 14422 5010
rect 14376 4622 14422 4634
rect 14494 5010 14540 5022
rect 14494 4634 14500 5010
rect 14534 4634 14540 5010
rect 14796 5010 14842 5022
rect 14796 4834 14802 5010
rect 14836 4834 14842 5010
rect 14796 4822 14842 4834
rect 14914 5010 14960 5022
rect 14914 4834 14920 5010
rect 14954 4834 14960 5010
rect 14914 4822 14960 4834
rect 14494 4622 14540 4634
rect 14146 4528 14180 4622
rect 14803 4528 14837 4822
rect 13623 4496 14837 4528
rect 14212 4474 14344 4496
rect 14212 4416 14248 4474
rect 14310 4416 14344 4474
rect 14212 4411 14344 4416
rect 15100 3642 15164 5634
rect 15394 5336 15520 5342
rect 15394 5234 15406 5336
rect 15508 5234 15520 5336
rect 15394 5228 15520 5234
rect 15572 5193 15606 5976
rect 16275 5914 16309 5976
rect 15674 5888 15752 5894
rect 15674 5834 15686 5888
rect 15740 5834 15752 5888
rect 15674 5828 15752 5834
rect 15978 5876 16720 5914
rect 15978 5752 16012 5876
rect 16214 5752 16248 5876
rect 16450 5752 16484 5876
rect 16686 5752 16720 5876
rect 15972 5740 16018 5752
rect 15972 5364 15978 5740
rect 16012 5364 16018 5740
rect 15972 5352 16018 5364
rect 16090 5740 16136 5752
rect 16090 5364 16096 5740
rect 16130 5364 16136 5740
rect 16090 5352 16136 5364
rect 16208 5740 16254 5752
rect 16208 5364 16214 5740
rect 16248 5364 16254 5740
rect 16208 5352 16254 5364
rect 16326 5740 16372 5752
rect 16326 5364 16332 5740
rect 16366 5364 16372 5740
rect 16326 5352 16372 5364
rect 16444 5740 16490 5752
rect 16444 5364 16450 5740
rect 16484 5364 16490 5740
rect 16444 5352 16490 5364
rect 16562 5740 16608 5752
rect 16562 5364 16568 5740
rect 16602 5364 16608 5740
rect 16562 5352 16608 5364
rect 16680 5740 16726 5752
rect 16680 5364 16686 5740
rect 16720 5364 16726 5740
rect 16680 5352 16726 5364
rect 15572 5192 15879 5193
rect 16988 5192 17022 5976
rect 17052 5828 17062 5894
rect 17128 5828 17202 5894
rect 17062 5698 17238 5704
rect 17062 5638 17074 5698
rect 17140 5638 17238 5698
rect 17062 5632 17238 5638
rect 15572 5187 15992 5192
rect 16706 5187 17022 5192
rect 15572 5176 16059 5187
rect 15572 5149 16008 5176
rect 15572 5148 15879 5149
rect 15572 5020 15606 5148
rect 15992 5142 16008 5149
rect 16042 5142 16059 5176
rect 15992 5136 16059 5142
rect 16639 5176 17022 5187
rect 16639 5142 16656 5176
rect 16690 5149 17022 5176
rect 16690 5142 16706 5149
rect 16639 5136 16706 5142
rect 15712 5108 15768 5120
rect 16825 5109 16881 5121
rect 16825 5108 16841 5109
rect 15712 5074 15718 5108
rect 15752 5093 16322 5108
rect 15752 5074 16272 5093
rect 15712 5059 16272 5074
rect 16306 5059 16322 5093
rect 15712 5058 15768 5059
rect 16255 5049 16322 5059
rect 16374 5092 16841 5108
rect 16374 5058 16390 5092
rect 16424 5075 16841 5092
rect 16875 5075 16881 5109
rect 16424 5059 16881 5075
rect 16424 5058 16440 5059
rect 16374 5051 16440 5058
rect 16988 5020 17022 5149
rect 15566 5008 15612 5020
rect 15566 4832 15572 5008
rect 15606 4832 15612 5008
rect 15566 4820 15612 4832
rect 15684 5008 15730 5020
rect 15684 4832 15690 5008
rect 15724 4832 15730 5008
rect 15684 4820 15730 4832
rect 16090 5008 16136 5020
rect 15691 4526 15724 4820
rect 16090 4632 16096 5008
rect 16130 4632 16136 5008
rect 16090 4620 16136 4632
rect 16208 5008 16254 5020
rect 16208 4632 16214 5008
rect 16248 4632 16254 5008
rect 16208 4620 16254 4632
rect 16326 5008 16372 5020
rect 16326 4632 16332 5008
rect 16366 4632 16372 5008
rect 16326 4620 16372 4632
rect 16444 5008 16490 5020
rect 16444 4632 16450 5008
rect 16484 4632 16490 5008
rect 16444 4620 16490 4632
rect 16562 5008 16608 5020
rect 16562 4632 16568 5008
rect 16602 4632 16608 5008
rect 16864 5008 16910 5020
rect 16864 4832 16870 5008
rect 16904 4832 16910 5008
rect 16864 4820 16910 4832
rect 16982 5008 17028 5020
rect 16982 4832 16988 5008
rect 17022 4832 17028 5008
rect 16982 4820 17028 4832
rect 16562 4620 16608 4632
rect 16214 4526 16248 4620
rect 16871 4526 16905 4820
rect 15691 4494 16905 4526
rect 16280 4472 16412 4494
rect 16280 4414 16316 4472
rect 16378 4414 16412 4472
rect 16280 4409 16412 4414
rect 17174 3749 17238 5632
rect 17463 5336 17589 5342
rect 17463 5234 17475 5336
rect 17577 5234 17589 5336
rect 17463 5228 17589 5234
rect 17641 5193 17675 5976
rect 18344 5914 18378 5976
rect 17743 5888 17821 5894
rect 17743 5834 17755 5888
rect 17809 5834 17821 5888
rect 17743 5828 17821 5834
rect 18047 5876 18789 5914
rect 18047 5752 18081 5876
rect 18283 5752 18317 5876
rect 18519 5752 18553 5876
rect 18755 5752 18789 5876
rect 18041 5740 18087 5752
rect 18041 5364 18047 5740
rect 18081 5364 18087 5740
rect 18041 5352 18087 5364
rect 18159 5740 18205 5752
rect 18159 5364 18165 5740
rect 18199 5364 18205 5740
rect 18159 5352 18205 5364
rect 18277 5740 18323 5752
rect 18277 5364 18283 5740
rect 18317 5364 18323 5740
rect 18277 5352 18323 5364
rect 18395 5740 18441 5752
rect 18395 5364 18401 5740
rect 18435 5364 18441 5740
rect 18395 5352 18441 5364
rect 18513 5740 18559 5752
rect 18513 5364 18519 5740
rect 18553 5364 18559 5740
rect 18513 5352 18559 5364
rect 18631 5740 18677 5752
rect 18631 5364 18637 5740
rect 18671 5364 18677 5740
rect 18631 5352 18677 5364
rect 18749 5740 18795 5752
rect 18749 5364 18755 5740
rect 18789 5364 18795 5740
rect 18749 5352 18795 5364
rect 17641 5192 17948 5193
rect 19057 5192 19091 5976
rect 19575 5974 19845 6009
rect 20412 6009 20446 6043
rect 20648 6009 20682 6043
rect 21250 6009 21284 6043
rect 20412 5974 20682 6009
rect 21125 5974 21284 6009
rect 21644 6011 21678 6045
rect 21880 6011 21914 6045
rect 21644 5976 21914 6011
rect 22481 6011 22515 6045
rect 22717 6011 22751 6045
rect 23319 6011 23353 6045
rect 23706 6043 23752 6055
rect 23824 6231 23870 6243
rect 23824 6055 23830 6231
rect 23864 6055 23870 6231
rect 23824 6043 23870 6055
rect 23942 6231 23988 6243
rect 23942 6055 23948 6231
rect 23982 6055 23988 6231
rect 23942 6043 23988 6055
rect 24060 6231 24106 6243
rect 24189 6231 24195 6431
rect 24060 6055 24066 6231
rect 24100 6055 24195 6231
rect 24229 6055 24235 6431
rect 24060 6043 24106 6055
rect 24189 6043 24235 6055
rect 24307 6431 24353 6443
rect 24307 6055 24313 6431
rect 24347 6055 24353 6431
rect 24307 6043 24353 6055
rect 24425 6431 24471 6443
rect 24425 6055 24431 6431
rect 24465 6055 24471 6431
rect 24425 6043 24471 6055
rect 24543 6431 24589 6443
rect 24543 6055 24549 6431
rect 24583 6055 24589 6431
rect 24543 6043 24589 6055
rect 24661 6431 24707 6443
rect 24661 6055 24667 6431
rect 24701 6055 24707 6431
rect 24661 6043 24707 6055
rect 24779 6431 24825 6443
rect 24779 6055 24785 6431
rect 24819 6055 24825 6431
rect 24779 6043 24825 6055
rect 24897 6431 24943 6443
rect 24897 6055 24903 6431
rect 24937 6231 24943 6431
rect 25269 6243 25303 6546
rect 25027 6231 25073 6243
rect 24937 6055 25033 6231
rect 25067 6055 25073 6231
rect 24897 6043 24943 6055
rect 25027 6043 25073 6055
rect 25145 6231 25191 6243
rect 25145 6055 25151 6231
rect 25185 6055 25191 6231
rect 25145 6043 25191 6055
rect 25263 6231 25309 6243
rect 25263 6055 25269 6231
rect 25303 6055 25309 6231
rect 25263 6043 25309 6055
rect 25381 6231 25427 6243
rect 25381 6055 25387 6231
rect 25421 6055 25427 6231
rect 25381 6043 25427 6055
rect 22481 5976 22751 6011
rect 23194 5976 23353 6011
rect 23712 6009 23746 6043
rect 23948 6009 23982 6043
rect 19121 5828 19131 5894
rect 19197 5828 19271 5894
rect 19131 5698 19328 5704
rect 19131 5638 19143 5698
rect 19209 5638 19328 5698
rect 19131 5632 19328 5638
rect 17641 5187 18061 5192
rect 18775 5187 19091 5192
rect 17641 5176 18128 5187
rect 17641 5149 18077 5176
rect 17641 5148 17948 5149
rect 17641 5020 17675 5148
rect 18061 5142 18077 5149
rect 18111 5142 18128 5176
rect 18061 5136 18128 5142
rect 18708 5176 19091 5187
rect 18708 5142 18725 5176
rect 18759 5149 19091 5176
rect 18759 5142 18775 5149
rect 18708 5136 18775 5142
rect 17781 5108 17837 5120
rect 18894 5109 18950 5121
rect 18894 5108 18910 5109
rect 17781 5074 17787 5108
rect 17821 5093 18391 5108
rect 17821 5074 18341 5093
rect 17781 5059 18341 5074
rect 18375 5059 18391 5093
rect 17781 5058 17837 5059
rect 18324 5049 18391 5059
rect 18443 5092 18910 5108
rect 18443 5058 18459 5092
rect 18493 5075 18910 5092
rect 18944 5075 18950 5109
rect 18493 5059 18950 5075
rect 18493 5058 18509 5059
rect 18443 5051 18509 5058
rect 19057 5020 19091 5149
rect 17635 5008 17681 5020
rect 17635 4832 17641 5008
rect 17675 4832 17681 5008
rect 17635 4820 17681 4832
rect 17753 5008 17799 5020
rect 17753 4832 17759 5008
rect 17793 4832 17799 5008
rect 17753 4820 17799 4832
rect 18159 5008 18205 5020
rect 17760 4526 17793 4820
rect 18159 4632 18165 5008
rect 18199 4632 18205 5008
rect 18159 4620 18205 4632
rect 18277 5008 18323 5020
rect 18277 4632 18283 5008
rect 18317 4632 18323 5008
rect 18277 4620 18323 4632
rect 18395 5008 18441 5020
rect 18395 4632 18401 5008
rect 18435 4632 18441 5008
rect 18395 4620 18441 4632
rect 18513 5008 18559 5020
rect 18513 4632 18519 5008
rect 18553 4632 18559 5008
rect 18513 4620 18559 4632
rect 18631 5008 18677 5020
rect 18631 4632 18637 5008
rect 18671 4632 18677 5008
rect 18933 5008 18979 5020
rect 18933 4832 18939 5008
rect 18973 4832 18979 5008
rect 18933 4820 18979 4832
rect 19051 5008 19097 5020
rect 19051 4832 19057 5008
rect 19091 4832 19097 5008
rect 19051 4820 19097 4832
rect 18631 4620 18677 4632
rect 18283 4526 18317 4620
rect 18940 4526 18974 4820
rect 17760 4494 18974 4526
rect 18349 4472 18481 4494
rect 18349 4414 18385 4472
rect 18447 4414 18481 4472
rect 18349 4409 18481 4414
rect 19264 3849 19328 5632
rect 19531 5334 19657 5340
rect 19531 5232 19543 5334
rect 19645 5232 19657 5334
rect 19531 5226 19657 5232
rect 19709 5191 19743 5974
rect 20412 5912 20446 5974
rect 19811 5886 19889 5892
rect 19811 5832 19823 5886
rect 19877 5832 19889 5886
rect 19811 5826 19889 5832
rect 20115 5874 20857 5912
rect 20115 5750 20149 5874
rect 20351 5750 20385 5874
rect 20587 5750 20621 5874
rect 20823 5750 20857 5874
rect 20109 5738 20155 5750
rect 20109 5362 20115 5738
rect 20149 5362 20155 5738
rect 20109 5350 20155 5362
rect 20227 5738 20273 5750
rect 20227 5362 20233 5738
rect 20267 5362 20273 5738
rect 20227 5350 20273 5362
rect 20345 5738 20391 5750
rect 20345 5362 20351 5738
rect 20385 5362 20391 5738
rect 20345 5350 20391 5362
rect 20463 5738 20509 5750
rect 20463 5362 20469 5738
rect 20503 5362 20509 5738
rect 20463 5350 20509 5362
rect 20581 5738 20627 5750
rect 20581 5362 20587 5738
rect 20621 5362 20627 5738
rect 20581 5350 20627 5362
rect 20699 5738 20745 5750
rect 20699 5362 20705 5738
rect 20739 5362 20745 5738
rect 20699 5350 20745 5362
rect 20817 5738 20863 5750
rect 20817 5362 20823 5738
rect 20857 5362 20863 5738
rect 20817 5350 20863 5362
rect 19709 5190 20016 5191
rect 21125 5190 21159 5974
rect 21189 5826 21199 5892
rect 21265 5826 21339 5892
rect 21199 5696 21374 5702
rect 21199 5636 21211 5696
rect 21277 5636 21374 5696
rect 21199 5630 21374 5636
rect 19709 5185 20129 5190
rect 20843 5185 21159 5190
rect 19709 5174 20196 5185
rect 19709 5147 20145 5174
rect 19709 5146 20016 5147
rect 19709 5018 19743 5146
rect 20129 5140 20145 5147
rect 20179 5140 20196 5174
rect 20129 5134 20196 5140
rect 20776 5174 21159 5185
rect 20776 5140 20793 5174
rect 20827 5147 21159 5174
rect 20827 5140 20843 5147
rect 20776 5134 20843 5140
rect 19849 5106 19905 5118
rect 20962 5107 21018 5119
rect 20962 5106 20978 5107
rect 19849 5072 19855 5106
rect 19889 5091 20459 5106
rect 19889 5072 20409 5091
rect 19849 5057 20409 5072
rect 20443 5057 20459 5091
rect 19849 5056 19905 5057
rect 20392 5047 20459 5057
rect 20511 5090 20978 5106
rect 20511 5056 20527 5090
rect 20561 5073 20978 5090
rect 21012 5073 21018 5107
rect 20561 5057 21018 5073
rect 20561 5056 20577 5057
rect 20511 5049 20577 5056
rect 21125 5018 21159 5147
rect 19703 5006 19749 5018
rect 19703 4830 19709 5006
rect 19743 4830 19749 5006
rect 19703 4818 19749 4830
rect 19821 5006 19867 5018
rect 19821 4830 19827 5006
rect 19861 4830 19867 5006
rect 19821 4818 19867 4830
rect 20227 5006 20273 5018
rect 19828 4524 19861 4818
rect 20227 4630 20233 5006
rect 20267 4630 20273 5006
rect 20227 4618 20273 4630
rect 20345 5006 20391 5018
rect 20345 4630 20351 5006
rect 20385 4630 20391 5006
rect 20345 4618 20391 4630
rect 20463 5006 20509 5018
rect 20463 4630 20469 5006
rect 20503 4630 20509 5006
rect 20463 4618 20509 4630
rect 20581 5006 20627 5018
rect 20581 4630 20587 5006
rect 20621 4630 20627 5006
rect 20581 4618 20627 4630
rect 20699 5006 20745 5018
rect 20699 4630 20705 5006
rect 20739 4630 20745 5006
rect 21001 5006 21047 5018
rect 21001 4830 21007 5006
rect 21041 4830 21047 5006
rect 21001 4818 21047 4830
rect 21119 5006 21165 5018
rect 21119 4830 21125 5006
rect 21159 4830 21165 5006
rect 21119 4818 21165 4830
rect 20699 4618 20745 4630
rect 20351 4524 20385 4618
rect 21008 4524 21042 4818
rect 19828 4492 21042 4524
rect 20417 4470 20549 4492
rect 20417 4412 20453 4470
rect 20515 4412 20549 4470
rect 20417 4407 20549 4412
rect 21310 3958 21374 5630
rect 21600 5336 21726 5342
rect 21600 5234 21612 5336
rect 21714 5234 21726 5336
rect 21600 5228 21726 5234
rect 21778 5193 21812 5976
rect 22481 5914 22515 5976
rect 21880 5888 21958 5894
rect 21880 5834 21892 5888
rect 21946 5834 21958 5888
rect 21880 5828 21958 5834
rect 22184 5876 22926 5914
rect 22184 5752 22218 5876
rect 22420 5752 22454 5876
rect 22656 5752 22690 5876
rect 22892 5752 22926 5876
rect 22178 5740 22224 5752
rect 22178 5364 22184 5740
rect 22218 5364 22224 5740
rect 22178 5352 22224 5364
rect 22296 5740 22342 5752
rect 22296 5364 22302 5740
rect 22336 5364 22342 5740
rect 22296 5352 22342 5364
rect 22414 5740 22460 5752
rect 22414 5364 22420 5740
rect 22454 5364 22460 5740
rect 22414 5352 22460 5364
rect 22532 5740 22578 5752
rect 22532 5364 22538 5740
rect 22572 5364 22578 5740
rect 22532 5352 22578 5364
rect 22650 5740 22696 5752
rect 22650 5364 22656 5740
rect 22690 5364 22696 5740
rect 22650 5352 22696 5364
rect 22768 5740 22814 5752
rect 22768 5364 22774 5740
rect 22808 5364 22814 5740
rect 22768 5352 22814 5364
rect 22886 5740 22932 5752
rect 22886 5364 22892 5740
rect 22926 5364 22932 5740
rect 22886 5352 22932 5364
rect 21778 5192 22085 5193
rect 23194 5192 23228 5976
rect 23712 5974 23982 6009
rect 24549 6009 24583 6043
rect 24785 6009 24819 6043
rect 25387 6009 25421 6043
rect 24549 5974 24819 6009
rect 25262 5974 25421 6009
rect 23258 5828 23268 5894
rect 23334 5828 23408 5894
rect 23268 5698 23408 5704
rect 23268 5638 23280 5698
rect 23346 5638 23408 5698
rect 23268 5632 23408 5638
rect 21778 5187 22198 5192
rect 22912 5187 23228 5192
rect 21778 5176 22265 5187
rect 21778 5149 22214 5176
rect 21778 5148 22085 5149
rect 21778 5020 21812 5148
rect 22198 5142 22214 5149
rect 22248 5142 22265 5176
rect 22198 5136 22265 5142
rect 22845 5176 23228 5187
rect 22845 5142 22862 5176
rect 22896 5149 23228 5176
rect 22896 5142 22912 5149
rect 22845 5136 22912 5142
rect 21918 5108 21974 5120
rect 23031 5109 23087 5121
rect 23031 5108 23047 5109
rect 21918 5074 21924 5108
rect 21958 5093 22528 5108
rect 21958 5074 22478 5093
rect 21918 5059 22478 5074
rect 22512 5059 22528 5093
rect 21918 5058 21974 5059
rect 22461 5049 22528 5059
rect 22580 5092 23047 5108
rect 22580 5058 22596 5092
rect 22630 5075 23047 5092
rect 23081 5075 23087 5109
rect 22630 5059 23087 5075
rect 22630 5058 22646 5059
rect 22580 5051 22646 5058
rect 23194 5020 23228 5149
rect 21772 5008 21818 5020
rect 21772 4832 21778 5008
rect 21812 4832 21818 5008
rect 21772 4820 21818 4832
rect 21890 5008 21936 5020
rect 21890 4832 21896 5008
rect 21930 4832 21936 5008
rect 21890 4820 21936 4832
rect 22296 5008 22342 5020
rect 21897 4526 21930 4820
rect 22296 4632 22302 5008
rect 22336 4632 22342 5008
rect 22296 4620 22342 4632
rect 22414 5008 22460 5020
rect 22414 4632 22420 5008
rect 22454 4632 22460 5008
rect 22414 4620 22460 4632
rect 22532 5008 22578 5020
rect 22532 4632 22538 5008
rect 22572 4632 22578 5008
rect 22532 4620 22578 4632
rect 22650 5008 22696 5020
rect 22650 4632 22656 5008
rect 22690 4632 22696 5008
rect 22650 4620 22696 4632
rect 22768 5008 22814 5020
rect 22768 4632 22774 5008
rect 22808 4632 22814 5008
rect 23070 5008 23116 5020
rect 23070 4832 23076 5008
rect 23110 4832 23116 5008
rect 23070 4820 23116 4832
rect 23188 5008 23234 5020
rect 23188 4832 23194 5008
rect 23228 4832 23234 5008
rect 23188 4820 23234 4832
rect 22768 4620 22814 4632
rect 22420 4526 22454 4620
rect 23077 4526 23111 4820
rect 21897 4494 23111 4526
rect 22486 4472 22618 4494
rect 22486 4414 22522 4472
rect 22584 4414 22618 4472
rect 22486 4409 22618 4414
rect 23344 4269 23408 5632
rect 23668 5334 23794 5340
rect 23668 5232 23680 5334
rect 23782 5232 23794 5334
rect 23668 5226 23794 5232
rect 23846 5191 23880 5974
rect 24549 5912 24583 5974
rect 23948 5886 24026 5892
rect 23948 5832 23960 5886
rect 24014 5832 24026 5886
rect 23948 5826 24026 5832
rect 24252 5874 24994 5912
rect 24252 5750 24286 5874
rect 24488 5750 24522 5874
rect 24724 5750 24758 5874
rect 24960 5750 24994 5874
rect 24246 5738 24292 5750
rect 24246 5362 24252 5738
rect 24286 5362 24292 5738
rect 24246 5350 24292 5362
rect 24364 5738 24410 5750
rect 24364 5362 24370 5738
rect 24404 5362 24410 5738
rect 24364 5350 24410 5362
rect 24482 5738 24528 5750
rect 24482 5362 24488 5738
rect 24522 5362 24528 5738
rect 24482 5350 24528 5362
rect 24600 5738 24646 5750
rect 24600 5362 24606 5738
rect 24640 5362 24646 5738
rect 24600 5350 24646 5362
rect 24718 5738 24764 5750
rect 24718 5362 24724 5738
rect 24758 5362 24764 5738
rect 24718 5350 24764 5362
rect 24836 5738 24882 5750
rect 24836 5362 24842 5738
rect 24876 5362 24882 5738
rect 24836 5350 24882 5362
rect 24954 5738 25000 5750
rect 24954 5362 24960 5738
rect 24994 5362 25000 5738
rect 24954 5350 25000 5362
rect 23846 5190 24153 5191
rect 25262 5190 25296 5974
rect 26047 5901 26111 17348
rect 26277 6085 26341 17543
rect 26464 6248 26538 17720
rect 26662 6398 26741 17909
rect 26849 6555 26913 18093
rect 27062 6863 27142 18278
rect 27316 7157 27395 18464
rect 28449 18446 28525 19292
rect 29568 18953 32760 19043
rect 27819 18436 28525 18446
rect 27819 18374 27829 18436
rect 27889 18374 28525 18436
rect 27819 18363 28525 18374
rect 28555 18854 32760 18953
rect 27819 18362 28438 18363
rect 28555 18256 28625 18854
rect 29565 18491 32623 18603
rect 27825 18252 28625 18256
rect 28662 18424 32623 18491
rect 28662 18420 29654 18424
rect 27825 18246 28564 18252
rect 27825 18184 27836 18246
rect 27896 18184 28564 18246
rect 27825 18177 28564 18184
rect 28616 18177 28626 18252
rect 27825 18170 28625 18177
rect 28662 18074 28732 18420
rect 29562 18080 32485 18178
rect 27826 18064 28732 18074
rect 27826 17995 27836 18064
rect 27896 17995 28461 18064
rect 27826 17987 28461 17995
rect 28515 17987 28732 18064
rect 27826 17980 28732 17987
rect 28840 18003 32485 18080
rect 28840 17888 28922 18003
rect 27836 17877 28922 17888
rect 27836 17814 27848 17877
rect 27909 17876 28922 17877
rect 27909 17814 28360 17876
rect 27836 17806 28360 17814
rect 28414 17824 28922 17876
rect 28414 17806 28921 17824
rect 27836 17798 28921 17806
rect 29565 17702 32343 17759
rect 27840 17686 32343 17702
rect 27840 17614 27851 17686
rect 27922 17675 32343 17686
rect 27922 17614 28258 17675
rect 27840 17600 28258 17614
rect 28311 17600 32343 17675
rect 27840 17574 32343 17600
rect 27840 17573 29649 17574
rect 29562 17223 32190 17328
rect 27841 17216 32190 17223
rect 27841 17209 28157 17216
rect 27841 17154 27851 17209
rect 27905 17154 28157 17209
rect 27841 17152 28157 17154
rect 28211 17152 32190 17216
rect 27841 17144 32190 17152
rect 30536 16922 30624 16924
rect 29559 16820 30624 16922
rect 27791 16807 30624 16820
rect 27791 16801 28052 16807
rect 27791 16747 27801 16801
rect 27857 16747 28052 16801
rect 27791 16731 28052 16747
rect 28118 16731 30624 16807
rect 27791 16723 30624 16731
rect 30503 13175 30624 16723
rect 30154 13168 30354 13174
rect 30154 13134 30166 13168
rect 30342 13134 30423 13168
rect 30154 13128 30354 13134
rect 30154 13050 30354 13056
rect 29808 13016 30166 13050
rect 30342 13016 30354 13050
rect 29808 12684 29851 13016
rect 30154 13010 30354 13016
rect 30388 13043 30423 13134
rect 30505 13149 30624 13175
rect 30695 13161 30767 13174
rect 30571 13128 30624 13149
rect 30691 13097 30701 13161
rect 30762 13097 30772 13161
rect 30695 13095 30701 13097
rect 30761 13095 30767 13097
rect 30695 13083 30767 13095
rect 30505 13073 30571 13083
rect 31379 13043 31579 13049
rect 30388 13009 31391 13043
rect 31567 13009 31579 13043
rect 30154 12932 30354 12938
rect 30154 12898 30166 12932
rect 30342 12898 30354 12932
rect 30154 12892 30354 12898
rect 30154 12814 30354 12820
rect 30154 12780 30166 12814
rect 30342 12780 30354 12814
rect 30154 12774 30354 12780
rect 30166 12690 30342 12774
rect 30647 12741 31047 12747
rect 30485 12707 30659 12741
rect 31035 12707 31047 12741
rect 31207 12727 31250 13009
rect 31379 13003 31579 13009
rect 31379 12926 31579 12931
rect 31379 12925 31905 12926
rect 31278 12896 31340 12902
rect 31278 12862 31290 12896
rect 31324 12862 31340 12896
rect 31379 12891 31391 12925
rect 31567 12892 31905 12925
rect 31567 12891 31579 12892
rect 31379 12885 31579 12891
rect 31278 12846 31340 12862
rect 29954 12684 30354 12690
rect 29808 12650 29966 12684
rect 30342 12650 30354 12684
rect 29808 12448 29851 12650
rect 29954 12644 30354 12650
rect 29954 12566 30354 12572
rect 29954 12532 29966 12566
rect 30342 12532 30423 12566
rect 29954 12526 30354 12532
rect 29954 12448 30354 12454
rect 29808 12414 29966 12448
rect 30342 12414 30354 12448
rect 29808 12379 29851 12414
rect 29954 12408 30354 12414
rect 29725 12351 29851 12379
rect 29703 12341 29851 12351
rect 29757 12287 29851 12341
rect 29954 12330 30354 12336
rect 30388 12330 30423 12532
rect 30485 12505 30523 12707
rect 30647 12701 31047 12707
rect 31212 12711 31263 12727
rect 31212 12677 31223 12711
rect 31257 12677 31263 12711
rect 31212 12660 31263 12677
rect 30647 12623 31047 12629
rect 30647 12589 30659 12623
rect 31035 12589 31047 12623
rect 30647 12583 31047 12589
rect 30647 12505 31047 12511
rect 30485 12471 30659 12505
rect 31035 12471 31047 12505
rect 30485 12330 30523 12471
rect 30647 12465 31047 12471
rect 31291 12461 31340 12846
rect 31379 12623 31779 12629
rect 31379 12589 31391 12623
rect 31767 12589 31779 12623
rect 31379 12583 31779 12589
rect 31379 12505 31779 12511
rect 31379 12471 31391 12505
rect 31767 12471 31779 12505
rect 31379 12465 31779 12471
rect 31291 12445 31348 12461
rect 31291 12411 31307 12445
rect 31341 12411 31348 12445
rect 31291 12395 31348 12411
rect 31873 12433 31905 12892
rect 31873 12399 31990 12433
rect 30647 12387 31047 12393
rect 30647 12353 30659 12387
rect 31035 12353 31047 12387
rect 30647 12347 31047 12353
rect 31379 12387 31779 12393
rect 31379 12353 31391 12387
rect 31767 12353 31779 12387
rect 31379 12347 31779 12353
rect 29954 12296 29966 12330
rect 30342 12296 30523 12330
rect 29954 12290 30354 12296
rect 29703 12277 29851 12287
rect 29725 12245 29851 12277
rect 29808 12212 29851 12245
rect 30485 12269 30523 12296
rect 31291 12327 31350 12343
rect 31291 12293 31306 12327
rect 31340 12293 31350 12327
rect 31291 12276 31350 12293
rect 31873 12337 31927 12399
rect 31985 12337 31990 12399
rect 31873 12301 31990 12337
rect 30647 12269 31047 12275
rect 30485 12235 30659 12269
rect 31035 12235 31047 12269
rect 29954 12212 30354 12218
rect 29808 12178 29966 12212
rect 30342 12178 30354 12212
rect 29808 11976 29851 12178
rect 29954 12172 30354 12178
rect 29954 12094 30354 12100
rect 29954 12060 29966 12094
rect 30342 12060 30354 12094
rect 29954 12054 30354 12060
rect 30485 12033 30523 12235
rect 30647 12229 31047 12235
rect 30647 12151 31047 12157
rect 30647 12117 30659 12151
rect 31035 12117 31047 12151
rect 30647 12111 31047 12117
rect 31212 12063 31263 12080
rect 30647 12033 31047 12039
rect 30485 11999 30659 12033
rect 31035 11999 31047 12033
rect 31212 12029 31223 12063
rect 31257 12029 31263 12063
rect 31212 12013 31263 12029
rect 30647 11993 31047 11999
rect 29954 11976 30354 11982
rect 29808 11942 29966 11976
rect 30342 11942 30354 11976
rect 29808 11611 29851 11942
rect 29954 11936 30354 11942
rect 30166 11853 30342 11936
rect 31207 11900 31250 12013
rect 30154 11847 30354 11853
rect 30154 11813 30166 11847
rect 30342 11813 30354 11847
rect 30154 11807 30354 11813
rect 30505 11761 30571 11773
rect 30154 11729 30354 11735
rect 30154 11695 30166 11729
rect 30342 11695 30423 11729
rect 30505 11707 30511 11761
rect 30565 11707 30571 11761
rect 30505 11695 30571 11707
rect 30154 11689 30354 11695
rect 30388 11627 30423 11695
rect 31206 11627 31251 11900
rect 31291 11789 31340 12276
rect 31379 12269 31779 12275
rect 31873 12269 31905 12301
rect 31379 12235 31391 12269
rect 31767 12235 31905 12269
rect 31379 12229 31779 12235
rect 31379 12151 31779 12157
rect 31379 12117 31391 12151
rect 31767 12117 31779 12151
rect 31379 12111 31779 12117
rect 31279 11773 31341 11789
rect 31279 11739 31291 11773
rect 31325 11739 31341 11773
rect 31279 11733 31341 11739
rect 31379 11745 31579 11751
rect 31873 11745 31905 12235
rect 31379 11711 31391 11745
rect 31567 11712 31905 11745
rect 31567 11711 31579 11712
rect 31379 11705 31579 11711
rect 31379 11627 31579 11633
rect 30154 11611 30354 11617
rect 29808 11577 30166 11611
rect 30342 11577 30354 11611
rect 30154 11571 30354 11577
rect 30388 11593 31391 11627
rect 31567 11593 31579 11627
rect 30154 11493 30354 11499
rect 30388 11493 30423 11593
rect 31379 11587 31579 11593
rect 30154 11459 30166 11493
rect 30342 11459 30423 11493
rect 31057 11529 31171 11541
rect 30154 11453 30354 11459
rect 31057 11427 31063 11529
rect 31165 11427 31171 11529
rect 31057 11415 31171 11427
rect 32101 11264 32190 17144
rect 30503 11178 32190 11264
rect 30503 11108 30570 11178
rect 30152 11100 30352 11106
rect 30152 11066 30164 11100
rect 30340 11066 30421 11100
rect 30152 11060 30352 11066
rect 30152 10982 30352 10988
rect 29806 10948 30164 10982
rect 30340 10948 30352 10982
rect 29806 10616 29849 10948
rect 30152 10942 30352 10948
rect 30386 10975 30421 11066
rect 30503 11081 30569 11108
rect 30692 11093 30765 11106
rect 30692 11028 30699 11093
rect 30693 11027 30699 11028
rect 30759 11027 30765 11093
rect 30693 11015 30765 11027
rect 30503 11005 30569 11015
rect 31377 10975 31577 10981
rect 30386 10941 31389 10975
rect 31565 10941 31577 10975
rect 30152 10864 30352 10870
rect 30152 10830 30164 10864
rect 30340 10830 30352 10864
rect 30152 10824 30352 10830
rect 30152 10746 30352 10752
rect 30152 10712 30164 10746
rect 30340 10712 30352 10746
rect 30152 10706 30352 10712
rect 30164 10622 30340 10706
rect 30645 10673 31045 10679
rect 30483 10639 30657 10673
rect 31033 10639 31045 10673
rect 31205 10659 31248 10941
rect 31377 10935 31577 10941
rect 31377 10858 31577 10863
rect 31377 10857 31903 10858
rect 31276 10828 31338 10834
rect 31276 10794 31288 10828
rect 31322 10794 31338 10828
rect 31377 10823 31389 10857
rect 31565 10824 31903 10857
rect 31565 10823 31577 10824
rect 31377 10817 31577 10823
rect 31276 10778 31338 10794
rect 29952 10616 30352 10622
rect 29806 10582 29964 10616
rect 30340 10582 30352 10616
rect 29806 10380 29849 10582
rect 29952 10576 30352 10582
rect 29952 10498 30352 10504
rect 29952 10464 29964 10498
rect 30340 10464 30421 10498
rect 29952 10458 30352 10464
rect 29952 10380 30352 10386
rect 29806 10346 29964 10380
rect 30340 10346 30352 10380
rect 29806 10311 29849 10346
rect 29952 10340 30352 10346
rect 29723 10283 29849 10311
rect 29701 10273 29849 10283
rect 29755 10219 29849 10273
rect 29952 10262 30352 10268
rect 30386 10262 30421 10464
rect 30483 10437 30521 10639
rect 30645 10633 31045 10639
rect 31210 10643 31261 10659
rect 31210 10609 31221 10643
rect 31255 10609 31261 10643
rect 31210 10592 31261 10609
rect 30645 10555 31045 10561
rect 30645 10521 30657 10555
rect 31033 10521 31045 10555
rect 30645 10515 31045 10521
rect 30645 10437 31045 10443
rect 30483 10403 30657 10437
rect 31033 10403 31045 10437
rect 30483 10262 30521 10403
rect 30645 10397 31045 10403
rect 31289 10393 31338 10778
rect 31377 10555 31777 10561
rect 31377 10521 31389 10555
rect 31765 10521 31777 10555
rect 31377 10515 31777 10521
rect 31377 10437 31777 10443
rect 31377 10403 31389 10437
rect 31765 10403 31777 10437
rect 31377 10397 31777 10403
rect 31289 10377 31346 10393
rect 31289 10343 31305 10377
rect 31339 10343 31346 10377
rect 31289 10327 31346 10343
rect 31871 10365 31903 10824
rect 31871 10331 31988 10365
rect 30645 10319 31045 10325
rect 30645 10285 30657 10319
rect 31033 10285 31045 10319
rect 30645 10279 31045 10285
rect 31377 10319 31777 10325
rect 31377 10285 31389 10319
rect 31765 10285 31777 10319
rect 31377 10279 31777 10285
rect 29952 10228 29964 10262
rect 30340 10228 30521 10262
rect 29952 10222 30352 10228
rect 29701 10209 29849 10219
rect 29723 10177 29849 10209
rect 29806 10144 29849 10177
rect 30483 10201 30521 10228
rect 31289 10259 31348 10275
rect 31289 10225 31304 10259
rect 31338 10225 31348 10259
rect 31289 10208 31348 10225
rect 31871 10269 31925 10331
rect 31983 10269 31988 10331
rect 31871 10233 31988 10269
rect 30645 10201 31045 10207
rect 30483 10167 30657 10201
rect 31033 10167 31045 10201
rect 29952 10144 30352 10150
rect 29806 10110 29964 10144
rect 30340 10110 30352 10144
rect 29806 9908 29849 10110
rect 29952 10104 30352 10110
rect 29952 10026 30352 10032
rect 29952 9992 29964 10026
rect 30340 9992 30352 10026
rect 29952 9986 30352 9992
rect 30483 9965 30521 10167
rect 30645 10161 31045 10167
rect 30645 10083 31045 10089
rect 30645 10049 30657 10083
rect 31033 10049 31045 10083
rect 30645 10043 31045 10049
rect 31210 9995 31261 10012
rect 30645 9965 31045 9971
rect 30483 9931 30657 9965
rect 31033 9931 31045 9965
rect 31210 9961 31221 9995
rect 31255 9961 31261 9995
rect 31210 9945 31261 9961
rect 30645 9925 31045 9931
rect 29952 9908 30352 9914
rect 29806 9874 29964 9908
rect 30340 9874 30352 9908
rect 29806 9543 29849 9874
rect 29952 9868 30352 9874
rect 30164 9785 30340 9868
rect 31205 9832 31248 9945
rect 30152 9779 30352 9785
rect 30152 9745 30164 9779
rect 30340 9745 30352 9779
rect 30152 9739 30352 9745
rect 30503 9693 30569 9705
rect 30152 9661 30352 9667
rect 30152 9627 30164 9661
rect 30340 9627 30421 9661
rect 30503 9639 30509 9693
rect 30563 9639 30569 9693
rect 30503 9627 30569 9639
rect 30152 9621 30352 9627
rect 30386 9559 30421 9627
rect 31204 9559 31249 9832
rect 31289 9721 31338 10208
rect 31377 10201 31777 10207
rect 31871 10201 31903 10233
rect 31377 10167 31389 10201
rect 31765 10167 31903 10201
rect 31377 10161 31777 10167
rect 31377 10083 31777 10089
rect 31377 10049 31389 10083
rect 31765 10049 31777 10083
rect 31377 10043 31777 10049
rect 31277 9705 31339 9721
rect 31277 9671 31289 9705
rect 31323 9671 31339 9705
rect 31277 9665 31339 9671
rect 31377 9677 31577 9683
rect 31871 9677 31903 10167
rect 31377 9643 31389 9677
rect 31565 9644 31903 9677
rect 31565 9643 31577 9644
rect 31377 9637 31577 9643
rect 31377 9559 31577 9565
rect 30152 9543 30352 9549
rect 29806 9509 30164 9543
rect 30340 9509 30352 9543
rect 30152 9503 30352 9509
rect 30386 9525 31389 9559
rect 31565 9525 31577 9559
rect 30152 9425 30352 9431
rect 30386 9425 30421 9525
rect 31377 9519 31577 9525
rect 30152 9391 30164 9425
rect 30340 9391 30421 9425
rect 31055 9461 31169 9473
rect 30152 9385 30352 9391
rect 31055 9359 31061 9461
rect 31163 9359 31169 9461
rect 31055 9347 31169 9359
rect 32264 9394 32343 17574
rect 32264 9209 32344 9394
rect 30504 9123 32344 9209
rect 30154 9031 30354 9037
rect 30154 8997 30166 9031
rect 30342 8997 30423 9031
rect 30504 9027 30571 9123
rect 30154 8991 30354 8997
rect 30154 8913 30354 8919
rect 29808 8879 30166 8913
rect 30342 8879 30354 8913
rect 29808 8547 29851 8879
rect 30154 8873 30354 8879
rect 30388 8906 30423 8997
rect 30505 9012 30571 9027
rect 30695 9024 30767 9038
rect 30695 8958 30701 9024
rect 30761 9021 30767 9024
rect 30762 8961 30767 9021
rect 30761 8958 30767 8961
rect 30695 8946 30767 8958
rect 30505 8936 30571 8946
rect 31379 8906 31579 8912
rect 30388 8872 31391 8906
rect 31567 8872 31579 8906
rect 30154 8795 30354 8801
rect 30154 8761 30166 8795
rect 30342 8761 30354 8795
rect 30154 8755 30354 8761
rect 30154 8677 30354 8683
rect 30154 8643 30166 8677
rect 30342 8643 30354 8677
rect 30154 8637 30354 8643
rect 30166 8553 30342 8637
rect 30647 8604 31047 8610
rect 30485 8570 30659 8604
rect 31035 8570 31047 8604
rect 31207 8590 31250 8872
rect 31379 8866 31579 8872
rect 31379 8789 31579 8794
rect 31379 8788 31905 8789
rect 31278 8759 31340 8765
rect 31278 8725 31290 8759
rect 31324 8725 31340 8759
rect 31379 8754 31391 8788
rect 31567 8755 31905 8788
rect 31567 8754 31579 8755
rect 31379 8748 31579 8754
rect 31278 8709 31340 8725
rect 29954 8547 30354 8553
rect 29808 8513 29966 8547
rect 30342 8513 30354 8547
rect 29808 8311 29851 8513
rect 29954 8507 30354 8513
rect 29954 8429 30354 8435
rect 29954 8395 29966 8429
rect 30342 8395 30423 8429
rect 29954 8389 30354 8395
rect 29954 8311 30354 8317
rect 29808 8277 29966 8311
rect 30342 8277 30354 8311
rect 29808 8242 29851 8277
rect 29954 8271 30354 8277
rect 29725 8214 29851 8242
rect 29703 8204 29851 8214
rect 29757 8150 29851 8204
rect 29954 8193 30354 8199
rect 30388 8193 30423 8395
rect 30485 8368 30523 8570
rect 30647 8564 31047 8570
rect 31212 8574 31263 8590
rect 31212 8540 31223 8574
rect 31257 8540 31263 8574
rect 31212 8523 31263 8540
rect 30647 8486 31047 8492
rect 30647 8452 30659 8486
rect 31035 8452 31047 8486
rect 30647 8446 31047 8452
rect 30647 8368 31047 8374
rect 30485 8334 30659 8368
rect 31035 8334 31047 8368
rect 30485 8193 30523 8334
rect 30647 8328 31047 8334
rect 31291 8324 31340 8709
rect 31379 8486 31779 8492
rect 31379 8452 31391 8486
rect 31767 8452 31779 8486
rect 31379 8446 31779 8452
rect 31379 8368 31779 8374
rect 31379 8334 31391 8368
rect 31767 8334 31779 8368
rect 31379 8328 31779 8334
rect 31291 8308 31348 8324
rect 31291 8274 31307 8308
rect 31341 8274 31348 8308
rect 31291 8258 31348 8274
rect 31873 8296 31905 8755
rect 31873 8262 31990 8296
rect 30647 8250 31047 8256
rect 30647 8216 30659 8250
rect 31035 8216 31047 8250
rect 30647 8210 31047 8216
rect 31379 8250 31779 8256
rect 31379 8216 31391 8250
rect 31767 8216 31779 8250
rect 31379 8210 31779 8216
rect 29954 8159 29966 8193
rect 30342 8159 30523 8193
rect 29954 8153 30354 8159
rect 29703 8140 29851 8150
rect 29725 8108 29851 8140
rect 29808 8075 29851 8108
rect 30485 8132 30523 8159
rect 31291 8190 31350 8206
rect 31291 8156 31306 8190
rect 31340 8156 31350 8190
rect 31291 8139 31350 8156
rect 31873 8200 31927 8262
rect 31985 8200 31990 8262
rect 31873 8164 31990 8200
rect 30647 8132 31047 8138
rect 30485 8098 30659 8132
rect 31035 8098 31047 8132
rect 29954 8075 30354 8081
rect 29808 8041 29966 8075
rect 30342 8041 30354 8075
rect 29808 7839 29851 8041
rect 29954 8035 30354 8041
rect 29954 7957 30354 7963
rect 29954 7923 29966 7957
rect 30342 7923 30354 7957
rect 29954 7917 30354 7923
rect 30485 7896 30523 8098
rect 30647 8092 31047 8098
rect 30647 8014 31047 8020
rect 30647 7980 30659 8014
rect 31035 7980 31047 8014
rect 30647 7974 31047 7980
rect 31212 7926 31263 7943
rect 30647 7896 31047 7902
rect 30485 7862 30659 7896
rect 31035 7862 31047 7896
rect 31212 7892 31223 7926
rect 31257 7892 31263 7926
rect 31212 7876 31263 7892
rect 30647 7856 31047 7862
rect 29954 7839 30354 7845
rect 29808 7805 29966 7839
rect 30342 7805 30354 7839
rect 29808 7474 29851 7805
rect 29954 7799 30354 7805
rect 30166 7716 30342 7799
rect 31207 7763 31250 7876
rect 30154 7710 30354 7716
rect 30154 7676 30166 7710
rect 30342 7676 30354 7710
rect 30154 7670 30354 7676
rect 30505 7624 30571 7636
rect 30154 7592 30354 7598
rect 30154 7558 30166 7592
rect 30342 7558 30423 7592
rect 30505 7570 30511 7624
rect 30565 7570 30571 7624
rect 30505 7558 30571 7570
rect 30154 7552 30354 7558
rect 30388 7490 30423 7558
rect 31206 7490 31251 7763
rect 31291 7652 31340 8139
rect 31379 8132 31779 8138
rect 31873 8132 31905 8164
rect 31379 8098 31391 8132
rect 31767 8098 31905 8132
rect 31379 8092 31779 8098
rect 31379 8014 31779 8020
rect 31379 7980 31391 8014
rect 31767 7980 31779 8014
rect 31379 7974 31779 7980
rect 31279 7636 31341 7652
rect 31279 7602 31291 7636
rect 31325 7602 31341 7636
rect 31279 7596 31341 7602
rect 31379 7608 31579 7614
rect 31873 7608 31905 8098
rect 31379 7574 31391 7608
rect 31567 7575 31905 7608
rect 31567 7574 31579 7575
rect 31379 7568 31579 7574
rect 31379 7490 31579 7496
rect 30154 7474 30354 7480
rect 29808 7440 30166 7474
rect 30342 7440 30354 7474
rect 30154 7434 30354 7440
rect 30388 7456 31391 7490
rect 31567 7456 31579 7490
rect 30154 7356 30354 7362
rect 30388 7356 30423 7456
rect 31379 7450 31579 7456
rect 30154 7322 30166 7356
rect 30342 7322 30423 7356
rect 31057 7392 31171 7404
rect 30154 7316 30354 7322
rect 31057 7290 31063 7392
rect 31165 7290 31171 7392
rect 31057 7278 31171 7290
rect 32408 7207 32485 18003
rect 32542 9302 32623 18424
rect 32539 9228 32549 9302
rect 32615 9228 32625 9302
rect 27311 7099 27321 7157
rect 27389 7099 27399 7157
rect 32408 7143 32416 7207
rect 32478 7143 32486 7207
rect 32408 7135 32485 7143
rect 27062 6806 27074 6863
rect 27130 6806 27142 6863
rect 26841 6502 26851 6555
rect 26912 6502 26922 6555
rect 26657 6340 26667 6398
rect 26737 6340 26747 6398
rect 26457 6190 26467 6248
rect 26535 6190 26545 6248
rect 26271 6031 26281 6085
rect 26339 6031 26349 6085
rect 25326 5826 25336 5892
rect 25402 5885 25692 5892
rect 25402 5832 25628 5885
rect 25688 5832 25698 5885
rect 26037 5841 26047 5901
rect 26111 5841 26121 5901
rect 25402 5826 25692 5832
rect 25336 5627 25346 5704
rect 25417 5702 25427 5704
rect 25417 5693 25692 5702
rect 25417 5635 25636 5693
rect 25688 5635 25698 5693
rect 25417 5630 25692 5635
rect 25417 5627 25427 5630
rect 23846 5185 24266 5190
rect 24980 5185 25296 5190
rect 23846 5174 24333 5185
rect 23846 5147 24282 5174
rect 23846 5146 24153 5147
rect 23846 5018 23880 5146
rect 24266 5140 24282 5147
rect 24316 5140 24333 5174
rect 24266 5134 24333 5140
rect 24913 5174 25296 5185
rect 24913 5140 24930 5174
rect 24964 5147 25296 5174
rect 24964 5140 24980 5147
rect 24913 5134 24980 5140
rect 23986 5106 24042 5118
rect 25099 5107 25155 5119
rect 25099 5106 25115 5107
rect 23986 5072 23992 5106
rect 24026 5091 24596 5106
rect 24026 5072 24546 5091
rect 23986 5057 24546 5072
rect 24580 5057 24596 5091
rect 23986 5056 24042 5057
rect 24529 5047 24596 5057
rect 24648 5090 25115 5106
rect 24648 5056 24664 5090
rect 24698 5073 25115 5090
rect 25149 5073 25155 5107
rect 24698 5057 25155 5073
rect 24698 5056 24714 5057
rect 24648 5049 24714 5056
rect 25262 5018 25296 5147
rect 23840 5006 23886 5018
rect 23840 4830 23846 5006
rect 23880 4830 23886 5006
rect 23840 4818 23886 4830
rect 23958 5006 24004 5018
rect 23958 4830 23964 5006
rect 23998 4830 24004 5006
rect 23958 4818 24004 4830
rect 24364 5006 24410 5018
rect 23965 4524 23998 4818
rect 24364 4630 24370 5006
rect 24404 4630 24410 5006
rect 24364 4618 24410 4630
rect 24482 5006 24528 5018
rect 24482 4630 24488 5006
rect 24522 4630 24528 5006
rect 24482 4618 24528 4630
rect 24600 5006 24646 5018
rect 24600 4630 24606 5006
rect 24640 4630 24646 5006
rect 24600 4618 24646 4630
rect 24718 5006 24764 5018
rect 24718 4630 24724 5006
rect 24758 4630 24764 5006
rect 24718 4618 24764 4630
rect 24836 5006 24882 5018
rect 24836 4630 24842 5006
rect 24876 4630 24882 5006
rect 25138 5006 25184 5018
rect 25138 4830 25144 5006
rect 25178 4830 25184 5006
rect 25138 4818 25184 4830
rect 25256 5006 25302 5018
rect 25256 4830 25262 5006
rect 25296 4830 25302 5006
rect 25256 4818 25302 4830
rect 24836 4618 24882 4630
rect 24488 4524 24522 4618
rect 25145 4524 25179 4818
rect 23965 4492 25179 4524
rect 24554 4470 24686 4492
rect 24554 4412 24590 4470
rect 24652 4412 24686 4470
rect 24554 4407 24686 4412
rect 26047 4269 26111 5841
rect 23343 4205 26111 4269
rect 23344 4061 23408 4205
rect 25806 4204 26111 4205
rect 23338 4055 23413 4061
rect 23338 4004 23350 4055
rect 23401 4004 23413 4055
rect 23338 3998 23413 4004
rect 26277 3958 26341 6031
rect 21310 3950 26341 3958
rect 21310 3896 21319 3950
rect 21366 3896 26341 3950
rect 21310 3877 26341 3896
rect 26464 3849 26538 6190
rect 19264 3847 26538 3849
rect 19264 3793 19272 3847
rect 19319 3793 26538 3847
rect 19264 3757 26538 3793
rect 17173 3737 17238 3749
rect 17173 3729 17179 3737
rect 17145 3686 17179 3729
rect 17229 3729 17238 3737
rect 26662 3730 26741 6340
rect 26578 3729 26741 3730
rect 17229 3686 26741 3729
rect 17145 3649 26741 3686
rect 26578 3648 26741 3649
rect 15100 3602 15107 3642
rect 15099 3589 15107 3602
rect 15158 3602 15164 3642
rect 26849 3602 26913 6502
rect 15158 3589 26913 3602
rect 15099 3534 26913 3589
rect 26849 3533 26913 3534
rect 27062 3503 27142 6806
rect 13000 3498 27142 3503
rect 13000 3447 13011 3498
rect 13055 3447 27142 3498
rect 13000 3436 27142 3447
rect 13001 3435 13065 3436
rect 27062 3435 27142 3436
rect 132 3348 142 3411
rect 221 3348 231 3411
rect 10928 3404 10994 3415
rect 27316 3404 27395 7099
rect 30503 7056 32485 7135
rect 30152 6963 30352 6969
rect 30152 6929 30164 6963
rect 30340 6929 30421 6963
rect 30152 6923 30352 6929
rect 30152 6845 30352 6851
rect 29806 6811 30164 6845
rect 30340 6811 30352 6845
rect 29806 6479 29849 6811
rect 30152 6805 30352 6811
rect 30386 6838 30421 6929
rect 30503 6944 30569 7056
rect 30693 6956 30765 6969
rect 30693 6890 30699 6956
rect 30759 6890 30765 6956
rect 30693 6878 30765 6890
rect 30503 6868 30569 6878
rect 31377 6838 31577 6844
rect 30386 6804 31389 6838
rect 31565 6804 31577 6838
rect 30152 6727 30352 6733
rect 30152 6693 30164 6727
rect 30340 6693 30352 6727
rect 30152 6687 30352 6693
rect 30152 6609 30352 6615
rect 30152 6575 30164 6609
rect 30340 6575 30352 6609
rect 30152 6569 30352 6575
rect 30164 6485 30340 6569
rect 30645 6536 31045 6542
rect 30483 6502 30657 6536
rect 31033 6502 31045 6536
rect 31205 6522 31248 6804
rect 31377 6798 31577 6804
rect 31377 6721 31577 6726
rect 31377 6720 31903 6721
rect 31276 6691 31338 6697
rect 31276 6657 31288 6691
rect 31322 6657 31338 6691
rect 31377 6686 31389 6720
rect 31565 6687 31903 6720
rect 31565 6686 31577 6687
rect 31377 6680 31577 6686
rect 31276 6641 31338 6657
rect 29952 6479 30352 6485
rect 29806 6445 29964 6479
rect 30340 6445 30352 6479
rect 29806 6243 29849 6445
rect 29952 6439 30352 6445
rect 29952 6361 30352 6367
rect 29952 6327 29964 6361
rect 30340 6327 30421 6361
rect 29952 6321 30352 6327
rect 29952 6243 30352 6249
rect 29806 6209 29964 6243
rect 30340 6209 30352 6243
rect 29806 6174 29849 6209
rect 29952 6203 30352 6209
rect 29723 6146 29849 6174
rect 29701 6136 29849 6146
rect 29755 6082 29849 6136
rect 29952 6125 30352 6131
rect 30386 6125 30421 6327
rect 30483 6300 30521 6502
rect 30645 6496 31045 6502
rect 31210 6506 31261 6522
rect 31210 6472 31221 6506
rect 31255 6472 31261 6506
rect 31210 6455 31261 6472
rect 30645 6418 31045 6424
rect 30645 6384 30657 6418
rect 31033 6384 31045 6418
rect 30645 6378 31045 6384
rect 30645 6300 31045 6306
rect 30483 6266 30657 6300
rect 31033 6266 31045 6300
rect 30483 6125 30521 6266
rect 30645 6260 31045 6266
rect 31289 6256 31338 6641
rect 31377 6418 31777 6424
rect 31377 6384 31389 6418
rect 31765 6384 31777 6418
rect 31377 6378 31777 6384
rect 31377 6300 31777 6306
rect 31377 6266 31389 6300
rect 31765 6266 31777 6300
rect 31377 6260 31777 6266
rect 31289 6240 31346 6256
rect 31289 6206 31305 6240
rect 31339 6206 31346 6240
rect 31289 6190 31346 6206
rect 31871 6228 31903 6687
rect 31871 6194 31988 6228
rect 30645 6182 31045 6188
rect 30645 6148 30657 6182
rect 31033 6148 31045 6182
rect 30645 6142 31045 6148
rect 31377 6182 31777 6188
rect 31377 6148 31389 6182
rect 31765 6148 31777 6182
rect 31377 6142 31777 6148
rect 29952 6091 29964 6125
rect 30340 6091 30521 6125
rect 29952 6085 30352 6091
rect 29701 6072 29849 6082
rect 29723 6040 29849 6072
rect 29806 6007 29849 6040
rect 30483 6064 30521 6091
rect 31289 6122 31348 6138
rect 31289 6088 31304 6122
rect 31338 6088 31348 6122
rect 31289 6071 31348 6088
rect 31871 6132 31925 6194
rect 31983 6132 31988 6194
rect 31871 6096 31988 6132
rect 30645 6064 31045 6070
rect 30483 6030 30657 6064
rect 31033 6030 31045 6064
rect 29952 6007 30352 6013
rect 29806 5973 29964 6007
rect 30340 5973 30352 6007
rect 29806 5771 29849 5973
rect 29952 5967 30352 5973
rect 29952 5889 30352 5895
rect 29952 5855 29964 5889
rect 30340 5855 30352 5889
rect 29952 5849 30352 5855
rect 30483 5828 30521 6030
rect 30645 6024 31045 6030
rect 30645 5946 31045 5952
rect 30645 5912 30657 5946
rect 31033 5912 31045 5946
rect 30645 5906 31045 5912
rect 31210 5858 31261 5875
rect 30645 5828 31045 5834
rect 30483 5794 30657 5828
rect 31033 5794 31045 5828
rect 31210 5824 31221 5858
rect 31255 5824 31261 5858
rect 31210 5808 31261 5824
rect 30645 5788 31045 5794
rect 29952 5771 30352 5777
rect 29806 5737 29964 5771
rect 30340 5737 30352 5771
rect 29806 5406 29849 5737
rect 29952 5731 30352 5737
rect 30164 5648 30340 5731
rect 31205 5695 31248 5808
rect 30152 5642 30352 5648
rect 30152 5608 30164 5642
rect 30340 5608 30352 5642
rect 30152 5602 30352 5608
rect 30503 5556 30569 5568
rect 30152 5524 30352 5530
rect 30152 5490 30164 5524
rect 30340 5490 30421 5524
rect 30503 5502 30509 5556
rect 30563 5502 30569 5556
rect 30503 5490 30569 5502
rect 30152 5484 30352 5490
rect 30386 5422 30421 5490
rect 31204 5422 31249 5695
rect 31289 5584 31338 6071
rect 31377 6064 31777 6070
rect 31871 6064 31903 6096
rect 31377 6030 31389 6064
rect 31765 6030 31903 6064
rect 31377 6024 31777 6030
rect 31377 5946 31777 5952
rect 31377 5912 31389 5946
rect 31765 5912 31777 5946
rect 31377 5906 31777 5912
rect 31277 5568 31339 5584
rect 31277 5534 31289 5568
rect 31323 5534 31339 5568
rect 31277 5528 31339 5534
rect 31377 5540 31577 5546
rect 31871 5540 31903 6030
rect 31377 5506 31389 5540
rect 31565 5507 31903 5540
rect 31565 5506 31577 5507
rect 31377 5500 31577 5506
rect 31377 5422 31577 5428
rect 30152 5406 30352 5412
rect 29806 5372 30164 5406
rect 30340 5372 30352 5406
rect 30152 5366 30352 5372
rect 30386 5388 31389 5422
rect 31565 5388 31577 5422
rect 30152 5288 30352 5294
rect 30386 5288 30421 5388
rect 31377 5382 31577 5388
rect 30152 5254 30164 5288
rect 30340 5254 30421 5288
rect 31055 5324 31169 5336
rect 30152 5248 30352 5254
rect 31055 5222 31061 5324
rect 31163 5222 31169 5324
rect 31055 5210 31169 5222
rect 32542 5066 32623 9228
rect 30503 4987 32623 5066
rect 30152 4894 30352 4900
rect 30152 4860 30164 4894
rect 30340 4860 30421 4894
rect 30152 4854 30352 4860
rect 30152 4776 30352 4782
rect 29806 4742 30164 4776
rect 30340 4742 30352 4776
rect 29806 4410 29849 4742
rect 30152 4736 30352 4742
rect 30386 4769 30421 4860
rect 30503 4886 30570 4987
rect 30693 4887 30765 4902
rect 30503 4875 30569 4886
rect 30693 4884 30699 4887
rect 30759 4884 30765 4887
rect 30690 4823 30699 4884
rect 30759 4823 30766 4884
rect 30693 4821 30699 4823
rect 30759 4821 30765 4823
rect 30693 4809 30765 4821
rect 30503 4799 30569 4809
rect 31377 4769 31577 4775
rect 30386 4735 31389 4769
rect 31565 4735 31577 4769
rect 30152 4658 30352 4664
rect 30152 4624 30164 4658
rect 30340 4624 30352 4658
rect 30152 4618 30352 4624
rect 30152 4540 30352 4546
rect 30152 4506 30164 4540
rect 30340 4506 30352 4540
rect 30152 4500 30352 4506
rect 30164 4416 30340 4500
rect 30645 4467 31045 4473
rect 30483 4433 30657 4467
rect 31033 4433 31045 4467
rect 31205 4453 31248 4735
rect 31377 4729 31577 4735
rect 31377 4652 31577 4657
rect 31377 4651 31903 4652
rect 31276 4622 31338 4628
rect 31276 4588 31288 4622
rect 31322 4588 31338 4622
rect 31377 4617 31389 4651
rect 31565 4618 31903 4651
rect 31565 4617 31577 4618
rect 31377 4611 31577 4617
rect 31276 4572 31338 4588
rect 29952 4410 30352 4416
rect 29806 4376 29964 4410
rect 30340 4376 30352 4410
rect 29806 4174 29849 4376
rect 29952 4370 30352 4376
rect 29952 4292 30352 4298
rect 29952 4258 29964 4292
rect 30340 4258 30421 4292
rect 29952 4252 30352 4258
rect 29952 4174 30352 4180
rect 29806 4140 29964 4174
rect 30340 4140 30352 4174
rect 29806 4105 29849 4140
rect 29952 4134 30352 4140
rect 29723 4077 29849 4105
rect 29701 4067 29849 4077
rect 29755 4013 29849 4067
rect 29952 4056 30352 4062
rect 30386 4056 30421 4258
rect 30483 4231 30521 4433
rect 30645 4427 31045 4433
rect 31210 4437 31261 4453
rect 31210 4403 31221 4437
rect 31255 4403 31261 4437
rect 31210 4386 31261 4403
rect 30645 4349 31045 4355
rect 30645 4315 30657 4349
rect 31033 4315 31045 4349
rect 30645 4309 31045 4315
rect 30645 4231 31045 4237
rect 30483 4197 30657 4231
rect 31033 4197 31045 4231
rect 30483 4056 30521 4197
rect 30645 4191 31045 4197
rect 31289 4187 31338 4572
rect 31377 4349 31777 4355
rect 31377 4315 31389 4349
rect 31765 4315 31777 4349
rect 31377 4309 31777 4315
rect 31377 4231 31777 4237
rect 31377 4197 31389 4231
rect 31765 4197 31777 4231
rect 31377 4191 31777 4197
rect 31289 4171 31346 4187
rect 31289 4137 31305 4171
rect 31339 4137 31346 4171
rect 31289 4121 31346 4137
rect 31871 4159 31903 4618
rect 31871 4125 31988 4159
rect 30645 4113 31045 4119
rect 30645 4079 30657 4113
rect 31033 4079 31045 4113
rect 30645 4073 31045 4079
rect 31377 4113 31777 4119
rect 31377 4079 31389 4113
rect 31765 4079 31777 4113
rect 31377 4073 31777 4079
rect 29952 4022 29964 4056
rect 30340 4022 30521 4056
rect 29952 4016 30352 4022
rect 29701 4003 29849 4013
rect 29723 3971 29849 4003
rect 10928 3403 27395 3404
rect 10928 3349 10934 3403
rect 10987 3349 27395 3403
rect 10928 3326 27395 3349
rect 29806 3938 29849 3971
rect 30483 3995 30521 4022
rect 31289 4053 31348 4069
rect 31289 4019 31304 4053
rect 31338 4019 31348 4053
rect 31289 4002 31348 4019
rect 31871 4063 31925 4125
rect 31983 4063 31988 4125
rect 31871 4027 31988 4063
rect 30645 3995 31045 4001
rect 30483 3961 30657 3995
rect 31033 3961 31045 3995
rect 29952 3938 30352 3944
rect 29806 3904 29964 3938
rect 30340 3904 30352 3938
rect 29806 3702 29849 3904
rect 29952 3898 30352 3904
rect 29952 3820 30352 3826
rect 29952 3786 29964 3820
rect 30340 3786 30352 3820
rect 29952 3780 30352 3786
rect 30483 3759 30521 3961
rect 30645 3955 31045 3961
rect 30645 3877 31045 3883
rect 30645 3843 30657 3877
rect 31033 3843 31045 3877
rect 30645 3837 31045 3843
rect 31210 3789 31261 3806
rect 30645 3759 31045 3765
rect 30483 3725 30657 3759
rect 31033 3725 31045 3759
rect 31210 3755 31221 3789
rect 31255 3755 31261 3789
rect 31210 3739 31261 3755
rect 30645 3719 31045 3725
rect 29952 3702 30352 3708
rect 29806 3668 29964 3702
rect 30340 3668 30352 3702
rect 29806 3337 29849 3668
rect 29952 3662 30352 3668
rect 30164 3579 30340 3662
rect 31205 3626 31248 3739
rect 30152 3573 30352 3579
rect 30152 3539 30164 3573
rect 30340 3539 30352 3573
rect 30152 3533 30352 3539
rect 30503 3487 30569 3499
rect 30152 3455 30352 3461
rect 30152 3421 30164 3455
rect 30340 3421 30421 3455
rect 30503 3433 30509 3487
rect 30563 3433 30569 3487
rect 30503 3421 30569 3433
rect 30152 3415 30352 3421
rect 30386 3353 30421 3421
rect 31204 3353 31249 3626
rect 31289 3515 31338 4002
rect 31377 3995 31777 4001
rect 31871 3995 31903 4027
rect 31377 3961 31389 3995
rect 31765 3961 31903 3995
rect 31377 3955 31777 3961
rect 31377 3877 31777 3883
rect 31377 3843 31389 3877
rect 31765 3843 31777 3877
rect 31377 3837 31777 3843
rect 31277 3499 31339 3515
rect 31277 3465 31289 3499
rect 31323 3465 31339 3499
rect 31277 3459 31339 3465
rect 31377 3471 31577 3477
rect 31871 3471 31903 3961
rect 31377 3437 31389 3471
rect 31565 3438 31903 3471
rect 31565 3437 31577 3438
rect 31377 3431 31577 3437
rect 31377 3353 31577 3359
rect 30152 3337 30352 3343
rect 29806 3303 30164 3337
rect 30340 3303 30352 3337
rect 30152 3297 30352 3303
rect 30386 3319 31389 3353
rect 31565 3319 31577 3353
rect -4 3285 815 3286
rect 22864 3285 29427 3287
rect -4 3221 29427 3285
rect -4 2655 65 3221
rect 789 3220 29427 3221
rect 29310 3194 29427 3220
rect 128 3098 138 3161
rect 217 3098 227 3161
rect 3136 3100 29266 3181
rect 126 2985 136 3048
rect 215 2985 225 3048
rect 137 2984 215 2985
rect 124 2860 134 2921
rect 211 2860 221 2921
rect 3138 2678 3209 3100
rect 22930 3099 29266 3100
rect 29141 3098 29266 3099
rect 6273 2993 29103 3071
rect 29149 3065 29266 3098
rect 6273 2992 22859 2993
rect 6273 2737 6342 2992
rect 9419 2949 22461 2951
rect 9419 2875 28942 2949
rect 6273 2711 6343 2737
rect -4 1334 64 2655
rect 1498 2324 1508 2384
rect 1588 2324 1598 2384
rect 1498 2284 1598 2324
rect 701 2227 2504 2284
rect 701 2140 735 2227
rect 1876 2140 1910 2227
rect 695 2128 741 2140
rect 695 1940 701 2128
rect 254 1928 300 1940
rect 254 1752 260 1928
rect 294 1752 300 1928
rect 254 1740 300 1752
rect 372 1928 418 1940
rect 372 1752 378 1928
rect 412 1752 418 1928
rect 372 1740 418 1752
rect 490 1928 536 1940
rect 490 1752 496 1928
rect 530 1752 536 1928
rect 490 1740 536 1752
rect 608 1928 701 1940
rect 608 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 741 2128
rect 608 1740 741 1752
rect 813 2128 859 2140
rect 813 1752 819 2128
rect 853 1752 859 2128
rect 813 1740 859 1752
rect 931 2128 977 2140
rect 931 1752 937 2128
rect 971 1752 977 2128
rect 931 1740 977 1752
rect 1049 2128 1095 2140
rect 1049 1752 1055 2128
rect 1089 1752 1095 2128
rect 1049 1740 1095 1752
rect 1162 2128 1208 2140
rect 1162 1752 1168 2128
rect 1202 1752 1208 2128
rect 1162 1740 1208 1752
rect 1280 2128 1326 2140
rect 1280 1752 1286 2128
rect 1320 1752 1326 2128
rect 1280 1740 1326 1752
rect 1398 2128 1444 2140
rect 1398 1752 1404 2128
rect 1438 1752 1444 2128
rect 1398 1740 1444 1752
rect 1516 2128 1562 2140
rect 1516 1752 1522 2128
rect 1556 1752 1562 2128
rect 1516 1740 1562 1752
rect 1634 2128 1680 2140
rect 1634 1752 1640 2128
rect 1674 1752 1680 2128
rect 1634 1740 1680 1752
rect 1752 2128 1798 2140
rect 1752 1752 1758 2128
rect 1792 1752 1798 2128
rect 1752 1740 1798 1752
rect 1870 2128 1916 2140
rect 1870 1752 1876 2128
rect 1910 1752 1916 2128
rect 1870 1740 1916 1752
rect 1989 2128 2035 2140
rect 1989 1752 1995 2128
rect 2029 1752 2035 2128
rect 1989 1740 2035 1752
rect 2107 2128 2153 2140
rect 2107 1752 2113 2128
rect 2147 1752 2153 2128
rect 2107 1740 2153 1752
rect 2225 2128 2271 2140
rect 2225 1752 2231 2128
rect 2265 1752 2271 2128
rect 2225 1740 2271 1752
rect 2343 2128 2389 2140
rect 2343 1752 2349 2128
rect 2383 1752 2389 2128
rect 2467 1940 2504 2227
rect 2343 1740 2389 1752
rect 2462 1928 2508 1940
rect 2462 1752 2468 1928
rect 2502 1752 2508 1928
rect 2462 1740 2508 1752
rect 2580 1928 2626 1940
rect 2580 1752 2586 1928
rect 2620 1752 2626 1928
rect 2580 1740 2626 1752
rect 2698 1928 2744 1940
rect 2698 1752 2704 1928
rect 2738 1752 2744 1928
rect 2698 1740 2744 1752
rect 2816 1928 2862 1940
rect 2816 1752 2822 1928
rect 2856 1752 2862 1928
rect 2816 1740 2862 1752
rect 259 1554 294 1740
rect 1168 1656 1202 1740
rect 2349 1656 2383 1740
rect 1168 1614 2383 1656
rect 2349 1594 2383 1614
rect 2349 1578 2706 1594
rect 259 1537 1396 1554
rect 259 1503 1346 1537
rect 1380 1503 1396 1537
rect 2349 1544 2656 1578
rect 2690 1544 2706 1578
rect 2349 1528 2706 1544
rect 259 1487 1396 1503
rect 101 1442 176 1450
rect 101 1374 117 1442
rect 174 1374 184 1442
rect 101 1366 176 1374
rect -4 1326 176 1334
rect -4 1258 117 1326
rect 174 1258 184 1326
rect -4 1250 176 1258
rect -4 1249 64 1250
rect 259 977 294 1487
rect 349 1441 441 1454
rect 349 1378 361 1441
rect 432 1378 441 1441
rect 349 1369 441 1378
rect 1434 1441 1526 1451
rect 1434 1379 1446 1441
rect 1516 1379 1526 1441
rect 1434 1366 1526 1379
rect 2822 1386 2857 1740
rect 1681 1324 1746 1327
rect 1681 1321 1750 1324
rect 1681 1261 1687 1321
rect 1746 1261 1756 1321
rect 1681 1257 1750 1261
rect 1681 1255 1746 1257
rect 1316 1158 1408 1166
rect 1316 1093 1328 1158
rect 1396 1093 1408 1158
rect 1316 1081 1408 1093
rect 2822 978 3003 1386
rect 3138 1334 3206 2678
rect 4642 2324 4652 2384
rect 4732 2324 4742 2384
rect 4642 2284 4742 2324
rect 3845 2227 5648 2284
rect 3845 2140 3879 2227
rect 5020 2140 5054 2227
rect 3839 2128 3885 2140
rect 3839 1940 3845 2128
rect 3398 1928 3444 1940
rect 3398 1752 3404 1928
rect 3438 1752 3444 1928
rect 3398 1740 3444 1752
rect 3516 1928 3562 1940
rect 3516 1752 3522 1928
rect 3556 1752 3562 1928
rect 3516 1740 3562 1752
rect 3634 1928 3680 1940
rect 3634 1752 3640 1928
rect 3674 1752 3680 1928
rect 3634 1740 3680 1752
rect 3752 1928 3845 1940
rect 3752 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3885 2128
rect 3752 1740 3885 1752
rect 3957 2128 4003 2140
rect 3957 1752 3963 2128
rect 3997 1752 4003 2128
rect 3957 1740 4003 1752
rect 4075 2128 4121 2140
rect 4075 1752 4081 2128
rect 4115 1752 4121 2128
rect 4075 1740 4121 1752
rect 4193 2128 4239 2140
rect 4193 1752 4199 2128
rect 4233 1752 4239 2128
rect 4193 1740 4239 1752
rect 4306 2128 4352 2140
rect 4306 1752 4312 2128
rect 4346 1752 4352 2128
rect 4306 1740 4352 1752
rect 4424 2128 4470 2140
rect 4424 1752 4430 2128
rect 4464 1752 4470 2128
rect 4424 1740 4470 1752
rect 4542 2128 4588 2140
rect 4542 1752 4548 2128
rect 4582 1752 4588 2128
rect 4542 1740 4588 1752
rect 4660 2128 4706 2140
rect 4660 1752 4666 2128
rect 4700 1752 4706 2128
rect 4660 1740 4706 1752
rect 4778 2128 4824 2140
rect 4778 1752 4784 2128
rect 4818 1752 4824 2128
rect 4778 1740 4824 1752
rect 4896 2128 4942 2140
rect 4896 1752 4902 2128
rect 4936 1752 4942 2128
rect 4896 1740 4942 1752
rect 5014 2128 5060 2140
rect 5014 1752 5020 2128
rect 5054 1752 5060 2128
rect 5014 1740 5060 1752
rect 5133 2128 5179 2140
rect 5133 1752 5139 2128
rect 5173 1752 5179 2128
rect 5133 1740 5179 1752
rect 5251 2128 5297 2140
rect 5251 1752 5257 2128
rect 5291 1752 5297 2128
rect 5251 1740 5297 1752
rect 5369 2128 5415 2140
rect 5369 1752 5375 2128
rect 5409 1752 5415 2128
rect 5369 1740 5415 1752
rect 5487 2128 5533 2140
rect 5487 1752 5493 2128
rect 5527 1752 5533 2128
rect 5611 1940 5648 2227
rect 5487 1740 5533 1752
rect 5606 1928 5652 1940
rect 5606 1752 5612 1928
rect 5646 1752 5652 1928
rect 5606 1740 5652 1752
rect 5724 1928 5770 1940
rect 5724 1752 5730 1928
rect 5764 1752 5770 1928
rect 5724 1740 5770 1752
rect 5842 1928 5888 1940
rect 5842 1752 5848 1928
rect 5882 1752 5888 1928
rect 5842 1740 5888 1752
rect 5960 1928 6006 1940
rect 5960 1752 5966 1928
rect 6000 1752 6006 1928
rect 5960 1740 6006 1752
rect 3403 1554 3438 1740
rect 4312 1656 4346 1740
rect 5493 1656 5527 1740
rect 4312 1614 5527 1656
rect 5493 1594 5527 1614
rect 5493 1578 5850 1594
rect 3403 1537 4540 1554
rect 3403 1503 4490 1537
rect 4524 1503 4540 1537
rect 5493 1544 5800 1578
rect 5834 1544 5850 1578
rect 5493 1528 5850 1544
rect 3403 1487 4540 1503
rect 3247 1442 3320 1450
rect 3247 1374 3261 1442
rect 3318 1374 3328 1442
rect 3247 1366 3320 1374
rect 3138 1326 3320 1334
rect 3138 1258 3261 1326
rect 3318 1258 3328 1326
rect 3138 1250 3320 1258
rect 3138 1247 3215 1250
rect 259 930 1631 977
rect 1953 931 3003 978
rect 1093 807 1127 930
rect 1565 917 1631 930
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1954 807 1988 931
rect 1088 795 1134 807
rect 1088 619 1094 795
rect 1128 619 1134 795
rect 1088 607 1134 619
rect 1206 795 1326 807
rect 1206 619 1212 795
rect 1246 619 1286 795
rect 1206 607 1286 619
rect 1212 240 1246 607
rect 1280 419 1286 607
rect 1320 419 1326 795
rect 1280 407 1326 419
rect 1398 795 1444 807
rect 1398 419 1404 795
rect 1438 419 1444 795
rect 1398 407 1444 419
rect 1516 795 1562 807
rect 1516 419 1522 795
rect 1556 419 1562 795
rect 1516 407 1562 419
rect 1634 795 1680 807
rect 1634 419 1640 795
rect 1674 419 1680 795
rect 1634 407 1680 419
rect 1752 795 1876 807
rect 1752 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1876 795
rect 1792 607 1876 619
rect 1948 795 1994 807
rect 1948 619 1954 795
rect 1988 619 1994 795
rect 1948 607 1994 619
rect 1792 419 1798 607
rect 1752 407 1798 419
rect 1522 334 1556 407
rect 1507 318 1573 334
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 1507 268 1573 284
rect 1836 240 1870 607
rect 1212 188 1870 240
rect 1510 166 1602 188
rect 1510 114 1522 166
rect 1588 114 1602 166
rect 1510 110 1602 114
rect -309 -317 -285 -155
rect -181 -317 -142 -155
rect -309 -346 -142 -317
rect -574 -498 -434 -479
rect -809 -766 -792 -604
rect -688 -766 -669 -604
rect -809 -781 -669 -766
rect 2857 -1063 3003 931
rect 3403 977 3438 1487
rect 3493 1441 3585 1454
rect 3493 1378 3505 1441
rect 3576 1378 3585 1441
rect 3493 1369 3585 1378
rect 4578 1441 4670 1451
rect 4578 1379 4590 1441
rect 4660 1379 4670 1441
rect 4578 1366 4670 1379
rect 5966 1386 6001 1740
rect 5966 1347 6147 1386
rect 4825 1324 4890 1327
rect 4825 1321 4894 1324
rect 4825 1261 4831 1321
rect 4890 1261 4900 1321
rect 4825 1257 4894 1261
rect 4825 1255 4890 1257
rect 4460 1158 4552 1166
rect 4460 1093 4472 1158
rect 4540 1093 4552 1158
rect 4460 1081 4552 1093
rect 5966 978 6149 1347
rect 6275 1338 6343 2711
rect 7774 2328 7784 2388
rect 7864 2328 7874 2388
rect 7774 2288 7874 2328
rect 6977 2231 8780 2288
rect 6977 2144 7011 2231
rect 8152 2144 8186 2231
rect 6971 2132 7017 2144
rect 6971 1944 6977 2132
rect 6530 1932 6576 1944
rect 6530 1756 6536 1932
rect 6570 1756 6576 1932
rect 6530 1744 6576 1756
rect 6648 1932 6694 1944
rect 6648 1756 6654 1932
rect 6688 1756 6694 1932
rect 6648 1744 6694 1756
rect 6766 1932 6812 1944
rect 6766 1756 6772 1932
rect 6806 1756 6812 1932
rect 6766 1744 6812 1756
rect 6884 1932 6977 1944
rect 6884 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7017 2132
rect 6884 1744 7017 1756
rect 7089 2132 7135 2144
rect 7089 1756 7095 2132
rect 7129 1756 7135 2132
rect 7089 1744 7135 1756
rect 7207 2132 7253 2144
rect 7207 1756 7213 2132
rect 7247 1756 7253 2132
rect 7207 1744 7253 1756
rect 7325 2132 7371 2144
rect 7325 1756 7331 2132
rect 7365 1756 7371 2132
rect 7325 1744 7371 1756
rect 7438 2132 7484 2144
rect 7438 1756 7444 2132
rect 7478 1756 7484 2132
rect 7438 1744 7484 1756
rect 7556 2132 7602 2144
rect 7556 1756 7562 2132
rect 7596 1756 7602 2132
rect 7556 1744 7602 1756
rect 7674 2132 7720 2144
rect 7674 1756 7680 2132
rect 7714 1756 7720 2132
rect 7674 1744 7720 1756
rect 7792 2132 7838 2144
rect 7792 1756 7798 2132
rect 7832 1756 7838 2132
rect 7792 1744 7838 1756
rect 7910 2132 7956 2144
rect 7910 1756 7916 2132
rect 7950 1756 7956 2132
rect 7910 1744 7956 1756
rect 8028 2132 8074 2144
rect 8028 1756 8034 2132
rect 8068 1756 8074 2132
rect 8028 1744 8074 1756
rect 8146 2132 8192 2144
rect 8146 1756 8152 2132
rect 8186 1756 8192 2132
rect 8146 1744 8192 1756
rect 8265 2132 8311 2144
rect 8265 1756 8271 2132
rect 8305 1756 8311 2132
rect 8265 1744 8311 1756
rect 8383 2132 8429 2144
rect 8383 1756 8389 2132
rect 8423 1756 8429 2132
rect 8383 1744 8429 1756
rect 8501 2132 8547 2144
rect 8501 1756 8507 2132
rect 8541 1756 8547 2132
rect 8501 1744 8547 1756
rect 8619 2132 8665 2144
rect 8619 1756 8625 2132
rect 8659 1756 8665 2132
rect 8743 1944 8780 2231
rect 8619 1744 8665 1756
rect 8738 1932 8784 1944
rect 8738 1756 8744 1932
rect 8778 1756 8784 1932
rect 8738 1744 8784 1756
rect 8856 1932 8902 1944
rect 8856 1756 8862 1932
rect 8896 1756 8902 1932
rect 8856 1744 8902 1756
rect 8974 1932 9020 1944
rect 8974 1756 8980 1932
rect 9014 1756 9020 1932
rect 8974 1744 9020 1756
rect 9092 1932 9138 1944
rect 9092 1756 9098 1932
rect 9132 1756 9138 1932
rect 9092 1744 9138 1756
rect 6535 1558 6570 1744
rect 7444 1660 7478 1744
rect 8625 1660 8659 1744
rect 7444 1618 8659 1660
rect 8625 1598 8659 1618
rect 8625 1582 8982 1598
rect 6535 1541 7672 1558
rect 6535 1507 7622 1541
rect 7656 1507 7672 1541
rect 8625 1548 8932 1582
rect 8966 1548 8982 1582
rect 8625 1532 8982 1548
rect 6535 1491 7672 1507
rect 6377 1446 6452 1454
rect 6377 1378 6393 1446
rect 6450 1378 6460 1446
rect 6377 1370 6452 1378
rect 6275 1330 6452 1338
rect 6275 1297 6393 1330
rect 6276 1262 6393 1297
rect 6450 1262 6460 1330
rect 6276 1254 6452 1262
rect 3403 930 4775 977
rect 5097 931 6149 978
rect 6535 981 6570 1491
rect 6625 1445 6717 1458
rect 6625 1382 6637 1445
rect 6708 1382 6717 1445
rect 6625 1373 6717 1382
rect 7710 1445 7802 1455
rect 7710 1383 7722 1445
rect 7792 1383 7802 1445
rect 7710 1370 7802 1383
rect 9098 1390 9133 1744
rect 9098 1352 9279 1390
rect 7957 1328 8022 1331
rect 7957 1325 8026 1328
rect 7957 1265 7963 1325
rect 8022 1265 8032 1325
rect 7957 1261 8026 1265
rect 7957 1259 8022 1261
rect 7592 1162 7684 1170
rect 7592 1097 7604 1162
rect 7672 1097 7684 1162
rect 7592 1085 7684 1097
rect 9098 982 9283 1352
rect 9419 1338 9487 2875
rect 28822 2856 28942 2875
rect 22290 2836 28557 2837
rect 12623 2772 28764 2836
rect 28826 2800 28942 2856
rect 12623 2767 28766 2772
rect 12623 2751 12690 2767
rect 12744 2766 28766 2767
rect 10918 2328 10928 2388
rect 11008 2328 11018 2388
rect 10918 2288 11018 2328
rect 10121 2231 11924 2288
rect 10121 2144 10155 2231
rect 11296 2144 11330 2231
rect 10115 2132 10161 2144
rect 10115 1944 10121 2132
rect 9674 1932 9720 1944
rect 9674 1756 9680 1932
rect 9714 1756 9720 1932
rect 9674 1744 9720 1756
rect 9792 1932 9838 1944
rect 9792 1756 9798 1932
rect 9832 1756 9838 1932
rect 9792 1744 9838 1756
rect 9910 1932 9956 1944
rect 9910 1756 9916 1932
rect 9950 1756 9956 1932
rect 9910 1744 9956 1756
rect 10028 1932 10121 1944
rect 10028 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10161 2132
rect 10028 1744 10161 1756
rect 10233 2132 10279 2144
rect 10233 1756 10239 2132
rect 10273 1756 10279 2132
rect 10233 1744 10279 1756
rect 10351 2132 10397 2144
rect 10351 1756 10357 2132
rect 10391 1756 10397 2132
rect 10351 1744 10397 1756
rect 10469 2132 10515 2144
rect 10469 1756 10475 2132
rect 10509 1756 10515 2132
rect 10469 1744 10515 1756
rect 10582 2132 10628 2144
rect 10582 1756 10588 2132
rect 10622 1756 10628 2132
rect 10582 1744 10628 1756
rect 10700 2132 10746 2144
rect 10700 1756 10706 2132
rect 10740 1756 10746 2132
rect 10700 1744 10746 1756
rect 10818 2132 10864 2144
rect 10818 1756 10824 2132
rect 10858 1756 10864 2132
rect 10818 1744 10864 1756
rect 10936 2132 10982 2144
rect 10936 1756 10942 2132
rect 10976 1756 10982 2132
rect 10936 1744 10982 1756
rect 11054 2132 11100 2144
rect 11054 1756 11060 2132
rect 11094 1756 11100 2132
rect 11054 1744 11100 1756
rect 11172 2132 11218 2144
rect 11172 1756 11178 2132
rect 11212 1756 11218 2132
rect 11172 1744 11218 1756
rect 11290 2132 11336 2144
rect 11290 1756 11296 2132
rect 11330 1756 11336 2132
rect 11290 1744 11336 1756
rect 11409 2132 11455 2144
rect 11409 1756 11415 2132
rect 11449 1756 11455 2132
rect 11409 1744 11455 1756
rect 11527 2132 11573 2144
rect 11527 1756 11533 2132
rect 11567 1756 11573 2132
rect 11527 1744 11573 1756
rect 11645 2132 11691 2144
rect 11645 1756 11651 2132
rect 11685 1756 11691 2132
rect 11645 1744 11691 1756
rect 11763 2132 11809 2144
rect 11763 1756 11769 2132
rect 11803 1756 11809 2132
rect 11887 1944 11924 2231
rect 11763 1744 11809 1756
rect 11882 1932 11928 1944
rect 11882 1756 11888 1932
rect 11922 1756 11928 1932
rect 11882 1744 11928 1756
rect 12000 1932 12046 1944
rect 12000 1756 12006 1932
rect 12040 1756 12046 1932
rect 12000 1744 12046 1756
rect 12118 1932 12164 1944
rect 12118 1756 12124 1932
rect 12158 1756 12164 1932
rect 12118 1744 12164 1756
rect 12236 1932 12282 1944
rect 12236 1756 12242 1932
rect 12276 1756 12282 1932
rect 12236 1744 12282 1756
rect 9679 1558 9714 1744
rect 10588 1660 10622 1744
rect 11769 1660 11803 1744
rect 10588 1618 11803 1660
rect 11769 1598 11803 1618
rect 11769 1582 12126 1598
rect 9679 1541 10816 1558
rect 9679 1507 10766 1541
rect 10800 1507 10816 1541
rect 11769 1548 12076 1582
rect 12110 1548 12126 1582
rect 11769 1532 12126 1548
rect 9679 1491 10816 1507
rect 9521 1446 9596 1454
rect 9521 1378 9537 1446
rect 9594 1378 9604 1446
rect 9521 1370 9596 1378
rect 9419 1330 9596 1338
rect 9419 1310 9537 1330
rect 9420 1262 9537 1310
rect 9594 1262 9604 1330
rect 9420 1254 9596 1262
rect 6535 934 7907 981
rect 8229 935 9283 982
rect 4237 807 4271 930
rect 4709 917 4775 930
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 5098 807 5132 931
rect 5980 925 6149 931
rect 4232 795 4278 807
rect 4232 619 4238 795
rect 4272 619 4278 795
rect 4232 607 4278 619
rect 4350 795 4470 807
rect 4350 619 4356 795
rect 4390 619 4430 795
rect 4350 607 4430 619
rect 4356 240 4390 607
rect 4424 419 4430 607
rect 4464 419 4470 795
rect 4424 407 4470 419
rect 4542 795 4588 807
rect 4542 419 4548 795
rect 4582 419 4588 795
rect 4542 407 4588 419
rect 4660 795 4706 807
rect 4660 419 4666 795
rect 4700 419 4706 795
rect 4660 407 4706 419
rect 4778 795 4824 807
rect 4778 419 4784 795
rect 4818 419 4824 795
rect 4778 407 4824 419
rect 4896 795 5020 807
rect 4896 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5020 795
rect 4936 607 5020 619
rect 5092 795 5138 807
rect 5092 619 5098 795
rect 5132 619 5138 795
rect 5092 607 5138 619
rect 4936 419 4942 607
rect 4896 407 4942 419
rect 4666 334 4700 407
rect 4651 318 4717 334
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 4651 268 4717 284
rect 4980 240 5014 607
rect 4356 188 5014 240
rect 4654 166 4746 188
rect 4654 114 4666 166
rect 4732 114 4746 166
rect 4654 110 4746 114
rect -64 -1188 3003 -1063
rect 3113 -1063 3215 -1062
rect 6003 -1063 6149 925
rect 7369 811 7403 934
rect 7841 921 7907 934
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 8230 811 8264 935
rect 7364 799 7410 811
rect 7364 623 7370 799
rect 7404 623 7410 799
rect 7364 611 7410 623
rect 7482 799 7602 811
rect 7482 623 7488 799
rect 7522 623 7562 799
rect 7482 611 7562 623
rect 7488 244 7522 611
rect 7556 423 7562 611
rect 7596 423 7602 799
rect 7556 411 7602 423
rect 7674 799 7720 811
rect 7674 423 7680 799
rect 7714 423 7720 799
rect 7674 411 7720 423
rect 7792 799 7838 811
rect 7792 423 7798 799
rect 7832 423 7838 799
rect 7792 411 7838 423
rect 7910 799 7956 811
rect 7910 423 7916 799
rect 7950 423 7956 799
rect 7910 411 7956 423
rect 8028 799 8152 811
rect 8028 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8152 799
rect 8068 611 8152 623
rect 8224 799 8270 811
rect 8224 623 8230 799
rect 8264 623 8270 799
rect 8224 611 8270 623
rect 8068 423 8074 611
rect 8028 411 8074 423
rect 7798 338 7832 411
rect 7783 322 7849 338
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 7783 272 7849 288
rect 8112 244 8146 611
rect 7488 192 8146 244
rect 7786 170 7878 192
rect 7786 118 7798 170
rect 7864 118 7878 170
rect 7786 114 7878 118
rect -63 -1192 2999 -1188
rect 3113 -1192 6149 -1063
rect 9137 -1066 9283 935
rect 9679 981 9714 1491
rect 9769 1445 9861 1458
rect 9769 1382 9781 1445
rect 9852 1382 9861 1445
rect 9769 1373 9861 1382
rect 10854 1445 10946 1455
rect 10854 1383 10866 1445
rect 10936 1383 10946 1445
rect 10854 1370 10946 1383
rect 12242 1390 12277 1744
rect 11101 1328 11166 1331
rect 11101 1325 11170 1328
rect 11101 1265 11107 1325
rect 11166 1265 11176 1325
rect 11101 1261 11170 1265
rect 11101 1259 11166 1261
rect 10736 1162 10828 1170
rect 10736 1097 10748 1162
rect 10816 1097 10828 1162
rect 10736 1085 10828 1097
rect 12242 982 12423 1390
rect 12622 1334 12690 2751
rect 15761 2735 21617 2736
rect 15761 2672 28582 2735
rect 14120 2324 14130 2384
rect 14210 2324 14220 2384
rect 14120 2284 14220 2324
rect 13323 2227 15126 2284
rect 13323 2140 13357 2227
rect 14498 2140 14532 2227
rect 13317 2128 13363 2140
rect 13317 1940 13323 2128
rect 12876 1928 12922 1940
rect 12876 1752 12882 1928
rect 12916 1752 12922 1928
rect 12876 1740 12922 1752
rect 12994 1928 13040 1940
rect 12994 1752 13000 1928
rect 13034 1752 13040 1928
rect 12994 1740 13040 1752
rect 13112 1928 13158 1940
rect 13112 1752 13118 1928
rect 13152 1752 13158 1928
rect 13112 1740 13158 1752
rect 13230 1928 13323 1940
rect 13230 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13363 2128
rect 13230 1740 13363 1752
rect 13435 2128 13481 2140
rect 13435 1752 13441 2128
rect 13475 1752 13481 2128
rect 13435 1740 13481 1752
rect 13553 2128 13599 2140
rect 13553 1752 13559 2128
rect 13593 1752 13599 2128
rect 13553 1740 13599 1752
rect 13671 2128 13717 2140
rect 13671 1752 13677 2128
rect 13711 1752 13717 2128
rect 13671 1740 13717 1752
rect 13784 2128 13830 2140
rect 13784 1752 13790 2128
rect 13824 1752 13830 2128
rect 13784 1740 13830 1752
rect 13902 2128 13948 2140
rect 13902 1752 13908 2128
rect 13942 1752 13948 2128
rect 13902 1740 13948 1752
rect 14020 2128 14066 2140
rect 14020 1752 14026 2128
rect 14060 1752 14066 2128
rect 14020 1740 14066 1752
rect 14138 2128 14184 2140
rect 14138 1752 14144 2128
rect 14178 1752 14184 2128
rect 14138 1740 14184 1752
rect 14256 2128 14302 2140
rect 14256 1752 14262 2128
rect 14296 1752 14302 2128
rect 14256 1740 14302 1752
rect 14374 2128 14420 2140
rect 14374 1752 14380 2128
rect 14414 1752 14420 2128
rect 14374 1740 14420 1752
rect 14492 2128 14538 2140
rect 14492 1752 14498 2128
rect 14532 1752 14538 2128
rect 14492 1740 14538 1752
rect 14611 2128 14657 2140
rect 14611 1752 14617 2128
rect 14651 1752 14657 2128
rect 14611 1740 14657 1752
rect 14729 2128 14775 2140
rect 14729 1752 14735 2128
rect 14769 1752 14775 2128
rect 14729 1740 14775 1752
rect 14847 2128 14893 2140
rect 14847 1752 14853 2128
rect 14887 1752 14893 2128
rect 14847 1740 14893 1752
rect 14965 2128 15011 2140
rect 14965 1752 14971 2128
rect 15005 1752 15011 2128
rect 15089 1940 15126 2227
rect 14965 1740 15011 1752
rect 15084 1928 15130 1940
rect 15084 1752 15090 1928
rect 15124 1752 15130 1928
rect 15084 1740 15130 1752
rect 15202 1928 15248 1940
rect 15202 1752 15208 1928
rect 15242 1752 15248 1928
rect 15202 1740 15248 1752
rect 15320 1928 15366 1940
rect 15320 1752 15326 1928
rect 15360 1752 15366 1928
rect 15320 1740 15366 1752
rect 15438 1928 15484 1940
rect 15438 1752 15444 1928
rect 15478 1752 15484 1928
rect 15438 1740 15484 1752
rect 12881 1554 12916 1740
rect 13790 1656 13824 1740
rect 14971 1656 15005 1740
rect 13790 1614 15005 1656
rect 14971 1594 15005 1614
rect 14971 1578 15328 1594
rect 12881 1537 14018 1554
rect 12881 1503 13968 1537
rect 14002 1503 14018 1537
rect 14971 1544 15278 1578
rect 15312 1544 15328 1578
rect 14971 1528 15328 1544
rect 12881 1487 14018 1503
rect 12725 1442 12798 1450
rect 12725 1374 12739 1442
rect 12796 1374 12806 1442
rect 12725 1366 12798 1374
rect 12622 1326 12798 1334
rect 12622 1258 12739 1326
rect 12796 1258 12806 1326
rect 12622 1250 12798 1258
rect 9679 934 11051 981
rect 11373 935 12423 982
rect 10513 811 10547 934
rect 10985 921 11051 934
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 11374 811 11408 935
rect 10508 799 10554 811
rect 10508 623 10514 799
rect 10548 623 10554 799
rect 10508 611 10554 623
rect 10626 799 10746 811
rect 10626 623 10632 799
rect 10666 623 10706 799
rect 10626 611 10706 623
rect 10632 244 10666 611
rect 10700 423 10706 611
rect 10740 423 10746 799
rect 10700 411 10746 423
rect 10818 799 10864 811
rect 10818 423 10824 799
rect 10858 423 10864 799
rect 10818 411 10864 423
rect 10936 799 10982 811
rect 10936 423 10942 799
rect 10976 423 10982 799
rect 10936 411 10982 423
rect 11054 799 11100 811
rect 11054 423 11060 799
rect 11094 423 11100 799
rect 11054 411 11100 423
rect 11172 799 11296 811
rect 11172 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11296 799
rect 11212 611 11296 623
rect 11368 799 11414 811
rect 11368 623 11374 799
rect 11408 623 11414 799
rect 11368 611 11414 623
rect 11212 423 11218 611
rect 11172 411 11218 423
rect 10942 338 10976 411
rect 10927 322 10993 338
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 10927 272 10993 288
rect 11256 244 11290 611
rect 10632 192 11290 244
rect 10930 170 11022 192
rect 10930 118 10942 170
rect 11008 118 11022 170
rect 10930 114 11022 118
rect 12277 -1060 12423 935
rect 12881 977 12916 1487
rect 12971 1441 13063 1454
rect 12971 1378 12983 1441
rect 13054 1378 13063 1441
rect 12971 1369 13063 1378
rect 14056 1441 14148 1451
rect 14056 1379 14068 1441
rect 14138 1379 14148 1441
rect 14056 1366 14148 1379
rect 15444 1386 15479 1740
rect 14303 1324 14368 1327
rect 14303 1321 14372 1324
rect 14303 1261 14309 1321
rect 14368 1261 14378 1321
rect 14303 1257 14372 1261
rect 14303 1255 14368 1257
rect 15444 1240 15625 1386
rect 15761 1334 15829 2672
rect 18896 2632 21309 2637
rect 18896 2621 28425 2632
rect 18895 2581 28425 2621
rect 18895 2550 18965 2581
rect 28308 2569 28425 2581
rect 17264 2324 17274 2384
rect 17354 2324 17364 2384
rect 17264 2284 17364 2324
rect 16467 2227 18270 2284
rect 16467 2140 16501 2227
rect 17642 2140 17676 2227
rect 16461 2128 16507 2140
rect 16461 1940 16467 2128
rect 16020 1928 16066 1940
rect 16020 1752 16026 1928
rect 16060 1752 16066 1928
rect 16020 1740 16066 1752
rect 16138 1928 16184 1940
rect 16138 1752 16144 1928
rect 16178 1752 16184 1928
rect 16138 1740 16184 1752
rect 16256 1928 16302 1940
rect 16256 1752 16262 1928
rect 16296 1752 16302 1928
rect 16256 1740 16302 1752
rect 16374 1928 16467 1940
rect 16374 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16507 2128
rect 16374 1740 16507 1752
rect 16579 2128 16625 2140
rect 16579 1752 16585 2128
rect 16619 1752 16625 2128
rect 16579 1740 16625 1752
rect 16697 2128 16743 2140
rect 16697 1752 16703 2128
rect 16737 1752 16743 2128
rect 16697 1740 16743 1752
rect 16815 2128 16861 2140
rect 16815 1752 16821 2128
rect 16855 1752 16861 2128
rect 16815 1740 16861 1752
rect 16928 2128 16974 2140
rect 16928 1752 16934 2128
rect 16968 1752 16974 2128
rect 16928 1740 16974 1752
rect 17046 2128 17092 2140
rect 17046 1752 17052 2128
rect 17086 1752 17092 2128
rect 17046 1740 17092 1752
rect 17164 2128 17210 2140
rect 17164 1752 17170 2128
rect 17204 1752 17210 2128
rect 17164 1740 17210 1752
rect 17282 2128 17328 2140
rect 17282 1752 17288 2128
rect 17322 1752 17328 2128
rect 17282 1740 17328 1752
rect 17400 2128 17446 2140
rect 17400 1752 17406 2128
rect 17440 1752 17446 2128
rect 17400 1740 17446 1752
rect 17518 2128 17564 2140
rect 17518 1752 17524 2128
rect 17558 1752 17564 2128
rect 17518 1740 17564 1752
rect 17636 2128 17682 2140
rect 17636 1752 17642 2128
rect 17676 1752 17682 2128
rect 17636 1740 17682 1752
rect 17755 2128 17801 2140
rect 17755 1752 17761 2128
rect 17795 1752 17801 2128
rect 17755 1740 17801 1752
rect 17873 2128 17919 2140
rect 17873 1752 17879 2128
rect 17913 1752 17919 2128
rect 17873 1740 17919 1752
rect 17991 2128 18037 2140
rect 17991 1752 17997 2128
rect 18031 1752 18037 2128
rect 17991 1740 18037 1752
rect 18109 2128 18155 2140
rect 18109 1752 18115 2128
rect 18149 1752 18155 2128
rect 18233 1940 18270 2227
rect 18109 1740 18155 1752
rect 18228 1928 18274 1940
rect 18228 1752 18234 1928
rect 18268 1752 18274 1928
rect 18228 1740 18274 1752
rect 18346 1928 18392 1940
rect 18346 1752 18352 1928
rect 18386 1752 18392 1928
rect 18346 1740 18392 1752
rect 18464 1928 18510 1940
rect 18464 1752 18470 1928
rect 18504 1752 18510 1928
rect 18464 1740 18510 1752
rect 18582 1928 18628 1940
rect 18582 1752 18588 1928
rect 18622 1752 18628 1928
rect 18582 1740 18628 1752
rect 16025 1554 16060 1740
rect 16934 1656 16968 1740
rect 18115 1656 18149 1740
rect 16934 1614 18149 1656
rect 18115 1594 18149 1614
rect 18115 1578 18472 1594
rect 16025 1537 17162 1554
rect 16025 1503 17112 1537
rect 17146 1503 17162 1537
rect 18115 1544 18422 1578
rect 18456 1544 18472 1578
rect 18115 1528 18472 1544
rect 16025 1487 17162 1503
rect 15868 1442 15942 1450
rect 15868 1374 15883 1442
rect 15940 1374 15950 1442
rect 15868 1366 15942 1374
rect 15761 1326 15942 1334
rect 15761 1258 15883 1326
rect 15940 1258 15950 1326
rect 15761 1250 15942 1258
rect 15761 1249 15795 1250
rect 13938 1158 14030 1166
rect 13938 1093 13950 1158
rect 14018 1093 14030 1158
rect 13938 1081 14030 1093
rect 15444 978 15620 1240
rect 12881 930 14253 977
rect 14575 931 15620 978
rect 13715 807 13749 930
rect 14187 917 14253 930
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14576 807 14610 931
rect 13710 795 13756 807
rect 13710 619 13716 795
rect 13750 619 13756 795
rect 13710 607 13756 619
rect 13828 795 13948 807
rect 13828 619 13834 795
rect 13868 619 13908 795
rect 13828 607 13908 619
rect 13834 240 13868 607
rect 13902 419 13908 607
rect 13942 419 13948 795
rect 13902 407 13948 419
rect 14020 795 14066 807
rect 14020 419 14026 795
rect 14060 419 14066 795
rect 14020 407 14066 419
rect 14138 795 14184 807
rect 14138 419 14144 795
rect 14178 419 14184 795
rect 14138 407 14184 419
rect 14256 795 14302 807
rect 14256 419 14262 795
rect 14296 419 14302 795
rect 14256 407 14302 419
rect 14374 795 14498 807
rect 14374 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14498 795
rect 14414 607 14498 619
rect 14570 795 14616 807
rect 14570 619 14576 795
rect 14610 619 14616 795
rect 14570 607 14616 619
rect 14414 419 14420 607
rect 14374 407 14420 419
rect 14144 334 14178 407
rect 14129 318 14195 334
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 14129 268 14195 284
rect 14458 240 14492 607
rect 13834 188 14492 240
rect 14132 166 14224 188
rect 14132 114 14144 166
rect 14210 114 14224 166
rect 14132 110 14224 114
rect -63 -2558 41 -1192
rect 1530 -1568 1540 -1508
rect 1620 -1568 1630 -1508
rect 1530 -1608 1630 -1568
rect 733 -1665 2536 -1608
rect 733 -1752 767 -1665
rect 1908 -1752 1942 -1665
rect 727 -1764 773 -1752
rect 727 -1952 733 -1764
rect 286 -1964 332 -1952
rect 286 -2140 292 -1964
rect 326 -2140 332 -1964
rect 286 -2152 332 -2140
rect 404 -1964 450 -1952
rect 404 -2140 410 -1964
rect 444 -2140 450 -1964
rect 404 -2152 450 -2140
rect 522 -1964 568 -1952
rect 522 -2140 528 -1964
rect 562 -2140 568 -1964
rect 522 -2152 568 -2140
rect 640 -1964 733 -1952
rect 640 -2140 646 -1964
rect 680 -2140 733 -1964
rect 767 -2140 773 -1764
rect 640 -2152 773 -2140
rect 845 -1764 891 -1752
rect 845 -2140 851 -1764
rect 885 -2140 891 -1764
rect 845 -2152 891 -2140
rect 963 -1764 1009 -1752
rect 963 -2140 969 -1764
rect 1003 -2140 1009 -1764
rect 963 -2152 1009 -2140
rect 1081 -1764 1127 -1752
rect 1081 -2140 1087 -1764
rect 1121 -2140 1127 -1764
rect 1081 -2152 1127 -2140
rect 1194 -1764 1240 -1752
rect 1194 -2140 1200 -1764
rect 1234 -2140 1240 -1764
rect 1194 -2152 1240 -2140
rect 1312 -1764 1358 -1752
rect 1312 -2140 1318 -1764
rect 1352 -2140 1358 -1764
rect 1312 -2152 1358 -2140
rect 1430 -1764 1476 -1752
rect 1430 -2140 1436 -1764
rect 1470 -2140 1476 -1764
rect 1430 -2152 1476 -2140
rect 1548 -1764 1594 -1752
rect 1548 -2140 1554 -1764
rect 1588 -2140 1594 -1764
rect 1548 -2152 1594 -2140
rect 1666 -1764 1712 -1752
rect 1666 -2140 1672 -1764
rect 1706 -2140 1712 -1764
rect 1666 -2152 1712 -2140
rect 1784 -1764 1830 -1752
rect 1784 -2140 1790 -1764
rect 1824 -2140 1830 -1764
rect 1784 -2152 1830 -2140
rect 1902 -1764 1948 -1752
rect 1902 -2140 1908 -1764
rect 1942 -2140 1948 -1764
rect 1902 -2152 1948 -2140
rect 2021 -1764 2067 -1752
rect 2021 -2140 2027 -1764
rect 2061 -2140 2067 -1764
rect 2021 -2152 2067 -2140
rect 2139 -1764 2185 -1752
rect 2139 -2140 2145 -1764
rect 2179 -2140 2185 -1764
rect 2139 -2152 2185 -2140
rect 2257 -1764 2303 -1752
rect 2257 -2140 2263 -1764
rect 2297 -2140 2303 -1764
rect 2257 -2152 2303 -2140
rect 2375 -1764 2421 -1752
rect 2375 -2140 2381 -1764
rect 2415 -2140 2421 -1764
rect 2499 -1952 2536 -1665
rect 2375 -2152 2421 -2140
rect 2494 -1964 2540 -1952
rect 2494 -2140 2500 -1964
rect 2534 -2140 2540 -1964
rect 2494 -2152 2540 -2140
rect 2612 -1964 2658 -1952
rect 2612 -2140 2618 -1964
rect 2652 -2140 2658 -1964
rect 2612 -2152 2658 -2140
rect 2730 -1964 2776 -1952
rect 2730 -2140 2736 -1964
rect 2770 -2140 2776 -1964
rect 2730 -2152 2776 -2140
rect 2848 -1964 2894 -1952
rect 2848 -2140 2854 -1964
rect 2888 -2140 2894 -1964
rect 2848 -2152 2894 -2140
rect 291 -2338 326 -2152
rect 1200 -2236 1234 -2152
rect 2381 -2236 2415 -2152
rect 1200 -2278 2415 -2236
rect 2381 -2298 2415 -2278
rect 2381 -2314 2738 -2298
rect 291 -2355 1428 -2338
rect 291 -2389 1378 -2355
rect 1412 -2389 1428 -2355
rect 2381 -2348 2688 -2314
rect 2722 -2348 2738 -2314
rect 2381 -2364 2738 -2348
rect 291 -2405 1428 -2389
rect 132 -2450 208 -2442
rect 132 -2518 149 -2450
rect 206 -2518 216 -2450
rect 132 -2526 208 -2518
rect -63 -2566 208 -2558
rect -63 -2634 149 -2566
rect 206 -2634 216 -2566
rect -63 -2642 208 -2634
rect -63 -2643 41 -2642
rect 291 -2915 326 -2405
rect 381 -2451 473 -2438
rect 381 -2514 393 -2451
rect 464 -2514 473 -2451
rect 381 -2523 473 -2514
rect 1466 -2451 1558 -2441
rect 1466 -2513 1478 -2451
rect 1548 -2513 1558 -2451
rect 1466 -2526 1558 -2513
rect 2854 -2506 2889 -2152
rect 2854 -2532 3035 -2506
rect 1713 -2568 1778 -2565
rect 1713 -2571 1782 -2568
rect 1713 -2631 1719 -2571
rect 1778 -2631 1788 -2571
rect 1713 -2635 1782 -2631
rect 1713 -2637 1778 -2635
rect 1348 -2734 1440 -2726
rect 1348 -2799 1360 -2734
rect 1428 -2799 1440 -2734
rect 1348 -2811 1440 -2799
rect 2854 -2914 3039 -2532
rect 3113 -2558 3217 -1192
rect 6003 -1198 6149 -1192
rect 6249 -1193 9283 -1066
rect 9374 -1189 12423 -1060
rect 6249 -1195 9275 -1193
rect 4674 -1568 4684 -1508
rect 4764 -1568 4774 -1508
rect 4674 -1608 4774 -1568
rect 3877 -1665 5680 -1608
rect 3877 -1752 3911 -1665
rect 5052 -1752 5086 -1665
rect 3871 -1764 3917 -1752
rect 3871 -1952 3877 -1764
rect 3430 -1964 3476 -1952
rect 3430 -2140 3436 -1964
rect 3470 -2140 3476 -1964
rect 3430 -2152 3476 -2140
rect 3548 -1964 3594 -1952
rect 3548 -2140 3554 -1964
rect 3588 -2140 3594 -1964
rect 3548 -2152 3594 -2140
rect 3666 -1964 3712 -1952
rect 3666 -2140 3672 -1964
rect 3706 -2140 3712 -1964
rect 3666 -2152 3712 -2140
rect 3784 -1964 3877 -1952
rect 3784 -2140 3790 -1964
rect 3824 -2140 3877 -1964
rect 3911 -2140 3917 -1764
rect 3784 -2152 3917 -2140
rect 3989 -1764 4035 -1752
rect 3989 -2140 3995 -1764
rect 4029 -2140 4035 -1764
rect 3989 -2152 4035 -2140
rect 4107 -1764 4153 -1752
rect 4107 -2140 4113 -1764
rect 4147 -2140 4153 -1764
rect 4107 -2152 4153 -2140
rect 4225 -1764 4271 -1752
rect 4225 -2140 4231 -1764
rect 4265 -2140 4271 -1764
rect 4225 -2152 4271 -2140
rect 4338 -1764 4384 -1752
rect 4338 -2140 4344 -1764
rect 4378 -2140 4384 -1764
rect 4338 -2152 4384 -2140
rect 4456 -1764 4502 -1752
rect 4456 -2140 4462 -1764
rect 4496 -2140 4502 -1764
rect 4456 -2152 4502 -2140
rect 4574 -1764 4620 -1752
rect 4574 -2140 4580 -1764
rect 4614 -2140 4620 -1764
rect 4574 -2152 4620 -2140
rect 4692 -1764 4738 -1752
rect 4692 -2140 4698 -1764
rect 4732 -2140 4738 -1764
rect 4692 -2152 4738 -2140
rect 4810 -1764 4856 -1752
rect 4810 -2140 4816 -1764
rect 4850 -2140 4856 -1764
rect 4810 -2152 4856 -2140
rect 4928 -1764 4974 -1752
rect 4928 -2140 4934 -1764
rect 4968 -2140 4974 -1764
rect 4928 -2152 4974 -2140
rect 5046 -1764 5092 -1752
rect 5046 -2140 5052 -1764
rect 5086 -2140 5092 -1764
rect 5046 -2152 5092 -2140
rect 5165 -1764 5211 -1752
rect 5165 -2140 5171 -1764
rect 5205 -2140 5211 -1764
rect 5165 -2152 5211 -2140
rect 5283 -1764 5329 -1752
rect 5283 -2140 5289 -1764
rect 5323 -2140 5329 -1764
rect 5283 -2152 5329 -2140
rect 5401 -1764 5447 -1752
rect 5401 -2140 5407 -1764
rect 5441 -2140 5447 -1764
rect 5401 -2152 5447 -2140
rect 5519 -1764 5565 -1752
rect 5519 -2140 5525 -1764
rect 5559 -2140 5565 -1764
rect 5643 -1952 5680 -1665
rect 5519 -2152 5565 -2140
rect 5638 -1964 5684 -1952
rect 5638 -2140 5644 -1964
rect 5678 -2140 5684 -1964
rect 5638 -2152 5684 -2140
rect 5756 -1964 5802 -1952
rect 5756 -2140 5762 -1964
rect 5796 -2140 5802 -1964
rect 5756 -2152 5802 -2140
rect 5874 -1964 5920 -1952
rect 5874 -2140 5880 -1964
rect 5914 -2140 5920 -1964
rect 5874 -2152 5920 -2140
rect 5992 -1964 6038 -1952
rect 5992 -2140 5998 -1964
rect 6032 -2140 6038 -1964
rect 5992 -2152 6038 -2140
rect 3435 -2338 3470 -2152
rect 4344 -2236 4378 -2152
rect 5525 -2236 5559 -2152
rect 4344 -2278 5559 -2236
rect 5525 -2298 5559 -2278
rect 5525 -2314 5882 -2298
rect 3435 -2355 4572 -2338
rect 3435 -2389 4522 -2355
rect 4556 -2389 4572 -2355
rect 5525 -2348 5832 -2314
rect 5866 -2348 5882 -2314
rect 5525 -2364 5882 -2348
rect 3435 -2405 4572 -2389
rect 3276 -2450 3352 -2442
rect 3276 -2518 3293 -2450
rect 3350 -2518 3360 -2450
rect 3276 -2526 3352 -2518
rect 3113 -2566 3352 -2558
rect 3113 -2634 3293 -2566
rect 3350 -2634 3360 -2566
rect 3113 -2641 3352 -2634
rect 3176 -2642 3352 -2641
rect 291 -2962 1663 -2915
rect 1985 -2961 3039 -2914
rect 1125 -3085 1159 -2962
rect 1597 -2975 1663 -2962
rect 1597 -3009 1613 -2975
rect 1647 -3009 1663 -2975
rect 1597 -3025 1663 -3009
rect 1986 -3085 2020 -2961
rect 1120 -3097 1166 -3085
rect 1120 -3273 1126 -3097
rect 1160 -3273 1166 -3097
rect 1120 -3285 1166 -3273
rect 1238 -3097 1358 -3085
rect 1238 -3273 1244 -3097
rect 1278 -3273 1318 -3097
rect 1238 -3285 1318 -3273
rect 1244 -3652 1278 -3285
rect 1312 -3473 1318 -3285
rect 1352 -3473 1358 -3097
rect 1312 -3485 1358 -3473
rect 1430 -3097 1476 -3085
rect 1430 -3473 1436 -3097
rect 1470 -3473 1476 -3097
rect 1430 -3485 1476 -3473
rect 1548 -3097 1594 -3085
rect 1548 -3473 1554 -3097
rect 1588 -3473 1594 -3097
rect 1548 -3485 1594 -3473
rect 1666 -3097 1712 -3085
rect 1666 -3473 1672 -3097
rect 1706 -3473 1712 -3097
rect 1666 -3485 1712 -3473
rect 1784 -3097 1908 -3085
rect 1784 -3473 1790 -3097
rect 1824 -3273 1868 -3097
rect 1902 -3273 1908 -3097
rect 1824 -3285 1908 -3273
rect 1980 -3097 2026 -3085
rect 1980 -3273 1986 -3097
rect 2020 -3273 2026 -3097
rect 1980 -3285 2026 -3273
rect 1824 -3473 1830 -3285
rect 1784 -3485 1830 -3473
rect 1554 -3558 1588 -3485
rect 1539 -3574 1605 -3558
rect 1539 -3608 1555 -3574
rect 1589 -3608 1605 -3574
rect 1539 -3624 1605 -3608
rect 1868 -3652 1902 -3285
rect 1244 -3704 1902 -3652
rect 1542 -3726 1634 -3704
rect 1542 -3778 1554 -3726
rect 1620 -3778 1634 -3726
rect 1542 -3782 1634 -3778
rect 2889 -4497 3039 -2961
rect 3435 -2915 3470 -2405
rect 3525 -2451 3617 -2438
rect 3525 -2514 3537 -2451
rect 3608 -2514 3617 -2451
rect 3525 -2523 3617 -2514
rect 4610 -2451 4702 -2441
rect 4610 -2513 4622 -2451
rect 4692 -2513 4702 -2451
rect 4610 -2526 4702 -2513
rect 5998 -2506 6033 -2152
rect 4857 -2568 4922 -2565
rect 4857 -2571 4926 -2568
rect 4857 -2631 4863 -2571
rect 4922 -2631 4932 -2571
rect 5998 -2596 6179 -2506
rect 6249 -2554 6353 -1195
rect 7806 -1564 7816 -1504
rect 7896 -1564 7906 -1504
rect 7806 -1604 7906 -1564
rect 7009 -1661 8812 -1604
rect 7009 -1748 7043 -1661
rect 8184 -1748 8218 -1661
rect 7003 -1760 7049 -1748
rect 7003 -1948 7009 -1760
rect 6562 -1960 6608 -1948
rect 6562 -2136 6568 -1960
rect 6602 -2136 6608 -1960
rect 6562 -2148 6608 -2136
rect 6680 -1960 6726 -1948
rect 6680 -2136 6686 -1960
rect 6720 -2136 6726 -1960
rect 6680 -2148 6726 -2136
rect 6798 -1960 6844 -1948
rect 6798 -2136 6804 -1960
rect 6838 -2136 6844 -1960
rect 6798 -2148 6844 -2136
rect 6916 -1960 7009 -1948
rect 6916 -2136 6922 -1960
rect 6956 -2136 7009 -1960
rect 7043 -2136 7049 -1760
rect 6916 -2148 7049 -2136
rect 7121 -1760 7167 -1748
rect 7121 -2136 7127 -1760
rect 7161 -2136 7167 -1760
rect 7121 -2148 7167 -2136
rect 7239 -1760 7285 -1748
rect 7239 -2136 7245 -1760
rect 7279 -2136 7285 -1760
rect 7239 -2148 7285 -2136
rect 7357 -1760 7403 -1748
rect 7357 -2136 7363 -1760
rect 7397 -2136 7403 -1760
rect 7357 -2148 7403 -2136
rect 7470 -1760 7516 -1748
rect 7470 -2136 7476 -1760
rect 7510 -2136 7516 -1760
rect 7470 -2148 7516 -2136
rect 7588 -1760 7634 -1748
rect 7588 -2136 7594 -1760
rect 7628 -2136 7634 -1760
rect 7588 -2148 7634 -2136
rect 7706 -1760 7752 -1748
rect 7706 -2136 7712 -1760
rect 7746 -2136 7752 -1760
rect 7706 -2148 7752 -2136
rect 7824 -1760 7870 -1748
rect 7824 -2136 7830 -1760
rect 7864 -2136 7870 -1760
rect 7824 -2148 7870 -2136
rect 7942 -1760 7988 -1748
rect 7942 -2136 7948 -1760
rect 7982 -2136 7988 -1760
rect 7942 -2148 7988 -2136
rect 8060 -1760 8106 -1748
rect 8060 -2136 8066 -1760
rect 8100 -2136 8106 -1760
rect 8060 -2148 8106 -2136
rect 8178 -1760 8224 -1748
rect 8178 -2136 8184 -1760
rect 8218 -2136 8224 -1760
rect 8178 -2148 8224 -2136
rect 8297 -1760 8343 -1748
rect 8297 -2136 8303 -1760
rect 8337 -2136 8343 -1760
rect 8297 -2148 8343 -2136
rect 8415 -1760 8461 -1748
rect 8415 -2136 8421 -1760
rect 8455 -2136 8461 -1760
rect 8415 -2148 8461 -2136
rect 8533 -1760 8579 -1748
rect 8533 -2136 8539 -1760
rect 8573 -2136 8579 -1760
rect 8533 -2148 8579 -2136
rect 8651 -1760 8697 -1748
rect 8651 -2136 8657 -1760
rect 8691 -2136 8697 -1760
rect 8775 -1948 8812 -1661
rect 8651 -2148 8697 -2136
rect 8770 -1960 8816 -1948
rect 8770 -2136 8776 -1960
rect 8810 -2136 8816 -1960
rect 8770 -2148 8816 -2136
rect 8888 -1960 8934 -1948
rect 8888 -2136 8894 -1960
rect 8928 -2136 8934 -1960
rect 8888 -2148 8934 -2136
rect 9006 -1960 9052 -1948
rect 9006 -2136 9012 -1960
rect 9046 -2136 9052 -1960
rect 9006 -2148 9052 -2136
rect 9124 -1960 9170 -1948
rect 9124 -2136 9130 -1960
rect 9164 -2136 9170 -1960
rect 9124 -2148 9170 -2136
rect 6567 -2334 6602 -2148
rect 7476 -2232 7510 -2148
rect 8657 -2232 8691 -2148
rect 7476 -2274 8691 -2232
rect 8657 -2294 8691 -2274
rect 8657 -2310 9014 -2294
rect 6567 -2351 7704 -2334
rect 6567 -2385 7654 -2351
rect 7688 -2385 7704 -2351
rect 8657 -2344 8964 -2310
rect 8998 -2344 9014 -2310
rect 8657 -2360 9014 -2344
rect 6567 -2401 7704 -2385
rect 6406 -2446 6484 -2438
rect 6406 -2514 6425 -2446
rect 6482 -2514 6492 -2446
rect 6406 -2522 6484 -2514
rect 6249 -2562 6484 -2554
rect 4857 -2635 4926 -2631
rect 4857 -2637 4922 -2635
rect 4492 -2734 4584 -2726
rect 4492 -2799 4504 -2734
rect 4572 -2799 4584 -2734
rect 4492 -2811 4584 -2799
rect 5998 -2914 6182 -2596
rect 6249 -2630 6425 -2562
rect 6482 -2630 6492 -2562
rect 6249 -2638 6484 -2630
rect 6249 -2641 6353 -2638
rect 3435 -2962 4807 -2915
rect 5129 -2961 6182 -2914
rect 6567 -2911 6602 -2401
rect 6657 -2447 6749 -2434
rect 6657 -2510 6669 -2447
rect 6740 -2510 6749 -2447
rect 6657 -2519 6749 -2510
rect 7742 -2447 7834 -2437
rect 7742 -2509 7754 -2447
rect 7824 -2509 7834 -2447
rect 7742 -2522 7834 -2509
rect 9130 -2502 9165 -2148
rect 7989 -2564 8054 -2561
rect 7989 -2567 8058 -2564
rect 7989 -2627 7995 -2567
rect 8054 -2627 8064 -2567
rect 9130 -2591 9311 -2502
rect 9374 -2554 9478 -1189
rect 12277 -1198 12423 -1189
rect 12585 -1060 12697 -1059
rect 15474 -1060 15620 931
rect 16025 977 16060 1487
rect 16115 1441 16207 1454
rect 16115 1378 16127 1441
rect 16198 1378 16207 1441
rect 16115 1369 16207 1378
rect 17200 1441 17292 1451
rect 17200 1379 17212 1441
rect 17282 1379 17292 1441
rect 17200 1366 17292 1379
rect 18588 1386 18623 1740
rect 18588 1352 18769 1386
rect 17447 1324 17512 1327
rect 17447 1321 17516 1324
rect 17447 1261 17453 1321
rect 17512 1261 17522 1321
rect 17447 1257 17516 1261
rect 17447 1255 17512 1257
rect 17082 1158 17174 1166
rect 17082 1093 17094 1158
rect 17162 1093 17174 1158
rect 17082 1081 17174 1093
rect 18588 978 18771 1352
rect 18895 1338 18966 2550
rect 22041 2495 28255 2547
rect 22041 2452 22116 2495
rect 28136 2493 28255 2495
rect 20396 2328 20406 2388
rect 20486 2328 20496 2388
rect 20396 2288 20496 2328
rect 19599 2231 21402 2288
rect 19599 2144 19633 2231
rect 20774 2144 20808 2231
rect 19593 2132 19639 2144
rect 19593 1944 19599 2132
rect 19152 1932 19198 1944
rect 19152 1756 19158 1932
rect 19192 1756 19198 1932
rect 19152 1744 19198 1756
rect 19270 1932 19316 1944
rect 19270 1756 19276 1932
rect 19310 1756 19316 1932
rect 19270 1744 19316 1756
rect 19388 1932 19434 1944
rect 19388 1756 19394 1932
rect 19428 1756 19434 1932
rect 19388 1744 19434 1756
rect 19506 1932 19599 1944
rect 19506 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19639 2132
rect 19506 1744 19639 1756
rect 19711 2132 19757 2144
rect 19711 1756 19717 2132
rect 19751 1756 19757 2132
rect 19711 1744 19757 1756
rect 19829 2132 19875 2144
rect 19829 1756 19835 2132
rect 19869 1756 19875 2132
rect 19829 1744 19875 1756
rect 19947 2132 19993 2144
rect 19947 1756 19953 2132
rect 19987 1756 19993 2132
rect 19947 1744 19993 1756
rect 20060 2132 20106 2144
rect 20060 1756 20066 2132
rect 20100 1756 20106 2132
rect 20060 1744 20106 1756
rect 20178 2132 20224 2144
rect 20178 1756 20184 2132
rect 20218 1756 20224 2132
rect 20178 1744 20224 1756
rect 20296 2132 20342 2144
rect 20296 1756 20302 2132
rect 20336 1756 20342 2132
rect 20296 1744 20342 1756
rect 20414 2132 20460 2144
rect 20414 1756 20420 2132
rect 20454 1756 20460 2132
rect 20414 1744 20460 1756
rect 20532 2132 20578 2144
rect 20532 1756 20538 2132
rect 20572 1756 20578 2132
rect 20532 1744 20578 1756
rect 20650 2132 20696 2144
rect 20650 1756 20656 2132
rect 20690 1756 20696 2132
rect 20650 1744 20696 1756
rect 20768 2132 20814 2144
rect 20768 1756 20774 2132
rect 20808 1756 20814 2132
rect 20768 1744 20814 1756
rect 20887 2132 20933 2144
rect 20887 1756 20893 2132
rect 20927 1756 20933 2132
rect 20887 1744 20933 1756
rect 21005 2132 21051 2144
rect 21005 1756 21011 2132
rect 21045 1756 21051 2132
rect 21005 1744 21051 1756
rect 21123 2132 21169 2144
rect 21123 1756 21129 2132
rect 21163 1756 21169 2132
rect 21123 1744 21169 1756
rect 21241 2132 21287 2144
rect 21241 1756 21247 2132
rect 21281 1756 21287 2132
rect 21365 1944 21402 2231
rect 21241 1744 21287 1756
rect 21360 1932 21406 1944
rect 21360 1756 21366 1932
rect 21400 1756 21406 1932
rect 21360 1744 21406 1756
rect 21478 1932 21524 1944
rect 21478 1756 21484 1932
rect 21518 1756 21524 1932
rect 21478 1744 21524 1756
rect 21596 1932 21642 1944
rect 21596 1756 21602 1932
rect 21636 1756 21642 1932
rect 21596 1744 21642 1756
rect 21714 1932 21760 1944
rect 21714 1756 21720 1932
rect 21754 1756 21760 1932
rect 21714 1744 21760 1756
rect 19157 1558 19192 1744
rect 20066 1660 20100 1744
rect 21247 1660 21281 1744
rect 20066 1618 21281 1660
rect 21247 1598 21281 1618
rect 21247 1582 21604 1598
rect 19157 1541 20294 1558
rect 19157 1507 20244 1541
rect 20278 1507 20294 1541
rect 21247 1548 21554 1582
rect 21588 1548 21604 1582
rect 21247 1532 21604 1548
rect 19157 1491 20294 1507
rect 18995 1446 19074 1454
rect 18995 1378 19015 1446
rect 19072 1378 19082 1446
rect 18995 1370 19074 1378
rect 18895 1330 19074 1338
rect 18895 1262 19015 1330
rect 19072 1262 19082 1330
rect 18895 1254 19074 1262
rect 16025 930 17397 977
rect 17719 931 18771 978
rect 19157 981 19192 1491
rect 19247 1445 19339 1458
rect 19247 1382 19259 1445
rect 19330 1382 19339 1445
rect 19247 1373 19339 1382
rect 20332 1445 20424 1455
rect 20332 1383 20344 1445
rect 20414 1383 20424 1445
rect 20332 1370 20424 1383
rect 21720 1390 21755 1744
rect 21720 1357 21901 1390
rect 20579 1328 20644 1331
rect 20579 1325 20648 1328
rect 20579 1265 20585 1325
rect 20644 1265 20654 1325
rect 20579 1261 20648 1265
rect 20579 1259 20644 1261
rect 20214 1162 20306 1170
rect 20214 1097 20226 1162
rect 20294 1097 20306 1162
rect 20214 1085 20306 1097
rect 21720 982 21905 1357
rect 22041 1339 22115 2452
rect 23540 2328 23550 2388
rect 23630 2328 23640 2388
rect 23540 2288 23640 2328
rect 22743 2231 24546 2288
rect 22743 2144 22777 2231
rect 23918 2144 23952 2231
rect 22737 2132 22783 2144
rect 22737 1944 22743 2132
rect 22296 1932 22342 1944
rect 22296 1756 22302 1932
rect 22336 1756 22342 1932
rect 22296 1744 22342 1756
rect 22414 1932 22460 1944
rect 22414 1756 22420 1932
rect 22454 1756 22460 1932
rect 22414 1744 22460 1756
rect 22532 1932 22578 1944
rect 22532 1756 22538 1932
rect 22572 1756 22578 1932
rect 22532 1744 22578 1756
rect 22650 1932 22743 1944
rect 22650 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22783 2132
rect 22650 1744 22783 1756
rect 22855 2132 22901 2144
rect 22855 1756 22861 2132
rect 22895 1756 22901 2132
rect 22855 1744 22901 1756
rect 22973 2132 23019 2144
rect 22973 1756 22979 2132
rect 23013 1756 23019 2132
rect 22973 1744 23019 1756
rect 23091 2132 23137 2144
rect 23091 1756 23097 2132
rect 23131 1756 23137 2132
rect 23091 1744 23137 1756
rect 23204 2132 23250 2144
rect 23204 1756 23210 2132
rect 23244 1756 23250 2132
rect 23204 1744 23250 1756
rect 23322 2132 23368 2144
rect 23322 1756 23328 2132
rect 23362 1756 23368 2132
rect 23322 1744 23368 1756
rect 23440 2132 23486 2144
rect 23440 1756 23446 2132
rect 23480 1756 23486 2132
rect 23440 1744 23486 1756
rect 23558 2132 23604 2144
rect 23558 1756 23564 2132
rect 23598 1756 23604 2132
rect 23558 1744 23604 1756
rect 23676 2132 23722 2144
rect 23676 1756 23682 2132
rect 23716 1756 23722 2132
rect 23676 1744 23722 1756
rect 23794 2132 23840 2144
rect 23794 1756 23800 2132
rect 23834 1756 23840 2132
rect 23794 1744 23840 1756
rect 23912 2132 23958 2144
rect 23912 1756 23918 2132
rect 23952 1756 23958 2132
rect 23912 1744 23958 1756
rect 24031 2132 24077 2144
rect 24031 1756 24037 2132
rect 24071 1756 24077 2132
rect 24031 1744 24077 1756
rect 24149 2132 24195 2144
rect 24149 1756 24155 2132
rect 24189 1756 24195 2132
rect 24149 1744 24195 1756
rect 24267 2132 24313 2144
rect 24267 1756 24273 2132
rect 24307 1756 24313 2132
rect 24267 1744 24313 1756
rect 24385 2132 24431 2144
rect 24385 1756 24391 2132
rect 24425 1756 24431 2132
rect 24509 1944 24546 2231
rect 28136 2079 28254 2493
rect 28308 2202 28426 2569
rect 28464 2382 28582 2672
rect 28648 2445 28766 2766
rect 28825 2473 28943 2800
rect 28987 2797 29103 2993
rect 29150 2819 29266 3065
rect 24385 1744 24431 1756
rect 24504 1932 24550 1944
rect 24504 1756 24510 1932
rect 24544 1756 24550 1932
rect 24504 1744 24550 1756
rect 24622 1932 24668 1944
rect 24622 1756 24628 1932
rect 24662 1756 24668 1932
rect 24622 1744 24668 1756
rect 24740 1932 24786 1944
rect 24740 1756 24746 1932
rect 24780 1756 24786 1932
rect 24740 1744 24786 1756
rect 24858 1932 24904 1944
rect 24858 1756 24864 1932
rect 24898 1756 24904 1932
rect 24858 1744 24904 1756
rect 22301 1558 22336 1744
rect 23210 1660 23244 1744
rect 24391 1660 24425 1744
rect 23210 1618 24425 1660
rect 24391 1598 24425 1618
rect 24391 1582 24748 1598
rect 22301 1541 23438 1558
rect 22301 1507 23388 1541
rect 23422 1507 23438 1541
rect 24391 1548 24698 1582
rect 24732 1548 24748 1582
rect 24391 1532 24748 1548
rect 22301 1491 23438 1507
rect 22143 1446 22218 1454
rect 22143 1378 22159 1446
rect 22216 1378 22226 1446
rect 22143 1370 22218 1378
rect 22041 1338 22126 1339
rect 22041 1330 22218 1338
rect 22041 1311 22159 1330
rect 22042 1262 22159 1311
rect 22216 1262 22226 1330
rect 22042 1254 22218 1262
rect 19157 934 20529 981
rect 20851 935 21905 982
rect 16859 807 16893 930
rect 17331 917 17397 930
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17720 807 17754 931
rect 18594 930 18771 931
rect 16854 795 16900 807
rect 16854 619 16860 795
rect 16894 619 16900 795
rect 16854 607 16900 619
rect 16972 795 17092 807
rect 16972 619 16978 795
rect 17012 619 17052 795
rect 16972 607 17052 619
rect 16978 240 17012 607
rect 17046 419 17052 607
rect 17086 419 17092 795
rect 17046 407 17092 419
rect 17164 795 17210 807
rect 17164 419 17170 795
rect 17204 419 17210 795
rect 17164 407 17210 419
rect 17282 795 17328 807
rect 17282 419 17288 795
rect 17322 419 17328 795
rect 17282 407 17328 419
rect 17400 795 17446 807
rect 17400 419 17406 795
rect 17440 419 17446 795
rect 17400 407 17446 419
rect 17518 795 17642 807
rect 17518 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17642 795
rect 17558 607 17642 619
rect 17714 795 17760 807
rect 17714 619 17720 795
rect 17754 619 17760 795
rect 17714 607 17760 619
rect 17558 419 17564 607
rect 17518 407 17564 419
rect 17288 334 17322 407
rect 17273 318 17339 334
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 17273 268 17339 284
rect 17602 240 17636 607
rect 16978 188 17636 240
rect 17276 166 17368 188
rect 17276 114 17288 166
rect 17354 114 17368 166
rect 17276 110 17368 114
rect 12585 -1189 15620 -1060
rect 10950 -1564 10960 -1504
rect 11040 -1564 11050 -1504
rect 10950 -1604 11050 -1564
rect 10153 -1661 11956 -1604
rect 10153 -1748 10187 -1661
rect 11328 -1748 11362 -1661
rect 10147 -1760 10193 -1748
rect 10147 -1948 10153 -1760
rect 9706 -1960 9752 -1948
rect 9706 -2136 9712 -1960
rect 9746 -2136 9752 -1960
rect 9706 -2148 9752 -2136
rect 9824 -1960 9870 -1948
rect 9824 -2136 9830 -1960
rect 9864 -2136 9870 -1960
rect 9824 -2148 9870 -2136
rect 9942 -1960 9988 -1948
rect 9942 -2136 9948 -1960
rect 9982 -2136 9988 -1960
rect 9942 -2148 9988 -2136
rect 10060 -1960 10153 -1948
rect 10060 -2136 10066 -1960
rect 10100 -2136 10153 -1960
rect 10187 -2136 10193 -1760
rect 10060 -2148 10193 -2136
rect 10265 -1760 10311 -1748
rect 10265 -2136 10271 -1760
rect 10305 -2136 10311 -1760
rect 10265 -2148 10311 -2136
rect 10383 -1760 10429 -1748
rect 10383 -2136 10389 -1760
rect 10423 -2136 10429 -1760
rect 10383 -2148 10429 -2136
rect 10501 -1760 10547 -1748
rect 10501 -2136 10507 -1760
rect 10541 -2136 10547 -1760
rect 10501 -2148 10547 -2136
rect 10614 -1760 10660 -1748
rect 10614 -2136 10620 -1760
rect 10654 -2136 10660 -1760
rect 10614 -2148 10660 -2136
rect 10732 -1760 10778 -1748
rect 10732 -2136 10738 -1760
rect 10772 -2136 10778 -1760
rect 10732 -2148 10778 -2136
rect 10850 -1760 10896 -1748
rect 10850 -2136 10856 -1760
rect 10890 -2136 10896 -1760
rect 10850 -2148 10896 -2136
rect 10968 -1760 11014 -1748
rect 10968 -2136 10974 -1760
rect 11008 -2136 11014 -1760
rect 10968 -2148 11014 -2136
rect 11086 -1760 11132 -1748
rect 11086 -2136 11092 -1760
rect 11126 -2136 11132 -1760
rect 11086 -2148 11132 -2136
rect 11204 -1760 11250 -1748
rect 11204 -2136 11210 -1760
rect 11244 -2136 11250 -1760
rect 11204 -2148 11250 -2136
rect 11322 -1760 11368 -1748
rect 11322 -2136 11328 -1760
rect 11362 -2136 11368 -1760
rect 11322 -2148 11368 -2136
rect 11441 -1760 11487 -1748
rect 11441 -2136 11447 -1760
rect 11481 -2136 11487 -1760
rect 11441 -2148 11487 -2136
rect 11559 -1760 11605 -1748
rect 11559 -2136 11565 -1760
rect 11599 -2136 11605 -1760
rect 11559 -2148 11605 -2136
rect 11677 -1760 11723 -1748
rect 11677 -2136 11683 -1760
rect 11717 -2136 11723 -1760
rect 11677 -2148 11723 -2136
rect 11795 -1760 11841 -1748
rect 11795 -2136 11801 -1760
rect 11835 -2136 11841 -1760
rect 11919 -1948 11956 -1661
rect 11795 -2148 11841 -2136
rect 11914 -1960 11960 -1948
rect 11914 -2136 11920 -1960
rect 11954 -2136 11960 -1960
rect 11914 -2148 11960 -2136
rect 12032 -1960 12078 -1948
rect 12032 -2136 12038 -1960
rect 12072 -2136 12078 -1960
rect 12032 -2148 12078 -2136
rect 12150 -1960 12196 -1948
rect 12150 -2136 12156 -1960
rect 12190 -2136 12196 -1960
rect 12150 -2148 12196 -2136
rect 12268 -1960 12314 -1948
rect 12268 -2136 12274 -1960
rect 12308 -2136 12314 -1960
rect 12268 -2148 12314 -2136
rect 9711 -2334 9746 -2148
rect 10620 -2232 10654 -2148
rect 11801 -2232 11835 -2148
rect 10620 -2274 11835 -2232
rect 11801 -2294 11835 -2274
rect 11801 -2310 12158 -2294
rect 9711 -2351 10848 -2334
rect 9711 -2385 10798 -2351
rect 10832 -2385 10848 -2351
rect 11801 -2344 12108 -2310
rect 12142 -2344 12158 -2310
rect 11801 -2360 12158 -2344
rect 9711 -2401 10848 -2385
rect 9553 -2446 9628 -2438
rect 9553 -2514 9569 -2446
rect 9626 -2514 9636 -2446
rect 9553 -2522 9628 -2514
rect 9374 -2562 9628 -2554
rect 7989 -2631 8058 -2627
rect 7989 -2633 8054 -2631
rect 7624 -2730 7716 -2722
rect 7624 -2795 7636 -2730
rect 7704 -2795 7716 -2730
rect 7624 -2807 7716 -2795
rect 9130 -2910 9317 -2591
rect 9374 -2630 9569 -2562
rect 9626 -2630 9636 -2562
rect 9374 -2638 9628 -2630
rect 6567 -2958 7939 -2911
rect 8261 -2957 9317 -2910
rect 4269 -3085 4303 -2962
rect 4741 -2975 4807 -2962
rect 4741 -3009 4757 -2975
rect 4791 -3009 4807 -2975
rect 4741 -3025 4807 -3009
rect 5130 -3085 5164 -2961
rect 4264 -3097 4310 -3085
rect 4264 -3273 4270 -3097
rect 4304 -3273 4310 -3097
rect 4264 -3285 4310 -3273
rect 4382 -3097 4502 -3085
rect 4382 -3273 4388 -3097
rect 4422 -3273 4462 -3097
rect 4382 -3285 4462 -3273
rect 4388 -3652 4422 -3285
rect 4456 -3473 4462 -3285
rect 4496 -3473 4502 -3097
rect 4456 -3485 4502 -3473
rect 4574 -3097 4620 -3085
rect 4574 -3473 4580 -3097
rect 4614 -3473 4620 -3097
rect 4574 -3485 4620 -3473
rect 4692 -3097 4738 -3085
rect 4692 -3473 4698 -3097
rect 4732 -3473 4738 -3097
rect 4692 -3485 4738 -3473
rect 4810 -3097 4856 -3085
rect 4810 -3473 4816 -3097
rect 4850 -3473 4856 -3097
rect 4810 -3485 4856 -3473
rect 4928 -3097 5052 -3085
rect 4928 -3473 4934 -3097
rect 4968 -3273 5012 -3097
rect 5046 -3273 5052 -3097
rect 4968 -3285 5052 -3273
rect 5124 -3097 5170 -3085
rect 5124 -3273 5130 -3097
rect 5164 -3273 5170 -3097
rect 5124 -3285 5170 -3273
rect 4968 -3473 4974 -3285
rect 4928 -3485 4974 -3473
rect 4698 -3558 4732 -3485
rect 4683 -3574 4749 -3558
rect 4683 -3608 4699 -3574
rect 4733 -3608 4749 -3574
rect 4683 -3624 4749 -3608
rect 5012 -3652 5046 -3285
rect 4388 -3704 5046 -3652
rect 4686 -3726 4778 -3704
rect 4686 -3778 4698 -3726
rect 4764 -3778 4778 -3726
rect 4686 -3782 4778 -3778
rect 6031 -4499 6182 -2961
rect 7401 -3081 7435 -2958
rect 7873 -2971 7939 -2958
rect 7873 -3005 7889 -2971
rect 7923 -3005 7939 -2971
rect 7873 -3021 7939 -3005
rect 8262 -3081 8296 -2957
rect 9133 -2960 9317 -2957
rect 9711 -2911 9746 -2401
rect 9801 -2447 9893 -2434
rect 9801 -2510 9813 -2447
rect 9884 -2510 9893 -2447
rect 9801 -2519 9893 -2510
rect 10886 -2447 10978 -2437
rect 10886 -2509 10898 -2447
rect 10968 -2509 10978 -2447
rect 10886 -2522 10978 -2509
rect 12274 -2502 12309 -2148
rect 11133 -2564 11198 -2561
rect 11133 -2567 11202 -2564
rect 11133 -2627 11139 -2567
rect 11198 -2627 11208 -2567
rect 12274 -2581 12455 -2502
rect 12585 -2558 12689 -1189
rect 15474 -1193 15620 -1189
rect 15744 -1060 15837 -1059
rect 18625 -1060 18771 930
rect 19991 811 20025 934
rect 20463 921 20529 934
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20852 811 20886 935
rect 21726 933 21905 935
rect 22301 981 22336 1491
rect 22391 1445 22483 1458
rect 22391 1382 22403 1445
rect 22474 1382 22483 1445
rect 22391 1373 22483 1382
rect 23476 1445 23568 1455
rect 23476 1383 23488 1445
rect 23558 1383 23568 1445
rect 23476 1370 23568 1383
rect 24864 1390 24899 1744
rect 23723 1328 23788 1331
rect 23723 1325 23792 1328
rect 23723 1265 23729 1325
rect 23788 1265 23798 1325
rect 23723 1261 23792 1265
rect 23723 1259 23788 1261
rect 23358 1162 23450 1170
rect 23358 1097 23370 1162
rect 23438 1097 23450 1162
rect 23358 1085 23450 1097
rect 24864 982 25045 1390
rect 22301 934 23673 981
rect 23995 935 25045 982
rect 19986 799 20032 811
rect 19986 623 19992 799
rect 20026 623 20032 799
rect 19986 611 20032 623
rect 20104 799 20224 811
rect 20104 623 20110 799
rect 20144 623 20184 799
rect 20104 611 20184 623
rect 20110 244 20144 611
rect 20178 423 20184 611
rect 20218 423 20224 799
rect 20178 411 20224 423
rect 20296 799 20342 811
rect 20296 423 20302 799
rect 20336 423 20342 799
rect 20296 411 20342 423
rect 20414 799 20460 811
rect 20414 423 20420 799
rect 20454 423 20460 799
rect 20414 411 20460 423
rect 20532 799 20578 811
rect 20532 423 20538 799
rect 20572 423 20578 799
rect 20532 411 20578 423
rect 20650 799 20774 811
rect 20650 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20774 799
rect 20690 611 20774 623
rect 20846 799 20892 811
rect 20846 623 20852 799
rect 20886 623 20892 799
rect 20846 611 20892 623
rect 20690 423 20696 611
rect 20650 411 20696 423
rect 20420 338 20454 411
rect 20405 322 20471 338
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 20405 272 20471 288
rect 20734 244 20768 611
rect 20110 192 20768 244
rect 20408 170 20500 192
rect 20408 118 20420 170
rect 20486 118 20500 170
rect 20408 114 20500 118
rect 21759 -1060 21905 933
rect 23135 811 23169 934
rect 23607 921 23673 934
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23996 811 24030 935
rect 23130 799 23176 811
rect 23130 623 23136 799
rect 23170 623 23176 799
rect 23130 611 23176 623
rect 23248 799 23368 811
rect 23248 623 23254 799
rect 23288 623 23328 799
rect 23248 611 23328 623
rect 23254 244 23288 611
rect 23322 423 23328 611
rect 23362 423 23368 799
rect 23322 411 23368 423
rect 23440 799 23486 811
rect 23440 423 23446 799
rect 23480 423 23486 799
rect 23440 411 23486 423
rect 23558 799 23604 811
rect 23558 423 23564 799
rect 23598 423 23604 799
rect 23558 411 23604 423
rect 23676 799 23722 811
rect 23676 423 23682 799
rect 23716 423 23722 799
rect 23676 411 23722 423
rect 23794 799 23918 811
rect 23794 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23918 799
rect 23834 611 23918 623
rect 23990 799 24036 811
rect 23990 623 23996 799
rect 24030 623 24036 799
rect 23990 611 24036 623
rect 23834 423 23840 611
rect 23794 411 23840 423
rect 23564 338 23598 411
rect 23549 322 23615 338
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 23549 272 23615 288
rect 23878 244 23912 611
rect 23254 192 23912 244
rect 23552 170 23644 192
rect 23552 118 23564 170
rect 23630 118 23644 170
rect 23552 114 23644 118
rect 15744 -1189 18771 -1060
rect 18885 -1165 21905 -1060
rect 24899 -1063 25045 935
rect 15744 -1199 15849 -1189
rect 18625 -1193 18771 -1189
rect 18884 -1188 21905 -1165
rect 18884 -1189 21898 -1188
rect 14152 -1568 14162 -1508
rect 14242 -1568 14252 -1508
rect 14152 -1608 14252 -1568
rect 13355 -1665 15158 -1608
rect 13355 -1752 13389 -1665
rect 14530 -1752 14564 -1665
rect 13349 -1764 13395 -1752
rect 13349 -1952 13355 -1764
rect 12908 -1964 12954 -1952
rect 12908 -2140 12914 -1964
rect 12948 -2140 12954 -1964
rect 12908 -2152 12954 -2140
rect 13026 -1964 13072 -1952
rect 13026 -2140 13032 -1964
rect 13066 -2140 13072 -1964
rect 13026 -2152 13072 -2140
rect 13144 -1964 13190 -1952
rect 13144 -2140 13150 -1964
rect 13184 -2140 13190 -1964
rect 13144 -2152 13190 -2140
rect 13262 -1964 13355 -1952
rect 13262 -2140 13268 -1964
rect 13302 -2140 13355 -1964
rect 13389 -2140 13395 -1764
rect 13262 -2152 13395 -2140
rect 13467 -1764 13513 -1752
rect 13467 -2140 13473 -1764
rect 13507 -2140 13513 -1764
rect 13467 -2152 13513 -2140
rect 13585 -1764 13631 -1752
rect 13585 -2140 13591 -1764
rect 13625 -2140 13631 -1764
rect 13585 -2152 13631 -2140
rect 13703 -1764 13749 -1752
rect 13703 -2140 13709 -1764
rect 13743 -2140 13749 -1764
rect 13703 -2152 13749 -2140
rect 13816 -1764 13862 -1752
rect 13816 -2140 13822 -1764
rect 13856 -2140 13862 -1764
rect 13816 -2152 13862 -2140
rect 13934 -1764 13980 -1752
rect 13934 -2140 13940 -1764
rect 13974 -2140 13980 -1764
rect 13934 -2152 13980 -2140
rect 14052 -1764 14098 -1752
rect 14052 -2140 14058 -1764
rect 14092 -2140 14098 -1764
rect 14052 -2152 14098 -2140
rect 14170 -1764 14216 -1752
rect 14170 -2140 14176 -1764
rect 14210 -2140 14216 -1764
rect 14170 -2152 14216 -2140
rect 14288 -1764 14334 -1752
rect 14288 -2140 14294 -1764
rect 14328 -2140 14334 -1764
rect 14288 -2152 14334 -2140
rect 14406 -1764 14452 -1752
rect 14406 -2140 14412 -1764
rect 14446 -2140 14452 -1764
rect 14406 -2152 14452 -2140
rect 14524 -1764 14570 -1752
rect 14524 -2140 14530 -1764
rect 14564 -2140 14570 -1764
rect 14524 -2152 14570 -2140
rect 14643 -1764 14689 -1752
rect 14643 -2140 14649 -1764
rect 14683 -2140 14689 -1764
rect 14643 -2152 14689 -2140
rect 14761 -1764 14807 -1752
rect 14761 -2140 14767 -1764
rect 14801 -2140 14807 -1764
rect 14761 -2152 14807 -2140
rect 14879 -1764 14925 -1752
rect 14879 -2140 14885 -1764
rect 14919 -2140 14925 -1764
rect 14879 -2152 14925 -2140
rect 14997 -1764 15043 -1752
rect 14997 -2140 15003 -1764
rect 15037 -2140 15043 -1764
rect 15121 -1952 15158 -1665
rect 14997 -2152 15043 -2140
rect 15116 -1964 15162 -1952
rect 15116 -2140 15122 -1964
rect 15156 -2140 15162 -1964
rect 15116 -2152 15162 -2140
rect 15234 -1964 15280 -1952
rect 15234 -2140 15240 -1964
rect 15274 -2140 15280 -1964
rect 15234 -2152 15280 -2140
rect 15352 -1964 15398 -1952
rect 15352 -2140 15358 -1964
rect 15392 -2140 15398 -1964
rect 15352 -2152 15398 -2140
rect 15470 -1964 15516 -1952
rect 15470 -2140 15476 -1964
rect 15510 -2140 15516 -1964
rect 15470 -2152 15516 -2140
rect 12913 -2338 12948 -2152
rect 13822 -2236 13856 -2152
rect 15003 -2236 15037 -2152
rect 13822 -2278 15037 -2236
rect 15003 -2298 15037 -2278
rect 15003 -2314 15360 -2298
rect 12913 -2355 14050 -2338
rect 12913 -2389 14000 -2355
rect 14034 -2389 14050 -2355
rect 15003 -2348 15310 -2314
rect 15344 -2348 15360 -2314
rect 15003 -2364 15360 -2348
rect 12913 -2405 14050 -2389
rect 12752 -2450 12830 -2442
rect 12752 -2518 12771 -2450
rect 12828 -2518 12838 -2450
rect 12752 -2526 12830 -2518
rect 12585 -2566 12830 -2558
rect 11133 -2631 11202 -2627
rect 11133 -2633 11198 -2631
rect 10768 -2730 10860 -2722
rect 10768 -2795 10780 -2730
rect 10848 -2795 10860 -2730
rect 10768 -2807 10860 -2795
rect 12274 -2910 12459 -2581
rect 12585 -2634 12771 -2566
rect 12828 -2634 12838 -2566
rect 12585 -2642 12830 -2634
rect 12585 -2643 12689 -2642
rect 9711 -2958 11083 -2911
rect 11405 -2957 12459 -2910
rect 7396 -3093 7442 -3081
rect 7396 -3269 7402 -3093
rect 7436 -3269 7442 -3093
rect 7396 -3281 7442 -3269
rect 7514 -3093 7634 -3081
rect 7514 -3269 7520 -3093
rect 7554 -3269 7594 -3093
rect 7514 -3281 7594 -3269
rect 7520 -3648 7554 -3281
rect 7588 -3469 7594 -3281
rect 7628 -3469 7634 -3093
rect 7588 -3481 7634 -3469
rect 7706 -3093 7752 -3081
rect 7706 -3469 7712 -3093
rect 7746 -3469 7752 -3093
rect 7706 -3481 7752 -3469
rect 7824 -3093 7870 -3081
rect 7824 -3469 7830 -3093
rect 7864 -3469 7870 -3093
rect 7824 -3481 7870 -3469
rect 7942 -3093 7988 -3081
rect 7942 -3469 7948 -3093
rect 7982 -3469 7988 -3093
rect 7942 -3481 7988 -3469
rect 8060 -3093 8184 -3081
rect 8060 -3469 8066 -3093
rect 8100 -3269 8144 -3093
rect 8178 -3269 8184 -3093
rect 8100 -3281 8184 -3269
rect 8256 -3093 8302 -3081
rect 8256 -3269 8262 -3093
rect 8296 -3269 8302 -3093
rect 8256 -3281 8302 -3269
rect 8100 -3469 8106 -3281
rect 8060 -3481 8106 -3469
rect 7830 -3554 7864 -3481
rect 7815 -3570 7881 -3554
rect 7815 -3604 7831 -3570
rect 7865 -3604 7881 -3570
rect 7815 -3620 7881 -3604
rect 8144 -3648 8178 -3281
rect 7520 -3700 8178 -3648
rect 7818 -3722 7910 -3700
rect 7818 -3774 7830 -3722
rect 7896 -3774 7910 -3722
rect 7818 -3778 7910 -3774
rect 9166 -4494 9317 -2960
rect 10545 -3081 10579 -2958
rect 11017 -2971 11083 -2958
rect 11017 -3005 11033 -2971
rect 11067 -3005 11083 -2971
rect 11017 -3021 11083 -3005
rect 11406 -3081 11440 -2957
rect 10540 -3093 10586 -3081
rect 10540 -3269 10546 -3093
rect 10580 -3269 10586 -3093
rect 10540 -3281 10586 -3269
rect 10658 -3093 10778 -3081
rect 10658 -3269 10664 -3093
rect 10698 -3269 10738 -3093
rect 10658 -3281 10738 -3269
rect 10664 -3648 10698 -3281
rect 10732 -3469 10738 -3281
rect 10772 -3469 10778 -3093
rect 10732 -3481 10778 -3469
rect 10850 -3093 10896 -3081
rect 10850 -3469 10856 -3093
rect 10890 -3469 10896 -3093
rect 10850 -3481 10896 -3469
rect 10968 -3093 11014 -3081
rect 10968 -3469 10974 -3093
rect 11008 -3469 11014 -3093
rect 10968 -3481 11014 -3469
rect 11086 -3093 11132 -3081
rect 11086 -3469 11092 -3093
rect 11126 -3469 11132 -3093
rect 11086 -3481 11132 -3469
rect 11204 -3093 11328 -3081
rect 11204 -3469 11210 -3093
rect 11244 -3269 11288 -3093
rect 11322 -3269 11328 -3093
rect 11244 -3281 11328 -3269
rect 11400 -3093 11446 -3081
rect 11400 -3269 11406 -3093
rect 11440 -3269 11446 -3093
rect 11400 -3281 11446 -3269
rect 11244 -3469 11250 -3281
rect 11204 -3481 11250 -3469
rect 10974 -3554 11008 -3481
rect 10959 -3570 11025 -3554
rect 10959 -3604 10975 -3570
rect 11009 -3604 11025 -3570
rect 10959 -3620 11025 -3604
rect 11288 -3648 11322 -3281
rect 10664 -3700 11322 -3648
rect 10962 -3722 11054 -3700
rect 10962 -3774 10974 -3722
rect 11040 -3774 11054 -3722
rect 10962 -3778 11054 -3774
rect 12308 -4484 12459 -2957
rect 12913 -2915 12948 -2405
rect 13003 -2451 13095 -2438
rect 13003 -2514 13015 -2451
rect 13086 -2514 13095 -2451
rect 13003 -2523 13095 -2514
rect 14088 -2451 14180 -2441
rect 14088 -2513 14100 -2451
rect 14170 -2513 14180 -2451
rect 14088 -2526 14180 -2513
rect 15476 -2506 15511 -2152
rect 14335 -2568 14400 -2565
rect 14335 -2571 14404 -2568
rect 14335 -2631 14341 -2571
rect 14400 -2631 14410 -2571
rect 15476 -2589 15657 -2506
rect 15745 -2558 15849 -1199
rect 17296 -1568 17306 -1508
rect 17386 -1568 17396 -1508
rect 17296 -1608 17396 -1568
rect 16499 -1665 18302 -1608
rect 16499 -1752 16533 -1665
rect 17674 -1752 17708 -1665
rect 16493 -1764 16539 -1752
rect 16493 -1952 16499 -1764
rect 16052 -1964 16098 -1952
rect 16052 -2140 16058 -1964
rect 16092 -2140 16098 -1964
rect 16052 -2152 16098 -2140
rect 16170 -1964 16216 -1952
rect 16170 -2140 16176 -1964
rect 16210 -2140 16216 -1964
rect 16170 -2152 16216 -2140
rect 16288 -1964 16334 -1952
rect 16288 -2140 16294 -1964
rect 16328 -2140 16334 -1964
rect 16288 -2152 16334 -2140
rect 16406 -1964 16499 -1952
rect 16406 -2140 16412 -1964
rect 16446 -2140 16499 -1964
rect 16533 -2140 16539 -1764
rect 16406 -2152 16539 -2140
rect 16611 -1764 16657 -1752
rect 16611 -2140 16617 -1764
rect 16651 -2140 16657 -1764
rect 16611 -2152 16657 -2140
rect 16729 -1764 16775 -1752
rect 16729 -2140 16735 -1764
rect 16769 -2140 16775 -1764
rect 16729 -2152 16775 -2140
rect 16847 -1764 16893 -1752
rect 16847 -2140 16853 -1764
rect 16887 -2140 16893 -1764
rect 16847 -2152 16893 -2140
rect 16960 -1764 17006 -1752
rect 16960 -2140 16966 -1764
rect 17000 -2140 17006 -1764
rect 16960 -2152 17006 -2140
rect 17078 -1764 17124 -1752
rect 17078 -2140 17084 -1764
rect 17118 -2140 17124 -1764
rect 17078 -2152 17124 -2140
rect 17196 -1764 17242 -1752
rect 17196 -2140 17202 -1764
rect 17236 -2140 17242 -1764
rect 17196 -2152 17242 -2140
rect 17314 -1764 17360 -1752
rect 17314 -2140 17320 -1764
rect 17354 -2140 17360 -1764
rect 17314 -2152 17360 -2140
rect 17432 -1764 17478 -1752
rect 17432 -2140 17438 -1764
rect 17472 -2140 17478 -1764
rect 17432 -2152 17478 -2140
rect 17550 -1764 17596 -1752
rect 17550 -2140 17556 -1764
rect 17590 -2140 17596 -1764
rect 17550 -2152 17596 -2140
rect 17668 -1764 17714 -1752
rect 17668 -2140 17674 -1764
rect 17708 -2140 17714 -1764
rect 17668 -2152 17714 -2140
rect 17787 -1764 17833 -1752
rect 17787 -2140 17793 -1764
rect 17827 -2140 17833 -1764
rect 17787 -2152 17833 -2140
rect 17905 -1764 17951 -1752
rect 17905 -2140 17911 -1764
rect 17945 -2140 17951 -1764
rect 17905 -2152 17951 -2140
rect 18023 -1764 18069 -1752
rect 18023 -2140 18029 -1764
rect 18063 -2140 18069 -1764
rect 18023 -2152 18069 -2140
rect 18141 -1764 18187 -1752
rect 18141 -2140 18147 -1764
rect 18181 -2140 18187 -1764
rect 18265 -1952 18302 -1665
rect 18141 -2152 18187 -2140
rect 18260 -1964 18306 -1952
rect 18260 -2140 18266 -1964
rect 18300 -2140 18306 -1964
rect 18260 -2152 18306 -2140
rect 18378 -1964 18424 -1952
rect 18378 -2140 18384 -1964
rect 18418 -2140 18424 -1964
rect 18378 -2152 18424 -2140
rect 18496 -1964 18542 -1952
rect 18496 -2140 18502 -1964
rect 18536 -2140 18542 -1964
rect 18496 -2152 18542 -2140
rect 18614 -1964 18660 -1952
rect 18614 -2140 18620 -1964
rect 18654 -2140 18660 -1964
rect 18614 -2152 18660 -2140
rect 16057 -2338 16092 -2152
rect 16966 -2236 17000 -2152
rect 18147 -2236 18181 -2152
rect 16966 -2278 18181 -2236
rect 18147 -2298 18181 -2278
rect 18147 -2314 18504 -2298
rect 16057 -2355 17194 -2338
rect 16057 -2389 17144 -2355
rect 17178 -2389 17194 -2355
rect 18147 -2348 18454 -2314
rect 18488 -2348 18504 -2314
rect 18147 -2364 18504 -2348
rect 16057 -2405 17194 -2389
rect 15899 -2450 15974 -2442
rect 15899 -2518 15915 -2450
rect 15972 -2518 15982 -2450
rect 15899 -2526 15974 -2518
rect 15745 -2566 15974 -2558
rect 14335 -2635 14404 -2631
rect 14335 -2637 14400 -2635
rect 13970 -2734 14062 -2726
rect 13970 -2799 13982 -2734
rect 14050 -2799 14062 -2734
rect 13970 -2811 14062 -2799
rect 15476 -2914 15660 -2589
rect 15745 -2634 15915 -2566
rect 15972 -2634 15982 -2566
rect 15745 -2641 15974 -2634
rect 15798 -2642 15974 -2641
rect 12913 -2962 14285 -2915
rect 14607 -2961 15660 -2914
rect 13747 -3085 13781 -2962
rect 14219 -2975 14285 -2962
rect 14219 -3009 14235 -2975
rect 14269 -3009 14285 -2975
rect 14219 -3025 14285 -3009
rect 14608 -3085 14642 -2961
rect 13742 -3097 13788 -3085
rect 13742 -3273 13748 -3097
rect 13782 -3273 13788 -3097
rect 13742 -3285 13788 -3273
rect 13860 -3097 13980 -3085
rect 13860 -3273 13866 -3097
rect 13900 -3273 13940 -3097
rect 13860 -3285 13940 -3273
rect 13866 -3652 13900 -3285
rect 13934 -3473 13940 -3285
rect 13974 -3473 13980 -3097
rect 13934 -3485 13980 -3473
rect 14052 -3097 14098 -3085
rect 14052 -3473 14058 -3097
rect 14092 -3473 14098 -3097
rect 14052 -3485 14098 -3473
rect 14170 -3097 14216 -3085
rect 14170 -3473 14176 -3097
rect 14210 -3473 14216 -3097
rect 14170 -3485 14216 -3473
rect 14288 -3097 14334 -3085
rect 14288 -3473 14294 -3097
rect 14328 -3473 14334 -3097
rect 14288 -3485 14334 -3473
rect 14406 -3097 14530 -3085
rect 14406 -3473 14412 -3097
rect 14446 -3273 14490 -3097
rect 14524 -3273 14530 -3097
rect 14446 -3285 14530 -3273
rect 14602 -3097 14648 -3085
rect 14602 -3273 14608 -3097
rect 14642 -3273 14648 -3097
rect 14602 -3285 14648 -3273
rect 14446 -3473 14452 -3285
rect 14406 -3485 14452 -3473
rect 14176 -3558 14210 -3485
rect 14161 -3574 14227 -3558
rect 14161 -3608 14177 -3574
rect 14211 -3608 14227 -3574
rect 14161 -3624 14227 -3608
rect 14490 -3652 14524 -3285
rect 13866 -3704 14524 -3652
rect 14164 -3726 14256 -3704
rect 14164 -3778 14176 -3726
rect 14242 -3778 14256 -3726
rect 14164 -3782 14256 -3778
rect 15509 -4492 15660 -2961
rect 16057 -2915 16092 -2405
rect 16147 -2451 16239 -2438
rect 16147 -2514 16159 -2451
rect 16230 -2514 16239 -2451
rect 16147 -2523 16239 -2514
rect 17232 -2451 17324 -2441
rect 17232 -2513 17244 -2451
rect 17314 -2513 17324 -2451
rect 17232 -2526 17324 -2513
rect 18620 -2482 18655 -2152
rect 18620 -2484 18693 -2482
rect 17479 -2568 17544 -2565
rect 17479 -2571 17548 -2568
rect 17479 -2631 17485 -2571
rect 17544 -2631 17554 -2571
rect 17479 -2635 17548 -2631
rect 17479 -2637 17544 -2635
rect 17114 -2734 17206 -2726
rect 17114 -2799 17126 -2734
rect 17194 -2799 17206 -2734
rect 17114 -2811 17206 -2799
rect 18620 -2914 18807 -2484
rect 18884 -2554 18988 -1189
rect 22004 -1192 25045 -1063
rect 20428 -1564 20438 -1504
rect 20518 -1564 20528 -1504
rect 20428 -1604 20528 -1564
rect 19631 -1661 21434 -1604
rect 19631 -1748 19665 -1661
rect 20806 -1748 20840 -1661
rect 19625 -1760 19671 -1748
rect 19625 -1948 19631 -1760
rect 19184 -1960 19230 -1948
rect 19184 -2136 19190 -1960
rect 19224 -2136 19230 -1960
rect 19184 -2148 19230 -2136
rect 19302 -1960 19348 -1948
rect 19302 -2136 19308 -1960
rect 19342 -2136 19348 -1960
rect 19302 -2148 19348 -2136
rect 19420 -1960 19466 -1948
rect 19420 -2136 19426 -1960
rect 19460 -2136 19466 -1960
rect 19420 -2148 19466 -2136
rect 19538 -1960 19631 -1948
rect 19538 -2136 19544 -1960
rect 19578 -2136 19631 -1960
rect 19665 -2136 19671 -1760
rect 19538 -2148 19671 -2136
rect 19743 -1760 19789 -1748
rect 19743 -2136 19749 -1760
rect 19783 -2136 19789 -1760
rect 19743 -2148 19789 -2136
rect 19861 -1760 19907 -1748
rect 19861 -2136 19867 -1760
rect 19901 -2136 19907 -1760
rect 19861 -2148 19907 -2136
rect 19979 -1760 20025 -1748
rect 19979 -2136 19985 -1760
rect 20019 -2136 20025 -1760
rect 19979 -2148 20025 -2136
rect 20092 -1760 20138 -1748
rect 20092 -2136 20098 -1760
rect 20132 -2136 20138 -1760
rect 20092 -2148 20138 -2136
rect 20210 -1760 20256 -1748
rect 20210 -2136 20216 -1760
rect 20250 -2136 20256 -1760
rect 20210 -2148 20256 -2136
rect 20328 -1760 20374 -1748
rect 20328 -2136 20334 -1760
rect 20368 -2136 20374 -1760
rect 20328 -2148 20374 -2136
rect 20446 -1760 20492 -1748
rect 20446 -2136 20452 -1760
rect 20486 -2136 20492 -1760
rect 20446 -2148 20492 -2136
rect 20564 -1760 20610 -1748
rect 20564 -2136 20570 -1760
rect 20604 -2136 20610 -1760
rect 20564 -2148 20610 -2136
rect 20682 -1760 20728 -1748
rect 20682 -2136 20688 -1760
rect 20722 -2136 20728 -1760
rect 20682 -2148 20728 -2136
rect 20800 -1760 20846 -1748
rect 20800 -2136 20806 -1760
rect 20840 -2136 20846 -1760
rect 20800 -2148 20846 -2136
rect 20919 -1760 20965 -1748
rect 20919 -2136 20925 -1760
rect 20959 -2136 20965 -1760
rect 20919 -2148 20965 -2136
rect 21037 -1760 21083 -1748
rect 21037 -2136 21043 -1760
rect 21077 -2136 21083 -1760
rect 21037 -2148 21083 -2136
rect 21155 -1760 21201 -1748
rect 21155 -2136 21161 -1760
rect 21195 -2136 21201 -1760
rect 21155 -2148 21201 -2136
rect 21273 -1760 21319 -1748
rect 21273 -2136 21279 -1760
rect 21313 -2136 21319 -1760
rect 21397 -1948 21434 -1661
rect 21273 -2148 21319 -2136
rect 21392 -1960 21438 -1948
rect 21392 -2136 21398 -1960
rect 21432 -2136 21438 -1960
rect 21392 -2148 21438 -2136
rect 21510 -1960 21556 -1948
rect 21510 -2136 21516 -1960
rect 21550 -2136 21556 -1960
rect 21510 -2148 21556 -2136
rect 21628 -1960 21674 -1948
rect 21628 -2136 21634 -1960
rect 21668 -2136 21674 -1960
rect 21628 -2148 21674 -2136
rect 21746 -1960 21792 -1948
rect 21746 -2136 21752 -1960
rect 21786 -2136 21792 -1960
rect 21746 -2148 21792 -2136
rect 19189 -2334 19224 -2148
rect 20098 -2232 20132 -2148
rect 21279 -2232 21313 -2148
rect 20098 -2274 21313 -2232
rect 21279 -2294 21313 -2274
rect 21279 -2310 21636 -2294
rect 19189 -2351 20326 -2334
rect 19189 -2385 20276 -2351
rect 20310 -2385 20326 -2351
rect 21279 -2344 21586 -2310
rect 21620 -2344 21636 -2310
rect 21279 -2360 21636 -2344
rect 19189 -2401 20326 -2385
rect 19029 -2446 19106 -2438
rect 19029 -2514 19047 -2446
rect 19104 -2514 19114 -2446
rect 19029 -2522 19106 -2514
rect 18884 -2562 19106 -2554
rect 18884 -2630 19047 -2562
rect 19104 -2630 19114 -2562
rect 18884 -2638 19106 -2630
rect 18884 -2641 18988 -2638
rect 16057 -2962 17429 -2915
rect 17751 -2961 18807 -2914
rect 19189 -2911 19224 -2401
rect 19279 -2447 19371 -2434
rect 19279 -2510 19291 -2447
rect 19362 -2510 19371 -2447
rect 19279 -2519 19371 -2510
rect 20364 -2447 20456 -2437
rect 20364 -2509 20376 -2447
rect 20446 -2509 20456 -2447
rect 20364 -2522 20456 -2509
rect 21752 -2502 21787 -2148
rect 20611 -2564 20676 -2561
rect 20611 -2567 20680 -2564
rect 20611 -2627 20617 -2567
rect 20676 -2627 20686 -2567
rect 20611 -2631 20680 -2627
rect 20611 -2633 20676 -2631
rect 21752 -2648 21933 -2502
rect 22004 -2554 22108 -1192
rect 24899 -1193 25045 -1192
rect 23572 -1564 23582 -1504
rect 23662 -1564 23672 -1504
rect 23572 -1604 23672 -1564
rect 22775 -1661 24578 -1604
rect 22775 -1748 22809 -1661
rect 23950 -1748 23984 -1661
rect 22769 -1760 22815 -1748
rect 22769 -1948 22775 -1760
rect 22328 -1960 22374 -1948
rect 22328 -2136 22334 -1960
rect 22368 -2136 22374 -1960
rect 22328 -2148 22374 -2136
rect 22446 -1960 22492 -1948
rect 22446 -2136 22452 -1960
rect 22486 -2136 22492 -1960
rect 22446 -2148 22492 -2136
rect 22564 -1960 22610 -1948
rect 22564 -2136 22570 -1960
rect 22604 -2136 22610 -1960
rect 22564 -2148 22610 -2136
rect 22682 -1960 22775 -1948
rect 22682 -2136 22688 -1960
rect 22722 -2136 22775 -1960
rect 22809 -2136 22815 -1760
rect 22682 -2148 22815 -2136
rect 22887 -1760 22933 -1748
rect 22887 -2136 22893 -1760
rect 22927 -2136 22933 -1760
rect 22887 -2148 22933 -2136
rect 23005 -1760 23051 -1748
rect 23005 -2136 23011 -1760
rect 23045 -2136 23051 -1760
rect 23005 -2148 23051 -2136
rect 23123 -1760 23169 -1748
rect 23123 -2136 23129 -1760
rect 23163 -2136 23169 -1760
rect 23123 -2148 23169 -2136
rect 23236 -1760 23282 -1748
rect 23236 -2136 23242 -1760
rect 23276 -2136 23282 -1760
rect 23236 -2148 23282 -2136
rect 23354 -1760 23400 -1748
rect 23354 -2136 23360 -1760
rect 23394 -2136 23400 -1760
rect 23354 -2148 23400 -2136
rect 23472 -1760 23518 -1748
rect 23472 -2136 23478 -1760
rect 23512 -2136 23518 -1760
rect 23472 -2148 23518 -2136
rect 23590 -1760 23636 -1748
rect 23590 -2136 23596 -1760
rect 23630 -2136 23636 -1760
rect 23590 -2148 23636 -2136
rect 23708 -1760 23754 -1748
rect 23708 -2136 23714 -1760
rect 23748 -2136 23754 -1760
rect 23708 -2148 23754 -2136
rect 23826 -1760 23872 -1748
rect 23826 -2136 23832 -1760
rect 23866 -2136 23872 -1760
rect 23826 -2148 23872 -2136
rect 23944 -1760 23990 -1748
rect 23944 -2136 23950 -1760
rect 23984 -2136 23990 -1760
rect 23944 -2148 23990 -2136
rect 24063 -1760 24109 -1748
rect 24063 -2136 24069 -1760
rect 24103 -2136 24109 -1760
rect 24063 -2148 24109 -2136
rect 24181 -1760 24227 -1748
rect 24181 -2136 24187 -1760
rect 24221 -2136 24227 -1760
rect 24181 -2148 24227 -2136
rect 24299 -1760 24345 -1748
rect 24299 -2136 24305 -1760
rect 24339 -2136 24345 -1760
rect 24299 -2148 24345 -2136
rect 24417 -1760 24463 -1748
rect 24417 -2136 24423 -1760
rect 24457 -2136 24463 -1760
rect 24541 -1948 24578 -1661
rect 24417 -2148 24463 -2136
rect 24536 -1960 24582 -1948
rect 24536 -2136 24542 -1960
rect 24576 -2136 24582 -1960
rect 24536 -2148 24582 -2136
rect 24654 -1960 24700 -1948
rect 24654 -2136 24660 -1960
rect 24694 -2136 24700 -1960
rect 24654 -2148 24700 -2136
rect 24772 -1960 24818 -1948
rect 24772 -2136 24778 -1960
rect 24812 -2136 24818 -1960
rect 24772 -2148 24818 -2136
rect 24890 -1960 24936 -1948
rect 24890 -2136 24896 -1960
rect 24930 -2136 24936 -1960
rect 24890 -2148 24936 -2136
rect 22333 -2334 22368 -2148
rect 23242 -2232 23276 -2148
rect 24423 -2232 24457 -2148
rect 23242 -2274 24457 -2232
rect 24423 -2294 24457 -2274
rect 24423 -2310 24780 -2294
rect 22333 -2351 23470 -2334
rect 22333 -2385 23420 -2351
rect 23454 -2385 23470 -2351
rect 24423 -2344 24730 -2310
rect 24764 -2344 24780 -2310
rect 24423 -2360 24780 -2344
rect 22333 -2401 23470 -2385
rect 22174 -2446 22250 -2438
rect 22174 -2514 22191 -2446
rect 22248 -2514 22258 -2446
rect 22174 -2522 22250 -2514
rect 22004 -2562 22250 -2554
rect 22004 -2630 22191 -2562
rect 22248 -2630 22258 -2562
rect 22004 -2638 22250 -2630
rect 22004 -2641 22108 -2638
rect 20246 -2730 20338 -2722
rect 20246 -2795 20258 -2730
rect 20326 -2795 20338 -2730
rect 20246 -2807 20338 -2795
rect 21752 -2910 21931 -2648
rect 19189 -2958 20561 -2911
rect 20883 -2957 21931 -2910
rect 16891 -3085 16925 -2962
rect 17363 -2975 17429 -2962
rect 17363 -3009 17379 -2975
rect 17413 -3009 17429 -2975
rect 17363 -3025 17429 -3009
rect 17752 -3085 17786 -2961
rect 18631 -2962 18807 -2961
rect 16886 -3097 16932 -3085
rect 16886 -3273 16892 -3097
rect 16926 -3273 16932 -3097
rect 16886 -3285 16932 -3273
rect 17004 -3097 17124 -3085
rect 17004 -3273 17010 -3097
rect 17044 -3273 17084 -3097
rect 17004 -3285 17084 -3273
rect 17010 -3652 17044 -3285
rect 17078 -3473 17084 -3285
rect 17118 -3473 17124 -3097
rect 17078 -3485 17124 -3473
rect 17196 -3097 17242 -3085
rect 17196 -3473 17202 -3097
rect 17236 -3473 17242 -3097
rect 17196 -3485 17242 -3473
rect 17314 -3097 17360 -3085
rect 17314 -3473 17320 -3097
rect 17354 -3473 17360 -3097
rect 17314 -3485 17360 -3473
rect 17432 -3097 17478 -3085
rect 17432 -3473 17438 -3097
rect 17472 -3473 17478 -3097
rect 17432 -3485 17478 -3473
rect 17550 -3097 17674 -3085
rect 17550 -3473 17556 -3097
rect 17590 -3273 17634 -3097
rect 17668 -3273 17674 -3097
rect 17590 -3285 17674 -3273
rect 17746 -3097 17792 -3085
rect 17746 -3273 17752 -3097
rect 17786 -3273 17792 -3097
rect 17746 -3285 17792 -3273
rect 17590 -3473 17596 -3285
rect 17550 -3485 17596 -3473
rect 17320 -3558 17354 -3485
rect 17305 -3574 17371 -3558
rect 17305 -3608 17321 -3574
rect 17355 -3608 17371 -3574
rect 17305 -3624 17371 -3608
rect 17634 -3652 17668 -3285
rect 17010 -3704 17668 -3652
rect 17308 -3726 17400 -3704
rect 17308 -3778 17320 -3726
rect 17386 -3778 17400 -3726
rect 17308 -3782 17400 -3778
rect 18656 -4476 18807 -2962
rect 20023 -3081 20057 -2958
rect 20495 -2971 20561 -2958
rect 20495 -3005 20511 -2971
rect 20545 -3005 20561 -2971
rect 20495 -3021 20561 -3005
rect 20884 -3081 20918 -2957
rect 20018 -3093 20064 -3081
rect 20018 -3269 20024 -3093
rect 20058 -3269 20064 -3093
rect 20018 -3281 20064 -3269
rect 20136 -3093 20256 -3081
rect 20136 -3269 20142 -3093
rect 20176 -3269 20216 -3093
rect 20136 -3281 20216 -3269
rect 20142 -3648 20176 -3281
rect 20210 -3469 20216 -3281
rect 20250 -3469 20256 -3093
rect 20210 -3481 20256 -3469
rect 20328 -3093 20374 -3081
rect 20328 -3469 20334 -3093
rect 20368 -3469 20374 -3093
rect 20328 -3481 20374 -3469
rect 20446 -3093 20492 -3081
rect 20446 -3469 20452 -3093
rect 20486 -3469 20492 -3093
rect 20446 -3481 20492 -3469
rect 20564 -3093 20610 -3081
rect 20564 -3469 20570 -3093
rect 20604 -3469 20610 -3093
rect 20564 -3481 20610 -3469
rect 20682 -3093 20806 -3081
rect 20682 -3469 20688 -3093
rect 20722 -3269 20766 -3093
rect 20800 -3269 20806 -3093
rect 20722 -3281 20806 -3269
rect 20878 -3093 20924 -3081
rect 20878 -3269 20884 -3093
rect 20918 -3269 20924 -3093
rect 20878 -3281 20924 -3269
rect 20722 -3469 20728 -3281
rect 20682 -3481 20728 -3469
rect 20452 -3554 20486 -3481
rect 20437 -3570 20503 -3554
rect 20437 -3604 20453 -3570
rect 20487 -3604 20503 -3570
rect 20437 -3620 20503 -3604
rect 20766 -3648 20800 -3281
rect 20142 -3700 20800 -3648
rect 20440 -3722 20532 -3700
rect 20440 -3774 20452 -3722
rect 20518 -3774 20532 -3722
rect 20440 -3778 20532 -3774
rect 21780 -4487 21931 -2957
rect 22333 -2911 22368 -2401
rect 22423 -2447 22515 -2434
rect 22423 -2510 22435 -2447
rect 22506 -2510 22515 -2447
rect 22423 -2519 22515 -2510
rect 23508 -2447 23600 -2437
rect 23508 -2509 23520 -2447
rect 23590 -2509 23600 -2447
rect 23508 -2522 23600 -2509
rect 24896 -2502 24931 -2148
rect 23755 -2564 23820 -2561
rect 23755 -2567 23824 -2564
rect 23755 -2627 23761 -2567
rect 23820 -2627 23830 -2567
rect 23755 -2631 23824 -2627
rect 23755 -2633 23820 -2631
rect 24896 -2648 25077 -2502
rect 23390 -2730 23482 -2722
rect 23390 -2795 23402 -2730
rect 23470 -2795 23482 -2730
rect 23390 -2807 23482 -2795
rect 24896 -2910 25076 -2648
rect 22333 -2958 23705 -2911
rect 24027 -2957 25076 -2910
rect 23167 -3081 23201 -2958
rect 23639 -2971 23705 -2958
rect 23639 -3005 23655 -2971
rect 23689 -3005 23705 -2971
rect 23639 -3021 23705 -3005
rect 24028 -3081 24062 -2957
rect 23162 -3093 23208 -3081
rect 23162 -3269 23168 -3093
rect 23202 -3269 23208 -3093
rect 23162 -3281 23208 -3269
rect 23280 -3093 23400 -3081
rect 23280 -3269 23286 -3093
rect 23320 -3269 23360 -3093
rect 23280 -3281 23360 -3269
rect 23286 -3648 23320 -3281
rect 23354 -3469 23360 -3281
rect 23394 -3469 23400 -3093
rect 23354 -3481 23400 -3469
rect 23472 -3093 23518 -3081
rect 23472 -3469 23478 -3093
rect 23512 -3469 23518 -3093
rect 23472 -3481 23518 -3469
rect 23590 -3093 23636 -3081
rect 23590 -3469 23596 -3093
rect 23630 -3469 23636 -3093
rect 23590 -3481 23636 -3469
rect 23708 -3093 23754 -3081
rect 23708 -3469 23714 -3093
rect 23748 -3469 23754 -3093
rect 23708 -3481 23754 -3469
rect 23826 -3093 23950 -3081
rect 23826 -3469 23832 -3093
rect 23866 -3269 23910 -3093
rect 23944 -3269 23950 -3093
rect 23866 -3281 23950 -3269
rect 24022 -3093 24068 -3081
rect 24022 -3269 24028 -3093
rect 24062 -3269 24068 -3093
rect 24022 -3281 24068 -3269
rect 23866 -3469 23872 -3281
rect 23826 -3481 23872 -3469
rect 23596 -3554 23630 -3481
rect 23581 -3570 23647 -3554
rect 23581 -3604 23597 -3570
rect 23631 -3604 23647 -3570
rect 23581 -3620 23647 -3604
rect 23910 -3648 23944 -3281
rect 23286 -3700 23944 -3648
rect 23584 -3722 23676 -3700
rect 23584 -3774 23596 -3722
rect 23662 -3774 23676 -3722
rect 23584 -3778 23676 -3774
rect 24925 -4479 25076 -2957
rect 28137 -4243 28253 2079
rect 28309 -4110 28425 2202
rect 28465 -3959 28581 2382
rect 28648 -3804 28764 2445
rect 28826 -3647 28942 2473
rect 28986 2470 29104 2797
rect 29148 2492 29266 2819
rect 29311 2807 29427 3194
rect 30152 3219 30352 3225
rect 30386 3219 30421 3319
rect 31377 3313 31577 3319
rect 30152 3185 30164 3219
rect 30340 3185 30421 3219
rect 31055 3255 31169 3267
rect 30152 3179 30352 3185
rect 31055 3153 31061 3255
rect 31163 3153 31169 3255
rect 31055 3141 31169 3153
rect 32681 3012 32760 18854
rect 30501 3000 32760 3012
rect 30501 2938 32681 3000
rect 32747 2938 32760 3000
rect 30501 2924 32760 2938
rect 30150 2826 30350 2832
rect 29310 2514 29428 2807
rect 30150 2792 30162 2826
rect 30338 2792 30419 2826
rect 30150 2786 30350 2792
rect 30150 2708 30350 2714
rect 28987 -3485 29103 2470
rect 29148 -3344 29264 2492
rect 29309 2480 29428 2514
rect 29804 2674 30162 2708
rect 30338 2674 30350 2708
rect 29309 -3179 29425 2480
rect 29804 2342 29847 2674
rect 30150 2668 30350 2674
rect 30384 2701 30419 2792
rect 30501 2807 30567 2924
rect 30691 2819 30763 2837
rect 30691 2817 30697 2819
rect 30757 2817 30763 2819
rect 30689 2755 30697 2817
rect 30757 2755 30765 2817
rect 30691 2753 30697 2755
rect 30757 2753 30763 2755
rect 30691 2741 30763 2753
rect 30501 2731 30567 2741
rect 31375 2701 31575 2707
rect 30384 2667 31387 2701
rect 31563 2667 31575 2701
rect 30150 2590 30350 2596
rect 30150 2556 30162 2590
rect 30338 2556 30350 2590
rect 30150 2550 30350 2556
rect 30150 2472 30350 2478
rect 30150 2438 30162 2472
rect 30338 2438 30350 2472
rect 30150 2432 30350 2438
rect 30162 2348 30338 2432
rect 30643 2399 31043 2405
rect 30481 2365 30655 2399
rect 31031 2365 31043 2399
rect 31203 2385 31246 2667
rect 31375 2661 31575 2667
rect 31375 2584 31575 2589
rect 31375 2583 31901 2584
rect 31274 2554 31336 2560
rect 31274 2520 31286 2554
rect 31320 2520 31336 2554
rect 31375 2549 31387 2583
rect 31563 2550 31901 2583
rect 31563 2549 31575 2550
rect 31375 2543 31575 2549
rect 31274 2504 31336 2520
rect 29950 2342 30350 2348
rect 29804 2308 29962 2342
rect 30338 2308 30350 2342
rect 29804 2106 29847 2308
rect 29950 2302 30350 2308
rect 29950 2224 30350 2230
rect 29950 2190 29962 2224
rect 30338 2190 30419 2224
rect 29950 2184 30350 2190
rect 29950 2106 30350 2112
rect 29804 2072 29962 2106
rect 30338 2072 30350 2106
rect 29804 2037 29847 2072
rect 29950 2066 30350 2072
rect 29721 2009 29847 2037
rect 29699 1999 29847 2009
rect 29753 1945 29847 1999
rect 29950 1988 30350 1994
rect 30384 1988 30419 2190
rect 30481 2163 30519 2365
rect 30643 2359 31043 2365
rect 31208 2369 31259 2385
rect 31208 2335 31219 2369
rect 31253 2335 31259 2369
rect 31208 2318 31259 2335
rect 30643 2281 31043 2287
rect 30643 2247 30655 2281
rect 31031 2247 31043 2281
rect 30643 2241 31043 2247
rect 30643 2163 31043 2169
rect 30481 2129 30655 2163
rect 31031 2129 31043 2163
rect 30481 1988 30519 2129
rect 30643 2123 31043 2129
rect 31287 2119 31336 2504
rect 31375 2281 31775 2287
rect 31375 2247 31387 2281
rect 31763 2247 31775 2281
rect 31375 2241 31775 2247
rect 31375 2163 31775 2169
rect 31375 2129 31387 2163
rect 31763 2129 31775 2163
rect 31375 2123 31775 2129
rect 31287 2103 31344 2119
rect 31287 2069 31303 2103
rect 31337 2069 31344 2103
rect 31287 2053 31344 2069
rect 31869 2091 31901 2550
rect 31869 2057 31986 2091
rect 30643 2045 31043 2051
rect 30643 2011 30655 2045
rect 31031 2011 31043 2045
rect 30643 2005 31043 2011
rect 31375 2045 31775 2051
rect 31375 2011 31387 2045
rect 31763 2011 31775 2045
rect 31375 2005 31775 2011
rect 29950 1954 29962 1988
rect 30338 1954 30519 1988
rect 29950 1948 30350 1954
rect 29699 1935 29847 1945
rect 29721 1903 29847 1935
rect 29804 1870 29847 1903
rect 30481 1927 30519 1954
rect 31287 1985 31346 2001
rect 31287 1951 31302 1985
rect 31336 1951 31346 1985
rect 31287 1934 31346 1951
rect 31869 1995 31923 2057
rect 31981 1995 31986 2057
rect 31869 1959 31986 1995
rect 30643 1927 31043 1933
rect 30481 1893 30655 1927
rect 31031 1893 31043 1927
rect 29950 1870 30350 1876
rect 29804 1836 29962 1870
rect 30338 1836 30350 1870
rect 29804 1634 29847 1836
rect 29950 1830 30350 1836
rect 29950 1752 30350 1758
rect 29950 1718 29962 1752
rect 30338 1718 30350 1752
rect 29950 1712 30350 1718
rect 30481 1691 30519 1893
rect 30643 1887 31043 1893
rect 30643 1809 31043 1815
rect 30643 1775 30655 1809
rect 31031 1775 31043 1809
rect 30643 1769 31043 1775
rect 31208 1721 31259 1738
rect 30643 1691 31043 1697
rect 30481 1657 30655 1691
rect 31031 1657 31043 1691
rect 31208 1687 31219 1721
rect 31253 1687 31259 1721
rect 31208 1671 31259 1687
rect 30643 1651 31043 1657
rect 29950 1634 30350 1640
rect 29804 1600 29962 1634
rect 30338 1600 30350 1634
rect 29804 1269 29847 1600
rect 29950 1594 30350 1600
rect 30162 1511 30338 1594
rect 31203 1558 31246 1671
rect 30150 1505 30350 1511
rect 30150 1471 30162 1505
rect 30338 1471 30350 1505
rect 30150 1465 30350 1471
rect 30501 1419 30567 1431
rect 30150 1387 30350 1393
rect 30150 1353 30162 1387
rect 30338 1353 30419 1387
rect 30501 1365 30507 1419
rect 30561 1365 30567 1419
rect 30501 1353 30567 1365
rect 30150 1347 30350 1353
rect 30384 1285 30419 1353
rect 31202 1285 31247 1558
rect 31287 1447 31336 1934
rect 31375 1927 31775 1933
rect 31869 1927 31901 1959
rect 31375 1893 31387 1927
rect 31763 1893 31901 1927
rect 31375 1887 31775 1893
rect 31375 1809 31775 1815
rect 31375 1775 31387 1809
rect 31763 1775 31775 1809
rect 31375 1769 31775 1775
rect 31275 1431 31337 1447
rect 31275 1397 31287 1431
rect 31321 1397 31337 1431
rect 31275 1391 31337 1397
rect 31375 1403 31575 1409
rect 31869 1403 31901 1893
rect 31375 1369 31387 1403
rect 31563 1370 31901 1403
rect 31563 1369 31575 1370
rect 31375 1363 31575 1369
rect 31375 1285 31575 1291
rect 30150 1269 30350 1275
rect 29804 1235 30162 1269
rect 30338 1235 30350 1269
rect 30150 1229 30350 1235
rect 30384 1251 31387 1285
rect 31563 1251 31575 1285
rect 30150 1151 30350 1157
rect 30384 1151 30419 1251
rect 31375 1245 31575 1251
rect 30150 1117 30162 1151
rect 30338 1117 30419 1151
rect 31053 1187 31167 1199
rect 30150 1111 30350 1117
rect 31053 1085 31059 1187
rect 31161 1085 31167 1187
rect 31053 1073 31167 1085
rect 32825 932 32900 19294
rect 30503 921 32900 932
rect 30503 866 32534 921
rect 32604 866 32900 921
rect 30503 854 32900 866
rect 30152 757 30352 763
rect 30152 723 30164 757
rect 30340 723 30421 757
rect 30152 717 30352 723
rect 30152 639 30352 645
rect 29806 605 30164 639
rect 30340 605 30352 639
rect 29806 273 29849 605
rect 30152 599 30352 605
rect 30386 632 30421 723
rect 30503 738 30569 854
rect 30693 750 30765 771
rect 30693 684 30699 750
rect 30759 684 30765 750
rect 30693 672 30765 684
rect 30503 662 30569 672
rect 31377 632 31577 638
rect 30386 598 31389 632
rect 31565 598 31577 632
rect 30152 521 30352 527
rect 30152 487 30164 521
rect 30340 487 30352 521
rect 30152 481 30352 487
rect 30152 403 30352 409
rect 30152 369 30164 403
rect 30340 369 30352 403
rect 30152 363 30352 369
rect 30164 279 30340 363
rect 30645 330 31045 336
rect 30483 296 30657 330
rect 31033 296 31045 330
rect 31205 316 31248 598
rect 31377 592 31577 598
rect 31377 515 31577 520
rect 31377 514 31903 515
rect 31276 485 31338 491
rect 31276 451 31288 485
rect 31322 451 31338 485
rect 31377 480 31389 514
rect 31565 481 31903 514
rect 31565 480 31577 481
rect 31377 474 31577 480
rect 31276 435 31338 451
rect 29952 273 30352 279
rect 29806 239 29964 273
rect 30340 239 30352 273
rect 29806 37 29849 239
rect 29952 233 30352 239
rect 29952 155 30352 161
rect 29952 121 29964 155
rect 30340 121 30421 155
rect 29952 115 30352 121
rect 29952 37 30352 43
rect 29806 3 29964 37
rect 30340 3 30352 37
rect 29806 -32 29849 3
rect 29952 -3 30352 3
rect 29723 -60 29849 -32
rect 29701 -70 29849 -60
rect 29755 -124 29849 -70
rect 29952 -81 30352 -75
rect 30386 -81 30421 121
rect 30483 94 30521 296
rect 30645 290 31045 296
rect 31210 300 31261 316
rect 31210 266 31221 300
rect 31255 266 31261 300
rect 31210 249 31261 266
rect 30645 212 31045 218
rect 30645 178 30657 212
rect 31033 178 31045 212
rect 30645 172 31045 178
rect 30645 94 31045 100
rect 30483 60 30657 94
rect 31033 60 31045 94
rect 30483 -81 30521 60
rect 30645 54 31045 60
rect 31289 50 31338 435
rect 31377 212 31777 218
rect 31377 178 31389 212
rect 31765 178 31777 212
rect 31377 172 31777 178
rect 31377 94 31777 100
rect 31377 60 31389 94
rect 31765 60 31777 94
rect 31377 54 31777 60
rect 31289 34 31346 50
rect 31289 0 31305 34
rect 31339 0 31346 34
rect 31289 -16 31346 0
rect 31871 22 31903 481
rect 31871 -12 31988 22
rect 30645 -24 31045 -18
rect 30645 -58 30657 -24
rect 31033 -58 31045 -24
rect 30645 -64 31045 -58
rect 31377 -24 31777 -18
rect 31377 -58 31389 -24
rect 31765 -58 31777 -24
rect 31377 -64 31777 -58
rect 29952 -115 29964 -81
rect 30340 -115 30521 -81
rect 29952 -121 30352 -115
rect 29701 -134 29849 -124
rect 29723 -166 29849 -134
rect 29806 -199 29849 -166
rect 30483 -142 30521 -115
rect 31289 -84 31348 -68
rect 31289 -118 31304 -84
rect 31338 -118 31348 -84
rect 31289 -135 31348 -118
rect 31871 -74 31925 -12
rect 31983 -74 31988 -12
rect 31871 -110 31988 -74
rect 30645 -142 31045 -136
rect 30483 -176 30657 -142
rect 31033 -176 31045 -142
rect 29952 -199 30352 -193
rect 29806 -233 29964 -199
rect 30340 -233 30352 -199
rect 29806 -435 29849 -233
rect 29952 -239 30352 -233
rect 29952 -317 30352 -311
rect 29952 -351 29964 -317
rect 30340 -351 30352 -317
rect 29952 -357 30352 -351
rect 30483 -378 30521 -176
rect 30645 -182 31045 -176
rect 30645 -260 31045 -254
rect 30645 -294 30657 -260
rect 31033 -294 31045 -260
rect 30645 -300 31045 -294
rect 31210 -348 31261 -331
rect 30645 -378 31045 -372
rect 30483 -412 30657 -378
rect 31033 -412 31045 -378
rect 31210 -382 31221 -348
rect 31255 -382 31261 -348
rect 31210 -398 31261 -382
rect 30645 -418 31045 -412
rect 29952 -435 30352 -429
rect 29806 -469 29964 -435
rect 30340 -469 30352 -435
rect 29806 -800 29849 -469
rect 29952 -475 30352 -469
rect 30164 -558 30340 -475
rect 31205 -511 31248 -398
rect 30152 -564 30352 -558
rect 30152 -598 30164 -564
rect 30340 -598 30352 -564
rect 30152 -604 30352 -598
rect 30503 -650 30569 -638
rect 30152 -682 30352 -676
rect 30152 -716 30164 -682
rect 30340 -716 30421 -682
rect 30503 -704 30509 -650
rect 30563 -704 30569 -650
rect 30503 -716 30569 -704
rect 30152 -722 30352 -716
rect 30386 -784 30421 -716
rect 31204 -784 31249 -511
rect 31289 -622 31338 -135
rect 31377 -142 31777 -136
rect 31871 -142 31903 -110
rect 31377 -176 31389 -142
rect 31765 -176 31903 -142
rect 31377 -182 31777 -176
rect 31377 -260 31777 -254
rect 31377 -294 31389 -260
rect 31765 -294 31777 -260
rect 31377 -300 31777 -294
rect 31277 -638 31339 -622
rect 31277 -672 31289 -638
rect 31323 -672 31339 -638
rect 31277 -678 31339 -672
rect 31377 -666 31577 -660
rect 31871 -666 31903 -176
rect 31377 -700 31389 -666
rect 31565 -699 31903 -666
rect 31565 -700 31577 -699
rect 31377 -706 31577 -700
rect 31377 -784 31577 -778
rect 30152 -800 30352 -794
rect 29806 -834 30164 -800
rect 30340 -834 30352 -800
rect 30152 -840 30352 -834
rect 30386 -818 31389 -784
rect 31565 -818 31577 -784
rect 30152 -918 30352 -912
rect 30386 -918 30421 -818
rect 31377 -824 31577 -818
rect 30152 -952 30164 -918
rect 30340 -952 30421 -918
rect 31055 -882 31169 -870
rect 30152 -958 30352 -952
rect 31055 -984 31061 -882
rect 31163 -984 31169 -882
rect 31055 -996 31169 -984
rect 32960 -1147 33035 19715
rect 33097 19906 33170 20145
rect 33097 13247 33172 19906
rect 33097 13195 33107 13247
rect 33168 13195 33178 13247
rect 33097 11159 33172 13195
rect 33244 12876 33329 20563
rect 33409 13053 33482 20986
rect 33542 13209 33615 21216
rect 33672 21529 33744 21868
rect 33672 13360 33745 21529
rect 33810 13512 33883 22289
rect 33952 19663 34046 22721
rect 34112 19853 34190 23140
rect 34249 19997 34330 23561
rect 39088 21693 39181 23587
rect 39244 23528 39710 23550
rect 39998 23528 40064 23624
rect 41829 23634 41835 23810
rect 41869 23634 41875 23810
rect 41829 23622 41875 23634
rect 41947 23810 41993 23822
rect 41947 23634 41953 23810
rect 41987 23634 41993 23810
rect 41947 23622 41993 23634
rect 42065 23810 42111 23822
rect 42065 23634 42071 23810
rect 42105 23634 42111 23810
rect 42065 23622 42111 23634
rect 42183 23810 42229 23822
rect 42183 23634 42189 23810
rect 42223 23755 42229 23810
rect 42348 23810 42394 23822
rect 42348 23755 42354 23810
rect 42223 23667 42354 23755
rect 42223 23634 42229 23667
rect 42183 23622 42229 23634
rect 42348 23634 42354 23667
rect 42388 23634 42394 23810
rect 42348 23622 42394 23634
rect 42466 23810 42512 23822
rect 42466 23634 42472 23810
rect 42506 23634 42512 23810
rect 42466 23622 42512 23634
rect 42584 23810 42630 23822
rect 42584 23634 42590 23810
rect 42624 23634 42630 23810
rect 42584 23622 42630 23634
rect 42702 23810 42748 23822
rect 42702 23634 42708 23810
rect 42742 23634 42748 23810
rect 42702 23622 42748 23634
rect 41835 23583 41869 23622
rect 42071 23583 42105 23622
rect 41835 23548 42105 23583
rect 42472 23584 42505 23622
rect 42708 23584 42741 23622
rect 42472 23548 42741 23584
rect 39244 23480 40064 23528
rect 41869 23547 42105 23548
rect 39244 23449 39710 23480
rect 41869 23473 42001 23547
rect 39244 23193 39349 23449
rect 41859 23365 41869 23473
rect 42001 23365 42011 23473
rect 39244 23087 39307 23193
rect 39419 23087 39429 23193
rect 40011 23169 40231 23189
rect 39244 23076 39393 23087
rect 39244 21899 39349 23076
rect 40011 23061 40055 23169
rect 40187 23061 40231 23169
rect 40011 23019 40231 23061
rect 42809 23034 42871 24605
rect 43061 24597 43107 24609
rect 43061 24221 43067 24597
rect 43101 24221 43107 24597
rect 43061 24209 43107 24221
rect 43179 24597 43225 24609
rect 43179 24221 43185 24597
rect 43219 24221 43225 24597
rect 43179 24209 43225 24221
rect 43297 24597 43343 24609
rect 43297 24221 43303 24597
rect 43337 24221 43343 24597
rect 43297 24209 43343 24221
rect 43415 24597 43461 24609
rect 43415 24221 43421 24597
rect 43455 24221 43461 24597
rect 43415 24209 43461 24221
rect 43533 24597 43579 24609
rect 43533 24221 43539 24597
rect 43573 24221 43579 24597
rect 43533 24209 43579 24221
rect 43651 24597 43697 24609
rect 43651 24221 43657 24597
rect 43691 24221 43697 24597
rect 43651 24209 43697 24221
rect 43769 24597 43815 24609
rect 43769 24221 43775 24597
rect 43809 24221 43815 24597
rect 46114 24636 47091 24666
rect 46114 24530 46146 24636
rect 46350 24530 46382 24636
rect 46586 24530 46618 24636
rect 46822 24530 46854 24636
rect 47057 24530 47091 24636
rect 46107 24518 46153 24530
rect 46107 24342 46113 24518
rect 46147 24342 46153 24518
rect 46107 24330 46153 24342
rect 46225 24518 46271 24530
rect 46225 24342 46231 24518
rect 46265 24342 46271 24518
rect 46225 24330 46271 24342
rect 46343 24518 46389 24530
rect 46343 24342 46349 24518
rect 46383 24342 46389 24518
rect 46343 24330 46389 24342
rect 46461 24518 46507 24530
rect 46461 24342 46467 24518
rect 46501 24342 46507 24518
rect 46461 24330 46507 24342
rect 46579 24518 46625 24530
rect 46579 24342 46585 24518
rect 46619 24342 46625 24518
rect 46579 24330 46625 24342
rect 46697 24518 46743 24530
rect 46697 24342 46703 24518
rect 46737 24342 46743 24518
rect 46697 24330 46743 24342
rect 46815 24518 46861 24530
rect 46815 24342 46821 24518
rect 46855 24342 46861 24518
rect 46815 24330 46861 24342
rect 46933 24518 46979 24530
rect 46933 24342 46939 24518
rect 46973 24342 46979 24518
rect 46933 24330 46979 24342
rect 47051 24518 47097 24530
rect 47051 24342 47057 24518
rect 47091 24342 47097 24518
rect 47051 24330 47097 24342
rect 47169 24518 47215 24530
rect 47169 24342 47175 24518
rect 47209 24342 47215 24518
rect 47169 24330 47215 24342
rect 43769 24209 43815 24221
rect 46230 24236 46266 24330
rect 46466 24236 46502 24330
rect 46702 24237 46738 24330
rect 46864 24282 46930 24289
rect 46864 24248 46880 24282
rect 46914 24248 46930 24282
rect 46864 24237 46930 24248
rect 46702 24236 46930 24237
rect 43067 24167 43101 24209
rect 43303 24167 43337 24209
rect 43067 24139 43337 24167
rect 43421 24168 43455 24209
rect 43657 24168 43691 24209
rect 43421 24139 43691 24168
rect 43067 24091 43101 24139
rect 43067 24061 43130 24091
rect 43095 23969 43130 24061
rect 43602 24031 43702 24052
rect 43602 23977 43616 24031
rect 43681 23977 43702 24031
rect 43602 23972 43702 23977
rect 43775 24026 43809 24209
rect 46230 24207 46930 24236
rect 46230 24206 46812 24207
rect 46350 24093 46384 24206
rect 46746 24165 46812 24206
rect 46746 24131 46762 24165
rect 46796 24131 46812 24165
rect 46746 24124 46812 24131
rect 47174 24125 47209 24330
rect 47381 24125 47448 24715
rect 49140 24692 49181 24724
rect 49427 24720 49437 24786
rect 49493 24720 49503 24786
rect 50173 24762 50183 24870
rect 50315 24807 50325 24870
rect 53044 24811 53264 24831
rect 50315 24796 50327 24807
rect 50315 24762 50328 24796
rect 50183 24724 50328 24762
rect 50287 24696 50328 24724
rect 48556 24664 48826 24692
rect 48297 24598 48307 24664
rect 48373 24598 48383 24664
rect 48556 24602 48590 24664
rect 48792 24602 48826 24664
rect 48910 24664 49181 24692
rect 49698 24668 49968 24696
rect 48910 24602 48944 24664
rect 49146 24602 49181 24664
rect 49322 24652 49493 24668
rect 49322 24618 49453 24652
rect 49487 24618 49493 24652
rect 49322 24602 49493 24618
rect 49698 24606 49732 24668
rect 49934 24606 49968 24668
rect 50052 24668 50328 24696
rect 50052 24606 50086 24668
rect 50288 24606 50328 24668
rect 53044 24703 53088 24811
rect 53220 24703 53264 24811
rect 54841 24769 54897 24777
rect 53044 24661 53264 24703
rect 53915 24761 54897 24769
rect 53915 24727 54857 24761
rect 54891 24727 54897 24761
rect 55560 24757 55570 24865
rect 55702 24802 55712 24865
rect 55702 24791 55714 24802
rect 55702 24757 55715 24791
rect 55971 24781 56027 24783
rect 53915 24711 54897 24727
rect 55570 24719 55715 24757
rect 53915 24710 54894 24711
rect 48432 24590 48478 24602
rect 48432 24214 48438 24590
rect 48472 24214 48478 24590
rect 48432 24202 48478 24214
rect 48550 24590 48596 24602
rect 48550 24214 48556 24590
rect 48590 24214 48596 24590
rect 48550 24202 48596 24214
rect 48668 24590 48714 24602
rect 48668 24214 48674 24590
rect 48708 24214 48714 24590
rect 48668 24202 48714 24214
rect 48786 24590 48832 24602
rect 48786 24214 48792 24590
rect 48826 24214 48832 24590
rect 48786 24202 48832 24214
rect 48904 24590 48950 24602
rect 48904 24214 48910 24590
rect 48944 24214 48950 24590
rect 48904 24202 48950 24214
rect 49022 24590 49068 24602
rect 49022 24214 49028 24590
rect 49062 24214 49068 24590
rect 49022 24202 49068 24214
rect 49140 24590 49186 24602
rect 49140 24214 49146 24590
rect 49180 24214 49186 24590
rect 49140 24202 49186 24214
rect 47174 24097 47448 24125
rect 46820 24093 47448 24097
rect 46344 24081 46390 24093
rect 44777 24040 44884 24042
rect 43775 23972 43884 24026
rect 43095 23933 43322 23969
rect 43095 23826 43130 23933
rect 43256 23899 43322 23933
rect 43256 23865 43272 23899
rect 43306 23865 43322 23899
rect 43603 23957 43700 23972
rect 43603 23890 43660 23957
rect 43256 23859 43322 23865
rect 43497 23854 43766 23890
rect 43497 23826 43530 23854
rect 43733 23826 43766 23854
rect 43850 23826 43884 23972
rect 44701 23965 44711 24040
rect 44779 23965 44884 24040
rect 44728 23964 44884 23965
rect 42971 23814 43017 23826
rect 42971 23638 42977 23814
rect 43011 23638 43017 23814
rect 42971 23626 43017 23638
rect 43089 23814 43135 23826
rect 43089 23638 43095 23814
rect 43129 23638 43135 23814
rect 43089 23626 43135 23638
rect 43207 23814 43253 23826
rect 43207 23638 43213 23814
rect 43247 23638 43253 23814
rect 43207 23626 43253 23638
rect 43325 23814 43371 23826
rect 43325 23638 43331 23814
rect 43365 23759 43371 23814
rect 43490 23814 43536 23826
rect 43490 23759 43496 23814
rect 43365 23671 43496 23759
rect 43365 23638 43371 23671
rect 43325 23626 43371 23638
rect 43490 23638 43496 23671
rect 43530 23638 43536 23814
rect 43490 23626 43536 23638
rect 43608 23814 43654 23826
rect 43608 23638 43614 23814
rect 43648 23638 43654 23814
rect 43608 23626 43654 23638
rect 43726 23814 43772 23826
rect 43726 23638 43732 23814
rect 43766 23638 43772 23814
rect 43726 23626 43772 23638
rect 43844 23814 43890 23826
rect 43844 23638 43850 23814
rect 43884 23638 43890 23814
rect 43844 23626 43890 23638
rect 42977 23587 43011 23626
rect 43213 23587 43247 23626
rect 42977 23551 43247 23587
rect 43614 23588 43647 23626
rect 43850 23588 43883 23626
rect 43614 23552 43883 23588
rect 42977 23550 43143 23551
rect 43011 23471 43143 23550
rect 43001 23363 43011 23471
rect 43143 23363 43153 23471
rect 39615 22989 40592 23019
rect 42809 23017 42872 23034
rect 42734 23013 42872 23017
rect 39615 22883 39647 22989
rect 39851 22883 39883 22989
rect 40087 22883 40119 22989
rect 40323 22883 40355 22989
rect 40558 22883 40592 22989
rect 40902 22979 42872 23013
rect 40900 22950 42872 22979
rect 40900 22934 40946 22950
rect 42734 22948 42872 22950
rect 39608 22871 39654 22883
rect 39608 22695 39614 22871
rect 39648 22695 39654 22871
rect 39608 22683 39654 22695
rect 39726 22871 39772 22883
rect 39726 22695 39732 22871
rect 39766 22695 39772 22871
rect 39726 22683 39772 22695
rect 39844 22871 39890 22883
rect 39844 22695 39850 22871
rect 39884 22695 39890 22871
rect 39844 22683 39890 22695
rect 39962 22871 40008 22883
rect 39962 22695 39968 22871
rect 40002 22695 40008 22871
rect 39962 22683 40008 22695
rect 40080 22871 40126 22883
rect 40080 22695 40086 22871
rect 40120 22695 40126 22871
rect 40080 22683 40126 22695
rect 40198 22871 40244 22883
rect 40198 22695 40204 22871
rect 40238 22695 40244 22871
rect 40198 22683 40244 22695
rect 40316 22871 40362 22883
rect 40316 22695 40322 22871
rect 40356 22695 40362 22871
rect 40316 22683 40362 22695
rect 40434 22871 40480 22883
rect 40434 22695 40440 22871
rect 40474 22695 40480 22871
rect 40434 22683 40480 22695
rect 40552 22871 40598 22883
rect 40552 22695 40558 22871
rect 40592 22695 40598 22871
rect 40552 22683 40598 22695
rect 40670 22871 40716 22883
rect 40670 22695 40676 22871
rect 40710 22695 40716 22871
rect 40670 22683 40716 22695
rect 39731 22589 39767 22683
rect 39967 22589 40003 22683
rect 40203 22590 40239 22683
rect 40365 22635 40431 22642
rect 40365 22601 40381 22635
rect 40415 22601 40431 22635
rect 40365 22590 40431 22601
rect 40203 22589 40431 22590
rect 39731 22560 40431 22589
rect 39731 22559 40313 22560
rect 39851 22446 39885 22559
rect 40247 22518 40313 22559
rect 40247 22484 40263 22518
rect 40297 22484 40313 22518
rect 40247 22477 40313 22484
rect 40675 22465 40710 22683
rect 40899 22482 40946 22934
rect 41858 22718 41868 22826
rect 42000 22718 42010 22826
rect 43756 22718 43766 22826
rect 43898 22718 43908 22826
rect 41868 22678 42000 22718
rect 43766 22678 43898 22718
rect 41867 22612 42000 22678
rect 43765 22612 43898 22678
rect 41196 22569 42669 22612
rect 40899 22466 40945 22482
rect 40864 22465 40945 22466
rect 40675 22450 40945 22465
rect 40321 22446 40945 22450
rect 39845 22434 39891 22446
rect 39580 21956 39590 22074
rect 39708 22042 39718 22074
rect 39845 22058 39851 22434
rect 39885 22058 39891 22434
rect 39845 22046 39891 22058
rect 39963 22434 40009 22446
rect 39963 22058 39969 22434
rect 40003 22058 40009 22434
rect 39963 22046 40009 22058
rect 40081 22434 40127 22446
rect 40081 22058 40087 22434
rect 40121 22082 40127 22434
rect 40198 22434 40244 22446
rect 40198 22258 40204 22434
rect 40238 22258 40244 22434
rect 40198 22246 40244 22258
rect 40316 22434 40945 22446
rect 40316 22258 40322 22434
rect 40356 22422 40945 22434
rect 40356 22421 40598 22422
rect 40356 22258 40362 22421
rect 40864 22420 40945 22422
rect 41196 22266 41230 22569
rect 41562 22466 41596 22569
rect 41798 22466 41832 22569
rect 42034 22466 42068 22569
rect 42270 22466 42304 22569
rect 41556 22454 41602 22466
rect 40316 22246 40362 22258
rect 41072 22254 41118 22266
rect 40204 22130 40239 22246
rect 40335 22130 40443 22140
rect 40204 22082 40335 22130
rect 40121 22058 40335 22082
rect 40081 22046 40335 22058
rect 40087 22042 40335 22046
rect 39708 22014 39723 22042
rect 39708 22008 39960 22014
rect 39708 21974 39910 22008
rect 39944 21974 39960 22008
rect 39708 21958 39960 21974
rect 40012 22008 40078 22014
rect 40012 21974 40028 22008
rect 40062 21974 40078 22008
rect 40261 21998 40335 22042
rect 41072 22078 41078 22254
rect 41112 22078 41118 22254
rect 41072 22066 41118 22078
rect 41190 22254 41236 22266
rect 41190 22078 41196 22254
rect 41230 22078 41236 22254
rect 41190 22066 41236 22078
rect 41308 22254 41354 22266
rect 41308 22078 41314 22254
rect 41348 22078 41354 22254
rect 41308 22066 41354 22078
rect 41426 22254 41472 22266
rect 41556 22254 41562 22454
rect 41426 22078 41432 22254
rect 41466 22078 41562 22254
rect 41596 22078 41602 22454
rect 41426 22066 41472 22078
rect 41556 22066 41602 22078
rect 41674 22454 41720 22466
rect 41674 22078 41680 22454
rect 41714 22078 41720 22454
rect 41674 22066 41720 22078
rect 41792 22454 41838 22466
rect 41792 22078 41798 22454
rect 41832 22078 41838 22454
rect 41792 22066 41838 22078
rect 41910 22454 41956 22466
rect 41910 22078 41916 22454
rect 41950 22078 41956 22454
rect 41910 22066 41956 22078
rect 42028 22454 42074 22466
rect 42028 22078 42034 22454
rect 42068 22078 42074 22454
rect 42028 22066 42074 22078
rect 42146 22454 42192 22466
rect 42146 22078 42152 22454
rect 42186 22078 42192 22454
rect 42146 22066 42192 22078
rect 42264 22454 42310 22466
rect 42264 22078 42270 22454
rect 42304 22254 42310 22454
rect 42635 22266 42669 22569
rect 43094 22569 44567 22612
rect 43094 22266 43128 22569
rect 43460 22466 43494 22569
rect 43696 22466 43730 22569
rect 43932 22466 43966 22569
rect 44168 22466 44202 22569
rect 43454 22454 43500 22466
rect 42393 22254 42439 22266
rect 42304 22078 42399 22254
rect 42433 22078 42439 22254
rect 42264 22066 42310 22078
rect 42393 22066 42439 22078
rect 42511 22254 42557 22266
rect 42511 22078 42517 22254
rect 42551 22078 42557 22254
rect 42511 22066 42557 22078
rect 42629 22254 42675 22266
rect 42629 22078 42635 22254
rect 42669 22078 42675 22254
rect 42629 22066 42675 22078
rect 42747 22254 42793 22266
rect 42747 22078 42753 22254
rect 42787 22078 42793 22254
rect 42747 22066 42793 22078
rect 42970 22254 43016 22266
rect 42970 22078 42976 22254
rect 43010 22078 43016 22254
rect 42970 22066 43016 22078
rect 43088 22254 43134 22266
rect 43088 22078 43094 22254
rect 43128 22078 43134 22254
rect 43088 22066 43134 22078
rect 43206 22254 43252 22266
rect 43206 22078 43212 22254
rect 43246 22078 43252 22254
rect 43206 22066 43252 22078
rect 43324 22254 43370 22266
rect 43454 22254 43460 22454
rect 43324 22078 43330 22254
rect 43364 22078 43460 22254
rect 43494 22078 43500 22454
rect 43324 22066 43370 22078
rect 43454 22066 43500 22078
rect 43572 22454 43618 22466
rect 43572 22078 43578 22454
rect 43612 22078 43618 22454
rect 43572 22066 43618 22078
rect 43690 22454 43736 22466
rect 43690 22078 43696 22454
rect 43730 22078 43736 22454
rect 43690 22066 43736 22078
rect 43808 22454 43854 22466
rect 43808 22078 43814 22454
rect 43848 22078 43854 22454
rect 43808 22066 43854 22078
rect 43926 22454 43972 22466
rect 43926 22078 43932 22454
rect 43966 22078 43972 22454
rect 43926 22066 43972 22078
rect 44044 22454 44090 22466
rect 44044 22078 44050 22454
rect 44084 22078 44090 22454
rect 44044 22066 44090 22078
rect 44162 22454 44208 22466
rect 44162 22078 44168 22454
rect 44202 22254 44208 22454
rect 44533 22266 44567 22569
rect 44291 22254 44337 22266
rect 44202 22078 44297 22254
rect 44331 22078 44337 22254
rect 44162 22066 44208 22078
rect 44291 22066 44337 22078
rect 44409 22254 44455 22266
rect 44409 22078 44415 22254
rect 44449 22078 44455 22254
rect 44409 22066 44455 22078
rect 44527 22254 44573 22266
rect 44527 22078 44533 22254
rect 44567 22078 44573 22254
rect 44527 22066 44573 22078
rect 44645 22254 44691 22266
rect 44645 22078 44651 22254
rect 44685 22078 44691 22254
rect 44777 22220 44884 23964
rect 45172 23751 45461 23777
rect 45172 23607 45190 23751
rect 45426 23688 45461 23751
rect 46344 23705 46350 24081
rect 46384 23705 46390 24081
rect 46344 23693 46390 23705
rect 46462 24081 46508 24093
rect 46462 23705 46468 24081
rect 46502 23705 46508 24081
rect 46462 23693 46508 23705
rect 46580 24081 46626 24093
rect 46580 23705 46586 24081
rect 46620 23729 46626 24081
rect 46697 24081 46743 24093
rect 46697 23905 46703 24081
rect 46737 23905 46743 24081
rect 46697 23893 46743 23905
rect 46815 24081 47448 24093
rect 46815 23905 46821 24081
rect 46855 24068 47448 24081
rect 48438 24160 48472 24202
rect 48674 24160 48708 24202
rect 48438 24132 48708 24160
rect 48792 24161 48826 24202
rect 49028 24161 49062 24202
rect 48792 24132 49062 24161
rect 48438 24084 48472 24132
rect 46855 23905 46861 24068
rect 48438 24054 48501 24084
rect 46815 23893 46861 23905
rect 48466 23962 48501 24054
rect 48466 23926 48693 23962
rect 48963 23951 48973 24048
rect 49072 23951 49082 24048
rect 49146 24019 49180 24202
rect 49146 23965 49255 24019
rect 46703 23777 46738 23893
rect 48466 23819 48501 23926
rect 48627 23892 48693 23926
rect 48627 23858 48643 23892
rect 48677 23858 48693 23892
rect 48974 23950 49071 23951
rect 48974 23883 49031 23950
rect 48627 23852 48693 23858
rect 48868 23847 49137 23883
rect 48868 23819 48901 23847
rect 49104 23819 49137 23847
rect 49221 23819 49255 23965
rect 48342 23807 48388 23819
rect 46834 23777 46942 23787
rect 46703 23729 46834 23777
rect 46620 23705 46834 23729
rect 46580 23693 46834 23705
rect 46586 23689 46834 23693
rect 45426 23661 46222 23688
rect 45426 23655 46459 23661
rect 45426 23621 46409 23655
rect 46443 23621 46459 23655
rect 45426 23607 46459 23621
rect 45172 23605 46459 23607
rect 46511 23655 46577 23661
rect 46511 23621 46527 23655
rect 46561 23621 46577 23655
rect 46760 23645 46834 23689
rect 46834 23635 46942 23645
rect 45172 23589 46222 23605
rect 45172 23588 46159 23589
rect 45172 23584 45694 23588
rect 45172 23583 45461 23584
rect 45189 22220 45477 22223
rect 44777 22104 45477 22220
rect 44777 22101 44884 22104
rect 44645 22066 44691 22078
rect 40335 21988 40443 21998
rect 41078 22032 41112 22066
rect 41680 22032 41714 22066
rect 41916 22032 41950 22066
rect 41078 21997 41237 22032
rect 41680 21997 41950 22032
rect 42517 22032 42551 22066
rect 42753 22032 42787 22066
rect 42517 21997 42787 22032
rect 42976 22032 43010 22066
rect 43578 22032 43612 22066
rect 43814 22032 43848 22066
rect 42976 21997 43135 22032
rect 43578 21997 43848 22032
rect 44415 22032 44449 22066
rect 44651 22032 44685 22066
rect 44415 21997 44685 22032
rect 45189 22061 45477 22104
rect 39708 21956 39723 21958
rect 39623 21942 39723 21956
rect 39623 21899 39723 21900
rect 39244 21878 39723 21899
rect 40012 21878 40078 21974
rect 39244 21830 40078 21878
rect 39244 21801 39723 21830
rect 39244 21799 39349 21801
rect 39623 21800 39723 21801
rect 39077 21614 39087 21693
rect 39180 21614 39190 21693
rect 39088 20440 39181 21614
rect 40006 21565 40226 21585
rect 40006 21457 40050 21565
rect 40182 21457 40226 21565
rect 40006 21415 40226 21457
rect 39610 21385 40587 21415
rect 39610 21279 39642 21385
rect 39846 21279 39878 21385
rect 40082 21279 40114 21385
rect 40318 21279 40350 21385
rect 40553 21279 40587 21385
rect 39603 21267 39649 21279
rect 39603 21091 39609 21267
rect 39643 21091 39649 21267
rect 39603 21079 39649 21091
rect 39721 21267 39767 21279
rect 39721 21091 39727 21267
rect 39761 21091 39767 21267
rect 39721 21079 39767 21091
rect 39839 21267 39885 21279
rect 39839 21091 39845 21267
rect 39879 21091 39885 21267
rect 39839 21079 39885 21091
rect 39957 21267 40003 21279
rect 39957 21091 39963 21267
rect 39997 21091 40003 21267
rect 39957 21079 40003 21091
rect 40075 21267 40121 21279
rect 40075 21091 40081 21267
rect 40115 21091 40121 21267
rect 40075 21079 40121 21091
rect 40193 21267 40239 21279
rect 40193 21091 40199 21267
rect 40233 21091 40239 21267
rect 40193 21079 40239 21091
rect 40311 21267 40357 21279
rect 40311 21091 40317 21267
rect 40351 21091 40357 21267
rect 40311 21079 40357 21091
rect 40429 21267 40475 21279
rect 40429 21091 40435 21267
rect 40469 21091 40475 21267
rect 40429 21079 40475 21091
rect 40547 21267 40593 21279
rect 40547 21091 40553 21267
rect 40587 21091 40593 21267
rect 40547 21079 40593 21091
rect 40665 21267 40711 21279
rect 40665 21091 40671 21267
rect 40705 21091 40711 21267
rect 40665 21079 40711 21091
rect 41203 21213 41237 21997
rect 41916 21935 41950 21997
rect 41505 21897 42247 21935
rect 41505 21773 41539 21897
rect 41741 21773 41775 21897
rect 41977 21773 42011 21897
rect 42213 21773 42247 21897
rect 42503 21790 42513 21856
rect 42576 21790 42586 21856
rect 41499 21761 41545 21773
rect 41499 21385 41505 21761
rect 41539 21385 41545 21761
rect 41499 21373 41545 21385
rect 41617 21761 41663 21773
rect 41617 21385 41623 21761
rect 41657 21385 41663 21761
rect 41617 21373 41663 21385
rect 41735 21761 41781 21773
rect 41735 21385 41741 21761
rect 41775 21385 41781 21761
rect 41735 21373 41781 21385
rect 41853 21761 41899 21773
rect 41853 21385 41859 21761
rect 41893 21385 41899 21761
rect 41853 21373 41899 21385
rect 41971 21761 42017 21773
rect 41971 21385 41977 21761
rect 42011 21385 42017 21761
rect 41971 21373 42017 21385
rect 42089 21761 42135 21773
rect 42089 21385 42095 21761
rect 42129 21385 42135 21761
rect 42089 21373 42135 21385
rect 42207 21761 42253 21773
rect 42207 21385 42213 21761
rect 42247 21385 42253 21761
rect 42207 21373 42253 21385
rect 42619 21214 42653 21997
rect 42346 21213 42653 21214
rect 41203 21208 41519 21213
rect 42233 21208 42653 21213
rect 41203 21197 41586 21208
rect 41203 21170 41535 21197
rect 39726 20985 39762 21079
rect 39962 20985 39998 21079
rect 40198 20986 40234 21079
rect 40360 21031 40426 21038
rect 40360 20997 40376 21031
rect 40410 20997 40426 21031
rect 40360 20986 40426 20997
rect 40198 20985 40426 20986
rect 39726 20956 40426 20985
rect 39726 20955 40308 20956
rect 39846 20842 39880 20955
rect 40242 20914 40308 20955
rect 40242 20880 40258 20914
rect 40292 20880 40308 20914
rect 40242 20873 40308 20880
rect 40670 20846 40705 21079
rect 41203 21041 41237 21170
rect 41519 21163 41535 21170
rect 41569 21163 41586 21197
rect 41519 21157 41586 21163
rect 42166 21197 42653 21208
rect 42166 21163 42183 21197
rect 42217 21170 42653 21197
rect 42217 21163 42233 21170
rect 42346 21169 42653 21170
rect 42166 21157 42233 21163
rect 41344 21130 41400 21142
rect 41344 21096 41350 21130
rect 41384 21129 41400 21130
rect 42457 21129 42513 21141
rect 41384 21113 41851 21129
rect 41384 21096 41801 21113
rect 41344 21080 41801 21096
rect 41785 21079 41801 21080
rect 41835 21079 41851 21113
rect 41785 21072 41851 21079
rect 41903 21114 42473 21129
rect 41903 21080 41919 21114
rect 41953 21095 42473 21114
rect 42507 21095 42513 21129
rect 41953 21080 42513 21095
rect 41903 21070 41970 21080
rect 42457 21079 42513 21080
rect 42619 21041 42653 21169
rect 43101 21213 43135 21997
rect 43814 21935 43848 21997
rect 43403 21897 44145 21935
rect 43403 21773 43437 21897
rect 43639 21773 43673 21897
rect 43875 21773 43909 21897
rect 44111 21773 44145 21897
rect 43397 21761 43443 21773
rect 43397 21385 43403 21761
rect 43437 21385 43443 21761
rect 43397 21373 43443 21385
rect 43515 21761 43561 21773
rect 43515 21385 43521 21761
rect 43555 21385 43561 21761
rect 43515 21373 43561 21385
rect 43633 21761 43679 21773
rect 43633 21385 43639 21761
rect 43673 21385 43679 21761
rect 43633 21373 43679 21385
rect 43751 21761 43797 21773
rect 43751 21385 43757 21761
rect 43791 21385 43797 21761
rect 43751 21373 43797 21385
rect 43869 21761 43915 21773
rect 43869 21385 43875 21761
rect 43909 21385 43915 21761
rect 43869 21373 43915 21385
rect 43987 21761 44033 21773
rect 43987 21385 43993 21761
rect 44027 21385 44033 21761
rect 43987 21373 44033 21385
rect 44105 21761 44151 21773
rect 44105 21385 44111 21761
rect 44145 21385 44151 21761
rect 44105 21373 44151 21385
rect 44517 21214 44551 21997
rect 45189 21955 45325 22061
rect 45437 22059 45477 22061
rect 45443 22048 45477 22059
rect 45189 21953 45331 21955
rect 45443 21953 45478 22048
rect 45189 21944 45478 21953
rect 45189 21943 45477 21944
rect 45189 21942 45445 21943
rect 44129 21213 44198 21214
rect 44244 21213 44551 21214
rect 43101 21208 43417 21213
rect 44129 21209 44551 21213
rect 43101 21197 43484 21208
rect 43101 21170 43433 21197
rect 43101 21041 43135 21170
rect 43417 21163 43433 21170
rect 43467 21163 43484 21197
rect 43417 21157 43484 21163
rect 44062 21198 44551 21209
rect 44062 21164 44079 21198
rect 44113 21170 44551 21198
rect 44113 21164 44129 21170
rect 44244 21169 44551 21170
rect 44062 21158 44129 21164
rect 43242 21130 43298 21142
rect 43242 21096 43248 21130
rect 43282 21129 43298 21130
rect 44355 21129 44411 21141
rect 43282 21113 43749 21129
rect 43282 21096 43699 21113
rect 43242 21080 43699 21096
rect 43683 21079 43699 21080
rect 43733 21079 43749 21113
rect 43683 21072 43749 21079
rect 43801 21114 44371 21129
rect 43801 21080 43817 21114
rect 43851 21095 44371 21114
rect 44405 21095 44411 21129
rect 43851 21080 44411 21095
rect 43801 21070 43868 21080
rect 44355 21079 44411 21080
rect 44517 21041 44551 21169
rect 44632 21819 44699 21843
rect 44632 21785 44649 21819
rect 44683 21785 44699 21819
rect 40316 20842 40705 20846
rect 39840 20830 39886 20842
rect 39840 20454 39846 20830
rect 39880 20454 39886 20830
rect 39840 20442 39886 20454
rect 39958 20830 40004 20842
rect 39958 20454 39964 20830
rect 39998 20454 40004 20830
rect 39958 20442 40004 20454
rect 40076 20830 40122 20842
rect 40076 20454 40082 20830
rect 40116 20478 40122 20830
rect 40193 20830 40239 20842
rect 40193 20654 40199 20830
rect 40233 20654 40239 20830
rect 40193 20642 40239 20654
rect 40311 20830 40705 20842
rect 41197 21029 41243 21041
rect 41197 20853 41203 21029
rect 41237 20853 41243 21029
rect 41197 20841 41243 20853
rect 41315 21029 41361 21041
rect 41315 20853 41321 21029
rect 41355 20853 41361 21029
rect 41315 20841 41361 20853
rect 41617 21029 41663 21041
rect 40311 20654 40317 20830
rect 40351 20817 40705 20830
rect 40351 20654 40357 20817
rect 40627 20814 40705 20817
rect 40627 20762 40637 20814
rect 40700 20762 40710 20814
rect 40632 20756 40705 20762
rect 40311 20642 40357 20654
rect 40199 20526 40234 20642
rect 41320 20547 41354 20841
rect 41617 20653 41623 21029
rect 41657 20653 41663 21029
rect 41617 20641 41663 20653
rect 41735 21029 41781 21041
rect 41735 20653 41741 21029
rect 41775 20653 41781 21029
rect 41735 20641 41781 20653
rect 41853 21029 41899 21041
rect 41853 20653 41859 21029
rect 41893 20653 41899 21029
rect 41853 20641 41899 20653
rect 41971 21029 42017 21041
rect 41971 20653 41977 21029
rect 42011 20653 42017 21029
rect 41971 20641 42017 20653
rect 42089 21029 42135 21041
rect 42089 20653 42095 21029
rect 42129 20653 42135 21029
rect 42495 21029 42541 21041
rect 42495 20853 42501 21029
rect 42535 20853 42541 21029
rect 42495 20841 42541 20853
rect 42613 21029 42659 21041
rect 42613 20853 42619 21029
rect 42653 20853 42659 21029
rect 42613 20841 42659 20853
rect 43095 21029 43141 21041
rect 43095 20853 43101 21029
rect 43135 20853 43141 21029
rect 43095 20841 43141 20853
rect 43213 21029 43259 21041
rect 43213 20853 43219 21029
rect 43253 20853 43259 21029
rect 43213 20841 43259 20853
rect 43515 21029 43561 21041
rect 42089 20641 42135 20653
rect 41977 20547 42011 20641
rect 42501 20547 42534 20841
rect 40330 20526 40438 20536
rect 40199 20478 40330 20526
rect 40116 20454 40330 20478
rect 40076 20442 40330 20454
rect 39088 20438 39673 20440
rect 40082 20438 40330 20442
rect 39088 20410 39718 20438
rect 39088 20404 39955 20410
rect 39088 20370 39905 20404
rect 39939 20370 39955 20404
rect 39088 20354 39955 20370
rect 40007 20404 40073 20410
rect 40007 20370 40023 20404
rect 40057 20370 40073 20404
rect 40256 20394 40330 20438
rect 41320 20515 42534 20547
rect 43218 20547 43252 20841
rect 43515 20653 43521 21029
rect 43555 20653 43561 21029
rect 43515 20641 43561 20653
rect 43633 21029 43679 21041
rect 43633 20653 43639 21029
rect 43673 20653 43679 21029
rect 43633 20641 43679 20653
rect 43751 21029 43797 21041
rect 43751 20653 43757 21029
rect 43791 20653 43797 21029
rect 43751 20641 43797 20653
rect 43869 21029 43915 21041
rect 43869 20653 43875 21029
rect 43909 20653 43915 21029
rect 43869 20641 43915 20653
rect 43987 21029 44033 21041
rect 43987 20653 43993 21029
rect 44027 20653 44033 21029
rect 44393 21029 44439 21041
rect 44393 20853 44399 21029
rect 44433 20853 44439 21029
rect 44393 20841 44439 20853
rect 44511 21029 44557 21041
rect 44511 20853 44517 21029
rect 44551 20853 44557 21029
rect 44511 20841 44557 20853
rect 43987 20641 44033 20653
rect 43875 20547 43909 20641
rect 44399 20547 44432 20841
rect 43218 20515 44432 20547
rect 41813 20430 41945 20515
rect 43711 20430 43843 20515
rect 40330 20384 40438 20394
rect 39088 20338 39718 20354
rect 39088 20334 39673 20338
rect 39088 20333 39189 20334
rect 39618 20285 39718 20296
rect 39582 20179 39592 20285
rect 39704 20274 39718 20285
rect 40007 20274 40073 20370
rect 41803 20322 41813 20430
rect 41945 20322 41955 20430
rect 43701 20322 43711 20430
rect 43843 20322 43853 20430
rect 44632 20402 44699 21785
rect 45601 21690 45694 23584
rect 45757 23525 46223 23547
rect 46511 23525 46577 23621
rect 48342 23631 48348 23807
rect 48382 23631 48388 23807
rect 48342 23619 48388 23631
rect 48460 23807 48506 23819
rect 48460 23631 48466 23807
rect 48500 23631 48506 23807
rect 48460 23619 48506 23631
rect 48578 23807 48624 23819
rect 48578 23631 48584 23807
rect 48618 23631 48624 23807
rect 48578 23619 48624 23631
rect 48696 23807 48742 23819
rect 48696 23631 48702 23807
rect 48736 23752 48742 23807
rect 48861 23807 48907 23819
rect 48861 23752 48867 23807
rect 48736 23664 48867 23752
rect 48736 23631 48742 23664
rect 48696 23619 48742 23631
rect 48861 23631 48867 23664
rect 48901 23631 48907 23807
rect 48861 23619 48907 23631
rect 48979 23807 49025 23819
rect 48979 23631 48985 23807
rect 49019 23631 49025 23807
rect 48979 23619 49025 23631
rect 49097 23807 49143 23819
rect 49097 23631 49103 23807
rect 49137 23631 49143 23807
rect 49097 23619 49143 23631
rect 49215 23807 49261 23819
rect 49215 23631 49221 23807
rect 49255 23631 49261 23807
rect 49215 23619 49261 23631
rect 48348 23580 48382 23619
rect 48584 23580 48618 23619
rect 48348 23545 48618 23580
rect 48985 23581 49018 23619
rect 49221 23581 49254 23619
rect 48985 23545 49254 23581
rect 45757 23477 46577 23525
rect 48382 23544 48618 23545
rect 45757 23446 46223 23477
rect 48382 23470 48514 23544
rect 45757 23190 45862 23446
rect 48372 23362 48382 23470
rect 48514 23362 48524 23470
rect 45757 23084 45820 23190
rect 45932 23084 45942 23190
rect 46524 23166 46744 23186
rect 45757 23073 45906 23084
rect 45757 21896 45862 23073
rect 46524 23058 46568 23166
rect 46700 23058 46744 23166
rect 46524 23016 46744 23058
rect 49322 23031 49384 24602
rect 49574 24594 49620 24606
rect 49574 24218 49580 24594
rect 49614 24218 49620 24594
rect 49574 24206 49620 24218
rect 49692 24594 49738 24606
rect 49692 24218 49698 24594
rect 49732 24218 49738 24594
rect 49692 24206 49738 24218
rect 49810 24594 49856 24606
rect 49810 24218 49816 24594
rect 49850 24218 49856 24594
rect 49810 24206 49856 24218
rect 49928 24594 49974 24606
rect 49928 24218 49934 24594
rect 49968 24218 49974 24594
rect 49928 24206 49974 24218
rect 50046 24594 50092 24606
rect 50046 24218 50052 24594
rect 50086 24218 50092 24594
rect 50046 24206 50092 24218
rect 50164 24594 50210 24606
rect 50164 24218 50170 24594
rect 50204 24218 50210 24594
rect 50164 24206 50210 24218
rect 50282 24594 50328 24606
rect 50282 24218 50288 24594
rect 50322 24218 50328 24594
rect 52648 24631 53625 24661
rect 52648 24525 52680 24631
rect 52884 24525 52916 24631
rect 53120 24525 53152 24631
rect 53356 24525 53388 24631
rect 53591 24525 53625 24631
rect 52641 24513 52687 24525
rect 52641 24337 52647 24513
rect 52681 24337 52687 24513
rect 52641 24325 52687 24337
rect 52759 24513 52805 24525
rect 52759 24337 52765 24513
rect 52799 24337 52805 24513
rect 52759 24325 52805 24337
rect 52877 24513 52923 24525
rect 52877 24337 52883 24513
rect 52917 24337 52923 24513
rect 52877 24325 52923 24337
rect 52995 24513 53041 24525
rect 52995 24337 53001 24513
rect 53035 24337 53041 24513
rect 52995 24325 53041 24337
rect 53113 24513 53159 24525
rect 53113 24337 53119 24513
rect 53153 24337 53159 24513
rect 53113 24325 53159 24337
rect 53231 24513 53277 24525
rect 53231 24337 53237 24513
rect 53271 24337 53277 24513
rect 53231 24325 53277 24337
rect 53349 24513 53395 24525
rect 53349 24337 53355 24513
rect 53389 24337 53395 24513
rect 53349 24325 53395 24337
rect 53467 24513 53513 24525
rect 53467 24337 53473 24513
rect 53507 24337 53513 24513
rect 53467 24325 53513 24337
rect 53585 24513 53631 24525
rect 53585 24337 53591 24513
rect 53625 24337 53631 24513
rect 53585 24325 53631 24337
rect 53703 24513 53749 24525
rect 53703 24337 53709 24513
rect 53743 24337 53749 24513
rect 53703 24325 53749 24337
rect 50282 24206 50328 24218
rect 52764 24231 52800 24325
rect 53000 24231 53036 24325
rect 53236 24232 53272 24325
rect 53398 24277 53464 24284
rect 53398 24243 53414 24277
rect 53448 24243 53464 24277
rect 53398 24232 53464 24243
rect 53236 24231 53464 24232
rect 49580 24164 49614 24206
rect 49816 24164 49850 24206
rect 49580 24136 49850 24164
rect 49934 24165 49968 24206
rect 50170 24165 50204 24206
rect 49934 24136 50204 24165
rect 49580 24088 49614 24136
rect 49580 24058 49643 24088
rect 49608 23966 49643 24058
rect 50115 24028 50215 24049
rect 50115 23974 50129 24028
rect 50194 23974 50215 24028
rect 50115 23969 50215 23974
rect 50288 24023 50322 24206
rect 52764 24202 53464 24231
rect 52764 24201 53346 24202
rect 52884 24088 52918 24201
rect 53280 24160 53346 24201
rect 53280 24126 53296 24160
rect 53330 24126 53346 24160
rect 53280 24119 53346 24126
rect 53708 24120 53743 24325
rect 53915 24120 53982 24710
rect 55674 24687 55715 24719
rect 55961 24715 55971 24781
rect 56027 24715 56037 24781
rect 56707 24757 56717 24865
rect 56849 24802 56859 24865
rect 59602 24815 59822 24835
rect 56849 24791 56861 24802
rect 56849 24757 56862 24791
rect 56717 24719 56862 24757
rect 56821 24691 56862 24719
rect 55090 24659 55360 24687
rect 54831 24593 54841 24659
rect 54907 24593 54917 24659
rect 55090 24597 55124 24659
rect 55326 24597 55360 24659
rect 55444 24659 55715 24687
rect 56232 24663 56502 24691
rect 55444 24597 55478 24659
rect 55680 24597 55715 24659
rect 55856 24647 56027 24663
rect 55856 24613 55987 24647
rect 56021 24613 56027 24647
rect 55856 24597 56027 24613
rect 56232 24601 56266 24663
rect 56468 24601 56502 24663
rect 56586 24663 56862 24691
rect 59602 24707 59646 24815
rect 59778 24707 59822 24815
rect 61399 24773 61455 24781
rect 59602 24665 59822 24707
rect 60473 24765 61455 24773
rect 60473 24731 61415 24765
rect 61449 24731 61455 24765
rect 62118 24761 62128 24869
rect 62260 24806 62270 24869
rect 62260 24795 62272 24806
rect 62260 24761 62273 24795
rect 62529 24785 62585 24787
rect 60473 24715 61455 24731
rect 62128 24723 62273 24761
rect 60473 24714 61452 24715
rect 56586 24601 56620 24663
rect 56822 24601 56862 24663
rect 54966 24585 55012 24597
rect 54966 24209 54972 24585
rect 55006 24209 55012 24585
rect 54966 24197 55012 24209
rect 55084 24585 55130 24597
rect 55084 24209 55090 24585
rect 55124 24209 55130 24585
rect 55084 24197 55130 24209
rect 55202 24585 55248 24597
rect 55202 24209 55208 24585
rect 55242 24209 55248 24585
rect 55202 24197 55248 24209
rect 55320 24585 55366 24597
rect 55320 24209 55326 24585
rect 55360 24209 55366 24585
rect 55320 24197 55366 24209
rect 55438 24585 55484 24597
rect 55438 24209 55444 24585
rect 55478 24209 55484 24585
rect 55438 24197 55484 24209
rect 55556 24585 55602 24597
rect 55556 24209 55562 24585
rect 55596 24209 55602 24585
rect 55556 24197 55602 24209
rect 55674 24585 55720 24597
rect 55674 24209 55680 24585
rect 55714 24209 55720 24585
rect 55674 24197 55720 24209
rect 53708 24092 53982 24120
rect 53354 24088 53982 24092
rect 52878 24076 52924 24088
rect 51297 24037 51396 24041
rect 50288 23969 50397 24023
rect 49608 23930 49835 23966
rect 49608 23823 49643 23930
rect 49769 23896 49835 23930
rect 49769 23862 49785 23896
rect 49819 23862 49835 23896
rect 50116 23954 50213 23969
rect 50116 23887 50173 23954
rect 49769 23856 49835 23862
rect 50010 23851 50279 23887
rect 50010 23823 50043 23851
rect 50246 23823 50279 23851
rect 50363 23823 50397 23969
rect 51214 23962 51224 24037
rect 51292 23962 51396 24037
rect 51241 23961 51396 23962
rect 49484 23811 49530 23823
rect 49484 23635 49490 23811
rect 49524 23635 49530 23811
rect 49484 23623 49530 23635
rect 49602 23811 49648 23823
rect 49602 23635 49608 23811
rect 49642 23635 49648 23811
rect 49602 23623 49648 23635
rect 49720 23811 49766 23823
rect 49720 23635 49726 23811
rect 49760 23635 49766 23811
rect 49720 23623 49766 23635
rect 49838 23811 49884 23823
rect 49838 23635 49844 23811
rect 49878 23756 49884 23811
rect 50003 23811 50049 23823
rect 50003 23756 50009 23811
rect 49878 23668 50009 23756
rect 49878 23635 49884 23668
rect 49838 23623 49884 23635
rect 50003 23635 50009 23668
rect 50043 23635 50049 23811
rect 50003 23623 50049 23635
rect 50121 23811 50167 23823
rect 50121 23635 50127 23811
rect 50161 23635 50167 23811
rect 50121 23623 50167 23635
rect 50239 23811 50285 23823
rect 50239 23635 50245 23811
rect 50279 23635 50285 23811
rect 50239 23623 50285 23635
rect 50357 23811 50403 23823
rect 50357 23635 50363 23811
rect 50397 23635 50403 23811
rect 50357 23623 50403 23635
rect 49490 23584 49524 23623
rect 49726 23584 49760 23623
rect 49490 23548 49760 23584
rect 50127 23585 50160 23623
rect 50363 23585 50396 23623
rect 50127 23549 50396 23585
rect 49490 23547 49656 23548
rect 49524 23468 49656 23547
rect 49514 23360 49524 23468
rect 49656 23360 49666 23468
rect 46128 22986 47105 23016
rect 49322 23014 49385 23031
rect 49247 23010 49385 23014
rect 46128 22880 46160 22986
rect 46364 22880 46396 22986
rect 46600 22880 46632 22986
rect 46836 22880 46868 22986
rect 47071 22880 47105 22986
rect 47415 22976 49385 23010
rect 47413 22947 49385 22976
rect 47413 22931 47459 22947
rect 49247 22945 49385 22947
rect 46121 22868 46167 22880
rect 46121 22692 46127 22868
rect 46161 22692 46167 22868
rect 46121 22680 46167 22692
rect 46239 22868 46285 22880
rect 46239 22692 46245 22868
rect 46279 22692 46285 22868
rect 46239 22680 46285 22692
rect 46357 22868 46403 22880
rect 46357 22692 46363 22868
rect 46397 22692 46403 22868
rect 46357 22680 46403 22692
rect 46475 22868 46521 22880
rect 46475 22692 46481 22868
rect 46515 22692 46521 22868
rect 46475 22680 46521 22692
rect 46593 22868 46639 22880
rect 46593 22692 46599 22868
rect 46633 22692 46639 22868
rect 46593 22680 46639 22692
rect 46711 22868 46757 22880
rect 46711 22692 46717 22868
rect 46751 22692 46757 22868
rect 46711 22680 46757 22692
rect 46829 22868 46875 22880
rect 46829 22692 46835 22868
rect 46869 22692 46875 22868
rect 46829 22680 46875 22692
rect 46947 22868 46993 22880
rect 46947 22692 46953 22868
rect 46987 22692 46993 22868
rect 46947 22680 46993 22692
rect 47065 22868 47111 22880
rect 47065 22692 47071 22868
rect 47105 22692 47111 22868
rect 47065 22680 47111 22692
rect 47183 22868 47229 22880
rect 47183 22692 47189 22868
rect 47223 22692 47229 22868
rect 47183 22680 47229 22692
rect 46244 22586 46280 22680
rect 46480 22586 46516 22680
rect 46716 22587 46752 22680
rect 46878 22632 46944 22639
rect 46878 22598 46894 22632
rect 46928 22598 46944 22632
rect 46878 22587 46944 22598
rect 46716 22586 46944 22587
rect 46244 22557 46944 22586
rect 46244 22556 46826 22557
rect 46364 22443 46398 22556
rect 46760 22515 46826 22556
rect 46760 22481 46776 22515
rect 46810 22481 46826 22515
rect 46760 22474 46826 22481
rect 47188 22462 47223 22680
rect 47412 22479 47459 22931
rect 48371 22715 48381 22823
rect 48513 22715 48523 22823
rect 50269 22715 50279 22823
rect 50411 22715 50421 22823
rect 48381 22675 48513 22715
rect 50279 22675 50411 22715
rect 48380 22609 48513 22675
rect 50278 22609 50411 22675
rect 47709 22566 49182 22609
rect 47412 22463 47458 22479
rect 47377 22462 47458 22463
rect 47188 22447 47458 22462
rect 46834 22443 47458 22447
rect 46358 22431 46404 22443
rect 46093 21953 46103 22071
rect 46221 22039 46231 22071
rect 46358 22055 46364 22431
rect 46398 22055 46404 22431
rect 46358 22043 46404 22055
rect 46476 22431 46522 22443
rect 46476 22055 46482 22431
rect 46516 22055 46522 22431
rect 46476 22043 46522 22055
rect 46594 22431 46640 22443
rect 46594 22055 46600 22431
rect 46634 22079 46640 22431
rect 46711 22431 46757 22443
rect 46711 22255 46717 22431
rect 46751 22255 46757 22431
rect 46711 22243 46757 22255
rect 46829 22431 47458 22443
rect 46829 22255 46835 22431
rect 46869 22419 47458 22431
rect 46869 22418 47111 22419
rect 46869 22255 46875 22418
rect 47377 22417 47458 22419
rect 47709 22263 47743 22566
rect 48075 22463 48109 22566
rect 48311 22463 48345 22566
rect 48547 22463 48581 22566
rect 48783 22463 48817 22566
rect 48069 22451 48115 22463
rect 46829 22243 46875 22255
rect 47585 22251 47631 22263
rect 46717 22127 46752 22243
rect 46848 22127 46956 22137
rect 46717 22079 46848 22127
rect 46634 22055 46848 22079
rect 46594 22043 46848 22055
rect 46600 22039 46848 22043
rect 46221 22011 46236 22039
rect 46221 22005 46473 22011
rect 46221 21971 46423 22005
rect 46457 21971 46473 22005
rect 46221 21955 46473 21971
rect 46525 22005 46591 22011
rect 46525 21971 46541 22005
rect 46575 21971 46591 22005
rect 46774 21995 46848 22039
rect 47585 22075 47591 22251
rect 47625 22075 47631 22251
rect 47585 22063 47631 22075
rect 47703 22251 47749 22263
rect 47703 22075 47709 22251
rect 47743 22075 47749 22251
rect 47703 22063 47749 22075
rect 47821 22251 47867 22263
rect 47821 22075 47827 22251
rect 47861 22075 47867 22251
rect 47821 22063 47867 22075
rect 47939 22251 47985 22263
rect 48069 22251 48075 22451
rect 47939 22075 47945 22251
rect 47979 22075 48075 22251
rect 48109 22075 48115 22451
rect 47939 22063 47985 22075
rect 48069 22063 48115 22075
rect 48187 22451 48233 22463
rect 48187 22075 48193 22451
rect 48227 22075 48233 22451
rect 48187 22063 48233 22075
rect 48305 22451 48351 22463
rect 48305 22075 48311 22451
rect 48345 22075 48351 22451
rect 48305 22063 48351 22075
rect 48423 22451 48469 22463
rect 48423 22075 48429 22451
rect 48463 22075 48469 22451
rect 48423 22063 48469 22075
rect 48541 22451 48587 22463
rect 48541 22075 48547 22451
rect 48581 22075 48587 22451
rect 48541 22063 48587 22075
rect 48659 22451 48705 22463
rect 48659 22075 48665 22451
rect 48699 22075 48705 22451
rect 48659 22063 48705 22075
rect 48777 22451 48823 22463
rect 48777 22075 48783 22451
rect 48817 22251 48823 22451
rect 49148 22263 49182 22566
rect 49607 22566 51080 22609
rect 49607 22263 49641 22566
rect 49973 22463 50007 22566
rect 50209 22463 50243 22566
rect 50445 22463 50479 22566
rect 50681 22463 50715 22566
rect 49967 22451 50013 22463
rect 48906 22251 48952 22263
rect 48817 22075 48912 22251
rect 48946 22075 48952 22251
rect 48777 22063 48823 22075
rect 48906 22063 48952 22075
rect 49024 22251 49070 22263
rect 49024 22075 49030 22251
rect 49064 22075 49070 22251
rect 49024 22063 49070 22075
rect 49142 22251 49188 22263
rect 49142 22075 49148 22251
rect 49182 22075 49188 22251
rect 49142 22063 49188 22075
rect 49260 22251 49306 22263
rect 49260 22075 49266 22251
rect 49300 22075 49306 22251
rect 49260 22063 49306 22075
rect 49483 22251 49529 22263
rect 49483 22075 49489 22251
rect 49523 22075 49529 22251
rect 49483 22063 49529 22075
rect 49601 22251 49647 22263
rect 49601 22075 49607 22251
rect 49641 22075 49647 22251
rect 49601 22063 49647 22075
rect 49719 22251 49765 22263
rect 49719 22075 49725 22251
rect 49759 22075 49765 22251
rect 49719 22063 49765 22075
rect 49837 22251 49883 22263
rect 49967 22251 49973 22451
rect 49837 22075 49843 22251
rect 49877 22075 49973 22251
rect 50007 22075 50013 22451
rect 49837 22063 49883 22075
rect 49967 22063 50013 22075
rect 50085 22451 50131 22463
rect 50085 22075 50091 22451
rect 50125 22075 50131 22451
rect 50085 22063 50131 22075
rect 50203 22451 50249 22463
rect 50203 22075 50209 22451
rect 50243 22075 50249 22451
rect 50203 22063 50249 22075
rect 50321 22451 50367 22463
rect 50321 22075 50327 22451
rect 50361 22075 50367 22451
rect 50321 22063 50367 22075
rect 50439 22451 50485 22463
rect 50439 22075 50445 22451
rect 50479 22075 50485 22451
rect 50439 22063 50485 22075
rect 50557 22451 50603 22463
rect 50557 22075 50563 22451
rect 50597 22075 50603 22451
rect 50557 22063 50603 22075
rect 50675 22451 50721 22463
rect 50675 22075 50681 22451
rect 50715 22251 50721 22451
rect 51046 22263 51080 22566
rect 50804 22251 50850 22263
rect 50715 22075 50810 22251
rect 50844 22075 50850 22251
rect 50675 22063 50721 22075
rect 50804 22063 50850 22075
rect 50922 22251 50968 22263
rect 50922 22075 50928 22251
rect 50962 22075 50968 22251
rect 50922 22063 50968 22075
rect 51040 22251 51086 22263
rect 51040 22075 51046 22251
rect 51080 22075 51086 22251
rect 51040 22063 51086 22075
rect 51158 22251 51204 22263
rect 51158 22075 51164 22251
rect 51198 22075 51204 22251
rect 51297 22215 51396 23961
rect 51706 23758 51995 23777
rect 51706 23601 51727 23758
rect 51960 23683 51995 23758
rect 52878 23700 52884 24076
rect 52918 23700 52924 24076
rect 52878 23688 52924 23700
rect 52996 24076 53042 24088
rect 52996 23700 53002 24076
rect 53036 23700 53042 24076
rect 52996 23688 53042 23700
rect 53114 24076 53160 24088
rect 53114 23700 53120 24076
rect 53154 23724 53160 24076
rect 53231 24076 53277 24088
rect 53231 23900 53237 24076
rect 53271 23900 53277 24076
rect 53231 23888 53277 23900
rect 53349 24076 53982 24088
rect 53349 23900 53355 24076
rect 53389 24063 53982 24076
rect 54972 24155 55006 24197
rect 55208 24155 55242 24197
rect 54972 24127 55242 24155
rect 55326 24156 55360 24197
rect 55562 24156 55596 24197
rect 55326 24127 55596 24156
rect 54972 24079 55006 24127
rect 53389 23900 53395 24063
rect 54972 24049 55035 24079
rect 53349 23888 53395 23900
rect 55000 23957 55035 24049
rect 55000 23921 55227 23957
rect 55497 23946 55507 24043
rect 55606 23946 55616 24043
rect 55680 24014 55714 24197
rect 55680 23960 55789 24014
rect 53237 23772 53272 23888
rect 55000 23814 55035 23921
rect 55161 23887 55227 23921
rect 55161 23853 55177 23887
rect 55211 23853 55227 23887
rect 55508 23945 55605 23946
rect 55508 23878 55565 23945
rect 55161 23847 55227 23853
rect 55402 23842 55671 23878
rect 55402 23814 55435 23842
rect 55638 23814 55671 23842
rect 55755 23814 55789 23960
rect 54876 23802 54922 23814
rect 53368 23772 53476 23782
rect 53237 23724 53368 23772
rect 53154 23700 53368 23724
rect 53114 23688 53368 23700
rect 53120 23684 53368 23688
rect 51960 23656 52756 23683
rect 51960 23650 52993 23656
rect 51960 23616 52943 23650
rect 52977 23616 52993 23650
rect 51960 23601 52993 23616
rect 51706 23600 52993 23601
rect 53045 23650 53111 23656
rect 53045 23616 53061 23650
rect 53095 23616 53111 23650
rect 53294 23640 53368 23684
rect 53368 23630 53476 23640
rect 51706 23584 52756 23600
rect 51706 23583 52693 23584
rect 51706 23579 52228 23583
rect 51706 23578 51995 23579
rect 51723 22215 52011 22218
rect 51297 22105 52011 22215
rect 51158 22063 51204 22075
rect 46848 21985 46956 21995
rect 47591 22029 47625 22063
rect 48193 22029 48227 22063
rect 48429 22029 48463 22063
rect 47591 21994 47750 22029
rect 48193 21994 48463 22029
rect 49030 22029 49064 22063
rect 49266 22029 49300 22063
rect 49030 21994 49300 22029
rect 49489 22029 49523 22063
rect 50091 22029 50125 22063
rect 50327 22029 50361 22063
rect 49489 21994 49648 22029
rect 50091 21994 50361 22029
rect 50928 22029 50962 22063
rect 51164 22029 51198 22063
rect 50928 21994 51198 22029
rect 51723 22056 52011 22105
rect 46221 21953 46236 21955
rect 46136 21939 46236 21953
rect 46136 21896 46236 21897
rect 45757 21875 46236 21896
rect 46525 21875 46591 21971
rect 45757 21827 46591 21875
rect 45757 21798 46236 21827
rect 45757 21796 45862 21798
rect 46136 21797 46236 21798
rect 45590 21611 45600 21690
rect 45693 21611 45703 21690
rect 45601 20437 45694 21611
rect 46519 21562 46739 21582
rect 46519 21454 46563 21562
rect 46695 21454 46739 21562
rect 46519 21412 46739 21454
rect 46123 21382 47100 21412
rect 46123 21276 46155 21382
rect 46359 21276 46391 21382
rect 46595 21276 46627 21382
rect 46831 21276 46863 21382
rect 47066 21276 47100 21382
rect 46116 21264 46162 21276
rect 46116 21088 46122 21264
rect 46156 21088 46162 21264
rect 46116 21076 46162 21088
rect 46234 21264 46280 21276
rect 46234 21088 46240 21264
rect 46274 21088 46280 21264
rect 46234 21076 46280 21088
rect 46352 21264 46398 21276
rect 46352 21088 46358 21264
rect 46392 21088 46398 21264
rect 46352 21076 46398 21088
rect 46470 21264 46516 21276
rect 46470 21088 46476 21264
rect 46510 21088 46516 21264
rect 46470 21076 46516 21088
rect 46588 21264 46634 21276
rect 46588 21088 46594 21264
rect 46628 21088 46634 21264
rect 46588 21076 46634 21088
rect 46706 21264 46752 21276
rect 46706 21088 46712 21264
rect 46746 21088 46752 21264
rect 46706 21076 46752 21088
rect 46824 21264 46870 21276
rect 46824 21088 46830 21264
rect 46864 21088 46870 21264
rect 46824 21076 46870 21088
rect 46942 21264 46988 21276
rect 46942 21088 46948 21264
rect 46982 21088 46988 21264
rect 46942 21076 46988 21088
rect 47060 21264 47106 21276
rect 47060 21088 47066 21264
rect 47100 21088 47106 21264
rect 47060 21076 47106 21088
rect 47178 21264 47224 21276
rect 47178 21088 47184 21264
rect 47218 21088 47224 21264
rect 47178 21076 47224 21088
rect 47716 21210 47750 21994
rect 48429 21932 48463 21994
rect 48018 21894 48760 21932
rect 48018 21770 48052 21894
rect 48254 21770 48288 21894
rect 48490 21770 48524 21894
rect 48726 21770 48760 21894
rect 49016 21787 49026 21853
rect 49089 21787 49099 21853
rect 48012 21758 48058 21770
rect 48012 21382 48018 21758
rect 48052 21382 48058 21758
rect 48012 21370 48058 21382
rect 48130 21758 48176 21770
rect 48130 21382 48136 21758
rect 48170 21382 48176 21758
rect 48130 21370 48176 21382
rect 48248 21758 48294 21770
rect 48248 21382 48254 21758
rect 48288 21382 48294 21758
rect 48248 21370 48294 21382
rect 48366 21758 48412 21770
rect 48366 21382 48372 21758
rect 48406 21382 48412 21758
rect 48366 21370 48412 21382
rect 48484 21758 48530 21770
rect 48484 21382 48490 21758
rect 48524 21382 48530 21758
rect 48484 21370 48530 21382
rect 48602 21758 48648 21770
rect 48602 21382 48608 21758
rect 48642 21382 48648 21758
rect 48602 21370 48648 21382
rect 48720 21758 48766 21770
rect 48720 21382 48726 21758
rect 48760 21382 48766 21758
rect 48720 21370 48766 21382
rect 49132 21211 49166 21994
rect 48859 21210 49166 21211
rect 47716 21205 48032 21210
rect 48746 21205 49166 21210
rect 47716 21194 48099 21205
rect 47716 21167 48048 21194
rect 46239 20982 46275 21076
rect 46475 20982 46511 21076
rect 46711 20983 46747 21076
rect 46873 21028 46939 21035
rect 46873 20994 46889 21028
rect 46923 20994 46939 21028
rect 46873 20983 46939 20994
rect 46711 20982 46939 20983
rect 46239 20953 46939 20982
rect 46239 20952 46821 20953
rect 46359 20839 46393 20952
rect 46755 20911 46821 20952
rect 46755 20877 46771 20911
rect 46805 20877 46821 20911
rect 46755 20870 46821 20877
rect 47183 20843 47218 21076
rect 47716 21038 47750 21167
rect 48032 21160 48048 21167
rect 48082 21160 48099 21194
rect 48032 21154 48099 21160
rect 48679 21194 49166 21205
rect 48679 21160 48696 21194
rect 48730 21167 49166 21194
rect 48730 21160 48746 21167
rect 48859 21166 49166 21167
rect 48679 21154 48746 21160
rect 47857 21127 47913 21139
rect 47857 21093 47863 21127
rect 47897 21126 47913 21127
rect 48970 21126 49026 21138
rect 47897 21110 48364 21126
rect 47897 21093 48314 21110
rect 47857 21077 48314 21093
rect 48298 21076 48314 21077
rect 48348 21076 48364 21110
rect 48298 21069 48364 21076
rect 48416 21111 48986 21126
rect 48416 21077 48432 21111
rect 48466 21092 48986 21111
rect 49020 21092 49026 21126
rect 48466 21077 49026 21092
rect 48416 21067 48483 21077
rect 48970 21076 49026 21077
rect 49132 21038 49166 21166
rect 49614 21210 49648 21994
rect 50327 21932 50361 21994
rect 49916 21894 50658 21932
rect 49916 21770 49950 21894
rect 50152 21770 50186 21894
rect 50388 21770 50422 21894
rect 50624 21770 50658 21894
rect 49910 21758 49956 21770
rect 49910 21382 49916 21758
rect 49950 21382 49956 21758
rect 49910 21370 49956 21382
rect 50028 21758 50074 21770
rect 50028 21382 50034 21758
rect 50068 21382 50074 21758
rect 50028 21370 50074 21382
rect 50146 21758 50192 21770
rect 50146 21382 50152 21758
rect 50186 21382 50192 21758
rect 50146 21370 50192 21382
rect 50264 21758 50310 21770
rect 50264 21382 50270 21758
rect 50304 21382 50310 21758
rect 50264 21370 50310 21382
rect 50382 21758 50428 21770
rect 50382 21382 50388 21758
rect 50422 21382 50428 21758
rect 50382 21370 50428 21382
rect 50500 21758 50546 21770
rect 50500 21382 50506 21758
rect 50540 21382 50546 21758
rect 50500 21370 50546 21382
rect 50618 21758 50664 21770
rect 50618 21382 50624 21758
rect 50658 21382 50664 21758
rect 50618 21370 50664 21382
rect 51030 21211 51064 21994
rect 51723 21950 51859 22056
rect 51971 22054 52011 22056
rect 51977 22043 52011 22054
rect 51723 21948 51865 21950
rect 51977 21948 52012 22043
rect 51723 21939 52012 21948
rect 51723 21938 52011 21939
rect 51723 21937 51979 21938
rect 50642 21210 50711 21211
rect 50757 21210 51064 21211
rect 49614 21205 49930 21210
rect 50642 21206 51064 21210
rect 49614 21194 49997 21205
rect 49614 21167 49946 21194
rect 49614 21038 49648 21167
rect 49930 21160 49946 21167
rect 49980 21160 49997 21194
rect 49930 21154 49997 21160
rect 50575 21195 51064 21206
rect 50575 21161 50592 21195
rect 50626 21167 51064 21195
rect 50626 21161 50642 21167
rect 50757 21166 51064 21167
rect 50575 21155 50642 21161
rect 49755 21127 49811 21139
rect 49755 21093 49761 21127
rect 49795 21126 49811 21127
rect 50868 21126 50924 21138
rect 49795 21110 50262 21126
rect 49795 21093 50212 21110
rect 49755 21077 50212 21093
rect 50196 21076 50212 21077
rect 50246 21076 50262 21110
rect 50196 21069 50262 21076
rect 50314 21111 50884 21126
rect 50314 21077 50330 21111
rect 50364 21092 50884 21111
rect 50918 21092 50924 21126
rect 50364 21077 50924 21092
rect 50314 21067 50381 21077
rect 50868 21076 50924 21077
rect 51030 21038 51064 21166
rect 51145 21816 51212 21840
rect 51145 21782 51162 21816
rect 51196 21782 51212 21816
rect 46829 20839 47218 20843
rect 46353 20827 46399 20839
rect 46353 20451 46359 20827
rect 46393 20451 46399 20827
rect 46353 20439 46399 20451
rect 46471 20827 46517 20839
rect 46471 20451 46477 20827
rect 46511 20451 46517 20827
rect 46471 20439 46517 20451
rect 46589 20827 46635 20839
rect 46589 20451 46595 20827
rect 46629 20475 46635 20827
rect 46706 20827 46752 20839
rect 46706 20651 46712 20827
rect 46746 20651 46752 20827
rect 46706 20639 46752 20651
rect 46824 20827 47218 20839
rect 47710 21026 47756 21038
rect 47710 20850 47716 21026
rect 47750 20850 47756 21026
rect 47710 20838 47756 20850
rect 47828 21026 47874 21038
rect 47828 20850 47834 21026
rect 47868 20850 47874 21026
rect 47828 20838 47874 20850
rect 48130 21026 48176 21038
rect 46824 20651 46830 20827
rect 46864 20814 47218 20827
rect 46864 20651 46870 20814
rect 47140 20811 47218 20814
rect 47140 20759 47150 20811
rect 47213 20759 47223 20811
rect 47145 20753 47218 20759
rect 46824 20639 46870 20651
rect 46712 20523 46747 20639
rect 47833 20544 47867 20838
rect 48130 20650 48136 21026
rect 48170 20650 48176 21026
rect 48130 20638 48176 20650
rect 48248 21026 48294 21038
rect 48248 20650 48254 21026
rect 48288 20650 48294 21026
rect 48248 20638 48294 20650
rect 48366 21026 48412 21038
rect 48366 20650 48372 21026
rect 48406 20650 48412 21026
rect 48366 20638 48412 20650
rect 48484 21026 48530 21038
rect 48484 20650 48490 21026
rect 48524 20650 48530 21026
rect 48484 20638 48530 20650
rect 48602 21026 48648 21038
rect 48602 20650 48608 21026
rect 48642 20650 48648 21026
rect 49008 21026 49054 21038
rect 49008 20850 49014 21026
rect 49048 20850 49054 21026
rect 49008 20838 49054 20850
rect 49126 21026 49172 21038
rect 49126 20850 49132 21026
rect 49166 20850 49172 21026
rect 49126 20838 49172 20850
rect 49608 21026 49654 21038
rect 49608 20850 49614 21026
rect 49648 20850 49654 21026
rect 49608 20838 49654 20850
rect 49726 21026 49772 21038
rect 49726 20850 49732 21026
rect 49766 20850 49772 21026
rect 49726 20838 49772 20850
rect 50028 21026 50074 21038
rect 48602 20638 48648 20650
rect 48490 20544 48524 20638
rect 49014 20544 49047 20838
rect 46843 20523 46951 20533
rect 46712 20475 46843 20523
rect 46629 20451 46843 20475
rect 46589 20439 46843 20451
rect 45601 20435 46186 20437
rect 46595 20435 46843 20439
rect 45601 20407 46231 20435
rect 39704 20226 40073 20274
rect 39704 20196 39718 20226
rect 39704 20179 39714 20196
rect 40006 20123 40072 20226
rect 44632 20123 44698 20402
rect 45601 20401 46468 20407
rect 45601 20367 46418 20401
rect 46452 20367 46468 20401
rect 45601 20351 46468 20367
rect 46520 20401 46586 20407
rect 46520 20367 46536 20401
rect 46570 20367 46586 20401
rect 46769 20391 46843 20435
rect 47833 20512 49047 20544
rect 49731 20544 49765 20838
rect 50028 20650 50034 21026
rect 50068 20650 50074 21026
rect 50028 20638 50074 20650
rect 50146 21026 50192 21038
rect 50146 20650 50152 21026
rect 50186 20650 50192 21026
rect 50146 20638 50192 20650
rect 50264 21026 50310 21038
rect 50264 20650 50270 21026
rect 50304 20650 50310 21026
rect 50264 20638 50310 20650
rect 50382 21026 50428 21038
rect 50382 20650 50388 21026
rect 50422 20650 50428 21026
rect 50382 20638 50428 20650
rect 50500 21026 50546 21038
rect 50500 20650 50506 21026
rect 50540 20650 50546 21026
rect 50906 21026 50952 21038
rect 50906 20850 50912 21026
rect 50946 20850 50952 21026
rect 50906 20838 50952 20850
rect 51024 21026 51070 21038
rect 51024 20850 51030 21026
rect 51064 20850 51070 21026
rect 51024 20838 51070 20850
rect 50500 20638 50546 20650
rect 50388 20544 50422 20638
rect 50912 20544 50945 20838
rect 49731 20512 50945 20544
rect 48326 20427 48458 20512
rect 50224 20427 50356 20512
rect 46843 20381 46951 20391
rect 45601 20335 46231 20351
rect 45601 20331 46186 20335
rect 45601 20330 45702 20331
rect 46131 20282 46231 20293
rect 46095 20176 46105 20282
rect 46217 20271 46231 20282
rect 46520 20271 46586 20367
rect 48316 20319 48326 20427
rect 48458 20319 48468 20427
rect 50214 20319 50224 20427
rect 50356 20319 50366 20427
rect 51145 20399 51212 21782
rect 52135 21685 52228 23579
rect 52291 23520 52757 23542
rect 53045 23520 53111 23616
rect 54876 23626 54882 23802
rect 54916 23626 54922 23802
rect 54876 23614 54922 23626
rect 54994 23802 55040 23814
rect 54994 23626 55000 23802
rect 55034 23626 55040 23802
rect 54994 23614 55040 23626
rect 55112 23802 55158 23814
rect 55112 23626 55118 23802
rect 55152 23626 55158 23802
rect 55112 23614 55158 23626
rect 55230 23802 55276 23814
rect 55230 23626 55236 23802
rect 55270 23747 55276 23802
rect 55395 23802 55441 23814
rect 55395 23747 55401 23802
rect 55270 23659 55401 23747
rect 55270 23626 55276 23659
rect 55230 23614 55276 23626
rect 55395 23626 55401 23659
rect 55435 23626 55441 23802
rect 55395 23614 55441 23626
rect 55513 23802 55559 23814
rect 55513 23626 55519 23802
rect 55553 23626 55559 23802
rect 55513 23614 55559 23626
rect 55631 23802 55677 23814
rect 55631 23626 55637 23802
rect 55671 23626 55677 23802
rect 55631 23614 55677 23626
rect 55749 23802 55795 23814
rect 55749 23626 55755 23802
rect 55789 23626 55795 23802
rect 55749 23614 55795 23626
rect 54882 23575 54916 23614
rect 55118 23575 55152 23614
rect 54882 23540 55152 23575
rect 55519 23576 55552 23614
rect 55755 23576 55788 23614
rect 55519 23540 55788 23576
rect 52291 23472 53111 23520
rect 54916 23539 55152 23540
rect 52291 23441 52757 23472
rect 54916 23465 55048 23539
rect 52291 23185 52396 23441
rect 54906 23357 54916 23465
rect 55048 23357 55058 23465
rect 52291 23079 52354 23185
rect 52466 23079 52476 23185
rect 53058 23161 53278 23181
rect 52291 23068 52440 23079
rect 52291 21891 52396 23068
rect 53058 23053 53102 23161
rect 53234 23053 53278 23161
rect 53058 23011 53278 23053
rect 55856 23026 55918 24597
rect 56108 24589 56154 24601
rect 56108 24213 56114 24589
rect 56148 24213 56154 24589
rect 56108 24201 56154 24213
rect 56226 24589 56272 24601
rect 56226 24213 56232 24589
rect 56266 24213 56272 24589
rect 56226 24201 56272 24213
rect 56344 24589 56390 24601
rect 56344 24213 56350 24589
rect 56384 24213 56390 24589
rect 56344 24201 56390 24213
rect 56462 24589 56508 24601
rect 56462 24213 56468 24589
rect 56502 24213 56508 24589
rect 56462 24201 56508 24213
rect 56580 24589 56626 24601
rect 56580 24213 56586 24589
rect 56620 24213 56626 24589
rect 56580 24201 56626 24213
rect 56698 24589 56744 24601
rect 56698 24213 56704 24589
rect 56738 24213 56744 24589
rect 56698 24201 56744 24213
rect 56816 24589 56862 24601
rect 56816 24213 56822 24589
rect 56856 24213 56862 24589
rect 59206 24635 60183 24665
rect 59206 24529 59238 24635
rect 59442 24529 59474 24635
rect 59678 24529 59710 24635
rect 59914 24529 59946 24635
rect 60149 24529 60183 24635
rect 59199 24517 59245 24529
rect 59199 24341 59205 24517
rect 59239 24341 59245 24517
rect 59199 24329 59245 24341
rect 59317 24517 59363 24529
rect 59317 24341 59323 24517
rect 59357 24341 59363 24517
rect 59317 24329 59363 24341
rect 59435 24517 59481 24529
rect 59435 24341 59441 24517
rect 59475 24341 59481 24517
rect 59435 24329 59481 24341
rect 59553 24517 59599 24529
rect 59553 24341 59559 24517
rect 59593 24341 59599 24517
rect 59553 24329 59599 24341
rect 59671 24517 59717 24529
rect 59671 24341 59677 24517
rect 59711 24341 59717 24517
rect 59671 24329 59717 24341
rect 59789 24517 59835 24529
rect 59789 24341 59795 24517
rect 59829 24341 59835 24517
rect 59789 24329 59835 24341
rect 59907 24517 59953 24529
rect 59907 24341 59913 24517
rect 59947 24341 59953 24517
rect 59907 24329 59953 24341
rect 60025 24517 60071 24529
rect 60025 24341 60031 24517
rect 60065 24341 60071 24517
rect 60025 24329 60071 24341
rect 60143 24517 60189 24529
rect 60143 24341 60149 24517
rect 60183 24341 60189 24517
rect 60143 24329 60189 24341
rect 60261 24517 60307 24529
rect 60261 24341 60267 24517
rect 60301 24341 60307 24517
rect 60261 24329 60307 24341
rect 56816 24201 56862 24213
rect 59322 24235 59358 24329
rect 59558 24235 59594 24329
rect 59794 24236 59830 24329
rect 59956 24281 60022 24288
rect 59956 24247 59972 24281
rect 60006 24247 60022 24281
rect 59956 24236 60022 24247
rect 59794 24235 60022 24236
rect 59322 24206 60022 24235
rect 59322 24205 59904 24206
rect 56114 24159 56148 24201
rect 56350 24159 56384 24201
rect 56114 24131 56384 24159
rect 56468 24160 56502 24201
rect 56704 24160 56738 24201
rect 56468 24131 56738 24160
rect 56114 24083 56148 24131
rect 56114 24053 56177 24083
rect 56142 23961 56177 24053
rect 56649 24023 56749 24044
rect 56649 23969 56663 24023
rect 56728 23969 56749 24023
rect 56649 23964 56749 23969
rect 56822 24018 56856 24201
rect 59442 24092 59476 24205
rect 59838 24164 59904 24205
rect 59838 24130 59854 24164
rect 59888 24130 59904 24164
rect 59838 24123 59904 24130
rect 60266 24124 60301 24329
rect 60473 24124 60540 24714
rect 62232 24691 62273 24723
rect 62519 24719 62529 24785
rect 62585 24719 62595 24785
rect 63265 24761 63275 24869
rect 63407 24806 63417 24869
rect 63407 24795 63419 24806
rect 63407 24761 63420 24795
rect 63275 24723 63420 24761
rect 63379 24695 63420 24723
rect 61648 24663 61918 24691
rect 61389 24597 61399 24663
rect 61465 24597 61475 24663
rect 61648 24601 61682 24663
rect 61884 24601 61918 24663
rect 62002 24663 62273 24691
rect 62790 24667 63060 24695
rect 62002 24601 62036 24663
rect 62238 24601 62273 24663
rect 62414 24651 62585 24667
rect 62414 24617 62545 24651
rect 62579 24617 62585 24651
rect 62414 24601 62585 24617
rect 62790 24605 62824 24667
rect 63026 24605 63060 24667
rect 63144 24667 63420 24695
rect 63144 24605 63178 24667
rect 63380 24605 63420 24667
rect 61524 24589 61570 24601
rect 61524 24213 61530 24589
rect 61564 24213 61570 24589
rect 61524 24201 61570 24213
rect 61642 24589 61688 24601
rect 61642 24213 61648 24589
rect 61682 24213 61688 24589
rect 61642 24201 61688 24213
rect 61760 24589 61806 24601
rect 61760 24213 61766 24589
rect 61800 24213 61806 24589
rect 61760 24201 61806 24213
rect 61878 24589 61924 24601
rect 61878 24213 61884 24589
rect 61918 24213 61924 24589
rect 61878 24201 61924 24213
rect 61996 24589 62042 24601
rect 61996 24213 62002 24589
rect 62036 24213 62042 24589
rect 61996 24201 62042 24213
rect 62114 24589 62160 24601
rect 62114 24213 62120 24589
rect 62154 24213 62160 24589
rect 62114 24201 62160 24213
rect 62232 24589 62278 24601
rect 62232 24213 62238 24589
rect 62272 24213 62278 24589
rect 62232 24201 62278 24213
rect 60266 24096 60540 24124
rect 59912 24092 60540 24096
rect 59436 24080 59482 24092
rect 57834 24032 57926 24035
rect 56822 23964 56931 24018
rect 56142 23925 56369 23961
rect 56142 23818 56177 23925
rect 56303 23891 56369 23925
rect 56303 23857 56319 23891
rect 56353 23857 56369 23891
rect 56650 23949 56747 23964
rect 56650 23882 56707 23949
rect 56303 23851 56369 23857
rect 56544 23846 56813 23882
rect 56544 23818 56577 23846
rect 56780 23818 56813 23846
rect 56897 23818 56931 23964
rect 57748 23957 57758 24032
rect 57826 23957 57926 24032
rect 57775 23956 57926 23957
rect 56018 23806 56064 23818
rect 56018 23630 56024 23806
rect 56058 23630 56064 23806
rect 56018 23618 56064 23630
rect 56136 23806 56182 23818
rect 56136 23630 56142 23806
rect 56176 23630 56182 23806
rect 56136 23618 56182 23630
rect 56254 23806 56300 23818
rect 56254 23630 56260 23806
rect 56294 23630 56300 23806
rect 56254 23618 56300 23630
rect 56372 23806 56418 23818
rect 56372 23630 56378 23806
rect 56412 23751 56418 23806
rect 56537 23806 56583 23818
rect 56537 23751 56543 23806
rect 56412 23663 56543 23751
rect 56412 23630 56418 23663
rect 56372 23618 56418 23630
rect 56537 23630 56543 23663
rect 56577 23630 56583 23806
rect 56537 23618 56583 23630
rect 56655 23806 56701 23818
rect 56655 23630 56661 23806
rect 56695 23630 56701 23806
rect 56655 23618 56701 23630
rect 56773 23806 56819 23818
rect 56773 23630 56779 23806
rect 56813 23630 56819 23806
rect 56773 23618 56819 23630
rect 56891 23806 56937 23818
rect 56891 23630 56897 23806
rect 56931 23630 56937 23806
rect 56891 23618 56937 23630
rect 56024 23579 56058 23618
rect 56260 23579 56294 23618
rect 56024 23543 56294 23579
rect 56661 23580 56694 23618
rect 56897 23580 56930 23618
rect 56661 23544 56930 23580
rect 56024 23542 56190 23543
rect 56058 23463 56190 23542
rect 56048 23355 56058 23463
rect 56190 23355 56200 23463
rect 52662 22981 53639 23011
rect 55856 23009 55919 23026
rect 55781 23005 55919 23009
rect 52662 22875 52694 22981
rect 52898 22875 52930 22981
rect 53134 22875 53166 22981
rect 53370 22875 53402 22981
rect 53605 22875 53639 22981
rect 53949 22971 55919 23005
rect 53947 22942 55919 22971
rect 53947 22926 53993 22942
rect 55781 22940 55919 22942
rect 52655 22863 52701 22875
rect 52655 22687 52661 22863
rect 52695 22687 52701 22863
rect 52655 22675 52701 22687
rect 52773 22863 52819 22875
rect 52773 22687 52779 22863
rect 52813 22687 52819 22863
rect 52773 22675 52819 22687
rect 52891 22863 52937 22875
rect 52891 22687 52897 22863
rect 52931 22687 52937 22863
rect 52891 22675 52937 22687
rect 53009 22863 53055 22875
rect 53009 22687 53015 22863
rect 53049 22687 53055 22863
rect 53009 22675 53055 22687
rect 53127 22863 53173 22875
rect 53127 22687 53133 22863
rect 53167 22687 53173 22863
rect 53127 22675 53173 22687
rect 53245 22863 53291 22875
rect 53245 22687 53251 22863
rect 53285 22687 53291 22863
rect 53245 22675 53291 22687
rect 53363 22863 53409 22875
rect 53363 22687 53369 22863
rect 53403 22687 53409 22863
rect 53363 22675 53409 22687
rect 53481 22863 53527 22875
rect 53481 22687 53487 22863
rect 53521 22687 53527 22863
rect 53481 22675 53527 22687
rect 53599 22863 53645 22875
rect 53599 22687 53605 22863
rect 53639 22687 53645 22863
rect 53599 22675 53645 22687
rect 53717 22863 53763 22875
rect 53717 22687 53723 22863
rect 53757 22687 53763 22863
rect 53717 22675 53763 22687
rect 52778 22581 52814 22675
rect 53014 22581 53050 22675
rect 53250 22582 53286 22675
rect 53412 22627 53478 22634
rect 53412 22593 53428 22627
rect 53462 22593 53478 22627
rect 53412 22582 53478 22593
rect 53250 22581 53478 22582
rect 52778 22552 53478 22581
rect 52778 22551 53360 22552
rect 52898 22438 52932 22551
rect 53294 22510 53360 22551
rect 53294 22476 53310 22510
rect 53344 22476 53360 22510
rect 53294 22469 53360 22476
rect 53722 22457 53757 22675
rect 53946 22474 53993 22926
rect 54905 22710 54915 22818
rect 55047 22710 55057 22818
rect 56803 22710 56813 22818
rect 56945 22710 56955 22818
rect 54915 22670 55047 22710
rect 56813 22670 56945 22710
rect 54914 22604 55047 22670
rect 56812 22604 56945 22670
rect 54243 22561 55716 22604
rect 53946 22458 53992 22474
rect 53911 22457 53992 22458
rect 53722 22442 53992 22457
rect 53368 22438 53992 22442
rect 52892 22426 52938 22438
rect 52627 21948 52637 22066
rect 52755 22034 52765 22066
rect 52892 22050 52898 22426
rect 52932 22050 52938 22426
rect 52892 22038 52938 22050
rect 53010 22426 53056 22438
rect 53010 22050 53016 22426
rect 53050 22050 53056 22426
rect 53010 22038 53056 22050
rect 53128 22426 53174 22438
rect 53128 22050 53134 22426
rect 53168 22074 53174 22426
rect 53245 22426 53291 22438
rect 53245 22250 53251 22426
rect 53285 22250 53291 22426
rect 53245 22238 53291 22250
rect 53363 22426 53992 22438
rect 53363 22250 53369 22426
rect 53403 22414 53992 22426
rect 53403 22413 53645 22414
rect 53403 22250 53409 22413
rect 53911 22412 53992 22414
rect 54243 22258 54277 22561
rect 54609 22458 54643 22561
rect 54845 22458 54879 22561
rect 55081 22458 55115 22561
rect 55317 22458 55351 22561
rect 54603 22446 54649 22458
rect 53363 22238 53409 22250
rect 54119 22246 54165 22258
rect 53251 22122 53286 22238
rect 53382 22122 53490 22132
rect 53251 22074 53382 22122
rect 53168 22050 53382 22074
rect 53128 22038 53382 22050
rect 53134 22034 53382 22038
rect 52755 22006 52770 22034
rect 52755 22000 53007 22006
rect 52755 21966 52957 22000
rect 52991 21966 53007 22000
rect 52755 21950 53007 21966
rect 53059 22000 53125 22006
rect 53059 21966 53075 22000
rect 53109 21966 53125 22000
rect 53308 21990 53382 22034
rect 54119 22070 54125 22246
rect 54159 22070 54165 22246
rect 54119 22058 54165 22070
rect 54237 22246 54283 22258
rect 54237 22070 54243 22246
rect 54277 22070 54283 22246
rect 54237 22058 54283 22070
rect 54355 22246 54401 22258
rect 54355 22070 54361 22246
rect 54395 22070 54401 22246
rect 54355 22058 54401 22070
rect 54473 22246 54519 22258
rect 54603 22246 54609 22446
rect 54473 22070 54479 22246
rect 54513 22070 54609 22246
rect 54643 22070 54649 22446
rect 54473 22058 54519 22070
rect 54603 22058 54649 22070
rect 54721 22446 54767 22458
rect 54721 22070 54727 22446
rect 54761 22070 54767 22446
rect 54721 22058 54767 22070
rect 54839 22446 54885 22458
rect 54839 22070 54845 22446
rect 54879 22070 54885 22446
rect 54839 22058 54885 22070
rect 54957 22446 55003 22458
rect 54957 22070 54963 22446
rect 54997 22070 55003 22446
rect 54957 22058 55003 22070
rect 55075 22446 55121 22458
rect 55075 22070 55081 22446
rect 55115 22070 55121 22446
rect 55075 22058 55121 22070
rect 55193 22446 55239 22458
rect 55193 22070 55199 22446
rect 55233 22070 55239 22446
rect 55193 22058 55239 22070
rect 55311 22446 55357 22458
rect 55311 22070 55317 22446
rect 55351 22246 55357 22446
rect 55682 22258 55716 22561
rect 56141 22561 57614 22604
rect 56141 22258 56175 22561
rect 56507 22458 56541 22561
rect 56743 22458 56777 22561
rect 56979 22458 57013 22561
rect 57215 22458 57249 22561
rect 56501 22446 56547 22458
rect 55440 22246 55486 22258
rect 55351 22070 55446 22246
rect 55480 22070 55486 22246
rect 55311 22058 55357 22070
rect 55440 22058 55486 22070
rect 55558 22246 55604 22258
rect 55558 22070 55564 22246
rect 55598 22070 55604 22246
rect 55558 22058 55604 22070
rect 55676 22246 55722 22258
rect 55676 22070 55682 22246
rect 55716 22070 55722 22246
rect 55676 22058 55722 22070
rect 55794 22246 55840 22258
rect 55794 22070 55800 22246
rect 55834 22070 55840 22246
rect 55794 22058 55840 22070
rect 56017 22246 56063 22258
rect 56017 22070 56023 22246
rect 56057 22070 56063 22246
rect 56017 22058 56063 22070
rect 56135 22246 56181 22258
rect 56135 22070 56141 22246
rect 56175 22070 56181 22246
rect 56135 22058 56181 22070
rect 56253 22246 56299 22258
rect 56253 22070 56259 22246
rect 56293 22070 56299 22246
rect 56253 22058 56299 22070
rect 56371 22246 56417 22258
rect 56501 22246 56507 22446
rect 56371 22070 56377 22246
rect 56411 22070 56507 22246
rect 56541 22070 56547 22446
rect 56371 22058 56417 22070
rect 56501 22058 56547 22070
rect 56619 22446 56665 22458
rect 56619 22070 56625 22446
rect 56659 22070 56665 22446
rect 56619 22058 56665 22070
rect 56737 22446 56783 22458
rect 56737 22070 56743 22446
rect 56777 22070 56783 22446
rect 56737 22058 56783 22070
rect 56855 22446 56901 22458
rect 56855 22070 56861 22446
rect 56895 22070 56901 22446
rect 56855 22058 56901 22070
rect 56973 22446 57019 22458
rect 56973 22070 56979 22446
rect 57013 22070 57019 22446
rect 56973 22058 57019 22070
rect 57091 22446 57137 22458
rect 57091 22070 57097 22446
rect 57131 22070 57137 22446
rect 57091 22058 57137 22070
rect 57209 22446 57255 22458
rect 57209 22070 57215 22446
rect 57249 22246 57255 22446
rect 57580 22258 57614 22561
rect 57338 22246 57384 22258
rect 57249 22070 57344 22246
rect 57378 22070 57384 22246
rect 57209 22058 57255 22070
rect 57338 22058 57384 22070
rect 57456 22246 57502 22258
rect 57456 22070 57462 22246
rect 57496 22070 57502 22246
rect 57456 22058 57502 22070
rect 57574 22246 57620 22258
rect 57574 22070 57580 22246
rect 57614 22070 57620 22246
rect 57574 22058 57620 22070
rect 57692 22246 57738 22258
rect 57692 22070 57698 22246
rect 57732 22070 57738 22246
rect 57834 22220 57926 23956
rect 58264 23759 58553 23778
rect 58264 23596 58287 23759
rect 58534 23687 58553 23759
rect 59436 23704 59442 24080
rect 59476 23704 59482 24080
rect 59436 23692 59482 23704
rect 59554 24080 59600 24092
rect 59554 23704 59560 24080
rect 59594 23704 59600 24080
rect 59554 23692 59600 23704
rect 59672 24080 59718 24092
rect 59672 23704 59678 24080
rect 59712 23728 59718 24080
rect 59789 24080 59835 24092
rect 59789 23904 59795 24080
rect 59829 23904 59835 24080
rect 59789 23892 59835 23904
rect 59907 24080 60540 24092
rect 59907 23904 59913 24080
rect 59947 24067 60540 24080
rect 61530 24159 61564 24201
rect 61766 24159 61800 24201
rect 61530 24131 61800 24159
rect 61884 24160 61918 24201
rect 62120 24160 62154 24201
rect 61884 24131 62154 24160
rect 61530 24083 61564 24131
rect 59947 23904 59953 24067
rect 61530 24053 61593 24083
rect 59907 23892 59953 23904
rect 61558 23961 61593 24053
rect 61558 23925 61785 23961
rect 62055 23950 62065 24047
rect 62164 23950 62174 24047
rect 62238 24018 62272 24201
rect 62238 23964 62347 24018
rect 59795 23776 59830 23892
rect 61558 23818 61593 23925
rect 61719 23891 61785 23925
rect 61719 23857 61735 23891
rect 61769 23857 61785 23891
rect 62066 23949 62163 23950
rect 62066 23882 62123 23949
rect 61719 23851 61785 23857
rect 61960 23846 62229 23882
rect 61960 23818 61993 23846
rect 62196 23818 62229 23846
rect 62313 23818 62347 23964
rect 61434 23806 61480 23818
rect 59926 23776 60034 23786
rect 59795 23728 59926 23776
rect 59712 23704 59926 23728
rect 59672 23692 59926 23704
rect 59678 23688 59926 23692
rect 58534 23660 59314 23687
rect 58534 23654 59551 23660
rect 58534 23620 59501 23654
rect 59535 23620 59551 23654
rect 58534 23604 59551 23620
rect 59603 23654 59669 23660
rect 59603 23620 59619 23654
rect 59653 23620 59669 23654
rect 59852 23644 59926 23688
rect 59926 23634 60034 23644
rect 58534 23596 59314 23604
rect 58264 23588 59314 23596
rect 58264 23587 59251 23588
rect 58264 23583 58786 23587
rect 58264 23582 58553 23583
rect 58281 22220 58569 22222
rect 57834 22104 58569 22220
rect 57692 22058 57738 22070
rect 58281 22060 58569 22104
rect 53382 21980 53490 21990
rect 54125 22024 54159 22058
rect 54727 22024 54761 22058
rect 54963 22024 54997 22058
rect 54125 21989 54284 22024
rect 54727 21989 54997 22024
rect 55564 22024 55598 22058
rect 55800 22024 55834 22058
rect 55564 21989 55834 22024
rect 56023 22024 56057 22058
rect 56625 22024 56659 22058
rect 56861 22024 56895 22058
rect 56023 21989 56182 22024
rect 56625 21989 56895 22024
rect 57462 22024 57496 22058
rect 57698 22024 57732 22058
rect 57462 21989 57732 22024
rect 52755 21948 52770 21950
rect 52670 21934 52770 21948
rect 52670 21891 52770 21892
rect 52291 21870 52770 21891
rect 53059 21870 53125 21966
rect 52291 21822 53125 21870
rect 52291 21793 52770 21822
rect 52291 21791 52396 21793
rect 52670 21792 52770 21793
rect 52124 21606 52134 21685
rect 52227 21606 52237 21685
rect 52135 20432 52228 21606
rect 53053 21557 53273 21577
rect 53053 21449 53097 21557
rect 53229 21449 53273 21557
rect 53053 21407 53273 21449
rect 52657 21377 53634 21407
rect 52657 21271 52689 21377
rect 52893 21271 52925 21377
rect 53129 21271 53161 21377
rect 53365 21271 53397 21377
rect 53600 21271 53634 21377
rect 52650 21259 52696 21271
rect 52650 21083 52656 21259
rect 52690 21083 52696 21259
rect 52650 21071 52696 21083
rect 52768 21259 52814 21271
rect 52768 21083 52774 21259
rect 52808 21083 52814 21259
rect 52768 21071 52814 21083
rect 52886 21259 52932 21271
rect 52886 21083 52892 21259
rect 52926 21083 52932 21259
rect 52886 21071 52932 21083
rect 53004 21259 53050 21271
rect 53004 21083 53010 21259
rect 53044 21083 53050 21259
rect 53004 21071 53050 21083
rect 53122 21259 53168 21271
rect 53122 21083 53128 21259
rect 53162 21083 53168 21259
rect 53122 21071 53168 21083
rect 53240 21259 53286 21271
rect 53240 21083 53246 21259
rect 53280 21083 53286 21259
rect 53240 21071 53286 21083
rect 53358 21259 53404 21271
rect 53358 21083 53364 21259
rect 53398 21083 53404 21259
rect 53358 21071 53404 21083
rect 53476 21259 53522 21271
rect 53476 21083 53482 21259
rect 53516 21083 53522 21259
rect 53476 21071 53522 21083
rect 53594 21259 53640 21271
rect 53594 21083 53600 21259
rect 53634 21083 53640 21259
rect 53594 21071 53640 21083
rect 53712 21259 53758 21271
rect 53712 21083 53718 21259
rect 53752 21083 53758 21259
rect 53712 21071 53758 21083
rect 54250 21205 54284 21989
rect 54963 21927 54997 21989
rect 54552 21889 55294 21927
rect 54552 21765 54586 21889
rect 54788 21765 54822 21889
rect 55024 21765 55058 21889
rect 55260 21765 55294 21889
rect 55550 21782 55560 21848
rect 55623 21782 55633 21848
rect 54546 21753 54592 21765
rect 54546 21377 54552 21753
rect 54586 21377 54592 21753
rect 54546 21365 54592 21377
rect 54664 21753 54710 21765
rect 54664 21377 54670 21753
rect 54704 21377 54710 21753
rect 54664 21365 54710 21377
rect 54782 21753 54828 21765
rect 54782 21377 54788 21753
rect 54822 21377 54828 21753
rect 54782 21365 54828 21377
rect 54900 21753 54946 21765
rect 54900 21377 54906 21753
rect 54940 21377 54946 21753
rect 54900 21365 54946 21377
rect 55018 21753 55064 21765
rect 55018 21377 55024 21753
rect 55058 21377 55064 21753
rect 55018 21365 55064 21377
rect 55136 21753 55182 21765
rect 55136 21377 55142 21753
rect 55176 21377 55182 21753
rect 55136 21365 55182 21377
rect 55254 21753 55300 21765
rect 55254 21377 55260 21753
rect 55294 21377 55300 21753
rect 55254 21365 55300 21377
rect 55666 21206 55700 21989
rect 55393 21205 55700 21206
rect 54250 21200 54566 21205
rect 55280 21200 55700 21205
rect 54250 21189 54633 21200
rect 54250 21162 54582 21189
rect 52773 20977 52809 21071
rect 53009 20977 53045 21071
rect 53245 20978 53281 21071
rect 53407 21023 53473 21030
rect 53407 20989 53423 21023
rect 53457 20989 53473 21023
rect 53407 20978 53473 20989
rect 53245 20977 53473 20978
rect 52773 20948 53473 20977
rect 52773 20947 53355 20948
rect 52893 20834 52927 20947
rect 53289 20906 53355 20947
rect 53289 20872 53305 20906
rect 53339 20872 53355 20906
rect 53289 20865 53355 20872
rect 53717 20838 53752 21071
rect 54250 21033 54284 21162
rect 54566 21155 54582 21162
rect 54616 21155 54633 21189
rect 54566 21149 54633 21155
rect 55213 21189 55700 21200
rect 55213 21155 55230 21189
rect 55264 21162 55700 21189
rect 55264 21155 55280 21162
rect 55393 21161 55700 21162
rect 55213 21149 55280 21155
rect 54391 21122 54447 21134
rect 54391 21088 54397 21122
rect 54431 21121 54447 21122
rect 55504 21121 55560 21133
rect 54431 21105 54898 21121
rect 54431 21088 54848 21105
rect 54391 21072 54848 21088
rect 54832 21071 54848 21072
rect 54882 21071 54898 21105
rect 54832 21064 54898 21071
rect 54950 21106 55520 21121
rect 54950 21072 54966 21106
rect 55000 21087 55520 21106
rect 55554 21087 55560 21121
rect 55000 21072 55560 21087
rect 54950 21062 55017 21072
rect 55504 21071 55560 21072
rect 55666 21033 55700 21161
rect 56148 21205 56182 21989
rect 56861 21927 56895 21989
rect 56450 21889 57192 21927
rect 56450 21765 56484 21889
rect 56686 21765 56720 21889
rect 56922 21765 56956 21889
rect 57158 21765 57192 21889
rect 56444 21753 56490 21765
rect 56444 21377 56450 21753
rect 56484 21377 56490 21753
rect 56444 21365 56490 21377
rect 56562 21753 56608 21765
rect 56562 21377 56568 21753
rect 56602 21377 56608 21753
rect 56562 21365 56608 21377
rect 56680 21753 56726 21765
rect 56680 21377 56686 21753
rect 56720 21377 56726 21753
rect 56680 21365 56726 21377
rect 56798 21753 56844 21765
rect 56798 21377 56804 21753
rect 56838 21377 56844 21753
rect 56798 21365 56844 21377
rect 56916 21753 56962 21765
rect 56916 21377 56922 21753
rect 56956 21377 56962 21753
rect 56916 21365 56962 21377
rect 57034 21753 57080 21765
rect 57034 21377 57040 21753
rect 57074 21377 57080 21753
rect 57034 21365 57080 21377
rect 57152 21753 57198 21765
rect 57152 21377 57158 21753
rect 57192 21377 57198 21753
rect 57152 21365 57198 21377
rect 57564 21206 57598 21989
rect 58281 21954 58417 22060
rect 58529 22058 58569 22060
rect 58535 22047 58569 22058
rect 58281 21952 58423 21954
rect 58535 21952 58570 22047
rect 58281 21943 58570 21952
rect 58281 21942 58569 21943
rect 58281 21941 58537 21942
rect 57176 21205 57245 21206
rect 57291 21205 57598 21206
rect 56148 21200 56464 21205
rect 57176 21201 57598 21205
rect 56148 21189 56531 21200
rect 56148 21162 56480 21189
rect 56148 21033 56182 21162
rect 56464 21155 56480 21162
rect 56514 21155 56531 21189
rect 56464 21149 56531 21155
rect 57109 21190 57598 21201
rect 57109 21156 57126 21190
rect 57160 21162 57598 21190
rect 57160 21156 57176 21162
rect 57291 21161 57598 21162
rect 57109 21150 57176 21156
rect 56289 21122 56345 21134
rect 56289 21088 56295 21122
rect 56329 21121 56345 21122
rect 57402 21121 57458 21133
rect 56329 21105 56796 21121
rect 56329 21088 56746 21105
rect 56289 21072 56746 21088
rect 56730 21071 56746 21072
rect 56780 21071 56796 21105
rect 56730 21064 56796 21071
rect 56848 21106 57418 21121
rect 56848 21072 56864 21106
rect 56898 21087 57418 21106
rect 57452 21087 57458 21121
rect 56898 21072 57458 21087
rect 56848 21062 56915 21072
rect 57402 21071 57458 21072
rect 57564 21033 57598 21161
rect 57679 21811 57746 21835
rect 57679 21777 57696 21811
rect 57730 21777 57746 21811
rect 53363 20834 53752 20838
rect 52887 20822 52933 20834
rect 52887 20446 52893 20822
rect 52927 20446 52933 20822
rect 52887 20434 52933 20446
rect 53005 20822 53051 20834
rect 53005 20446 53011 20822
rect 53045 20446 53051 20822
rect 53005 20434 53051 20446
rect 53123 20822 53169 20834
rect 53123 20446 53129 20822
rect 53163 20470 53169 20822
rect 53240 20822 53286 20834
rect 53240 20646 53246 20822
rect 53280 20646 53286 20822
rect 53240 20634 53286 20646
rect 53358 20822 53752 20834
rect 54244 21021 54290 21033
rect 54244 20845 54250 21021
rect 54284 20845 54290 21021
rect 54244 20833 54290 20845
rect 54362 21021 54408 21033
rect 54362 20845 54368 21021
rect 54402 20845 54408 21021
rect 54362 20833 54408 20845
rect 54664 21021 54710 21033
rect 53358 20646 53364 20822
rect 53398 20809 53752 20822
rect 53398 20646 53404 20809
rect 53674 20806 53752 20809
rect 53674 20754 53684 20806
rect 53747 20754 53757 20806
rect 53679 20748 53752 20754
rect 53358 20634 53404 20646
rect 53246 20518 53281 20634
rect 54367 20539 54401 20833
rect 54664 20645 54670 21021
rect 54704 20645 54710 21021
rect 54664 20633 54710 20645
rect 54782 21021 54828 21033
rect 54782 20645 54788 21021
rect 54822 20645 54828 21021
rect 54782 20633 54828 20645
rect 54900 21021 54946 21033
rect 54900 20645 54906 21021
rect 54940 20645 54946 21021
rect 54900 20633 54946 20645
rect 55018 21021 55064 21033
rect 55018 20645 55024 21021
rect 55058 20645 55064 21021
rect 55018 20633 55064 20645
rect 55136 21021 55182 21033
rect 55136 20645 55142 21021
rect 55176 20645 55182 21021
rect 55542 21021 55588 21033
rect 55542 20845 55548 21021
rect 55582 20845 55588 21021
rect 55542 20833 55588 20845
rect 55660 21021 55706 21033
rect 55660 20845 55666 21021
rect 55700 20845 55706 21021
rect 55660 20833 55706 20845
rect 56142 21021 56188 21033
rect 56142 20845 56148 21021
rect 56182 20845 56188 21021
rect 56142 20833 56188 20845
rect 56260 21021 56306 21033
rect 56260 20845 56266 21021
rect 56300 20845 56306 21021
rect 56260 20833 56306 20845
rect 56562 21021 56608 21033
rect 55136 20633 55182 20645
rect 55024 20539 55058 20633
rect 55548 20539 55581 20833
rect 53377 20518 53485 20528
rect 53246 20470 53377 20518
rect 53163 20446 53377 20470
rect 53123 20434 53377 20446
rect 52135 20430 52720 20432
rect 53129 20430 53377 20434
rect 52135 20402 52765 20430
rect 46217 20223 46586 20271
rect 46217 20193 46231 20223
rect 46217 20176 46227 20193
rect 40004 20043 44698 20123
rect 46519 20120 46585 20223
rect 51145 20120 51211 20399
rect 52135 20396 53002 20402
rect 52135 20362 52952 20396
rect 52986 20362 53002 20396
rect 52135 20346 53002 20362
rect 53054 20396 53120 20402
rect 53054 20362 53070 20396
rect 53104 20362 53120 20396
rect 53303 20386 53377 20430
rect 54367 20507 55581 20539
rect 56265 20539 56299 20833
rect 56562 20645 56568 21021
rect 56602 20645 56608 21021
rect 56562 20633 56608 20645
rect 56680 21021 56726 21033
rect 56680 20645 56686 21021
rect 56720 20645 56726 21021
rect 56680 20633 56726 20645
rect 56798 21021 56844 21033
rect 56798 20645 56804 21021
rect 56838 20645 56844 21021
rect 56798 20633 56844 20645
rect 56916 21021 56962 21033
rect 56916 20645 56922 21021
rect 56956 20645 56962 21021
rect 56916 20633 56962 20645
rect 57034 21021 57080 21033
rect 57034 20645 57040 21021
rect 57074 20645 57080 21021
rect 57440 21021 57486 21033
rect 57440 20845 57446 21021
rect 57480 20845 57486 21021
rect 57440 20833 57486 20845
rect 57558 21021 57604 21033
rect 57558 20845 57564 21021
rect 57598 20845 57604 21021
rect 57558 20833 57604 20845
rect 57034 20633 57080 20645
rect 56922 20539 56956 20633
rect 57446 20539 57479 20833
rect 56265 20507 57479 20539
rect 54860 20422 54992 20507
rect 56758 20422 56890 20507
rect 53377 20376 53485 20386
rect 52135 20330 52765 20346
rect 52135 20326 52720 20330
rect 52135 20325 52236 20326
rect 52665 20277 52765 20288
rect 52629 20171 52639 20277
rect 52751 20266 52765 20277
rect 53054 20266 53120 20362
rect 54850 20314 54860 20422
rect 54992 20314 55002 20422
rect 56748 20314 56758 20422
rect 56890 20314 56900 20422
rect 57679 20394 57746 21777
rect 58693 21689 58786 23583
rect 58849 23524 59315 23546
rect 59603 23524 59669 23620
rect 61434 23630 61440 23806
rect 61474 23630 61480 23806
rect 61434 23618 61480 23630
rect 61552 23806 61598 23818
rect 61552 23630 61558 23806
rect 61592 23630 61598 23806
rect 61552 23618 61598 23630
rect 61670 23806 61716 23818
rect 61670 23630 61676 23806
rect 61710 23630 61716 23806
rect 61670 23618 61716 23630
rect 61788 23806 61834 23818
rect 61788 23630 61794 23806
rect 61828 23751 61834 23806
rect 61953 23806 61999 23818
rect 61953 23751 61959 23806
rect 61828 23663 61959 23751
rect 61828 23630 61834 23663
rect 61788 23618 61834 23630
rect 61953 23630 61959 23663
rect 61993 23630 61999 23806
rect 61953 23618 61999 23630
rect 62071 23806 62117 23818
rect 62071 23630 62077 23806
rect 62111 23630 62117 23806
rect 62071 23618 62117 23630
rect 62189 23806 62235 23818
rect 62189 23630 62195 23806
rect 62229 23630 62235 23806
rect 62189 23618 62235 23630
rect 62307 23806 62353 23818
rect 62307 23630 62313 23806
rect 62347 23630 62353 23806
rect 62307 23618 62353 23630
rect 61440 23579 61474 23618
rect 61676 23579 61710 23618
rect 61440 23544 61710 23579
rect 62077 23580 62110 23618
rect 62313 23580 62346 23618
rect 62077 23544 62346 23580
rect 58849 23476 59669 23524
rect 61474 23543 61710 23544
rect 58849 23445 59315 23476
rect 61474 23469 61606 23543
rect 58849 23189 58954 23445
rect 61464 23361 61474 23469
rect 61606 23361 61616 23469
rect 58849 23083 58912 23189
rect 59024 23083 59034 23189
rect 59616 23165 59836 23185
rect 58849 23072 58998 23083
rect 58849 21895 58954 23072
rect 59616 23057 59660 23165
rect 59792 23057 59836 23165
rect 59616 23015 59836 23057
rect 62414 23030 62476 24601
rect 62666 24593 62712 24605
rect 62666 24217 62672 24593
rect 62706 24217 62712 24593
rect 62666 24205 62712 24217
rect 62784 24593 62830 24605
rect 62784 24217 62790 24593
rect 62824 24217 62830 24593
rect 62784 24205 62830 24217
rect 62902 24593 62948 24605
rect 62902 24217 62908 24593
rect 62942 24217 62948 24593
rect 62902 24205 62948 24217
rect 63020 24593 63066 24605
rect 63020 24217 63026 24593
rect 63060 24217 63066 24593
rect 63020 24205 63066 24217
rect 63138 24593 63184 24605
rect 63138 24217 63144 24593
rect 63178 24217 63184 24593
rect 63138 24205 63184 24217
rect 63256 24593 63302 24605
rect 63256 24217 63262 24593
rect 63296 24217 63302 24593
rect 63256 24205 63302 24217
rect 63374 24593 63420 24605
rect 63374 24217 63380 24593
rect 63414 24217 63420 24593
rect 63374 24205 63420 24217
rect 62672 24163 62706 24205
rect 62908 24163 62942 24205
rect 62672 24135 62942 24163
rect 63026 24164 63060 24205
rect 63262 24164 63296 24205
rect 63026 24135 63296 24164
rect 62672 24087 62706 24135
rect 62672 24057 62735 24087
rect 62700 23965 62735 24057
rect 63207 24027 63307 24048
rect 63207 23973 63221 24027
rect 63286 23973 63307 24027
rect 63207 23968 63307 23973
rect 63380 24022 63414 24205
rect 64414 24036 64780 24038
rect 63380 23968 63489 24022
rect 62700 23929 62927 23965
rect 62700 23822 62735 23929
rect 62861 23895 62927 23929
rect 62861 23861 62877 23895
rect 62911 23861 62927 23895
rect 63208 23953 63305 23968
rect 63208 23886 63265 23953
rect 62861 23855 62927 23861
rect 63102 23850 63371 23886
rect 63102 23822 63135 23850
rect 63338 23822 63371 23850
rect 63455 23822 63489 23968
rect 64306 23961 64316 24036
rect 64384 23961 64780 24036
rect 64333 23960 64780 23961
rect 64379 23956 64780 23960
rect 62576 23810 62622 23822
rect 62576 23634 62582 23810
rect 62616 23634 62622 23810
rect 62576 23622 62622 23634
rect 62694 23810 62740 23822
rect 62694 23634 62700 23810
rect 62734 23634 62740 23810
rect 62694 23622 62740 23634
rect 62812 23810 62858 23822
rect 62812 23634 62818 23810
rect 62852 23634 62858 23810
rect 62812 23622 62858 23634
rect 62930 23810 62976 23822
rect 62930 23634 62936 23810
rect 62970 23755 62976 23810
rect 63095 23810 63141 23822
rect 63095 23755 63101 23810
rect 62970 23667 63101 23755
rect 62970 23634 62976 23667
rect 62930 23622 62976 23634
rect 63095 23634 63101 23667
rect 63135 23634 63141 23810
rect 63095 23622 63141 23634
rect 63213 23810 63259 23822
rect 63213 23634 63219 23810
rect 63253 23634 63259 23810
rect 63213 23622 63259 23634
rect 63331 23810 63377 23822
rect 63331 23634 63337 23810
rect 63371 23634 63377 23810
rect 63331 23622 63377 23634
rect 63449 23810 63495 23822
rect 63449 23634 63455 23810
rect 63489 23634 63495 23810
rect 63449 23622 63495 23634
rect 62582 23583 62616 23622
rect 62818 23583 62852 23622
rect 62582 23547 62852 23583
rect 63219 23584 63252 23622
rect 63455 23584 63488 23622
rect 63219 23548 63488 23584
rect 62582 23546 62748 23547
rect 62616 23467 62748 23546
rect 62606 23359 62616 23467
rect 62748 23359 62758 23467
rect 64653 23038 64780 23956
rect 59220 22985 60197 23015
rect 62414 23013 62477 23030
rect 62339 23009 62477 23013
rect 59220 22879 59252 22985
rect 59456 22879 59488 22985
rect 59692 22879 59724 22985
rect 59928 22879 59960 22985
rect 60163 22879 60197 22985
rect 60507 22975 62477 23009
rect 60505 22946 62477 22975
rect 60505 22930 60551 22946
rect 62339 22944 62477 22946
rect 64655 22931 64778 23038
rect 59213 22867 59259 22879
rect 59213 22691 59219 22867
rect 59253 22691 59259 22867
rect 59213 22679 59259 22691
rect 59331 22867 59377 22879
rect 59331 22691 59337 22867
rect 59371 22691 59377 22867
rect 59331 22679 59377 22691
rect 59449 22867 59495 22879
rect 59449 22691 59455 22867
rect 59489 22691 59495 22867
rect 59449 22679 59495 22691
rect 59567 22867 59613 22879
rect 59567 22691 59573 22867
rect 59607 22691 59613 22867
rect 59567 22679 59613 22691
rect 59685 22867 59731 22879
rect 59685 22691 59691 22867
rect 59725 22691 59731 22867
rect 59685 22679 59731 22691
rect 59803 22867 59849 22879
rect 59803 22691 59809 22867
rect 59843 22691 59849 22867
rect 59803 22679 59849 22691
rect 59921 22867 59967 22879
rect 59921 22691 59927 22867
rect 59961 22691 59967 22867
rect 59921 22679 59967 22691
rect 60039 22867 60085 22879
rect 60039 22691 60045 22867
rect 60079 22691 60085 22867
rect 60039 22679 60085 22691
rect 60157 22867 60203 22879
rect 60157 22691 60163 22867
rect 60197 22691 60203 22867
rect 60157 22679 60203 22691
rect 60275 22867 60321 22879
rect 60275 22691 60281 22867
rect 60315 22691 60321 22867
rect 60275 22679 60321 22691
rect 59336 22585 59372 22679
rect 59572 22585 59608 22679
rect 59808 22586 59844 22679
rect 59970 22631 60036 22638
rect 59970 22597 59986 22631
rect 60020 22597 60036 22631
rect 59970 22586 60036 22597
rect 59808 22585 60036 22586
rect 59336 22556 60036 22585
rect 59336 22555 59918 22556
rect 59456 22442 59490 22555
rect 59852 22514 59918 22555
rect 59852 22480 59868 22514
rect 59902 22480 59918 22514
rect 59852 22473 59918 22480
rect 60280 22461 60315 22679
rect 60504 22478 60551 22930
rect 61463 22714 61473 22822
rect 61605 22714 61615 22822
rect 63361 22714 63371 22822
rect 63503 22714 63513 22822
rect 61473 22674 61605 22714
rect 63371 22674 63503 22714
rect 61472 22608 61605 22674
rect 63370 22608 63503 22674
rect 60801 22565 62274 22608
rect 60504 22462 60550 22478
rect 60469 22461 60550 22462
rect 60280 22446 60550 22461
rect 59926 22442 60550 22446
rect 59450 22430 59496 22442
rect 59185 21952 59195 22070
rect 59313 22038 59323 22070
rect 59450 22054 59456 22430
rect 59490 22054 59496 22430
rect 59450 22042 59496 22054
rect 59568 22430 59614 22442
rect 59568 22054 59574 22430
rect 59608 22054 59614 22430
rect 59568 22042 59614 22054
rect 59686 22430 59732 22442
rect 59686 22054 59692 22430
rect 59726 22078 59732 22430
rect 59803 22430 59849 22442
rect 59803 22254 59809 22430
rect 59843 22254 59849 22430
rect 59803 22242 59849 22254
rect 59921 22430 60550 22442
rect 59921 22254 59927 22430
rect 59961 22418 60550 22430
rect 59961 22417 60203 22418
rect 59961 22254 59967 22417
rect 60469 22416 60550 22418
rect 60801 22262 60835 22565
rect 61167 22462 61201 22565
rect 61403 22462 61437 22565
rect 61639 22462 61673 22565
rect 61875 22462 61909 22565
rect 61161 22450 61207 22462
rect 59921 22242 59967 22254
rect 60677 22250 60723 22262
rect 59809 22126 59844 22242
rect 59940 22126 60048 22136
rect 59809 22078 59940 22126
rect 59726 22054 59940 22078
rect 59686 22042 59940 22054
rect 59692 22038 59940 22042
rect 59313 22010 59328 22038
rect 59313 22004 59565 22010
rect 59313 21970 59515 22004
rect 59549 21970 59565 22004
rect 59313 21954 59565 21970
rect 59617 22004 59683 22010
rect 59617 21970 59633 22004
rect 59667 21970 59683 22004
rect 59866 21994 59940 22038
rect 60677 22074 60683 22250
rect 60717 22074 60723 22250
rect 60677 22062 60723 22074
rect 60795 22250 60841 22262
rect 60795 22074 60801 22250
rect 60835 22074 60841 22250
rect 60795 22062 60841 22074
rect 60913 22250 60959 22262
rect 60913 22074 60919 22250
rect 60953 22074 60959 22250
rect 60913 22062 60959 22074
rect 61031 22250 61077 22262
rect 61161 22250 61167 22450
rect 61031 22074 61037 22250
rect 61071 22074 61167 22250
rect 61201 22074 61207 22450
rect 61031 22062 61077 22074
rect 61161 22062 61207 22074
rect 61279 22450 61325 22462
rect 61279 22074 61285 22450
rect 61319 22074 61325 22450
rect 61279 22062 61325 22074
rect 61397 22450 61443 22462
rect 61397 22074 61403 22450
rect 61437 22074 61443 22450
rect 61397 22062 61443 22074
rect 61515 22450 61561 22462
rect 61515 22074 61521 22450
rect 61555 22074 61561 22450
rect 61515 22062 61561 22074
rect 61633 22450 61679 22462
rect 61633 22074 61639 22450
rect 61673 22074 61679 22450
rect 61633 22062 61679 22074
rect 61751 22450 61797 22462
rect 61751 22074 61757 22450
rect 61791 22074 61797 22450
rect 61751 22062 61797 22074
rect 61869 22450 61915 22462
rect 61869 22074 61875 22450
rect 61909 22250 61915 22450
rect 62240 22262 62274 22565
rect 62699 22565 64172 22608
rect 62699 22262 62733 22565
rect 63065 22462 63099 22565
rect 63301 22462 63335 22565
rect 63537 22462 63571 22565
rect 63773 22462 63807 22565
rect 63059 22450 63105 22462
rect 61998 22250 62044 22262
rect 61909 22074 62004 22250
rect 62038 22074 62044 22250
rect 61869 22062 61915 22074
rect 61998 22062 62044 22074
rect 62116 22250 62162 22262
rect 62116 22074 62122 22250
rect 62156 22074 62162 22250
rect 62116 22062 62162 22074
rect 62234 22250 62280 22262
rect 62234 22074 62240 22250
rect 62274 22074 62280 22250
rect 62234 22062 62280 22074
rect 62352 22250 62398 22262
rect 62352 22074 62358 22250
rect 62392 22074 62398 22250
rect 62352 22062 62398 22074
rect 62575 22250 62621 22262
rect 62575 22074 62581 22250
rect 62615 22074 62621 22250
rect 62575 22062 62621 22074
rect 62693 22250 62739 22262
rect 62693 22074 62699 22250
rect 62733 22074 62739 22250
rect 62693 22062 62739 22074
rect 62811 22250 62857 22262
rect 62811 22074 62817 22250
rect 62851 22074 62857 22250
rect 62811 22062 62857 22074
rect 62929 22250 62975 22262
rect 63059 22250 63065 22450
rect 62929 22074 62935 22250
rect 62969 22074 63065 22250
rect 63099 22074 63105 22450
rect 62929 22062 62975 22074
rect 63059 22062 63105 22074
rect 63177 22450 63223 22462
rect 63177 22074 63183 22450
rect 63217 22074 63223 22450
rect 63177 22062 63223 22074
rect 63295 22450 63341 22462
rect 63295 22074 63301 22450
rect 63335 22074 63341 22450
rect 63295 22062 63341 22074
rect 63413 22450 63459 22462
rect 63413 22074 63419 22450
rect 63453 22074 63459 22450
rect 63413 22062 63459 22074
rect 63531 22450 63577 22462
rect 63531 22074 63537 22450
rect 63571 22074 63577 22450
rect 63531 22062 63577 22074
rect 63649 22450 63695 22462
rect 63649 22074 63655 22450
rect 63689 22074 63695 22450
rect 63649 22062 63695 22074
rect 63767 22450 63813 22462
rect 63767 22074 63773 22450
rect 63807 22250 63813 22450
rect 64138 22262 64172 22565
rect 63896 22250 63942 22262
rect 63807 22074 63902 22250
rect 63936 22074 63942 22250
rect 63767 22062 63813 22074
rect 63896 22062 63942 22074
rect 64014 22250 64060 22262
rect 64014 22074 64020 22250
rect 64054 22074 64060 22250
rect 64014 22062 64060 22074
rect 64132 22250 64178 22262
rect 64132 22074 64138 22250
rect 64172 22074 64178 22250
rect 64132 22062 64178 22074
rect 64250 22250 64296 22262
rect 64250 22074 64256 22250
rect 64290 22074 64296 22250
rect 64250 22062 64296 22074
rect 59940 21984 60048 21994
rect 60683 22028 60717 22062
rect 61285 22028 61319 22062
rect 61521 22028 61555 22062
rect 60683 21993 60842 22028
rect 61285 21993 61555 22028
rect 62122 22028 62156 22062
rect 62358 22028 62392 22062
rect 62122 21993 62392 22028
rect 62581 22028 62615 22062
rect 63183 22028 63217 22062
rect 63419 22028 63453 22062
rect 62581 21993 62740 22028
rect 63183 21993 63453 22028
rect 64020 22028 64054 22062
rect 64256 22028 64290 22062
rect 64020 21993 64290 22028
rect 59313 21952 59328 21954
rect 59228 21938 59328 21952
rect 59228 21895 59328 21896
rect 58849 21874 59328 21895
rect 59617 21874 59683 21970
rect 58849 21826 59683 21874
rect 58849 21797 59328 21826
rect 58849 21795 58954 21797
rect 59228 21796 59328 21797
rect 58682 21610 58692 21689
rect 58785 21610 58795 21689
rect 58693 20436 58786 21610
rect 59611 21561 59831 21581
rect 59611 21453 59655 21561
rect 59787 21453 59831 21561
rect 59611 21411 59831 21453
rect 59215 21381 60192 21411
rect 59215 21275 59247 21381
rect 59451 21275 59483 21381
rect 59687 21275 59719 21381
rect 59923 21275 59955 21381
rect 60158 21275 60192 21381
rect 59208 21263 59254 21275
rect 59208 21087 59214 21263
rect 59248 21087 59254 21263
rect 59208 21075 59254 21087
rect 59326 21263 59372 21275
rect 59326 21087 59332 21263
rect 59366 21087 59372 21263
rect 59326 21075 59372 21087
rect 59444 21263 59490 21275
rect 59444 21087 59450 21263
rect 59484 21087 59490 21263
rect 59444 21075 59490 21087
rect 59562 21263 59608 21275
rect 59562 21087 59568 21263
rect 59602 21087 59608 21263
rect 59562 21075 59608 21087
rect 59680 21263 59726 21275
rect 59680 21087 59686 21263
rect 59720 21087 59726 21263
rect 59680 21075 59726 21087
rect 59798 21263 59844 21275
rect 59798 21087 59804 21263
rect 59838 21087 59844 21263
rect 59798 21075 59844 21087
rect 59916 21263 59962 21275
rect 59916 21087 59922 21263
rect 59956 21087 59962 21263
rect 59916 21075 59962 21087
rect 60034 21263 60080 21275
rect 60034 21087 60040 21263
rect 60074 21087 60080 21263
rect 60034 21075 60080 21087
rect 60152 21263 60198 21275
rect 60152 21087 60158 21263
rect 60192 21087 60198 21263
rect 60152 21075 60198 21087
rect 60270 21263 60316 21275
rect 60270 21087 60276 21263
rect 60310 21087 60316 21263
rect 60270 21075 60316 21087
rect 60808 21209 60842 21993
rect 61521 21931 61555 21993
rect 61110 21893 61852 21931
rect 61110 21769 61144 21893
rect 61346 21769 61380 21893
rect 61582 21769 61616 21893
rect 61818 21769 61852 21893
rect 62108 21786 62118 21852
rect 62181 21786 62191 21852
rect 61104 21757 61150 21769
rect 61104 21381 61110 21757
rect 61144 21381 61150 21757
rect 61104 21369 61150 21381
rect 61222 21757 61268 21769
rect 61222 21381 61228 21757
rect 61262 21381 61268 21757
rect 61222 21369 61268 21381
rect 61340 21757 61386 21769
rect 61340 21381 61346 21757
rect 61380 21381 61386 21757
rect 61340 21369 61386 21381
rect 61458 21757 61504 21769
rect 61458 21381 61464 21757
rect 61498 21381 61504 21757
rect 61458 21369 61504 21381
rect 61576 21757 61622 21769
rect 61576 21381 61582 21757
rect 61616 21381 61622 21757
rect 61576 21369 61622 21381
rect 61694 21757 61740 21769
rect 61694 21381 61700 21757
rect 61734 21381 61740 21757
rect 61694 21369 61740 21381
rect 61812 21757 61858 21769
rect 61812 21381 61818 21757
rect 61852 21381 61858 21757
rect 61812 21369 61858 21381
rect 62224 21210 62258 21993
rect 61951 21209 62258 21210
rect 60808 21204 61124 21209
rect 61838 21204 62258 21209
rect 60808 21193 61191 21204
rect 60808 21166 61140 21193
rect 59331 20981 59367 21075
rect 59567 20981 59603 21075
rect 59803 20982 59839 21075
rect 59965 21027 60031 21034
rect 59965 20993 59981 21027
rect 60015 20993 60031 21027
rect 59965 20982 60031 20993
rect 59803 20981 60031 20982
rect 59331 20952 60031 20981
rect 59331 20951 59913 20952
rect 59451 20838 59485 20951
rect 59847 20910 59913 20951
rect 59847 20876 59863 20910
rect 59897 20876 59913 20910
rect 59847 20869 59913 20876
rect 60275 20842 60310 21075
rect 60808 21037 60842 21166
rect 61124 21159 61140 21166
rect 61174 21159 61191 21193
rect 61124 21153 61191 21159
rect 61771 21193 62258 21204
rect 61771 21159 61788 21193
rect 61822 21166 62258 21193
rect 61822 21159 61838 21166
rect 61951 21165 62258 21166
rect 61771 21153 61838 21159
rect 60949 21126 61005 21138
rect 60949 21092 60955 21126
rect 60989 21125 61005 21126
rect 62062 21125 62118 21137
rect 60989 21109 61456 21125
rect 60989 21092 61406 21109
rect 60949 21076 61406 21092
rect 61390 21075 61406 21076
rect 61440 21075 61456 21109
rect 61390 21068 61456 21075
rect 61508 21110 62078 21125
rect 61508 21076 61524 21110
rect 61558 21091 62078 21110
rect 62112 21091 62118 21125
rect 61558 21076 62118 21091
rect 61508 21066 61575 21076
rect 62062 21075 62118 21076
rect 62224 21037 62258 21165
rect 62706 21209 62740 21993
rect 63419 21931 63453 21993
rect 63008 21893 63750 21931
rect 63008 21769 63042 21893
rect 63244 21769 63278 21893
rect 63480 21769 63514 21893
rect 63716 21769 63750 21893
rect 63002 21757 63048 21769
rect 63002 21381 63008 21757
rect 63042 21381 63048 21757
rect 63002 21369 63048 21381
rect 63120 21757 63166 21769
rect 63120 21381 63126 21757
rect 63160 21381 63166 21757
rect 63120 21369 63166 21381
rect 63238 21757 63284 21769
rect 63238 21381 63244 21757
rect 63278 21381 63284 21757
rect 63238 21369 63284 21381
rect 63356 21757 63402 21769
rect 63356 21381 63362 21757
rect 63396 21381 63402 21757
rect 63356 21369 63402 21381
rect 63474 21757 63520 21769
rect 63474 21381 63480 21757
rect 63514 21381 63520 21757
rect 63474 21369 63520 21381
rect 63592 21757 63638 21769
rect 63592 21381 63598 21757
rect 63632 21381 63638 21757
rect 63592 21369 63638 21381
rect 63710 21757 63756 21769
rect 63710 21381 63716 21757
rect 63750 21381 63756 21757
rect 63710 21369 63756 21381
rect 64122 21210 64156 21993
rect 63734 21209 63803 21210
rect 63849 21209 64156 21210
rect 62706 21204 63022 21209
rect 63734 21205 64156 21209
rect 62706 21193 63089 21204
rect 62706 21166 63038 21193
rect 62706 21037 62740 21166
rect 63022 21159 63038 21166
rect 63072 21159 63089 21193
rect 63022 21153 63089 21159
rect 63667 21194 64156 21205
rect 63667 21160 63684 21194
rect 63718 21166 64156 21194
rect 63718 21160 63734 21166
rect 63849 21165 64156 21166
rect 63667 21154 63734 21160
rect 62847 21126 62903 21138
rect 62847 21092 62853 21126
rect 62887 21125 62903 21126
rect 63960 21125 64016 21137
rect 62887 21109 63354 21125
rect 62887 21092 63304 21109
rect 62847 21076 63304 21092
rect 63288 21075 63304 21076
rect 63338 21075 63354 21109
rect 63288 21068 63354 21075
rect 63406 21110 63976 21125
rect 63406 21076 63422 21110
rect 63456 21091 63976 21110
rect 64010 21091 64016 21125
rect 63456 21076 64016 21091
rect 63406 21066 63473 21076
rect 63960 21075 64016 21076
rect 64122 21037 64156 21165
rect 64237 21815 64304 21839
rect 64237 21781 64254 21815
rect 64288 21781 64304 21815
rect 59921 20838 60310 20842
rect 59445 20826 59491 20838
rect 59445 20450 59451 20826
rect 59485 20450 59491 20826
rect 59445 20438 59491 20450
rect 59563 20826 59609 20838
rect 59563 20450 59569 20826
rect 59603 20450 59609 20826
rect 59563 20438 59609 20450
rect 59681 20826 59727 20838
rect 59681 20450 59687 20826
rect 59721 20474 59727 20826
rect 59798 20826 59844 20838
rect 59798 20650 59804 20826
rect 59838 20650 59844 20826
rect 59798 20638 59844 20650
rect 59916 20826 60310 20838
rect 60802 21025 60848 21037
rect 60802 20849 60808 21025
rect 60842 20849 60848 21025
rect 60802 20837 60848 20849
rect 60920 21025 60966 21037
rect 60920 20849 60926 21025
rect 60960 20849 60966 21025
rect 60920 20837 60966 20849
rect 61222 21025 61268 21037
rect 59916 20650 59922 20826
rect 59956 20813 60310 20826
rect 59956 20650 59962 20813
rect 60232 20810 60310 20813
rect 60232 20758 60242 20810
rect 60305 20758 60315 20810
rect 60237 20752 60310 20758
rect 59916 20638 59962 20650
rect 59804 20522 59839 20638
rect 60925 20543 60959 20837
rect 61222 20649 61228 21025
rect 61262 20649 61268 21025
rect 61222 20637 61268 20649
rect 61340 21025 61386 21037
rect 61340 20649 61346 21025
rect 61380 20649 61386 21025
rect 61340 20637 61386 20649
rect 61458 21025 61504 21037
rect 61458 20649 61464 21025
rect 61498 20649 61504 21025
rect 61458 20637 61504 20649
rect 61576 21025 61622 21037
rect 61576 20649 61582 21025
rect 61616 20649 61622 21025
rect 61576 20637 61622 20649
rect 61694 21025 61740 21037
rect 61694 20649 61700 21025
rect 61734 20649 61740 21025
rect 62100 21025 62146 21037
rect 62100 20849 62106 21025
rect 62140 20849 62146 21025
rect 62100 20837 62146 20849
rect 62218 21025 62264 21037
rect 62218 20849 62224 21025
rect 62258 20849 62264 21025
rect 62218 20837 62264 20849
rect 62700 21025 62746 21037
rect 62700 20849 62706 21025
rect 62740 20849 62746 21025
rect 62700 20837 62746 20849
rect 62818 21025 62864 21037
rect 62818 20849 62824 21025
rect 62858 20849 62864 21025
rect 62818 20837 62864 20849
rect 63120 21025 63166 21037
rect 61694 20637 61740 20649
rect 61582 20543 61616 20637
rect 62106 20543 62139 20837
rect 59935 20522 60043 20532
rect 59804 20474 59935 20522
rect 59721 20450 59935 20474
rect 59681 20438 59935 20450
rect 58693 20434 59278 20436
rect 59687 20434 59935 20438
rect 58693 20406 59323 20434
rect 58693 20400 59560 20406
rect 52751 20218 53120 20266
rect 52751 20188 52765 20218
rect 52751 20171 52761 20188
rect 46517 20040 51211 20120
rect 53053 20115 53119 20218
rect 57679 20115 57745 20394
rect 58693 20366 59510 20400
rect 59544 20366 59560 20400
rect 58693 20350 59560 20366
rect 59612 20400 59678 20406
rect 59612 20366 59628 20400
rect 59662 20366 59678 20400
rect 59861 20390 59935 20434
rect 60925 20511 62139 20543
rect 62823 20543 62857 20837
rect 63120 20649 63126 21025
rect 63160 20649 63166 21025
rect 63120 20637 63166 20649
rect 63238 21025 63284 21037
rect 63238 20649 63244 21025
rect 63278 20649 63284 21025
rect 63238 20637 63284 20649
rect 63356 21025 63402 21037
rect 63356 20649 63362 21025
rect 63396 20649 63402 21025
rect 63356 20637 63402 20649
rect 63474 21025 63520 21037
rect 63474 20649 63480 21025
rect 63514 20649 63520 21025
rect 63474 20637 63520 20649
rect 63592 21025 63638 21037
rect 63592 20649 63598 21025
rect 63632 20649 63638 21025
rect 63998 21025 64044 21037
rect 63998 20849 64004 21025
rect 64038 20849 64044 21025
rect 63998 20837 64044 20849
rect 64116 21025 64162 21037
rect 64116 20849 64122 21025
rect 64156 20849 64162 21025
rect 64116 20837 64162 20849
rect 63592 20637 63638 20649
rect 63480 20543 63514 20637
rect 64004 20543 64037 20837
rect 62823 20511 64037 20543
rect 61418 20426 61550 20511
rect 63316 20426 63448 20511
rect 59935 20380 60043 20390
rect 58693 20334 59323 20350
rect 58693 20330 59278 20334
rect 58693 20329 58794 20330
rect 59223 20281 59323 20292
rect 59187 20175 59197 20281
rect 59309 20270 59323 20281
rect 59612 20270 59678 20366
rect 61408 20318 61418 20426
rect 61550 20318 61560 20426
rect 63306 20318 63316 20426
rect 63448 20318 63458 20426
rect 64237 20398 64304 21781
rect 59309 20222 59678 20270
rect 59309 20192 59323 20222
rect 59309 20175 59319 20192
rect 59611 20119 59677 20222
rect 64237 20119 64303 20398
rect 53051 20035 57745 20115
rect 59609 20039 64303 20119
rect 34249 19996 34648 19997
rect 34249 19985 45170 19996
rect 34249 19907 45026 19985
rect 45154 19907 45170 19985
rect 34249 19893 45170 19907
rect 34112 19834 51673 19853
rect 34112 19723 51539 19834
rect 51650 19723 51673 19834
rect 34112 19710 51673 19723
rect 34112 19709 51461 19710
rect 33952 19651 58274 19663
rect 33952 19533 58127 19651
rect 58261 19533 58274 19651
rect 33952 19519 58274 19533
rect 39608 19202 39618 19265
rect 39606 19191 39618 19202
rect 39605 19157 39618 19191
rect 39750 19157 39760 19265
rect 40755 19202 40765 19265
rect 40753 19191 40765 19202
rect 40440 19181 40496 19183
rect 39605 19119 39750 19157
rect 39605 19091 39646 19119
rect 40430 19115 40440 19181
rect 40496 19115 40506 19181
rect 40752 19157 40765 19191
rect 40897 19157 40907 19265
rect 43203 19211 43423 19231
rect 41570 19169 41626 19177
rect 41570 19161 42552 19169
rect 40752 19119 40897 19157
rect 41570 19127 41576 19161
rect 41610 19127 42552 19161
rect 39605 19063 39881 19091
rect 39605 19001 39645 19063
rect 39847 19001 39881 19063
rect 39965 19063 40235 19091
rect 40752 19087 40793 19119
rect 41570 19111 42552 19127
rect 41573 19110 42552 19111
rect 39965 19001 39999 19063
rect 40201 19001 40235 19063
rect 40440 19047 40611 19063
rect 40440 19013 40446 19047
rect 40480 19013 40611 19047
rect 39605 18989 39651 19001
rect 39605 18613 39611 18989
rect 39645 18613 39651 18989
rect 39605 18601 39651 18613
rect 39723 18989 39769 19001
rect 39723 18613 39729 18989
rect 39763 18613 39769 18989
rect 39723 18601 39769 18613
rect 39841 18989 39887 19001
rect 39841 18613 39847 18989
rect 39881 18613 39887 18989
rect 39841 18601 39887 18613
rect 39959 18989 40005 19001
rect 39959 18613 39965 18989
rect 39999 18613 40005 18989
rect 39959 18601 40005 18613
rect 40077 18989 40123 19001
rect 40077 18613 40083 18989
rect 40117 18613 40123 18989
rect 40077 18601 40123 18613
rect 40195 18989 40241 19001
rect 40195 18613 40201 18989
rect 40235 18613 40241 18989
rect 40195 18601 40241 18613
rect 40313 18989 40359 19001
rect 40440 18997 40611 19013
rect 40752 19059 41023 19087
rect 40752 18997 40787 19059
rect 40989 18997 41023 19059
rect 41107 19059 41377 19087
rect 41107 18997 41141 19059
rect 41343 18997 41377 19059
rect 40313 18613 40319 18989
rect 40353 18613 40359 18989
rect 40313 18601 40359 18613
rect 39611 18418 39645 18601
rect 39729 18560 39763 18601
rect 39965 18560 39999 18601
rect 39729 18531 39999 18560
rect 40083 18559 40117 18601
rect 40319 18559 40353 18601
rect 40083 18531 40353 18559
rect 40319 18483 40353 18531
rect 40290 18453 40353 18483
rect 39536 18364 39645 18418
rect 39718 18423 39818 18444
rect 39718 18369 39739 18423
rect 39804 18369 39818 18423
rect 39718 18364 39818 18369
rect 39536 18218 39570 18364
rect 39720 18349 39817 18364
rect 40290 18361 40325 18453
rect 39760 18282 39817 18349
rect 40098 18325 40325 18361
rect 40098 18291 40164 18325
rect 39654 18246 39923 18282
rect 40098 18257 40114 18291
rect 40148 18257 40164 18291
rect 40098 18251 40164 18257
rect 39654 18218 39687 18246
rect 39890 18218 39923 18246
rect 40290 18218 40325 18325
rect 39530 18206 39576 18218
rect 39530 18030 39536 18206
rect 39570 18030 39576 18206
rect 39530 18018 39576 18030
rect 39648 18206 39694 18218
rect 39648 18030 39654 18206
rect 39688 18030 39694 18206
rect 39648 18018 39694 18030
rect 39766 18206 39812 18218
rect 39766 18030 39772 18206
rect 39806 18030 39812 18206
rect 39766 18018 39812 18030
rect 39884 18206 39930 18218
rect 39884 18030 39890 18206
rect 39924 18151 39930 18206
rect 40049 18206 40095 18218
rect 40049 18151 40055 18206
rect 39924 18063 40055 18151
rect 39924 18030 39930 18063
rect 39884 18018 39930 18030
rect 40049 18030 40055 18063
rect 40089 18030 40095 18206
rect 40049 18018 40095 18030
rect 40167 18206 40213 18218
rect 40167 18030 40173 18206
rect 40207 18030 40213 18206
rect 40167 18018 40213 18030
rect 40285 18206 40331 18218
rect 40285 18030 40291 18206
rect 40325 18030 40331 18206
rect 40285 18018 40331 18030
rect 40403 18206 40449 18218
rect 40403 18030 40409 18206
rect 40443 18030 40449 18206
rect 40403 18018 40449 18030
rect 39537 17980 39570 18018
rect 39773 17980 39806 18018
rect 39537 17944 39806 17980
rect 40173 17979 40207 18018
rect 40409 17979 40443 18018
rect 40173 17943 40443 17979
rect 40277 17942 40443 17943
rect 40277 17863 40409 17942
rect 40267 17755 40277 17863
rect 40409 17755 40419 17863
rect 40549 17426 40611 18997
rect 40747 18985 40793 18997
rect 40747 18609 40753 18985
rect 40787 18609 40793 18985
rect 40747 18597 40793 18609
rect 40865 18985 40911 18997
rect 40865 18609 40871 18985
rect 40905 18609 40911 18985
rect 40865 18597 40911 18609
rect 40983 18985 41029 18997
rect 40983 18609 40989 18985
rect 41023 18609 41029 18985
rect 40983 18597 41029 18609
rect 41101 18985 41147 18997
rect 41101 18609 41107 18985
rect 41141 18609 41147 18985
rect 41101 18597 41147 18609
rect 41219 18985 41265 18997
rect 41219 18609 41225 18985
rect 41259 18609 41265 18985
rect 41219 18597 41265 18609
rect 41337 18985 41383 18997
rect 41337 18609 41343 18985
rect 41377 18609 41383 18985
rect 41337 18597 41383 18609
rect 41455 18985 41501 18997
rect 41550 18993 41560 19059
rect 41626 18993 41636 19059
rect 41455 18609 41461 18985
rect 41495 18609 41501 18985
rect 41455 18597 41501 18609
rect 40753 18414 40787 18597
rect 40871 18556 40905 18597
rect 41107 18556 41141 18597
rect 40871 18527 41141 18556
rect 41225 18555 41259 18597
rect 41461 18555 41495 18597
rect 41225 18527 41495 18555
rect 41461 18479 41495 18527
rect 41432 18449 41495 18479
rect 42485 18520 42552 19110
rect 43203 19103 43247 19211
rect 43379 19103 43423 19211
rect 46166 19198 46176 19261
rect 46164 19187 46176 19198
rect 43203 19061 43423 19103
rect 46163 19153 46176 19187
rect 46308 19153 46318 19261
rect 47313 19198 47323 19261
rect 47311 19187 47323 19198
rect 46998 19177 47054 19179
rect 46163 19115 46308 19153
rect 46163 19087 46204 19115
rect 46988 19111 46998 19177
rect 47054 19111 47064 19177
rect 47310 19153 47323 19187
rect 47455 19153 47465 19261
rect 49761 19207 49981 19227
rect 48128 19165 48184 19173
rect 48128 19157 49110 19165
rect 47310 19115 47455 19153
rect 48128 19123 48134 19157
rect 48168 19123 49110 19157
rect 42842 19031 43819 19061
rect 42842 18925 42876 19031
rect 43079 18925 43111 19031
rect 43315 18925 43347 19031
rect 43551 18925 43583 19031
rect 43787 18925 43819 19031
rect 46163 19059 46439 19087
rect 46163 18997 46203 19059
rect 46405 18997 46439 19059
rect 46523 19059 46793 19087
rect 47310 19083 47351 19115
rect 48128 19107 49110 19123
rect 48131 19106 49110 19107
rect 46523 18997 46557 19059
rect 46759 18997 46793 19059
rect 46998 19043 47169 19059
rect 46998 19009 47004 19043
rect 47038 19009 47169 19043
rect 46163 18985 46209 18997
rect 42718 18913 42764 18925
rect 42718 18737 42724 18913
rect 42758 18737 42764 18913
rect 42718 18725 42764 18737
rect 42836 18913 42882 18925
rect 42836 18737 42842 18913
rect 42876 18737 42882 18913
rect 42836 18725 42882 18737
rect 42954 18913 43000 18925
rect 42954 18737 42960 18913
rect 42994 18737 43000 18913
rect 42954 18725 43000 18737
rect 43072 18913 43118 18925
rect 43072 18737 43078 18913
rect 43112 18737 43118 18913
rect 43072 18725 43118 18737
rect 43190 18913 43236 18925
rect 43190 18737 43196 18913
rect 43230 18737 43236 18913
rect 43190 18725 43236 18737
rect 43308 18913 43354 18925
rect 43308 18737 43314 18913
rect 43348 18737 43354 18913
rect 43308 18725 43354 18737
rect 43426 18913 43472 18925
rect 43426 18737 43432 18913
rect 43466 18737 43472 18913
rect 43426 18725 43472 18737
rect 43544 18913 43590 18925
rect 43544 18737 43550 18913
rect 43584 18737 43590 18913
rect 43544 18725 43590 18737
rect 43662 18913 43708 18925
rect 43662 18737 43668 18913
rect 43702 18737 43708 18913
rect 43662 18725 43708 18737
rect 43780 18913 43826 18925
rect 43780 18737 43786 18913
rect 43820 18737 43826 18913
rect 43780 18725 43826 18737
rect 42724 18520 42759 18725
rect 43003 18677 43069 18684
rect 43003 18643 43019 18677
rect 43053 18643 43069 18677
rect 43003 18632 43069 18643
rect 43195 18632 43231 18725
rect 43003 18631 43231 18632
rect 43431 18631 43467 18725
rect 43667 18631 43703 18725
rect 43003 18602 43703 18631
rect 42485 18492 42759 18520
rect 43121 18601 43703 18602
rect 46163 18609 46169 18985
rect 46203 18609 46209 18985
rect 43121 18560 43187 18601
rect 43121 18526 43137 18560
rect 43171 18526 43187 18560
rect 43121 18519 43187 18526
rect 42485 18488 43113 18492
rect 43549 18488 43583 18601
rect 46163 18597 46209 18609
rect 46281 18985 46327 18997
rect 46281 18609 46287 18985
rect 46321 18609 46327 18985
rect 46281 18597 46327 18609
rect 46399 18985 46445 18997
rect 46399 18609 46405 18985
rect 46439 18609 46445 18985
rect 46399 18597 46445 18609
rect 46517 18985 46563 18997
rect 46517 18609 46523 18985
rect 46557 18609 46563 18985
rect 46517 18597 46563 18609
rect 46635 18985 46681 18997
rect 46635 18609 46641 18985
rect 46675 18609 46681 18985
rect 46635 18597 46681 18609
rect 46753 18985 46799 18997
rect 46753 18609 46759 18985
rect 46793 18609 46799 18985
rect 46753 18597 46799 18609
rect 46871 18985 46917 18997
rect 46998 18993 47169 19009
rect 47310 19055 47581 19083
rect 47310 18993 47345 19055
rect 47547 18993 47581 19055
rect 47665 19055 47935 19083
rect 47665 18993 47699 19055
rect 47901 18993 47935 19055
rect 46871 18609 46877 18985
rect 46911 18609 46917 18985
rect 46871 18597 46917 18609
rect 42485 18476 43118 18488
rect 42485 18463 43078 18476
rect 40678 18360 40787 18414
rect 40678 18214 40712 18360
rect 40851 18346 40861 18443
rect 40960 18346 40970 18443
rect 41432 18357 41467 18449
rect 40862 18345 40959 18346
rect 40902 18278 40959 18345
rect 41240 18321 41467 18357
rect 41240 18287 41306 18321
rect 40796 18242 41065 18278
rect 41240 18253 41256 18287
rect 41290 18253 41306 18287
rect 41240 18247 41306 18253
rect 40796 18214 40829 18242
rect 41032 18214 41065 18242
rect 41432 18214 41467 18321
rect 43072 18300 43078 18463
rect 43112 18300 43118 18476
rect 43072 18288 43118 18300
rect 43190 18476 43236 18488
rect 43190 18300 43196 18476
rect 43230 18300 43236 18476
rect 43190 18288 43236 18300
rect 43307 18476 43353 18488
rect 40672 18202 40718 18214
rect 40672 18026 40678 18202
rect 40712 18026 40718 18202
rect 40672 18014 40718 18026
rect 40790 18202 40836 18214
rect 40790 18026 40796 18202
rect 40830 18026 40836 18202
rect 40790 18014 40836 18026
rect 40908 18202 40954 18214
rect 40908 18026 40914 18202
rect 40948 18026 40954 18202
rect 40908 18014 40954 18026
rect 41026 18202 41072 18214
rect 41026 18026 41032 18202
rect 41066 18147 41072 18202
rect 41191 18202 41237 18214
rect 41191 18147 41197 18202
rect 41066 18059 41197 18147
rect 41066 18026 41072 18059
rect 41026 18014 41072 18026
rect 41191 18026 41197 18059
rect 41231 18026 41237 18202
rect 41191 18014 41237 18026
rect 41309 18202 41355 18214
rect 41309 18026 41315 18202
rect 41349 18026 41355 18202
rect 41309 18014 41355 18026
rect 41427 18202 41473 18214
rect 41427 18026 41433 18202
rect 41467 18026 41473 18202
rect 41427 18014 41473 18026
rect 41545 18202 41591 18214
rect 41545 18026 41551 18202
rect 41585 18026 41591 18202
rect 42991 18172 43099 18182
rect 43195 18172 43230 18288
rect 43099 18124 43230 18172
rect 43307 18124 43313 18476
rect 43099 18100 43313 18124
rect 43347 18100 43353 18476
rect 43099 18088 43353 18100
rect 43425 18476 43471 18488
rect 43425 18100 43431 18476
rect 43465 18100 43471 18476
rect 43425 18088 43471 18100
rect 43543 18476 43589 18488
rect 43543 18100 43549 18476
rect 43583 18100 43589 18476
rect 45099 18428 45198 18430
rect 45099 18353 45199 18428
rect 45267 18353 45277 18428
rect 46169 18414 46203 18597
rect 46287 18556 46321 18597
rect 46523 18556 46557 18597
rect 46287 18527 46557 18556
rect 46641 18555 46675 18597
rect 46877 18555 46911 18597
rect 46641 18527 46911 18555
rect 46877 18479 46911 18527
rect 46848 18449 46911 18479
rect 46094 18360 46203 18414
rect 46276 18419 46376 18440
rect 46276 18365 46297 18419
rect 46362 18365 46376 18419
rect 46276 18360 46376 18365
rect 45099 18352 45250 18353
rect 43543 18088 43589 18100
rect 44472 18132 44761 18151
rect 43099 18084 43347 18088
rect 43099 18040 43173 18084
rect 44472 18083 44513 18132
rect 43711 18056 44513 18083
rect 43356 18050 43422 18056
rect 42991 18030 43099 18040
rect 41545 18014 41591 18026
rect 43356 18016 43372 18050
rect 43406 18016 43422 18050
rect 40679 17976 40712 18014
rect 40915 17976 40948 18014
rect 40679 17940 40948 17976
rect 41315 17975 41349 18014
rect 41551 17975 41585 18014
rect 41315 17940 41585 17975
rect 41315 17939 41551 17940
rect 41419 17865 41551 17939
rect 43356 17920 43422 18016
rect 43474 18050 44513 18056
rect 43474 18016 43490 18050
rect 43524 18016 44513 18050
rect 43474 18000 44513 18016
rect 43711 17996 44513 18000
rect 44737 17996 44761 18132
rect 43711 17984 44761 17996
rect 43774 17983 44761 17984
rect 44239 17979 44761 17983
rect 43710 17920 44176 17942
rect 43356 17872 44176 17920
rect 41409 17757 41419 17865
rect 41551 17757 41561 17865
rect 43710 17841 44176 17872
rect 44071 17585 44176 17841
rect 40548 17409 40611 17426
rect 43189 17561 43409 17581
rect 43189 17453 43233 17561
rect 43365 17453 43409 17561
rect 43991 17479 44001 17585
rect 44113 17479 44176 17585
rect 44027 17468 44176 17479
rect 43189 17411 43409 17453
rect 40548 17405 40686 17409
rect 40548 17371 42518 17405
rect 42828 17381 43805 17411
rect 40548 17342 42520 17371
rect 40548 17340 40686 17342
rect 42474 17326 42520 17342
rect 39512 17110 39522 17218
rect 39654 17110 39664 17218
rect 41410 17110 41420 17218
rect 41552 17110 41562 17218
rect 39522 17070 39654 17110
rect 41420 17070 41552 17110
rect 39522 17004 39655 17070
rect 41420 17004 41553 17070
rect 38853 16961 40326 17004
rect 38853 16658 38887 16961
rect 39218 16858 39252 16961
rect 39454 16858 39488 16961
rect 39690 16858 39724 16961
rect 39926 16858 39960 16961
rect 39212 16846 39258 16858
rect 38729 16646 38775 16658
rect 38729 16470 38735 16646
rect 38769 16470 38775 16646
rect 38729 16458 38775 16470
rect 38847 16646 38893 16658
rect 38847 16470 38853 16646
rect 38887 16470 38893 16646
rect 38847 16458 38893 16470
rect 38965 16646 39011 16658
rect 38965 16470 38971 16646
rect 39005 16470 39011 16646
rect 38965 16458 39011 16470
rect 39083 16646 39129 16658
rect 39212 16646 39218 16846
rect 39083 16470 39089 16646
rect 39123 16470 39218 16646
rect 39252 16470 39258 16846
rect 39083 16458 39129 16470
rect 39212 16458 39258 16470
rect 39330 16846 39376 16858
rect 39330 16470 39336 16846
rect 39370 16470 39376 16846
rect 39330 16458 39376 16470
rect 39448 16846 39494 16858
rect 39448 16470 39454 16846
rect 39488 16470 39494 16846
rect 39448 16458 39494 16470
rect 39566 16846 39612 16858
rect 39566 16470 39572 16846
rect 39606 16470 39612 16846
rect 39566 16458 39612 16470
rect 39684 16846 39730 16858
rect 39684 16470 39690 16846
rect 39724 16470 39730 16846
rect 39684 16458 39730 16470
rect 39802 16846 39848 16858
rect 39802 16470 39808 16846
rect 39842 16470 39848 16846
rect 39802 16458 39848 16470
rect 39920 16846 39966 16858
rect 39920 16470 39926 16846
rect 39960 16646 39966 16846
rect 40292 16658 40326 16961
rect 40751 16961 42224 17004
rect 40751 16658 40785 16961
rect 41116 16858 41150 16961
rect 41352 16858 41386 16961
rect 41588 16858 41622 16961
rect 41824 16858 41858 16961
rect 41110 16846 41156 16858
rect 40050 16646 40096 16658
rect 39960 16470 40056 16646
rect 40090 16470 40096 16646
rect 39920 16458 39966 16470
rect 40050 16458 40096 16470
rect 40168 16646 40214 16658
rect 40168 16470 40174 16646
rect 40208 16470 40214 16646
rect 40168 16458 40214 16470
rect 40286 16646 40332 16658
rect 40286 16470 40292 16646
rect 40326 16470 40332 16646
rect 40286 16458 40332 16470
rect 40404 16646 40450 16658
rect 40404 16470 40410 16646
rect 40444 16470 40450 16646
rect 40404 16458 40450 16470
rect 40627 16646 40673 16658
rect 40627 16470 40633 16646
rect 40667 16470 40673 16646
rect 40627 16458 40673 16470
rect 40745 16646 40791 16658
rect 40745 16470 40751 16646
rect 40785 16470 40791 16646
rect 40745 16458 40791 16470
rect 40863 16646 40909 16658
rect 40863 16470 40869 16646
rect 40903 16470 40909 16646
rect 40863 16458 40909 16470
rect 40981 16646 41027 16658
rect 41110 16646 41116 16846
rect 40981 16470 40987 16646
rect 41021 16470 41116 16646
rect 41150 16470 41156 16846
rect 40981 16458 41027 16470
rect 41110 16458 41156 16470
rect 41228 16846 41274 16858
rect 41228 16470 41234 16846
rect 41268 16470 41274 16846
rect 41228 16458 41274 16470
rect 41346 16846 41392 16858
rect 41346 16470 41352 16846
rect 41386 16470 41392 16846
rect 41346 16458 41392 16470
rect 41464 16846 41510 16858
rect 41464 16470 41470 16846
rect 41504 16470 41510 16846
rect 41464 16458 41510 16470
rect 41582 16846 41628 16858
rect 41582 16470 41588 16846
rect 41622 16470 41628 16846
rect 41582 16458 41628 16470
rect 41700 16846 41746 16858
rect 41700 16470 41706 16846
rect 41740 16470 41746 16846
rect 41700 16458 41746 16470
rect 41818 16846 41864 16858
rect 41818 16470 41824 16846
rect 41858 16646 41864 16846
rect 42190 16658 42224 16961
rect 42474 16874 42521 17326
rect 42828 17275 42862 17381
rect 43065 17275 43097 17381
rect 43301 17275 43333 17381
rect 43537 17275 43569 17381
rect 43773 17275 43805 17381
rect 42704 17263 42750 17275
rect 42704 17087 42710 17263
rect 42744 17087 42750 17263
rect 42704 17075 42750 17087
rect 42822 17263 42868 17275
rect 42822 17087 42828 17263
rect 42862 17087 42868 17263
rect 42822 17075 42868 17087
rect 42940 17263 42986 17275
rect 42940 17087 42946 17263
rect 42980 17087 42986 17263
rect 42940 17075 42986 17087
rect 43058 17263 43104 17275
rect 43058 17087 43064 17263
rect 43098 17087 43104 17263
rect 43058 17075 43104 17087
rect 43176 17263 43222 17275
rect 43176 17087 43182 17263
rect 43216 17087 43222 17263
rect 43176 17075 43222 17087
rect 43294 17263 43340 17275
rect 43294 17087 43300 17263
rect 43334 17087 43340 17263
rect 43294 17075 43340 17087
rect 43412 17263 43458 17275
rect 43412 17087 43418 17263
rect 43452 17087 43458 17263
rect 43412 17075 43458 17087
rect 43530 17263 43576 17275
rect 43530 17087 43536 17263
rect 43570 17087 43576 17263
rect 43530 17075 43576 17087
rect 43648 17263 43694 17275
rect 43648 17087 43654 17263
rect 43688 17087 43694 17263
rect 43648 17075 43694 17087
rect 43766 17263 43812 17275
rect 43766 17087 43772 17263
rect 43806 17087 43812 17263
rect 43766 17075 43812 17087
rect 42475 16858 42521 16874
rect 42475 16857 42556 16858
rect 42710 16857 42745 17075
rect 42989 17027 43055 17034
rect 42989 16993 43005 17027
rect 43039 16993 43055 17027
rect 42989 16982 43055 16993
rect 43181 16982 43217 17075
rect 42989 16981 43217 16982
rect 43417 16981 43453 17075
rect 43653 16981 43689 17075
rect 42989 16952 43689 16981
rect 43107 16951 43689 16952
rect 43107 16910 43173 16951
rect 43107 16876 43123 16910
rect 43157 16876 43173 16910
rect 43107 16869 43173 16876
rect 42475 16842 42745 16857
rect 42475 16838 43099 16842
rect 43535 16838 43569 16951
rect 42475 16826 43104 16838
rect 42475 16814 43064 16826
rect 42475 16812 42556 16814
rect 42822 16813 43064 16814
rect 41948 16646 41994 16658
rect 41858 16470 41954 16646
rect 41988 16470 41994 16646
rect 41818 16458 41864 16470
rect 41948 16458 41994 16470
rect 42066 16646 42112 16658
rect 42066 16470 42072 16646
rect 42106 16470 42112 16646
rect 42066 16458 42112 16470
rect 42184 16646 42230 16658
rect 42184 16470 42190 16646
rect 42224 16470 42230 16646
rect 42184 16458 42230 16470
rect 42302 16646 42348 16658
rect 42302 16470 42308 16646
rect 42342 16470 42348 16646
rect 43058 16650 43064 16813
rect 43098 16650 43104 16826
rect 43058 16638 43104 16650
rect 43176 16826 43222 16838
rect 43176 16650 43182 16826
rect 43216 16650 43222 16826
rect 43176 16638 43222 16650
rect 43293 16826 43339 16838
rect 42302 16458 42348 16470
rect 42977 16522 43085 16532
rect 43181 16522 43216 16638
rect 38735 16424 38769 16458
rect 38971 16424 39005 16458
rect 38735 16389 39005 16424
rect 39572 16424 39606 16458
rect 39808 16424 39842 16458
rect 40410 16424 40444 16458
rect 39572 16389 39842 16424
rect 40285 16389 40444 16424
rect 40633 16424 40667 16458
rect 40869 16424 40903 16458
rect 40633 16389 40903 16424
rect 41470 16424 41504 16458
rect 41706 16424 41740 16458
rect 42308 16424 42342 16458
rect 41470 16389 41740 16424
rect 42183 16389 42342 16424
rect 43085 16474 43216 16522
rect 43293 16474 43299 16826
rect 43085 16450 43299 16474
rect 43333 16450 43339 16826
rect 43085 16438 43339 16450
rect 43411 16826 43457 16838
rect 43411 16450 43417 16826
rect 43451 16450 43457 16826
rect 43411 16438 43457 16450
rect 43529 16826 43575 16838
rect 43529 16450 43535 16826
rect 43569 16450 43575 16826
rect 43529 16438 43575 16450
rect 43085 16434 43333 16438
rect 43702 16434 43712 16466
rect 43085 16390 43159 16434
rect 43697 16406 43712 16434
rect 43342 16400 43408 16406
rect 38721 16211 38788 16235
rect 38721 16177 38737 16211
rect 38771 16177 38788 16211
rect 38505 15754 38660 15762
rect 38504 15748 38660 15754
rect 38504 15650 38516 15748
rect 38648 15650 38660 15748
rect 38504 13652 38660 15650
rect 38721 14794 38788 16177
rect 38869 15606 38903 16389
rect 39572 16327 39606 16389
rect 39275 16289 40017 16327
rect 39275 16165 39309 16289
rect 39511 16165 39545 16289
rect 39747 16165 39781 16289
rect 39983 16165 40017 16289
rect 39269 16153 39315 16165
rect 39269 15777 39275 16153
rect 39309 15777 39315 16153
rect 39269 15765 39315 15777
rect 39387 16153 39433 16165
rect 39387 15777 39393 16153
rect 39427 15777 39433 16153
rect 39387 15765 39433 15777
rect 39505 16153 39551 16165
rect 39505 15777 39511 16153
rect 39545 15777 39551 16153
rect 39505 15765 39551 15777
rect 39623 16153 39669 16165
rect 39623 15777 39629 16153
rect 39663 15777 39669 16153
rect 39623 15765 39669 15777
rect 39741 16153 39787 16165
rect 39741 15777 39747 16153
rect 39781 15777 39787 16153
rect 39741 15765 39787 15777
rect 39859 16153 39905 16165
rect 39859 15777 39865 16153
rect 39899 15777 39905 16153
rect 39859 15765 39905 15777
rect 39977 16153 40023 16165
rect 39977 15777 39983 16153
rect 40017 15777 40023 16153
rect 39977 15765 40023 15777
rect 38869 15605 39176 15606
rect 39222 15605 39291 15606
rect 40285 15605 40319 16389
rect 38869 15601 39291 15605
rect 38869 15590 39358 15601
rect 40003 15600 40319 15605
rect 38869 15562 39307 15590
rect 38869 15561 39176 15562
rect 38869 15433 38903 15561
rect 39291 15556 39307 15562
rect 39341 15556 39358 15590
rect 39291 15550 39358 15556
rect 39936 15589 40319 15600
rect 39936 15555 39953 15589
rect 39987 15562 40319 15589
rect 39987 15555 40003 15562
rect 39936 15549 40003 15555
rect 39009 15521 39065 15533
rect 40122 15522 40178 15534
rect 40122 15521 40138 15522
rect 39009 15487 39015 15521
rect 39049 15506 39619 15521
rect 39049 15487 39569 15506
rect 39009 15472 39569 15487
rect 39603 15472 39619 15506
rect 39009 15471 39065 15472
rect 39552 15462 39619 15472
rect 39671 15505 40138 15521
rect 39671 15471 39687 15505
rect 39721 15488 40138 15505
rect 40172 15488 40178 15522
rect 39721 15472 40178 15488
rect 39721 15471 39737 15472
rect 39671 15464 39737 15471
rect 40285 15433 40319 15562
rect 40767 15606 40801 16389
rect 41470 16327 41504 16389
rect 41173 16289 41915 16327
rect 40834 16182 40844 16248
rect 40907 16182 40917 16248
rect 41173 16165 41207 16289
rect 41409 16165 41443 16289
rect 41645 16165 41679 16289
rect 41881 16165 41915 16289
rect 41167 16153 41213 16165
rect 41167 15777 41173 16153
rect 41207 15777 41213 16153
rect 41167 15765 41213 15777
rect 41285 16153 41331 16165
rect 41285 15777 41291 16153
rect 41325 15777 41331 16153
rect 41285 15765 41331 15777
rect 41403 16153 41449 16165
rect 41403 15777 41409 16153
rect 41443 15777 41449 16153
rect 41403 15765 41449 15777
rect 41521 16153 41567 16165
rect 41521 15777 41527 16153
rect 41561 15777 41567 16153
rect 41521 15765 41567 15777
rect 41639 16153 41685 16165
rect 41639 15777 41645 16153
rect 41679 15777 41685 16153
rect 41639 15765 41685 15777
rect 41757 16153 41803 16165
rect 41757 15777 41763 16153
rect 41797 15777 41803 16153
rect 41757 15765 41803 15777
rect 41875 16153 41921 16165
rect 41875 15777 41881 16153
rect 41915 15777 41921 16153
rect 41875 15765 41921 15777
rect 40767 15605 41074 15606
rect 42183 15605 42217 16389
rect 42977 16380 43085 16390
rect 43342 16366 43358 16400
rect 43392 16366 43408 16400
rect 43342 16270 43408 16366
rect 43460 16400 43712 16406
rect 43460 16366 43476 16400
rect 43510 16366 43712 16400
rect 43460 16350 43712 16366
rect 43697 16348 43712 16350
rect 43830 16348 43840 16466
rect 43697 16334 43797 16348
rect 43697 16291 43797 16292
rect 44071 16291 44176 17468
rect 43697 16270 44176 16291
rect 43342 16222 44176 16270
rect 43697 16193 44176 16222
rect 43697 16192 43797 16193
rect 44071 16191 44176 16193
rect 44239 16085 44332 17979
rect 44472 17978 44761 17979
rect 44455 17571 44622 17618
rect 44455 17568 44496 17571
rect 44455 17555 44495 17568
rect 44453 17462 44495 17555
rect 44607 17462 44622 17571
rect 44453 17451 44622 17462
rect 44455 17450 44622 17451
rect 45099 16618 45198 18352
rect 46094 18214 46128 18360
rect 46278 18345 46375 18360
rect 46848 18357 46883 18449
rect 46318 18278 46375 18345
rect 46656 18321 46883 18357
rect 46656 18287 46722 18321
rect 46212 18242 46481 18278
rect 46656 18253 46672 18287
rect 46706 18253 46722 18287
rect 46656 18247 46722 18253
rect 46212 18214 46245 18242
rect 46448 18214 46481 18242
rect 46848 18214 46883 18321
rect 46088 18202 46134 18214
rect 46088 18026 46094 18202
rect 46128 18026 46134 18202
rect 46088 18014 46134 18026
rect 46206 18202 46252 18214
rect 46206 18026 46212 18202
rect 46246 18026 46252 18202
rect 46206 18014 46252 18026
rect 46324 18202 46370 18214
rect 46324 18026 46330 18202
rect 46364 18026 46370 18202
rect 46324 18014 46370 18026
rect 46442 18202 46488 18214
rect 46442 18026 46448 18202
rect 46482 18147 46488 18202
rect 46607 18202 46653 18214
rect 46607 18147 46613 18202
rect 46482 18059 46613 18147
rect 46482 18026 46488 18059
rect 46442 18014 46488 18026
rect 46607 18026 46613 18059
rect 46647 18026 46653 18202
rect 46607 18014 46653 18026
rect 46725 18202 46771 18214
rect 46725 18026 46731 18202
rect 46765 18026 46771 18202
rect 46725 18014 46771 18026
rect 46843 18202 46889 18214
rect 46843 18026 46849 18202
rect 46883 18026 46889 18202
rect 46843 18014 46889 18026
rect 46961 18202 47007 18214
rect 46961 18026 46967 18202
rect 47001 18026 47007 18202
rect 46961 18014 47007 18026
rect 46095 17976 46128 18014
rect 46331 17976 46364 18014
rect 46095 17940 46364 17976
rect 46731 17975 46765 18014
rect 46967 17975 47001 18014
rect 46731 17939 47001 17975
rect 46835 17938 47001 17939
rect 46835 17859 46967 17938
rect 46825 17751 46835 17859
rect 46967 17751 46977 17859
rect 47107 17422 47169 18993
rect 47305 18981 47351 18993
rect 47305 18605 47311 18981
rect 47345 18605 47351 18981
rect 47305 18593 47351 18605
rect 47423 18981 47469 18993
rect 47423 18605 47429 18981
rect 47463 18605 47469 18981
rect 47423 18593 47469 18605
rect 47541 18981 47587 18993
rect 47541 18605 47547 18981
rect 47581 18605 47587 18981
rect 47541 18593 47587 18605
rect 47659 18981 47705 18993
rect 47659 18605 47665 18981
rect 47699 18605 47705 18981
rect 47659 18593 47705 18605
rect 47777 18981 47823 18993
rect 47777 18605 47783 18981
rect 47817 18605 47823 18981
rect 47777 18593 47823 18605
rect 47895 18981 47941 18993
rect 47895 18605 47901 18981
rect 47935 18605 47941 18981
rect 47895 18593 47941 18605
rect 48013 18981 48059 18993
rect 48108 18989 48118 19055
rect 48184 18989 48194 19055
rect 48013 18605 48019 18981
rect 48053 18605 48059 18981
rect 48013 18593 48059 18605
rect 47311 18410 47345 18593
rect 47429 18552 47463 18593
rect 47665 18552 47699 18593
rect 47429 18523 47699 18552
rect 47783 18551 47817 18593
rect 48019 18551 48053 18593
rect 47783 18523 48053 18551
rect 48019 18475 48053 18523
rect 47990 18445 48053 18475
rect 49043 18516 49110 19106
rect 49761 19099 49805 19207
rect 49937 19099 49981 19207
rect 52700 19203 52710 19266
rect 52698 19192 52710 19203
rect 49761 19057 49981 19099
rect 52697 19158 52710 19192
rect 52842 19158 52852 19266
rect 53847 19203 53857 19266
rect 53845 19192 53857 19203
rect 53532 19182 53588 19184
rect 52697 19120 52842 19158
rect 52697 19092 52738 19120
rect 53522 19116 53532 19182
rect 53588 19116 53598 19182
rect 53844 19158 53857 19192
rect 53989 19158 53999 19266
rect 56295 19212 56515 19232
rect 54662 19170 54718 19178
rect 54662 19162 55644 19170
rect 53844 19120 53989 19158
rect 54662 19128 54668 19162
rect 54702 19128 55644 19162
rect 52697 19064 52973 19092
rect 49400 19027 50377 19057
rect 49400 18921 49434 19027
rect 49637 18921 49669 19027
rect 49873 18921 49905 19027
rect 50109 18921 50141 19027
rect 50345 18921 50377 19027
rect 52697 19002 52737 19064
rect 52939 19002 52973 19064
rect 53057 19064 53327 19092
rect 53844 19088 53885 19120
rect 54662 19112 55644 19128
rect 54665 19111 55644 19112
rect 53057 19002 53091 19064
rect 53293 19002 53327 19064
rect 53532 19048 53703 19064
rect 53532 19014 53538 19048
rect 53572 19014 53703 19048
rect 52697 18990 52743 19002
rect 49276 18909 49322 18921
rect 49276 18733 49282 18909
rect 49316 18733 49322 18909
rect 49276 18721 49322 18733
rect 49394 18909 49440 18921
rect 49394 18733 49400 18909
rect 49434 18733 49440 18909
rect 49394 18721 49440 18733
rect 49512 18909 49558 18921
rect 49512 18733 49518 18909
rect 49552 18733 49558 18909
rect 49512 18721 49558 18733
rect 49630 18909 49676 18921
rect 49630 18733 49636 18909
rect 49670 18733 49676 18909
rect 49630 18721 49676 18733
rect 49748 18909 49794 18921
rect 49748 18733 49754 18909
rect 49788 18733 49794 18909
rect 49748 18721 49794 18733
rect 49866 18909 49912 18921
rect 49866 18733 49872 18909
rect 49906 18733 49912 18909
rect 49866 18721 49912 18733
rect 49984 18909 50030 18921
rect 49984 18733 49990 18909
rect 50024 18733 50030 18909
rect 49984 18721 50030 18733
rect 50102 18909 50148 18921
rect 50102 18733 50108 18909
rect 50142 18733 50148 18909
rect 50102 18721 50148 18733
rect 50220 18909 50266 18921
rect 50220 18733 50226 18909
rect 50260 18733 50266 18909
rect 50220 18721 50266 18733
rect 50338 18909 50384 18921
rect 50338 18733 50344 18909
rect 50378 18733 50384 18909
rect 50338 18721 50384 18733
rect 49282 18516 49317 18721
rect 49561 18673 49627 18680
rect 49561 18639 49577 18673
rect 49611 18639 49627 18673
rect 49561 18628 49627 18639
rect 49753 18628 49789 18721
rect 49561 18627 49789 18628
rect 49989 18627 50025 18721
rect 50225 18627 50261 18721
rect 49561 18598 50261 18627
rect 52697 18614 52703 18990
rect 52737 18614 52743 18990
rect 52697 18602 52743 18614
rect 52815 18990 52861 19002
rect 52815 18614 52821 18990
rect 52855 18614 52861 18990
rect 52815 18602 52861 18614
rect 52933 18990 52979 19002
rect 52933 18614 52939 18990
rect 52973 18614 52979 18990
rect 52933 18602 52979 18614
rect 53051 18990 53097 19002
rect 53051 18614 53057 18990
rect 53091 18614 53097 18990
rect 53051 18602 53097 18614
rect 53169 18990 53215 19002
rect 53169 18614 53175 18990
rect 53209 18614 53215 18990
rect 53169 18602 53215 18614
rect 53287 18990 53333 19002
rect 53287 18614 53293 18990
rect 53327 18614 53333 18990
rect 53287 18602 53333 18614
rect 53405 18990 53451 19002
rect 53532 18998 53703 19014
rect 53844 19060 54115 19088
rect 53844 18998 53879 19060
rect 54081 18998 54115 19060
rect 54199 19060 54469 19088
rect 54199 18998 54233 19060
rect 54435 18998 54469 19060
rect 53405 18614 53411 18990
rect 53445 18614 53451 18990
rect 53405 18602 53451 18614
rect 49043 18488 49317 18516
rect 49679 18597 50261 18598
rect 49679 18556 49745 18597
rect 49679 18522 49695 18556
rect 49729 18522 49745 18556
rect 49679 18515 49745 18522
rect 49043 18484 49671 18488
rect 50107 18484 50141 18597
rect 49043 18472 49676 18484
rect 49043 18459 49636 18472
rect 47236 18356 47345 18410
rect 47236 18210 47270 18356
rect 47409 18342 47419 18439
rect 47518 18342 47528 18439
rect 47990 18353 48025 18445
rect 47420 18341 47517 18342
rect 47460 18274 47517 18341
rect 47798 18317 48025 18353
rect 47798 18283 47864 18317
rect 47354 18238 47623 18274
rect 47798 18249 47814 18283
rect 47848 18249 47864 18283
rect 47798 18243 47864 18249
rect 47354 18210 47387 18238
rect 47590 18210 47623 18238
rect 47990 18210 48025 18317
rect 49630 18296 49636 18459
rect 49670 18296 49676 18472
rect 49630 18284 49676 18296
rect 49748 18472 49794 18484
rect 49748 18296 49754 18472
rect 49788 18296 49794 18472
rect 49748 18284 49794 18296
rect 49865 18472 49911 18484
rect 47230 18198 47276 18210
rect 47230 18022 47236 18198
rect 47270 18022 47276 18198
rect 47230 18010 47276 18022
rect 47348 18198 47394 18210
rect 47348 18022 47354 18198
rect 47388 18022 47394 18198
rect 47348 18010 47394 18022
rect 47466 18198 47512 18210
rect 47466 18022 47472 18198
rect 47506 18022 47512 18198
rect 47466 18010 47512 18022
rect 47584 18198 47630 18210
rect 47584 18022 47590 18198
rect 47624 18143 47630 18198
rect 47749 18198 47795 18210
rect 47749 18143 47755 18198
rect 47624 18055 47755 18143
rect 47624 18022 47630 18055
rect 47584 18010 47630 18022
rect 47749 18022 47755 18055
rect 47789 18022 47795 18198
rect 47749 18010 47795 18022
rect 47867 18198 47913 18210
rect 47867 18022 47873 18198
rect 47907 18022 47913 18198
rect 47867 18010 47913 18022
rect 47985 18198 48031 18210
rect 47985 18022 47991 18198
rect 48025 18022 48031 18198
rect 47985 18010 48031 18022
rect 48103 18198 48149 18210
rect 48103 18022 48109 18198
rect 48143 18022 48149 18198
rect 49549 18168 49657 18178
rect 49753 18168 49788 18284
rect 49657 18120 49788 18168
rect 49865 18120 49871 18472
rect 49657 18096 49871 18120
rect 49905 18096 49911 18472
rect 49657 18084 49911 18096
rect 49983 18472 50029 18484
rect 49983 18096 49989 18472
rect 50023 18096 50029 18472
rect 49983 18084 50029 18096
rect 50101 18472 50147 18484
rect 50101 18096 50107 18472
rect 50141 18096 50147 18472
rect 51633 18416 51733 18433
rect 51631 18358 51733 18416
rect 51801 18358 51811 18433
rect 52703 18419 52737 18602
rect 52821 18561 52855 18602
rect 53057 18561 53091 18602
rect 52821 18532 53091 18561
rect 53175 18560 53209 18602
rect 53411 18560 53445 18602
rect 53175 18532 53445 18560
rect 53411 18484 53445 18532
rect 53382 18454 53445 18484
rect 52628 18365 52737 18419
rect 52810 18424 52910 18445
rect 52810 18370 52831 18424
rect 52896 18370 52910 18424
rect 52810 18365 52910 18370
rect 51631 18357 51784 18358
rect 50101 18084 50147 18096
rect 51030 18146 51319 18158
rect 49657 18080 49905 18084
rect 49657 18036 49731 18080
rect 51030 18079 51056 18146
rect 50269 18052 51056 18079
rect 49914 18046 49980 18052
rect 49549 18026 49657 18036
rect 48103 18010 48149 18022
rect 49914 18012 49930 18046
rect 49964 18012 49980 18046
rect 47237 17972 47270 18010
rect 47473 17972 47506 18010
rect 47237 17936 47506 17972
rect 47873 17971 47907 18010
rect 48109 17971 48143 18010
rect 47873 17936 48143 17971
rect 47873 17935 48109 17936
rect 47977 17861 48109 17935
rect 49914 17916 49980 18012
rect 50032 18046 51056 18052
rect 50032 18012 50048 18046
rect 50082 18012 51056 18046
rect 50032 17996 51056 18012
rect 50269 17990 51056 17996
rect 51306 17990 51319 18146
rect 50269 17980 51319 17990
rect 50332 17979 51319 17980
rect 50797 17975 51319 17979
rect 50268 17916 50734 17938
rect 49914 17868 50734 17916
rect 47967 17753 47977 17861
rect 48109 17753 48119 17861
rect 50268 17837 50734 17868
rect 50629 17581 50734 17837
rect 47106 17405 47169 17422
rect 49747 17557 49967 17577
rect 49747 17449 49791 17557
rect 49923 17449 49967 17557
rect 50549 17475 50559 17581
rect 50671 17475 50734 17581
rect 50585 17464 50734 17475
rect 49747 17407 49967 17449
rect 47106 17401 47244 17405
rect 47106 17367 49076 17401
rect 49386 17377 50363 17407
rect 47106 17338 49078 17367
rect 47106 17336 47244 17338
rect 49032 17322 49078 17338
rect 46070 17106 46080 17214
rect 46212 17106 46222 17214
rect 47968 17106 47978 17214
rect 48110 17106 48120 17214
rect 46080 17066 46212 17106
rect 47978 17066 48110 17106
rect 46080 17000 46213 17066
rect 47978 17000 48111 17066
rect 45411 16957 46884 17000
rect 45411 16654 45445 16957
rect 45776 16854 45810 16957
rect 46012 16854 46046 16957
rect 46248 16854 46282 16957
rect 46484 16854 46518 16957
rect 45770 16842 45816 16854
rect 44456 16515 45198 16618
rect 45287 16642 45333 16654
rect 44456 16456 44744 16515
rect 44456 16454 44496 16456
rect 44456 16443 44490 16454
rect 44455 16348 44490 16443
rect 44608 16350 44744 16456
rect 45287 16466 45293 16642
rect 45327 16466 45333 16642
rect 45287 16454 45333 16466
rect 45405 16642 45451 16654
rect 45405 16466 45411 16642
rect 45445 16466 45451 16642
rect 45405 16454 45451 16466
rect 45523 16642 45569 16654
rect 45523 16466 45529 16642
rect 45563 16466 45569 16642
rect 45523 16454 45569 16466
rect 45641 16642 45687 16654
rect 45770 16642 45776 16842
rect 45641 16466 45647 16642
rect 45681 16466 45776 16642
rect 45810 16466 45816 16842
rect 45641 16454 45687 16466
rect 45770 16454 45816 16466
rect 45888 16842 45934 16854
rect 45888 16466 45894 16842
rect 45928 16466 45934 16842
rect 45888 16454 45934 16466
rect 46006 16842 46052 16854
rect 46006 16466 46012 16842
rect 46046 16466 46052 16842
rect 46006 16454 46052 16466
rect 46124 16842 46170 16854
rect 46124 16466 46130 16842
rect 46164 16466 46170 16842
rect 46124 16454 46170 16466
rect 46242 16842 46288 16854
rect 46242 16466 46248 16842
rect 46282 16466 46288 16842
rect 46242 16454 46288 16466
rect 46360 16842 46406 16854
rect 46360 16466 46366 16842
rect 46400 16466 46406 16842
rect 46360 16454 46406 16466
rect 46478 16842 46524 16854
rect 46478 16466 46484 16842
rect 46518 16642 46524 16842
rect 46850 16654 46884 16957
rect 47309 16957 48782 17000
rect 47309 16654 47343 16957
rect 47674 16854 47708 16957
rect 47910 16854 47944 16957
rect 48146 16854 48180 16957
rect 48382 16854 48416 16957
rect 47668 16842 47714 16854
rect 46608 16642 46654 16654
rect 46518 16466 46614 16642
rect 46648 16466 46654 16642
rect 46478 16454 46524 16466
rect 46608 16454 46654 16466
rect 46726 16642 46772 16654
rect 46726 16466 46732 16642
rect 46766 16466 46772 16642
rect 46726 16454 46772 16466
rect 46844 16642 46890 16654
rect 46844 16466 46850 16642
rect 46884 16466 46890 16642
rect 46844 16454 46890 16466
rect 46962 16642 47008 16654
rect 46962 16466 46968 16642
rect 47002 16466 47008 16642
rect 46962 16454 47008 16466
rect 47185 16642 47231 16654
rect 47185 16466 47191 16642
rect 47225 16466 47231 16642
rect 47185 16454 47231 16466
rect 47303 16642 47349 16654
rect 47303 16466 47309 16642
rect 47343 16466 47349 16642
rect 47303 16454 47349 16466
rect 47421 16642 47467 16654
rect 47421 16466 47427 16642
rect 47461 16466 47467 16642
rect 47421 16454 47467 16466
rect 47539 16642 47585 16654
rect 47668 16642 47674 16842
rect 47539 16466 47545 16642
rect 47579 16466 47674 16642
rect 47708 16466 47714 16842
rect 47539 16454 47585 16466
rect 47668 16454 47714 16466
rect 47786 16842 47832 16854
rect 47786 16466 47792 16842
rect 47826 16466 47832 16842
rect 47786 16454 47832 16466
rect 47904 16842 47950 16854
rect 47904 16466 47910 16842
rect 47944 16466 47950 16842
rect 47904 16454 47950 16466
rect 48022 16842 48068 16854
rect 48022 16466 48028 16842
rect 48062 16466 48068 16842
rect 48022 16454 48068 16466
rect 48140 16842 48186 16854
rect 48140 16466 48146 16842
rect 48180 16466 48186 16842
rect 48140 16454 48186 16466
rect 48258 16842 48304 16854
rect 48258 16466 48264 16842
rect 48298 16466 48304 16842
rect 48258 16454 48304 16466
rect 48376 16842 48422 16854
rect 48376 16466 48382 16842
rect 48416 16642 48422 16842
rect 48748 16654 48782 16957
rect 49032 16870 49079 17322
rect 49386 17271 49420 17377
rect 49623 17271 49655 17377
rect 49859 17271 49891 17377
rect 50095 17271 50127 17377
rect 50331 17271 50363 17377
rect 49262 17259 49308 17271
rect 49262 17083 49268 17259
rect 49302 17083 49308 17259
rect 49262 17071 49308 17083
rect 49380 17259 49426 17271
rect 49380 17083 49386 17259
rect 49420 17083 49426 17259
rect 49380 17071 49426 17083
rect 49498 17259 49544 17271
rect 49498 17083 49504 17259
rect 49538 17083 49544 17259
rect 49498 17071 49544 17083
rect 49616 17259 49662 17271
rect 49616 17083 49622 17259
rect 49656 17083 49662 17259
rect 49616 17071 49662 17083
rect 49734 17259 49780 17271
rect 49734 17083 49740 17259
rect 49774 17083 49780 17259
rect 49734 17071 49780 17083
rect 49852 17259 49898 17271
rect 49852 17083 49858 17259
rect 49892 17083 49898 17259
rect 49852 17071 49898 17083
rect 49970 17259 50016 17271
rect 49970 17083 49976 17259
rect 50010 17083 50016 17259
rect 49970 17071 50016 17083
rect 50088 17259 50134 17271
rect 50088 17083 50094 17259
rect 50128 17083 50134 17259
rect 50088 17071 50134 17083
rect 50206 17259 50252 17271
rect 50206 17083 50212 17259
rect 50246 17083 50252 17259
rect 50206 17071 50252 17083
rect 50324 17259 50370 17271
rect 50324 17083 50330 17259
rect 50364 17083 50370 17259
rect 50324 17071 50370 17083
rect 49033 16854 49079 16870
rect 49033 16853 49114 16854
rect 49268 16853 49303 17071
rect 49547 17023 49613 17030
rect 49547 16989 49563 17023
rect 49597 16989 49613 17023
rect 49547 16978 49613 16989
rect 49739 16978 49775 17071
rect 49547 16977 49775 16978
rect 49975 16977 50011 17071
rect 50211 16977 50247 17071
rect 49547 16948 50247 16977
rect 49665 16947 50247 16948
rect 49665 16906 49731 16947
rect 49665 16872 49681 16906
rect 49715 16872 49731 16906
rect 49665 16865 49731 16872
rect 49033 16838 49303 16853
rect 49033 16834 49657 16838
rect 50093 16834 50127 16947
rect 49033 16822 49662 16834
rect 49033 16810 49622 16822
rect 49033 16808 49114 16810
rect 49380 16809 49622 16810
rect 48506 16642 48552 16654
rect 48416 16466 48512 16642
rect 48546 16466 48552 16642
rect 48376 16454 48422 16466
rect 48506 16454 48552 16466
rect 48624 16642 48670 16654
rect 48624 16466 48630 16642
rect 48664 16466 48670 16642
rect 48624 16454 48670 16466
rect 48742 16642 48788 16654
rect 48742 16466 48748 16642
rect 48782 16466 48788 16642
rect 48742 16454 48788 16466
rect 48860 16642 48906 16654
rect 48860 16466 48866 16642
rect 48900 16466 48906 16642
rect 49616 16646 49622 16809
rect 49656 16646 49662 16822
rect 49616 16634 49662 16646
rect 49734 16822 49780 16834
rect 49734 16646 49740 16822
rect 49774 16646 49780 16822
rect 49734 16634 49780 16646
rect 49851 16822 49897 16834
rect 48860 16454 48906 16466
rect 49535 16518 49643 16528
rect 49739 16518 49774 16634
rect 45293 16420 45327 16454
rect 45529 16420 45563 16454
rect 45293 16385 45563 16420
rect 46130 16420 46164 16454
rect 46366 16420 46400 16454
rect 46968 16420 47002 16454
rect 46130 16385 46400 16420
rect 46843 16385 47002 16420
rect 47191 16420 47225 16454
rect 47427 16420 47461 16454
rect 47191 16385 47461 16420
rect 48028 16420 48062 16454
rect 48264 16420 48298 16454
rect 48866 16420 48900 16454
rect 48028 16385 48298 16420
rect 48741 16385 48900 16420
rect 49643 16470 49774 16518
rect 49851 16470 49857 16822
rect 49643 16446 49857 16470
rect 49891 16446 49897 16822
rect 49643 16434 49897 16446
rect 49969 16822 50015 16834
rect 49969 16446 49975 16822
rect 50009 16446 50015 16822
rect 49969 16434 50015 16446
rect 50087 16822 50133 16834
rect 50087 16446 50093 16822
rect 50127 16446 50133 16822
rect 50087 16434 50133 16446
rect 49643 16430 49891 16434
rect 50260 16430 50270 16462
rect 49643 16386 49717 16430
rect 50255 16402 50270 16430
rect 49900 16396 49966 16402
rect 44602 16348 44744 16350
rect 44455 16339 44744 16348
rect 44456 16338 44744 16339
rect 44488 16337 44744 16338
rect 45279 16207 45346 16231
rect 45279 16173 45295 16207
rect 45329 16173 45346 16207
rect 44230 16006 44240 16085
rect 44333 16006 44343 16085
rect 43194 15957 43414 15977
rect 43194 15849 43238 15957
rect 43370 15849 43414 15957
rect 43194 15807 43414 15849
rect 42833 15777 43810 15807
rect 42833 15671 42867 15777
rect 43070 15671 43102 15777
rect 43306 15671 43338 15777
rect 43542 15671 43574 15777
rect 43778 15671 43810 15777
rect 40767 15600 41187 15605
rect 41901 15600 42217 15605
rect 40767 15589 41254 15600
rect 40767 15562 41203 15589
rect 40767 15561 41074 15562
rect 40767 15433 40801 15561
rect 41187 15555 41203 15562
rect 41237 15555 41254 15589
rect 41187 15549 41254 15555
rect 41834 15589 42217 15600
rect 41834 15555 41851 15589
rect 41885 15562 42217 15589
rect 41885 15555 41901 15562
rect 41834 15549 41901 15555
rect 40907 15521 40963 15533
rect 42020 15522 42076 15534
rect 42020 15521 42036 15522
rect 40907 15487 40913 15521
rect 40947 15506 41517 15521
rect 40947 15487 41467 15506
rect 40907 15472 41467 15487
rect 41501 15472 41517 15506
rect 40907 15471 40963 15472
rect 41450 15462 41517 15472
rect 41569 15505 42036 15521
rect 41569 15471 41585 15505
rect 41619 15488 42036 15505
rect 42070 15488 42076 15522
rect 41619 15472 42076 15488
rect 41619 15471 41635 15472
rect 41569 15464 41635 15471
rect 42183 15433 42217 15562
rect 42709 15659 42755 15671
rect 42709 15483 42715 15659
rect 42749 15483 42755 15659
rect 42709 15471 42755 15483
rect 42827 15659 42873 15671
rect 42827 15483 42833 15659
rect 42867 15483 42873 15659
rect 42827 15471 42873 15483
rect 42945 15659 42991 15671
rect 42945 15483 42951 15659
rect 42985 15483 42991 15659
rect 42945 15471 42991 15483
rect 43063 15659 43109 15671
rect 43063 15483 43069 15659
rect 43103 15483 43109 15659
rect 43063 15471 43109 15483
rect 43181 15659 43227 15671
rect 43181 15483 43187 15659
rect 43221 15483 43227 15659
rect 43181 15471 43227 15483
rect 43299 15659 43345 15671
rect 43299 15483 43305 15659
rect 43339 15483 43345 15659
rect 43299 15471 43345 15483
rect 43417 15659 43463 15671
rect 43417 15483 43423 15659
rect 43457 15483 43463 15659
rect 43417 15471 43463 15483
rect 43535 15659 43581 15671
rect 43535 15483 43541 15659
rect 43575 15483 43581 15659
rect 43535 15471 43581 15483
rect 43653 15659 43699 15671
rect 43653 15483 43659 15659
rect 43693 15483 43699 15659
rect 43653 15471 43699 15483
rect 43771 15659 43817 15671
rect 43771 15483 43777 15659
rect 43811 15483 43817 15659
rect 43771 15471 43817 15483
rect 38863 15421 38909 15433
rect 38863 15245 38869 15421
rect 38903 15245 38909 15421
rect 38863 15233 38909 15245
rect 38981 15421 39027 15433
rect 38981 15245 38987 15421
rect 39021 15245 39027 15421
rect 38981 15233 39027 15245
rect 39387 15421 39433 15433
rect 38988 14939 39021 15233
rect 39387 15045 39393 15421
rect 39427 15045 39433 15421
rect 39387 15033 39433 15045
rect 39505 15421 39551 15433
rect 39505 15045 39511 15421
rect 39545 15045 39551 15421
rect 39505 15033 39551 15045
rect 39623 15421 39669 15433
rect 39623 15045 39629 15421
rect 39663 15045 39669 15421
rect 39623 15033 39669 15045
rect 39741 15421 39787 15433
rect 39741 15045 39747 15421
rect 39781 15045 39787 15421
rect 39741 15033 39787 15045
rect 39859 15421 39905 15433
rect 39859 15045 39865 15421
rect 39899 15045 39905 15421
rect 40161 15421 40207 15433
rect 40161 15245 40167 15421
rect 40201 15245 40207 15421
rect 40161 15233 40207 15245
rect 40279 15421 40325 15433
rect 40279 15245 40285 15421
rect 40319 15245 40325 15421
rect 40279 15233 40325 15245
rect 40761 15421 40807 15433
rect 40761 15245 40767 15421
rect 40801 15245 40807 15421
rect 40761 15233 40807 15245
rect 40879 15421 40925 15433
rect 40879 15245 40885 15421
rect 40919 15245 40925 15421
rect 40879 15233 40925 15245
rect 41285 15421 41331 15433
rect 39859 15033 39905 15045
rect 39511 14939 39545 15033
rect 40168 14939 40202 15233
rect 38988 14907 40202 14939
rect 40886 14939 40919 15233
rect 41285 15045 41291 15421
rect 41325 15045 41331 15421
rect 41285 15033 41331 15045
rect 41403 15421 41449 15433
rect 41403 15045 41409 15421
rect 41443 15045 41449 15421
rect 41403 15033 41449 15045
rect 41521 15421 41567 15433
rect 41521 15045 41527 15421
rect 41561 15045 41567 15421
rect 41521 15033 41567 15045
rect 41639 15421 41685 15433
rect 41639 15045 41645 15421
rect 41679 15045 41685 15421
rect 41639 15033 41685 15045
rect 41757 15421 41803 15433
rect 41757 15045 41763 15421
rect 41797 15045 41803 15421
rect 42059 15421 42105 15433
rect 42059 15245 42065 15421
rect 42099 15245 42105 15421
rect 42059 15233 42105 15245
rect 42177 15421 42223 15433
rect 42177 15245 42183 15421
rect 42217 15245 42223 15421
rect 42177 15233 42223 15245
rect 42715 15238 42750 15471
rect 42994 15423 43060 15430
rect 42994 15389 43010 15423
rect 43044 15389 43060 15423
rect 42994 15378 43060 15389
rect 43186 15378 43222 15471
rect 42994 15377 43222 15378
rect 43422 15377 43458 15471
rect 43658 15377 43694 15471
rect 42994 15348 43694 15377
rect 43112 15347 43694 15348
rect 43112 15306 43178 15347
rect 43112 15272 43128 15306
rect 43162 15272 43178 15306
rect 43112 15265 43178 15272
rect 42715 15234 43104 15238
rect 43540 15234 43574 15347
rect 41757 15033 41803 15045
rect 41409 14939 41443 15033
rect 42066 14939 42100 15233
rect 42715 15222 43109 15234
rect 42715 15209 43069 15222
rect 42715 15206 42793 15209
rect 42710 15154 42720 15206
rect 42783 15154 42793 15206
rect 42715 15148 42788 15154
rect 43063 15046 43069 15209
rect 43103 15046 43109 15222
rect 43063 15034 43109 15046
rect 43181 15222 43227 15234
rect 43181 15046 43187 15222
rect 43221 15046 43227 15222
rect 43181 15034 43227 15046
rect 43298 15222 43344 15234
rect 40886 14907 42100 14939
rect 42982 14918 43090 14928
rect 43186 14918 43221 15034
rect 39577 14822 39709 14907
rect 41475 14822 41607 14907
rect 38722 14515 38788 14794
rect 39567 14714 39577 14822
rect 39709 14714 39719 14822
rect 41465 14714 41475 14822
rect 41607 14714 41617 14822
rect 43090 14870 43221 14918
rect 43298 14870 43304 15222
rect 43090 14846 43304 14870
rect 43338 14846 43344 15222
rect 43090 14834 43344 14846
rect 43416 15222 43462 15234
rect 43416 14846 43422 15222
rect 43456 14846 43462 15222
rect 43416 14834 43462 14846
rect 43534 15222 43580 15234
rect 43534 14846 43540 15222
rect 43574 14846 43580 15222
rect 43534 14834 43580 14846
rect 43090 14830 43338 14834
rect 44239 14832 44332 16006
rect 43747 14830 44332 14832
rect 43090 14786 43164 14830
rect 43702 14802 44332 14830
rect 43347 14796 43413 14802
rect 42982 14776 43090 14786
rect 43347 14762 43363 14796
rect 43397 14762 43413 14796
rect 43347 14666 43413 14762
rect 43465 14796 44332 14802
rect 43465 14762 43481 14796
rect 43515 14762 44332 14796
rect 43465 14746 44332 14762
rect 43702 14730 44332 14746
rect 43747 14726 44332 14730
rect 44231 14725 44332 14726
rect 45062 15744 45218 15750
rect 45062 15646 45074 15744
rect 45206 15646 45218 15744
rect 43702 14677 43802 14688
rect 43702 14666 43716 14677
rect 43347 14618 43716 14666
rect 43348 14515 43414 14618
rect 43702 14588 43716 14618
rect 43706 14571 43716 14588
rect 43828 14571 43838 14677
rect 38722 14435 43416 14515
rect 45062 13755 45218 15646
rect 45279 14790 45346 16173
rect 45427 15602 45461 16385
rect 46130 16323 46164 16385
rect 45833 16285 46575 16323
rect 45833 16161 45867 16285
rect 46069 16161 46103 16285
rect 46305 16161 46339 16285
rect 46541 16161 46575 16285
rect 45827 16149 45873 16161
rect 45827 15773 45833 16149
rect 45867 15773 45873 16149
rect 45827 15761 45873 15773
rect 45945 16149 45991 16161
rect 45945 15773 45951 16149
rect 45985 15773 45991 16149
rect 45945 15761 45991 15773
rect 46063 16149 46109 16161
rect 46063 15773 46069 16149
rect 46103 15773 46109 16149
rect 46063 15761 46109 15773
rect 46181 16149 46227 16161
rect 46181 15773 46187 16149
rect 46221 15773 46227 16149
rect 46181 15761 46227 15773
rect 46299 16149 46345 16161
rect 46299 15773 46305 16149
rect 46339 15773 46345 16149
rect 46299 15761 46345 15773
rect 46417 16149 46463 16161
rect 46417 15773 46423 16149
rect 46457 15773 46463 16149
rect 46417 15761 46463 15773
rect 46535 16149 46581 16161
rect 46535 15773 46541 16149
rect 46575 15773 46581 16149
rect 46535 15761 46581 15773
rect 45427 15601 45734 15602
rect 45780 15601 45849 15602
rect 46843 15601 46877 16385
rect 45427 15597 45849 15601
rect 45427 15586 45916 15597
rect 46561 15596 46877 15601
rect 45427 15558 45865 15586
rect 45427 15557 45734 15558
rect 45427 15429 45461 15557
rect 45849 15552 45865 15558
rect 45899 15552 45916 15586
rect 45849 15546 45916 15552
rect 46494 15585 46877 15596
rect 46494 15551 46511 15585
rect 46545 15558 46877 15585
rect 46545 15551 46561 15558
rect 46494 15545 46561 15551
rect 45567 15517 45623 15529
rect 46680 15518 46736 15530
rect 46680 15517 46696 15518
rect 45567 15483 45573 15517
rect 45607 15502 46177 15517
rect 45607 15483 46127 15502
rect 45567 15468 46127 15483
rect 46161 15468 46177 15502
rect 45567 15467 45623 15468
rect 46110 15458 46177 15468
rect 46229 15501 46696 15517
rect 46229 15467 46245 15501
rect 46279 15484 46696 15501
rect 46730 15484 46736 15518
rect 46279 15468 46736 15484
rect 46279 15467 46295 15468
rect 46229 15460 46295 15467
rect 46843 15429 46877 15558
rect 47325 15602 47359 16385
rect 48028 16323 48062 16385
rect 47731 16285 48473 16323
rect 47392 16178 47402 16244
rect 47465 16178 47475 16244
rect 47731 16161 47765 16285
rect 47967 16161 48001 16285
rect 48203 16161 48237 16285
rect 48439 16161 48473 16285
rect 47725 16149 47771 16161
rect 47725 15773 47731 16149
rect 47765 15773 47771 16149
rect 47725 15761 47771 15773
rect 47843 16149 47889 16161
rect 47843 15773 47849 16149
rect 47883 15773 47889 16149
rect 47843 15761 47889 15773
rect 47961 16149 48007 16161
rect 47961 15773 47967 16149
rect 48001 15773 48007 16149
rect 47961 15761 48007 15773
rect 48079 16149 48125 16161
rect 48079 15773 48085 16149
rect 48119 15773 48125 16149
rect 48079 15761 48125 15773
rect 48197 16149 48243 16161
rect 48197 15773 48203 16149
rect 48237 15773 48243 16149
rect 48197 15761 48243 15773
rect 48315 16149 48361 16161
rect 48315 15773 48321 16149
rect 48355 15773 48361 16149
rect 48315 15761 48361 15773
rect 48433 16149 48479 16161
rect 48433 15773 48439 16149
rect 48473 15773 48479 16149
rect 48433 15761 48479 15773
rect 47325 15601 47632 15602
rect 48741 15601 48775 16385
rect 49535 16376 49643 16386
rect 49900 16362 49916 16396
rect 49950 16362 49966 16396
rect 49900 16266 49966 16362
rect 50018 16396 50270 16402
rect 50018 16362 50034 16396
rect 50068 16362 50270 16396
rect 50018 16346 50270 16362
rect 50255 16344 50270 16346
rect 50388 16344 50398 16462
rect 50255 16330 50355 16344
rect 50255 16287 50355 16288
rect 50629 16287 50734 17464
rect 50255 16266 50734 16287
rect 49900 16218 50734 16266
rect 50255 16189 50734 16218
rect 50255 16188 50355 16189
rect 50629 16187 50734 16189
rect 50797 16081 50890 17975
rect 51030 17974 51319 17975
rect 51013 17564 51183 17617
rect 51013 17551 51053 17564
rect 51011 17458 51053 17551
rect 51165 17458 51183 17564
rect 51011 17447 51183 17458
rect 51013 17446 51183 17447
rect 51631 16617 51731 18357
rect 52628 18219 52662 18365
rect 52812 18350 52909 18365
rect 53382 18362 53417 18454
rect 52852 18283 52909 18350
rect 53190 18326 53417 18362
rect 53190 18292 53256 18326
rect 52746 18247 53015 18283
rect 53190 18258 53206 18292
rect 53240 18258 53256 18292
rect 53190 18252 53256 18258
rect 52746 18219 52779 18247
rect 52982 18219 53015 18247
rect 53382 18219 53417 18326
rect 52622 18207 52668 18219
rect 52622 18031 52628 18207
rect 52662 18031 52668 18207
rect 52622 18019 52668 18031
rect 52740 18207 52786 18219
rect 52740 18031 52746 18207
rect 52780 18031 52786 18207
rect 52740 18019 52786 18031
rect 52858 18207 52904 18219
rect 52858 18031 52864 18207
rect 52898 18031 52904 18207
rect 52858 18019 52904 18031
rect 52976 18207 53022 18219
rect 52976 18031 52982 18207
rect 53016 18152 53022 18207
rect 53141 18207 53187 18219
rect 53141 18152 53147 18207
rect 53016 18064 53147 18152
rect 53016 18031 53022 18064
rect 52976 18019 53022 18031
rect 53141 18031 53147 18064
rect 53181 18031 53187 18207
rect 53141 18019 53187 18031
rect 53259 18207 53305 18219
rect 53259 18031 53265 18207
rect 53299 18031 53305 18207
rect 53259 18019 53305 18031
rect 53377 18207 53423 18219
rect 53377 18031 53383 18207
rect 53417 18031 53423 18207
rect 53377 18019 53423 18031
rect 53495 18207 53541 18219
rect 53495 18031 53501 18207
rect 53535 18031 53541 18207
rect 53495 18019 53541 18031
rect 52629 17981 52662 18019
rect 52865 17981 52898 18019
rect 52629 17945 52898 17981
rect 53265 17980 53299 18019
rect 53501 17980 53535 18019
rect 53265 17944 53535 17980
rect 53369 17943 53535 17944
rect 53369 17864 53501 17943
rect 53359 17756 53369 17864
rect 53501 17756 53511 17864
rect 53641 17427 53703 18998
rect 53839 18986 53885 18998
rect 53839 18610 53845 18986
rect 53879 18610 53885 18986
rect 53839 18598 53885 18610
rect 53957 18986 54003 18998
rect 53957 18610 53963 18986
rect 53997 18610 54003 18986
rect 53957 18598 54003 18610
rect 54075 18986 54121 18998
rect 54075 18610 54081 18986
rect 54115 18610 54121 18986
rect 54075 18598 54121 18610
rect 54193 18986 54239 18998
rect 54193 18610 54199 18986
rect 54233 18610 54239 18986
rect 54193 18598 54239 18610
rect 54311 18986 54357 18998
rect 54311 18610 54317 18986
rect 54351 18610 54357 18986
rect 54311 18598 54357 18610
rect 54429 18986 54475 18998
rect 54429 18610 54435 18986
rect 54469 18610 54475 18986
rect 54429 18598 54475 18610
rect 54547 18986 54593 18998
rect 54642 18994 54652 19060
rect 54718 18994 54728 19060
rect 54547 18610 54553 18986
rect 54587 18610 54593 18986
rect 54547 18598 54593 18610
rect 53845 18415 53879 18598
rect 53963 18557 53997 18598
rect 54199 18557 54233 18598
rect 53963 18528 54233 18557
rect 54317 18556 54351 18598
rect 54553 18556 54587 18598
rect 54317 18528 54587 18556
rect 54553 18480 54587 18528
rect 54524 18450 54587 18480
rect 55577 18521 55644 19111
rect 56295 19104 56339 19212
rect 56471 19104 56515 19212
rect 59213 19206 59223 19269
rect 59211 19195 59223 19206
rect 56295 19062 56515 19104
rect 59210 19161 59223 19195
rect 59355 19161 59365 19269
rect 60360 19206 60370 19269
rect 60358 19195 60370 19206
rect 60045 19185 60101 19187
rect 59210 19123 59355 19161
rect 59210 19095 59251 19123
rect 60035 19119 60045 19185
rect 60101 19119 60111 19185
rect 60357 19161 60370 19195
rect 60502 19161 60512 19269
rect 62808 19215 63028 19235
rect 61175 19173 61231 19181
rect 61175 19165 62157 19173
rect 60357 19123 60502 19161
rect 61175 19131 61181 19165
rect 61215 19131 62157 19165
rect 59210 19067 59486 19095
rect 55934 19032 56911 19062
rect 55934 18926 55968 19032
rect 56171 18926 56203 19032
rect 56407 18926 56439 19032
rect 56643 18926 56675 19032
rect 56879 18926 56911 19032
rect 59210 19005 59250 19067
rect 59452 19005 59486 19067
rect 59570 19067 59840 19095
rect 60357 19091 60398 19123
rect 61175 19115 62157 19131
rect 61178 19114 62157 19115
rect 59570 19005 59604 19067
rect 59806 19005 59840 19067
rect 60045 19051 60216 19067
rect 60045 19017 60051 19051
rect 60085 19017 60216 19051
rect 59210 18993 59256 19005
rect 55810 18914 55856 18926
rect 55810 18738 55816 18914
rect 55850 18738 55856 18914
rect 55810 18726 55856 18738
rect 55928 18914 55974 18926
rect 55928 18738 55934 18914
rect 55968 18738 55974 18914
rect 55928 18726 55974 18738
rect 56046 18914 56092 18926
rect 56046 18738 56052 18914
rect 56086 18738 56092 18914
rect 56046 18726 56092 18738
rect 56164 18914 56210 18926
rect 56164 18738 56170 18914
rect 56204 18738 56210 18914
rect 56164 18726 56210 18738
rect 56282 18914 56328 18926
rect 56282 18738 56288 18914
rect 56322 18738 56328 18914
rect 56282 18726 56328 18738
rect 56400 18914 56446 18926
rect 56400 18738 56406 18914
rect 56440 18738 56446 18914
rect 56400 18726 56446 18738
rect 56518 18914 56564 18926
rect 56518 18738 56524 18914
rect 56558 18738 56564 18914
rect 56518 18726 56564 18738
rect 56636 18914 56682 18926
rect 56636 18738 56642 18914
rect 56676 18738 56682 18914
rect 56636 18726 56682 18738
rect 56754 18914 56800 18926
rect 56754 18738 56760 18914
rect 56794 18738 56800 18914
rect 56754 18726 56800 18738
rect 56872 18914 56918 18926
rect 56872 18738 56878 18914
rect 56912 18738 56918 18914
rect 56872 18726 56918 18738
rect 55816 18521 55851 18726
rect 56095 18678 56161 18685
rect 56095 18644 56111 18678
rect 56145 18644 56161 18678
rect 56095 18633 56161 18644
rect 56287 18633 56323 18726
rect 56095 18632 56323 18633
rect 56523 18632 56559 18726
rect 56759 18632 56795 18726
rect 56095 18603 56795 18632
rect 59210 18617 59216 18993
rect 59250 18617 59256 18993
rect 59210 18605 59256 18617
rect 59328 18993 59374 19005
rect 59328 18617 59334 18993
rect 59368 18617 59374 18993
rect 59328 18605 59374 18617
rect 59446 18993 59492 19005
rect 59446 18617 59452 18993
rect 59486 18617 59492 18993
rect 59446 18605 59492 18617
rect 59564 18993 59610 19005
rect 59564 18617 59570 18993
rect 59604 18617 59610 18993
rect 59564 18605 59610 18617
rect 59682 18993 59728 19005
rect 59682 18617 59688 18993
rect 59722 18617 59728 18993
rect 59682 18605 59728 18617
rect 59800 18993 59846 19005
rect 59800 18617 59806 18993
rect 59840 18617 59846 18993
rect 59800 18605 59846 18617
rect 59918 18993 59964 19005
rect 60045 19001 60216 19017
rect 60357 19063 60628 19091
rect 60357 19001 60392 19063
rect 60594 19001 60628 19063
rect 60712 19063 60982 19091
rect 60712 19001 60746 19063
rect 60948 19001 60982 19063
rect 59918 18617 59924 18993
rect 59958 18617 59964 18993
rect 59918 18605 59964 18617
rect 55577 18493 55851 18521
rect 56213 18602 56795 18603
rect 56213 18561 56279 18602
rect 56213 18527 56229 18561
rect 56263 18527 56279 18561
rect 56213 18520 56279 18527
rect 55577 18489 56205 18493
rect 56641 18489 56675 18602
rect 55577 18477 56210 18489
rect 55577 18464 56170 18477
rect 53770 18361 53879 18415
rect 53770 18215 53804 18361
rect 53943 18347 53953 18444
rect 54052 18347 54062 18444
rect 54524 18358 54559 18450
rect 53954 18346 54051 18347
rect 53994 18279 54051 18346
rect 54332 18322 54559 18358
rect 54332 18288 54398 18322
rect 53888 18243 54157 18279
rect 54332 18254 54348 18288
rect 54382 18254 54398 18288
rect 54332 18248 54398 18254
rect 53888 18215 53921 18243
rect 54124 18215 54157 18243
rect 54524 18215 54559 18322
rect 56164 18301 56170 18464
rect 56204 18301 56210 18477
rect 56164 18289 56210 18301
rect 56282 18477 56328 18489
rect 56282 18301 56288 18477
rect 56322 18301 56328 18477
rect 56282 18289 56328 18301
rect 56399 18477 56445 18489
rect 53764 18203 53810 18215
rect 53764 18027 53770 18203
rect 53804 18027 53810 18203
rect 53764 18015 53810 18027
rect 53882 18203 53928 18215
rect 53882 18027 53888 18203
rect 53922 18027 53928 18203
rect 53882 18015 53928 18027
rect 54000 18203 54046 18215
rect 54000 18027 54006 18203
rect 54040 18027 54046 18203
rect 54000 18015 54046 18027
rect 54118 18203 54164 18215
rect 54118 18027 54124 18203
rect 54158 18148 54164 18203
rect 54283 18203 54329 18215
rect 54283 18148 54289 18203
rect 54158 18060 54289 18148
rect 54158 18027 54164 18060
rect 54118 18015 54164 18027
rect 54283 18027 54289 18060
rect 54323 18027 54329 18203
rect 54283 18015 54329 18027
rect 54401 18203 54447 18215
rect 54401 18027 54407 18203
rect 54441 18027 54447 18203
rect 54401 18015 54447 18027
rect 54519 18203 54565 18215
rect 54519 18027 54525 18203
rect 54559 18027 54565 18203
rect 54519 18015 54565 18027
rect 54637 18203 54683 18215
rect 54637 18027 54643 18203
rect 54677 18027 54683 18203
rect 56083 18173 56191 18183
rect 56287 18173 56322 18289
rect 56191 18125 56322 18173
rect 56399 18125 56405 18477
rect 56191 18101 56405 18125
rect 56439 18101 56445 18477
rect 56191 18089 56445 18101
rect 56517 18477 56563 18489
rect 56517 18101 56523 18477
rect 56557 18101 56563 18477
rect 56517 18089 56563 18101
rect 56635 18477 56681 18489
rect 56635 18101 56641 18477
rect 56675 18101 56681 18477
rect 58146 18361 58246 18436
rect 58314 18361 58324 18436
rect 59216 18422 59250 18605
rect 59334 18564 59368 18605
rect 59570 18564 59604 18605
rect 59334 18535 59604 18564
rect 59688 18563 59722 18605
rect 59924 18563 59958 18605
rect 59688 18535 59958 18563
rect 59924 18487 59958 18535
rect 59895 18457 59958 18487
rect 59141 18368 59250 18422
rect 59323 18427 59423 18448
rect 59323 18373 59344 18427
rect 59409 18373 59423 18427
rect 59323 18368 59423 18373
rect 58146 18360 58297 18361
rect 56635 18089 56681 18101
rect 57564 18135 57853 18153
rect 56191 18085 56439 18089
rect 56191 18041 56265 18085
rect 57564 18084 57605 18135
rect 56803 18057 57605 18084
rect 56448 18051 56514 18057
rect 56083 18031 56191 18041
rect 54637 18015 54683 18027
rect 56448 18017 56464 18051
rect 56498 18017 56514 18051
rect 53771 17977 53804 18015
rect 54007 17977 54040 18015
rect 53771 17941 54040 17977
rect 54407 17976 54441 18015
rect 54643 17976 54677 18015
rect 54407 17941 54677 17976
rect 54407 17940 54643 17941
rect 54511 17866 54643 17940
rect 56448 17921 56514 18017
rect 56566 18051 57605 18057
rect 56566 18017 56582 18051
rect 56616 18017 57605 18051
rect 56566 18001 57605 18017
rect 56803 17998 57605 18001
rect 57833 17998 57853 18135
rect 56803 17985 57853 17998
rect 56866 17984 57853 17985
rect 57331 17980 57853 17984
rect 56802 17921 57268 17943
rect 56448 17873 57268 17921
rect 54501 17758 54511 17866
rect 54643 17758 54653 17866
rect 56802 17842 57268 17873
rect 57163 17586 57268 17842
rect 53640 17410 53703 17427
rect 56281 17562 56501 17582
rect 56281 17454 56325 17562
rect 56457 17454 56501 17562
rect 57083 17480 57093 17586
rect 57205 17480 57268 17586
rect 57119 17469 57268 17480
rect 56281 17412 56501 17454
rect 53640 17406 53778 17410
rect 53640 17372 55610 17406
rect 55920 17382 56897 17412
rect 53640 17343 55612 17372
rect 53640 17341 53778 17343
rect 55566 17327 55612 17343
rect 52604 17111 52614 17219
rect 52746 17111 52756 17219
rect 54502 17111 54512 17219
rect 54644 17111 54654 17219
rect 52614 17071 52746 17111
rect 54512 17071 54644 17111
rect 52614 17005 52747 17071
rect 54512 17005 54645 17071
rect 51945 16962 53418 17005
rect 51945 16659 51979 16962
rect 52310 16859 52344 16962
rect 52546 16859 52580 16962
rect 52782 16859 52816 16962
rect 53018 16859 53052 16962
rect 52304 16847 52350 16859
rect 51046 16614 51731 16617
rect 51014 16516 51731 16614
rect 51821 16647 51867 16659
rect 51014 16515 51489 16516
rect 51014 16452 51302 16515
rect 51821 16471 51827 16647
rect 51861 16471 51867 16647
rect 51821 16459 51867 16471
rect 51939 16647 51985 16659
rect 51939 16471 51945 16647
rect 51979 16471 51985 16647
rect 51939 16459 51985 16471
rect 52057 16647 52103 16659
rect 52057 16471 52063 16647
rect 52097 16471 52103 16647
rect 52057 16459 52103 16471
rect 52175 16647 52221 16659
rect 52304 16647 52310 16847
rect 52175 16471 52181 16647
rect 52215 16471 52310 16647
rect 52344 16471 52350 16847
rect 52175 16459 52221 16471
rect 52304 16459 52350 16471
rect 52422 16847 52468 16859
rect 52422 16471 52428 16847
rect 52462 16471 52468 16847
rect 52422 16459 52468 16471
rect 52540 16847 52586 16859
rect 52540 16471 52546 16847
rect 52580 16471 52586 16847
rect 52540 16459 52586 16471
rect 52658 16847 52704 16859
rect 52658 16471 52664 16847
rect 52698 16471 52704 16847
rect 52658 16459 52704 16471
rect 52776 16847 52822 16859
rect 52776 16471 52782 16847
rect 52816 16471 52822 16847
rect 52776 16459 52822 16471
rect 52894 16847 52940 16859
rect 52894 16471 52900 16847
rect 52934 16471 52940 16847
rect 52894 16459 52940 16471
rect 53012 16847 53058 16859
rect 53012 16471 53018 16847
rect 53052 16647 53058 16847
rect 53384 16659 53418 16962
rect 53843 16962 55316 17005
rect 53843 16659 53877 16962
rect 54208 16859 54242 16962
rect 54444 16859 54478 16962
rect 54680 16859 54714 16962
rect 54916 16859 54950 16962
rect 54202 16847 54248 16859
rect 53142 16647 53188 16659
rect 53052 16471 53148 16647
rect 53182 16471 53188 16647
rect 53012 16459 53058 16471
rect 53142 16459 53188 16471
rect 53260 16647 53306 16659
rect 53260 16471 53266 16647
rect 53300 16471 53306 16647
rect 53260 16459 53306 16471
rect 53378 16647 53424 16659
rect 53378 16471 53384 16647
rect 53418 16471 53424 16647
rect 53378 16459 53424 16471
rect 53496 16647 53542 16659
rect 53496 16471 53502 16647
rect 53536 16471 53542 16647
rect 53496 16459 53542 16471
rect 53719 16647 53765 16659
rect 53719 16471 53725 16647
rect 53759 16471 53765 16647
rect 53719 16459 53765 16471
rect 53837 16647 53883 16659
rect 53837 16471 53843 16647
rect 53877 16471 53883 16647
rect 53837 16459 53883 16471
rect 53955 16647 54001 16659
rect 53955 16471 53961 16647
rect 53995 16471 54001 16647
rect 53955 16459 54001 16471
rect 54073 16647 54119 16659
rect 54202 16647 54208 16847
rect 54073 16471 54079 16647
rect 54113 16471 54208 16647
rect 54242 16471 54248 16847
rect 54073 16459 54119 16471
rect 54202 16459 54248 16471
rect 54320 16847 54366 16859
rect 54320 16471 54326 16847
rect 54360 16471 54366 16847
rect 54320 16459 54366 16471
rect 54438 16847 54484 16859
rect 54438 16471 54444 16847
rect 54478 16471 54484 16847
rect 54438 16459 54484 16471
rect 54556 16847 54602 16859
rect 54556 16471 54562 16847
rect 54596 16471 54602 16847
rect 54556 16459 54602 16471
rect 54674 16847 54720 16859
rect 54674 16471 54680 16847
rect 54714 16471 54720 16847
rect 54674 16459 54720 16471
rect 54792 16847 54838 16859
rect 54792 16471 54798 16847
rect 54832 16471 54838 16847
rect 54792 16459 54838 16471
rect 54910 16847 54956 16859
rect 54910 16471 54916 16847
rect 54950 16647 54956 16847
rect 55282 16659 55316 16962
rect 55566 16875 55613 17327
rect 55920 17276 55954 17382
rect 56157 17276 56189 17382
rect 56393 17276 56425 17382
rect 56629 17276 56661 17382
rect 56865 17276 56897 17382
rect 55796 17264 55842 17276
rect 55796 17088 55802 17264
rect 55836 17088 55842 17264
rect 55796 17076 55842 17088
rect 55914 17264 55960 17276
rect 55914 17088 55920 17264
rect 55954 17088 55960 17264
rect 55914 17076 55960 17088
rect 56032 17264 56078 17276
rect 56032 17088 56038 17264
rect 56072 17088 56078 17264
rect 56032 17076 56078 17088
rect 56150 17264 56196 17276
rect 56150 17088 56156 17264
rect 56190 17088 56196 17264
rect 56150 17076 56196 17088
rect 56268 17264 56314 17276
rect 56268 17088 56274 17264
rect 56308 17088 56314 17264
rect 56268 17076 56314 17088
rect 56386 17264 56432 17276
rect 56386 17088 56392 17264
rect 56426 17088 56432 17264
rect 56386 17076 56432 17088
rect 56504 17264 56550 17276
rect 56504 17088 56510 17264
rect 56544 17088 56550 17264
rect 56504 17076 56550 17088
rect 56622 17264 56668 17276
rect 56622 17088 56628 17264
rect 56662 17088 56668 17264
rect 56622 17076 56668 17088
rect 56740 17264 56786 17276
rect 56740 17088 56746 17264
rect 56780 17088 56786 17264
rect 56740 17076 56786 17088
rect 56858 17264 56904 17276
rect 56858 17088 56864 17264
rect 56898 17088 56904 17264
rect 56858 17076 56904 17088
rect 55567 16859 55613 16875
rect 55567 16858 55648 16859
rect 55802 16858 55837 17076
rect 56081 17028 56147 17035
rect 56081 16994 56097 17028
rect 56131 16994 56147 17028
rect 56081 16983 56147 16994
rect 56273 16983 56309 17076
rect 56081 16982 56309 16983
rect 56509 16982 56545 17076
rect 56745 16982 56781 17076
rect 56081 16953 56781 16982
rect 56199 16952 56781 16953
rect 56199 16911 56265 16952
rect 56199 16877 56215 16911
rect 56249 16877 56265 16911
rect 56199 16870 56265 16877
rect 55567 16843 55837 16858
rect 55567 16839 56191 16843
rect 56627 16839 56661 16952
rect 55567 16827 56196 16839
rect 55567 16815 56156 16827
rect 55567 16813 55648 16815
rect 55914 16814 56156 16815
rect 55040 16647 55086 16659
rect 54950 16471 55046 16647
rect 55080 16471 55086 16647
rect 54910 16459 54956 16471
rect 55040 16459 55086 16471
rect 55158 16647 55204 16659
rect 55158 16471 55164 16647
rect 55198 16471 55204 16647
rect 55158 16459 55204 16471
rect 55276 16647 55322 16659
rect 55276 16471 55282 16647
rect 55316 16471 55322 16647
rect 55276 16459 55322 16471
rect 55394 16647 55440 16659
rect 55394 16471 55400 16647
rect 55434 16471 55440 16647
rect 56150 16651 56156 16814
rect 56190 16651 56196 16827
rect 56150 16639 56196 16651
rect 56268 16827 56314 16839
rect 56268 16651 56274 16827
rect 56308 16651 56314 16827
rect 56268 16639 56314 16651
rect 56385 16827 56431 16839
rect 55394 16459 55440 16471
rect 56069 16523 56177 16533
rect 56273 16523 56308 16639
rect 51014 16450 51054 16452
rect 51014 16439 51048 16450
rect 51013 16344 51048 16439
rect 51166 16346 51302 16452
rect 51827 16425 51861 16459
rect 52063 16425 52097 16459
rect 51827 16390 52097 16425
rect 52664 16425 52698 16459
rect 52900 16425 52934 16459
rect 53502 16425 53536 16459
rect 52664 16390 52934 16425
rect 53377 16390 53536 16425
rect 53725 16425 53759 16459
rect 53961 16425 53995 16459
rect 53725 16390 53995 16425
rect 54562 16425 54596 16459
rect 54798 16425 54832 16459
rect 55400 16425 55434 16459
rect 54562 16390 54832 16425
rect 55275 16390 55434 16425
rect 56177 16475 56308 16523
rect 56385 16475 56391 16827
rect 56177 16451 56391 16475
rect 56425 16451 56431 16827
rect 56177 16439 56431 16451
rect 56503 16827 56549 16839
rect 56503 16451 56509 16827
rect 56543 16451 56549 16827
rect 56503 16439 56549 16451
rect 56621 16827 56667 16839
rect 56621 16451 56627 16827
rect 56661 16451 56667 16827
rect 56621 16439 56667 16451
rect 56177 16435 56425 16439
rect 56794 16435 56804 16467
rect 56177 16391 56251 16435
rect 56789 16407 56804 16435
rect 56434 16401 56500 16407
rect 51160 16344 51302 16346
rect 51013 16335 51302 16344
rect 51014 16334 51302 16335
rect 51046 16333 51302 16334
rect 51813 16212 51880 16236
rect 51813 16178 51829 16212
rect 51863 16178 51880 16212
rect 50788 16002 50798 16081
rect 50891 16002 50901 16081
rect 49752 15953 49972 15973
rect 49752 15845 49796 15953
rect 49928 15845 49972 15953
rect 49752 15803 49972 15845
rect 49391 15773 50368 15803
rect 49391 15667 49425 15773
rect 49628 15667 49660 15773
rect 49864 15667 49896 15773
rect 50100 15667 50132 15773
rect 50336 15667 50368 15773
rect 47325 15596 47745 15601
rect 48459 15596 48775 15601
rect 47325 15585 47812 15596
rect 47325 15558 47761 15585
rect 47325 15557 47632 15558
rect 47325 15429 47359 15557
rect 47745 15551 47761 15558
rect 47795 15551 47812 15585
rect 47745 15545 47812 15551
rect 48392 15585 48775 15596
rect 48392 15551 48409 15585
rect 48443 15558 48775 15585
rect 48443 15551 48459 15558
rect 48392 15545 48459 15551
rect 47465 15517 47521 15529
rect 48578 15518 48634 15530
rect 48578 15517 48594 15518
rect 47465 15483 47471 15517
rect 47505 15502 48075 15517
rect 47505 15483 48025 15502
rect 47465 15468 48025 15483
rect 48059 15468 48075 15502
rect 47465 15467 47521 15468
rect 48008 15458 48075 15468
rect 48127 15501 48594 15517
rect 48127 15467 48143 15501
rect 48177 15484 48594 15501
rect 48628 15484 48634 15518
rect 48177 15468 48634 15484
rect 48177 15467 48193 15468
rect 48127 15460 48193 15467
rect 48741 15429 48775 15558
rect 49267 15655 49313 15667
rect 49267 15479 49273 15655
rect 49307 15479 49313 15655
rect 49267 15467 49313 15479
rect 49385 15655 49431 15667
rect 49385 15479 49391 15655
rect 49425 15479 49431 15655
rect 49385 15467 49431 15479
rect 49503 15655 49549 15667
rect 49503 15479 49509 15655
rect 49543 15479 49549 15655
rect 49503 15467 49549 15479
rect 49621 15655 49667 15667
rect 49621 15479 49627 15655
rect 49661 15479 49667 15655
rect 49621 15467 49667 15479
rect 49739 15655 49785 15667
rect 49739 15479 49745 15655
rect 49779 15479 49785 15655
rect 49739 15467 49785 15479
rect 49857 15655 49903 15667
rect 49857 15479 49863 15655
rect 49897 15479 49903 15655
rect 49857 15467 49903 15479
rect 49975 15655 50021 15667
rect 49975 15479 49981 15655
rect 50015 15479 50021 15655
rect 49975 15467 50021 15479
rect 50093 15655 50139 15667
rect 50093 15479 50099 15655
rect 50133 15479 50139 15655
rect 50093 15467 50139 15479
rect 50211 15655 50257 15667
rect 50211 15479 50217 15655
rect 50251 15479 50257 15655
rect 50211 15467 50257 15479
rect 50329 15655 50375 15667
rect 50329 15479 50335 15655
rect 50369 15479 50375 15655
rect 50329 15467 50375 15479
rect 45421 15417 45467 15429
rect 45421 15241 45427 15417
rect 45461 15241 45467 15417
rect 45421 15229 45467 15241
rect 45539 15417 45585 15429
rect 45539 15241 45545 15417
rect 45579 15241 45585 15417
rect 45539 15229 45585 15241
rect 45945 15417 45991 15429
rect 45546 14935 45579 15229
rect 45945 15041 45951 15417
rect 45985 15041 45991 15417
rect 45945 15029 45991 15041
rect 46063 15417 46109 15429
rect 46063 15041 46069 15417
rect 46103 15041 46109 15417
rect 46063 15029 46109 15041
rect 46181 15417 46227 15429
rect 46181 15041 46187 15417
rect 46221 15041 46227 15417
rect 46181 15029 46227 15041
rect 46299 15417 46345 15429
rect 46299 15041 46305 15417
rect 46339 15041 46345 15417
rect 46299 15029 46345 15041
rect 46417 15417 46463 15429
rect 46417 15041 46423 15417
rect 46457 15041 46463 15417
rect 46719 15417 46765 15429
rect 46719 15241 46725 15417
rect 46759 15241 46765 15417
rect 46719 15229 46765 15241
rect 46837 15417 46883 15429
rect 46837 15241 46843 15417
rect 46877 15241 46883 15417
rect 46837 15229 46883 15241
rect 47319 15417 47365 15429
rect 47319 15241 47325 15417
rect 47359 15241 47365 15417
rect 47319 15229 47365 15241
rect 47437 15417 47483 15429
rect 47437 15241 47443 15417
rect 47477 15241 47483 15417
rect 47437 15229 47483 15241
rect 47843 15417 47889 15429
rect 46417 15029 46463 15041
rect 46069 14935 46103 15029
rect 46726 14935 46760 15229
rect 45546 14903 46760 14935
rect 47444 14935 47477 15229
rect 47843 15041 47849 15417
rect 47883 15041 47889 15417
rect 47843 15029 47889 15041
rect 47961 15417 48007 15429
rect 47961 15041 47967 15417
rect 48001 15041 48007 15417
rect 47961 15029 48007 15041
rect 48079 15417 48125 15429
rect 48079 15041 48085 15417
rect 48119 15041 48125 15417
rect 48079 15029 48125 15041
rect 48197 15417 48243 15429
rect 48197 15041 48203 15417
rect 48237 15041 48243 15417
rect 48197 15029 48243 15041
rect 48315 15417 48361 15429
rect 48315 15041 48321 15417
rect 48355 15041 48361 15417
rect 48617 15417 48663 15429
rect 48617 15241 48623 15417
rect 48657 15241 48663 15417
rect 48617 15229 48663 15241
rect 48735 15417 48781 15429
rect 48735 15241 48741 15417
rect 48775 15241 48781 15417
rect 48735 15229 48781 15241
rect 49273 15234 49308 15467
rect 49552 15419 49618 15426
rect 49552 15385 49568 15419
rect 49602 15385 49618 15419
rect 49552 15374 49618 15385
rect 49744 15374 49780 15467
rect 49552 15373 49780 15374
rect 49980 15373 50016 15467
rect 50216 15373 50252 15467
rect 49552 15344 50252 15373
rect 49670 15343 50252 15344
rect 49670 15302 49736 15343
rect 49670 15268 49686 15302
rect 49720 15268 49736 15302
rect 49670 15261 49736 15268
rect 49273 15230 49662 15234
rect 50098 15230 50132 15343
rect 48315 15029 48361 15041
rect 47967 14935 48001 15029
rect 48624 14935 48658 15229
rect 49273 15218 49667 15230
rect 49273 15205 49627 15218
rect 49273 15202 49351 15205
rect 49268 15150 49278 15202
rect 49341 15150 49351 15202
rect 49273 15144 49346 15150
rect 49621 15042 49627 15205
rect 49661 15042 49667 15218
rect 49621 15030 49667 15042
rect 49739 15218 49785 15230
rect 49739 15042 49745 15218
rect 49779 15042 49785 15218
rect 49739 15030 49785 15042
rect 49856 15218 49902 15230
rect 47444 14903 48658 14935
rect 49540 14914 49648 14924
rect 49744 14914 49779 15030
rect 46135 14818 46267 14903
rect 48033 14818 48165 14903
rect 45280 14511 45346 14790
rect 46125 14710 46135 14818
rect 46267 14710 46277 14818
rect 48023 14710 48033 14818
rect 48165 14710 48175 14818
rect 49648 14866 49779 14914
rect 49856 14866 49862 15218
rect 49648 14842 49862 14866
rect 49896 14842 49902 15218
rect 49648 14830 49902 14842
rect 49974 15218 50020 15230
rect 49974 14842 49980 15218
rect 50014 14842 50020 15218
rect 49974 14830 50020 14842
rect 50092 15218 50138 15230
rect 50092 14842 50098 15218
rect 50132 14842 50138 15218
rect 50092 14830 50138 14842
rect 49648 14826 49896 14830
rect 50797 14828 50890 16002
rect 50305 14826 50890 14828
rect 49648 14782 49722 14826
rect 50260 14798 50890 14826
rect 49905 14792 49971 14798
rect 49540 14772 49648 14782
rect 49905 14758 49921 14792
rect 49955 14758 49971 14792
rect 49905 14662 49971 14758
rect 50023 14792 50890 14798
rect 50023 14758 50039 14792
rect 50073 14758 50890 14792
rect 50023 14742 50890 14758
rect 50260 14726 50890 14742
rect 50305 14722 50890 14726
rect 50789 14721 50890 14722
rect 51596 15749 51752 15755
rect 51596 15651 51608 15749
rect 51740 15706 51752 15749
rect 51740 15651 51753 15706
rect 50260 14673 50360 14684
rect 50260 14662 50274 14673
rect 49905 14614 50274 14662
rect 49906 14511 49972 14614
rect 50260 14584 50274 14614
rect 50264 14567 50274 14584
rect 50386 14567 50396 14673
rect 45280 14431 49974 14511
rect 51596 13866 51753 15651
rect 51813 14795 51880 16178
rect 51961 15607 51995 16390
rect 52664 16328 52698 16390
rect 52367 16290 53109 16328
rect 52367 16166 52401 16290
rect 52603 16166 52637 16290
rect 52839 16166 52873 16290
rect 53075 16166 53109 16290
rect 52361 16154 52407 16166
rect 52361 15778 52367 16154
rect 52401 15778 52407 16154
rect 52361 15766 52407 15778
rect 52479 16154 52525 16166
rect 52479 15778 52485 16154
rect 52519 15778 52525 16154
rect 52479 15766 52525 15778
rect 52597 16154 52643 16166
rect 52597 15778 52603 16154
rect 52637 15778 52643 16154
rect 52597 15766 52643 15778
rect 52715 16154 52761 16166
rect 52715 15778 52721 16154
rect 52755 15778 52761 16154
rect 52715 15766 52761 15778
rect 52833 16154 52879 16166
rect 52833 15778 52839 16154
rect 52873 15778 52879 16154
rect 52833 15766 52879 15778
rect 52951 16154 52997 16166
rect 52951 15778 52957 16154
rect 52991 15778 52997 16154
rect 52951 15766 52997 15778
rect 53069 16154 53115 16166
rect 53069 15778 53075 16154
rect 53109 15778 53115 16154
rect 53069 15766 53115 15778
rect 51961 15606 52268 15607
rect 52314 15606 52383 15607
rect 53377 15606 53411 16390
rect 51961 15602 52383 15606
rect 51961 15591 52450 15602
rect 53095 15601 53411 15606
rect 51961 15563 52399 15591
rect 51961 15562 52268 15563
rect 51961 15434 51995 15562
rect 52383 15557 52399 15563
rect 52433 15557 52450 15591
rect 52383 15551 52450 15557
rect 53028 15590 53411 15601
rect 53028 15556 53045 15590
rect 53079 15563 53411 15590
rect 53079 15556 53095 15563
rect 53028 15550 53095 15556
rect 52101 15522 52157 15534
rect 53214 15523 53270 15535
rect 53214 15522 53230 15523
rect 52101 15488 52107 15522
rect 52141 15507 52711 15522
rect 52141 15488 52661 15507
rect 52101 15473 52661 15488
rect 52695 15473 52711 15507
rect 52101 15472 52157 15473
rect 52644 15463 52711 15473
rect 52763 15506 53230 15522
rect 52763 15472 52779 15506
rect 52813 15489 53230 15506
rect 53264 15489 53270 15523
rect 52813 15473 53270 15489
rect 52813 15472 52829 15473
rect 52763 15465 52829 15472
rect 53377 15434 53411 15563
rect 53859 15607 53893 16390
rect 54562 16328 54596 16390
rect 54265 16290 55007 16328
rect 53926 16183 53936 16249
rect 53999 16183 54009 16249
rect 54265 16166 54299 16290
rect 54501 16166 54535 16290
rect 54737 16166 54771 16290
rect 54973 16166 55007 16290
rect 54259 16154 54305 16166
rect 54259 15778 54265 16154
rect 54299 15778 54305 16154
rect 54259 15766 54305 15778
rect 54377 16154 54423 16166
rect 54377 15778 54383 16154
rect 54417 15778 54423 16154
rect 54377 15766 54423 15778
rect 54495 16154 54541 16166
rect 54495 15778 54501 16154
rect 54535 15778 54541 16154
rect 54495 15766 54541 15778
rect 54613 16154 54659 16166
rect 54613 15778 54619 16154
rect 54653 15778 54659 16154
rect 54613 15766 54659 15778
rect 54731 16154 54777 16166
rect 54731 15778 54737 16154
rect 54771 15778 54777 16154
rect 54731 15766 54777 15778
rect 54849 16154 54895 16166
rect 54849 15778 54855 16154
rect 54889 15778 54895 16154
rect 54849 15766 54895 15778
rect 54967 16154 55013 16166
rect 54967 15778 54973 16154
rect 55007 15778 55013 16154
rect 54967 15766 55013 15778
rect 53859 15606 54166 15607
rect 55275 15606 55309 16390
rect 56069 16381 56177 16391
rect 56434 16367 56450 16401
rect 56484 16367 56500 16401
rect 56434 16271 56500 16367
rect 56552 16401 56804 16407
rect 56552 16367 56568 16401
rect 56602 16367 56804 16401
rect 56552 16351 56804 16367
rect 56789 16349 56804 16351
rect 56922 16349 56932 16467
rect 56789 16335 56889 16349
rect 56789 16292 56889 16293
rect 57163 16292 57268 17469
rect 56789 16271 57268 16292
rect 56434 16223 57268 16271
rect 56789 16194 57268 16223
rect 56789 16193 56889 16194
rect 57163 16192 57268 16194
rect 57331 16086 57424 17980
rect 57564 17979 57853 17980
rect 57547 17569 57724 17616
rect 57547 17556 57587 17569
rect 57545 17463 57587 17556
rect 57699 17463 57724 17569
rect 57545 17452 57724 17463
rect 57547 17451 57724 17452
rect 58146 16619 58247 18360
rect 59141 18222 59175 18368
rect 59325 18353 59422 18368
rect 59895 18365 59930 18457
rect 59365 18286 59422 18353
rect 59703 18329 59930 18365
rect 59703 18295 59769 18329
rect 59259 18250 59528 18286
rect 59703 18261 59719 18295
rect 59753 18261 59769 18295
rect 59703 18255 59769 18261
rect 59259 18222 59292 18250
rect 59495 18222 59528 18250
rect 59895 18222 59930 18329
rect 59135 18210 59181 18222
rect 59135 18034 59141 18210
rect 59175 18034 59181 18210
rect 59135 18022 59181 18034
rect 59253 18210 59299 18222
rect 59253 18034 59259 18210
rect 59293 18034 59299 18210
rect 59253 18022 59299 18034
rect 59371 18210 59417 18222
rect 59371 18034 59377 18210
rect 59411 18034 59417 18210
rect 59371 18022 59417 18034
rect 59489 18210 59535 18222
rect 59489 18034 59495 18210
rect 59529 18155 59535 18210
rect 59654 18210 59700 18222
rect 59654 18155 59660 18210
rect 59529 18067 59660 18155
rect 59529 18034 59535 18067
rect 59489 18022 59535 18034
rect 59654 18034 59660 18067
rect 59694 18034 59700 18210
rect 59654 18022 59700 18034
rect 59772 18210 59818 18222
rect 59772 18034 59778 18210
rect 59812 18034 59818 18210
rect 59772 18022 59818 18034
rect 59890 18210 59936 18222
rect 59890 18034 59896 18210
rect 59930 18034 59936 18210
rect 59890 18022 59936 18034
rect 60008 18210 60054 18222
rect 60008 18034 60014 18210
rect 60048 18034 60054 18210
rect 60008 18022 60054 18034
rect 59142 17984 59175 18022
rect 59378 17984 59411 18022
rect 59142 17948 59411 17984
rect 59778 17983 59812 18022
rect 60014 17983 60048 18022
rect 59778 17947 60048 17983
rect 59882 17946 60048 17947
rect 59882 17867 60014 17946
rect 59872 17759 59882 17867
rect 60014 17759 60024 17867
rect 60154 17430 60216 19001
rect 60352 18989 60398 19001
rect 60352 18613 60358 18989
rect 60392 18613 60398 18989
rect 60352 18601 60398 18613
rect 60470 18989 60516 19001
rect 60470 18613 60476 18989
rect 60510 18613 60516 18989
rect 60470 18601 60516 18613
rect 60588 18989 60634 19001
rect 60588 18613 60594 18989
rect 60628 18613 60634 18989
rect 60588 18601 60634 18613
rect 60706 18989 60752 19001
rect 60706 18613 60712 18989
rect 60746 18613 60752 18989
rect 60706 18601 60752 18613
rect 60824 18989 60870 19001
rect 60824 18613 60830 18989
rect 60864 18613 60870 18989
rect 60824 18601 60870 18613
rect 60942 18989 60988 19001
rect 60942 18613 60948 18989
rect 60982 18613 60988 18989
rect 60942 18601 60988 18613
rect 61060 18989 61106 19001
rect 61155 18997 61165 19063
rect 61231 18997 61241 19063
rect 61060 18613 61066 18989
rect 61100 18613 61106 18989
rect 61060 18601 61106 18613
rect 60358 18418 60392 18601
rect 60476 18560 60510 18601
rect 60712 18560 60746 18601
rect 60476 18531 60746 18560
rect 60830 18559 60864 18601
rect 61066 18559 61100 18601
rect 60830 18531 61100 18559
rect 61066 18483 61100 18531
rect 61037 18453 61100 18483
rect 62090 18524 62157 19114
rect 62808 19107 62852 19215
rect 62984 19107 63028 19215
rect 62808 19065 63028 19107
rect 62447 19035 63424 19065
rect 62447 18929 62481 19035
rect 62684 18929 62716 19035
rect 62920 18929 62952 19035
rect 63156 18929 63188 19035
rect 63392 18929 63424 19035
rect 62323 18917 62369 18929
rect 62323 18741 62329 18917
rect 62363 18741 62369 18917
rect 62323 18729 62369 18741
rect 62441 18917 62487 18929
rect 62441 18741 62447 18917
rect 62481 18741 62487 18917
rect 62441 18729 62487 18741
rect 62559 18917 62605 18929
rect 62559 18741 62565 18917
rect 62599 18741 62605 18917
rect 62559 18729 62605 18741
rect 62677 18917 62723 18929
rect 62677 18741 62683 18917
rect 62717 18741 62723 18917
rect 62677 18729 62723 18741
rect 62795 18917 62841 18929
rect 62795 18741 62801 18917
rect 62835 18741 62841 18917
rect 62795 18729 62841 18741
rect 62913 18917 62959 18929
rect 62913 18741 62919 18917
rect 62953 18741 62959 18917
rect 62913 18729 62959 18741
rect 63031 18917 63077 18929
rect 63031 18741 63037 18917
rect 63071 18741 63077 18917
rect 63031 18729 63077 18741
rect 63149 18917 63195 18929
rect 63149 18741 63155 18917
rect 63189 18741 63195 18917
rect 63149 18729 63195 18741
rect 63267 18917 63313 18929
rect 63267 18741 63273 18917
rect 63307 18741 63313 18917
rect 63267 18729 63313 18741
rect 63385 18917 63431 18929
rect 63385 18741 63391 18917
rect 63425 18741 63431 18917
rect 63385 18729 63431 18741
rect 62329 18524 62364 18729
rect 62608 18681 62674 18688
rect 62608 18647 62624 18681
rect 62658 18647 62674 18681
rect 62608 18636 62674 18647
rect 62800 18636 62836 18729
rect 62608 18635 62836 18636
rect 63036 18635 63072 18729
rect 63272 18635 63308 18729
rect 62608 18606 63308 18635
rect 62090 18496 62364 18524
rect 62726 18605 63308 18606
rect 62726 18564 62792 18605
rect 62726 18530 62742 18564
rect 62776 18530 62792 18564
rect 62726 18523 62792 18530
rect 62090 18492 62718 18496
rect 63154 18492 63188 18605
rect 62090 18480 62723 18492
rect 62090 18467 62683 18480
rect 60283 18364 60392 18418
rect 60283 18218 60317 18364
rect 60456 18350 60466 18447
rect 60565 18350 60575 18447
rect 61037 18361 61072 18453
rect 60467 18349 60564 18350
rect 60507 18282 60564 18349
rect 60845 18325 61072 18361
rect 60845 18291 60911 18325
rect 60401 18246 60670 18282
rect 60845 18257 60861 18291
rect 60895 18257 60911 18291
rect 60845 18251 60911 18257
rect 60401 18218 60434 18246
rect 60637 18218 60670 18246
rect 61037 18218 61072 18325
rect 62677 18304 62683 18467
rect 62717 18304 62723 18480
rect 62677 18292 62723 18304
rect 62795 18480 62841 18492
rect 62795 18304 62801 18480
rect 62835 18304 62841 18480
rect 62795 18292 62841 18304
rect 62912 18480 62958 18492
rect 60277 18206 60323 18218
rect 60277 18030 60283 18206
rect 60317 18030 60323 18206
rect 60277 18018 60323 18030
rect 60395 18206 60441 18218
rect 60395 18030 60401 18206
rect 60435 18030 60441 18206
rect 60395 18018 60441 18030
rect 60513 18206 60559 18218
rect 60513 18030 60519 18206
rect 60553 18030 60559 18206
rect 60513 18018 60559 18030
rect 60631 18206 60677 18218
rect 60631 18030 60637 18206
rect 60671 18151 60677 18206
rect 60796 18206 60842 18218
rect 60796 18151 60802 18206
rect 60671 18063 60802 18151
rect 60671 18030 60677 18063
rect 60631 18018 60677 18030
rect 60796 18030 60802 18063
rect 60836 18030 60842 18206
rect 60796 18018 60842 18030
rect 60914 18206 60960 18218
rect 60914 18030 60920 18206
rect 60954 18030 60960 18206
rect 60914 18018 60960 18030
rect 61032 18206 61078 18218
rect 61032 18030 61038 18206
rect 61072 18030 61078 18206
rect 61032 18018 61078 18030
rect 61150 18206 61196 18218
rect 61150 18030 61156 18206
rect 61190 18030 61196 18206
rect 62596 18176 62704 18186
rect 62800 18176 62835 18292
rect 62704 18128 62835 18176
rect 62912 18128 62918 18480
rect 62704 18104 62918 18128
rect 62952 18104 62958 18480
rect 62704 18092 62958 18104
rect 63030 18480 63076 18492
rect 63030 18104 63036 18480
rect 63070 18104 63076 18480
rect 63030 18092 63076 18104
rect 63148 18480 63194 18492
rect 63148 18104 63154 18480
rect 63188 18104 63194 18480
rect 63148 18092 63194 18104
rect 64077 18129 64366 18150
rect 62704 18088 62952 18092
rect 62704 18044 62778 18088
rect 64077 18087 64118 18129
rect 63316 18060 64118 18087
rect 62961 18054 63027 18060
rect 62596 18034 62704 18044
rect 61150 18018 61196 18030
rect 62961 18020 62977 18054
rect 63011 18020 63027 18054
rect 60284 17980 60317 18018
rect 60520 17980 60553 18018
rect 60284 17944 60553 17980
rect 60920 17979 60954 18018
rect 61156 17979 61190 18018
rect 60920 17944 61190 17979
rect 60920 17943 61156 17944
rect 61024 17869 61156 17943
rect 62961 17924 63027 18020
rect 63079 18054 64118 18060
rect 63079 18020 63095 18054
rect 63129 18020 64118 18054
rect 63079 18004 64118 18020
rect 63316 17998 64118 18004
rect 64350 17998 64366 18129
rect 63316 17988 64366 17998
rect 63379 17987 64366 17988
rect 63844 17983 64366 17987
rect 63315 17924 63781 17946
rect 62961 17876 63781 17924
rect 61014 17761 61024 17869
rect 61156 17761 61166 17869
rect 63315 17845 63781 17876
rect 63676 17589 63781 17845
rect 60153 17413 60216 17430
rect 62794 17565 63014 17585
rect 62794 17457 62838 17565
rect 62970 17457 63014 17565
rect 63596 17483 63606 17589
rect 63718 17483 63781 17589
rect 63632 17472 63781 17483
rect 62794 17415 63014 17457
rect 60153 17409 60291 17413
rect 60153 17375 62123 17409
rect 62433 17385 63410 17415
rect 60153 17346 62125 17375
rect 60153 17344 60291 17346
rect 62079 17330 62125 17346
rect 59117 17114 59127 17222
rect 59259 17114 59269 17222
rect 61015 17114 61025 17222
rect 61157 17114 61167 17222
rect 59127 17074 59259 17114
rect 61025 17074 61157 17114
rect 59127 17008 59260 17074
rect 61025 17008 61158 17074
rect 58458 16965 59931 17008
rect 58458 16662 58492 16965
rect 58823 16862 58857 16965
rect 59059 16862 59093 16965
rect 59295 16862 59329 16965
rect 59531 16862 59565 16965
rect 58817 16850 58863 16862
rect 57548 16517 58247 16619
rect 58334 16650 58380 16662
rect 57548 16457 57836 16517
rect 58334 16474 58340 16650
rect 58374 16474 58380 16650
rect 58334 16462 58380 16474
rect 58452 16650 58498 16662
rect 58452 16474 58458 16650
rect 58492 16474 58498 16650
rect 58452 16462 58498 16474
rect 58570 16650 58616 16662
rect 58570 16474 58576 16650
rect 58610 16474 58616 16650
rect 58570 16462 58616 16474
rect 58688 16650 58734 16662
rect 58817 16650 58823 16850
rect 58688 16474 58694 16650
rect 58728 16474 58823 16650
rect 58857 16474 58863 16850
rect 58688 16462 58734 16474
rect 58817 16462 58863 16474
rect 58935 16850 58981 16862
rect 58935 16474 58941 16850
rect 58975 16474 58981 16850
rect 58935 16462 58981 16474
rect 59053 16850 59099 16862
rect 59053 16474 59059 16850
rect 59093 16474 59099 16850
rect 59053 16462 59099 16474
rect 59171 16850 59217 16862
rect 59171 16474 59177 16850
rect 59211 16474 59217 16850
rect 59171 16462 59217 16474
rect 59289 16850 59335 16862
rect 59289 16474 59295 16850
rect 59329 16474 59335 16850
rect 59289 16462 59335 16474
rect 59407 16850 59453 16862
rect 59407 16474 59413 16850
rect 59447 16474 59453 16850
rect 59407 16462 59453 16474
rect 59525 16850 59571 16862
rect 59525 16474 59531 16850
rect 59565 16650 59571 16850
rect 59897 16662 59931 16965
rect 60356 16965 61829 17008
rect 60356 16662 60390 16965
rect 60721 16862 60755 16965
rect 60957 16862 60991 16965
rect 61193 16862 61227 16965
rect 61429 16862 61463 16965
rect 60715 16850 60761 16862
rect 59655 16650 59701 16662
rect 59565 16474 59661 16650
rect 59695 16474 59701 16650
rect 59525 16462 59571 16474
rect 59655 16462 59701 16474
rect 59773 16650 59819 16662
rect 59773 16474 59779 16650
rect 59813 16474 59819 16650
rect 59773 16462 59819 16474
rect 59891 16650 59937 16662
rect 59891 16474 59897 16650
rect 59931 16474 59937 16650
rect 59891 16462 59937 16474
rect 60009 16650 60055 16662
rect 60009 16474 60015 16650
rect 60049 16474 60055 16650
rect 60009 16462 60055 16474
rect 60232 16650 60278 16662
rect 60232 16474 60238 16650
rect 60272 16474 60278 16650
rect 60232 16462 60278 16474
rect 60350 16650 60396 16662
rect 60350 16474 60356 16650
rect 60390 16474 60396 16650
rect 60350 16462 60396 16474
rect 60468 16650 60514 16662
rect 60468 16474 60474 16650
rect 60508 16474 60514 16650
rect 60468 16462 60514 16474
rect 60586 16650 60632 16662
rect 60715 16650 60721 16850
rect 60586 16474 60592 16650
rect 60626 16474 60721 16650
rect 60755 16474 60761 16850
rect 60586 16462 60632 16474
rect 60715 16462 60761 16474
rect 60833 16850 60879 16862
rect 60833 16474 60839 16850
rect 60873 16474 60879 16850
rect 60833 16462 60879 16474
rect 60951 16850 60997 16862
rect 60951 16474 60957 16850
rect 60991 16474 60997 16850
rect 60951 16462 60997 16474
rect 61069 16850 61115 16862
rect 61069 16474 61075 16850
rect 61109 16474 61115 16850
rect 61069 16462 61115 16474
rect 61187 16850 61233 16862
rect 61187 16474 61193 16850
rect 61227 16474 61233 16850
rect 61187 16462 61233 16474
rect 61305 16850 61351 16862
rect 61305 16474 61311 16850
rect 61345 16474 61351 16850
rect 61305 16462 61351 16474
rect 61423 16850 61469 16862
rect 61423 16474 61429 16850
rect 61463 16650 61469 16850
rect 61795 16662 61829 16965
rect 62079 16878 62126 17330
rect 62433 17279 62467 17385
rect 62670 17279 62702 17385
rect 62906 17279 62938 17385
rect 63142 17279 63174 17385
rect 63378 17279 63410 17385
rect 62309 17267 62355 17279
rect 62309 17091 62315 17267
rect 62349 17091 62355 17267
rect 62309 17079 62355 17091
rect 62427 17267 62473 17279
rect 62427 17091 62433 17267
rect 62467 17091 62473 17267
rect 62427 17079 62473 17091
rect 62545 17267 62591 17279
rect 62545 17091 62551 17267
rect 62585 17091 62591 17267
rect 62545 17079 62591 17091
rect 62663 17267 62709 17279
rect 62663 17091 62669 17267
rect 62703 17091 62709 17267
rect 62663 17079 62709 17091
rect 62781 17267 62827 17279
rect 62781 17091 62787 17267
rect 62821 17091 62827 17267
rect 62781 17079 62827 17091
rect 62899 17267 62945 17279
rect 62899 17091 62905 17267
rect 62939 17091 62945 17267
rect 62899 17079 62945 17091
rect 63017 17267 63063 17279
rect 63017 17091 63023 17267
rect 63057 17091 63063 17267
rect 63017 17079 63063 17091
rect 63135 17267 63181 17279
rect 63135 17091 63141 17267
rect 63175 17091 63181 17267
rect 63135 17079 63181 17091
rect 63253 17267 63299 17279
rect 63253 17091 63259 17267
rect 63293 17091 63299 17267
rect 63253 17079 63299 17091
rect 63371 17267 63417 17279
rect 63371 17091 63377 17267
rect 63411 17091 63417 17267
rect 63371 17079 63417 17091
rect 62080 16862 62126 16878
rect 62080 16861 62161 16862
rect 62315 16861 62350 17079
rect 62594 17031 62660 17038
rect 62594 16997 62610 17031
rect 62644 16997 62660 17031
rect 62594 16986 62660 16997
rect 62786 16986 62822 17079
rect 62594 16985 62822 16986
rect 63022 16985 63058 17079
rect 63258 16985 63294 17079
rect 62594 16956 63294 16985
rect 62712 16955 63294 16956
rect 62712 16914 62778 16955
rect 62712 16880 62728 16914
rect 62762 16880 62778 16914
rect 62712 16873 62778 16880
rect 62080 16846 62350 16861
rect 62080 16842 62704 16846
rect 63140 16842 63174 16955
rect 62080 16830 62709 16842
rect 62080 16818 62669 16830
rect 62080 16816 62161 16818
rect 62427 16817 62669 16818
rect 61553 16650 61599 16662
rect 61463 16474 61559 16650
rect 61593 16474 61599 16650
rect 61423 16462 61469 16474
rect 61553 16462 61599 16474
rect 61671 16650 61717 16662
rect 61671 16474 61677 16650
rect 61711 16474 61717 16650
rect 61671 16462 61717 16474
rect 61789 16650 61835 16662
rect 61789 16474 61795 16650
rect 61829 16474 61835 16650
rect 61789 16462 61835 16474
rect 61907 16650 61953 16662
rect 61907 16474 61913 16650
rect 61947 16474 61953 16650
rect 62663 16654 62669 16817
rect 62703 16654 62709 16830
rect 62663 16642 62709 16654
rect 62781 16830 62827 16842
rect 62781 16654 62787 16830
rect 62821 16654 62827 16830
rect 62781 16642 62827 16654
rect 62898 16830 62944 16842
rect 61907 16462 61953 16474
rect 62582 16526 62690 16536
rect 62786 16526 62821 16642
rect 57548 16455 57588 16457
rect 57548 16444 57582 16455
rect 57547 16349 57582 16444
rect 57700 16351 57836 16457
rect 58340 16428 58374 16462
rect 58576 16428 58610 16462
rect 58340 16393 58610 16428
rect 59177 16428 59211 16462
rect 59413 16428 59447 16462
rect 60015 16428 60049 16462
rect 59177 16393 59447 16428
rect 59890 16393 60049 16428
rect 60238 16428 60272 16462
rect 60474 16428 60508 16462
rect 60238 16393 60508 16428
rect 61075 16428 61109 16462
rect 61311 16428 61345 16462
rect 61913 16428 61947 16462
rect 61075 16393 61345 16428
rect 61788 16393 61947 16428
rect 62690 16478 62821 16526
rect 62898 16478 62904 16830
rect 62690 16454 62904 16478
rect 62938 16454 62944 16830
rect 62690 16442 62944 16454
rect 63016 16830 63062 16842
rect 63016 16454 63022 16830
rect 63056 16454 63062 16830
rect 63016 16442 63062 16454
rect 63134 16830 63180 16842
rect 63134 16454 63140 16830
rect 63174 16454 63180 16830
rect 63134 16442 63180 16454
rect 62690 16438 62938 16442
rect 63307 16438 63317 16470
rect 62690 16394 62764 16438
rect 63302 16410 63317 16438
rect 62947 16404 63013 16410
rect 57694 16349 57836 16351
rect 57547 16340 57836 16349
rect 57548 16339 57836 16340
rect 57580 16338 57836 16339
rect 58326 16215 58393 16239
rect 58326 16181 58342 16215
rect 58376 16181 58393 16215
rect 57322 16007 57332 16086
rect 57425 16007 57435 16086
rect 56286 15958 56506 15978
rect 56286 15850 56330 15958
rect 56462 15850 56506 15958
rect 56286 15808 56506 15850
rect 55925 15778 56902 15808
rect 55925 15672 55959 15778
rect 56162 15672 56194 15778
rect 56398 15672 56430 15778
rect 56634 15672 56666 15778
rect 56870 15672 56902 15778
rect 53859 15601 54279 15606
rect 54993 15601 55309 15606
rect 53859 15590 54346 15601
rect 53859 15563 54295 15590
rect 53859 15562 54166 15563
rect 53859 15434 53893 15562
rect 54279 15556 54295 15563
rect 54329 15556 54346 15590
rect 54279 15550 54346 15556
rect 54926 15590 55309 15601
rect 54926 15556 54943 15590
rect 54977 15563 55309 15590
rect 54977 15556 54993 15563
rect 54926 15550 54993 15556
rect 53999 15522 54055 15534
rect 55112 15523 55168 15535
rect 55112 15522 55128 15523
rect 53999 15488 54005 15522
rect 54039 15507 54609 15522
rect 54039 15488 54559 15507
rect 53999 15473 54559 15488
rect 54593 15473 54609 15507
rect 53999 15472 54055 15473
rect 54542 15463 54609 15473
rect 54661 15506 55128 15522
rect 54661 15472 54677 15506
rect 54711 15489 55128 15506
rect 55162 15489 55168 15523
rect 54711 15473 55168 15489
rect 54711 15472 54727 15473
rect 54661 15465 54727 15472
rect 55275 15434 55309 15563
rect 55801 15660 55847 15672
rect 55801 15484 55807 15660
rect 55841 15484 55847 15660
rect 55801 15472 55847 15484
rect 55919 15660 55965 15672
rect 55919 15484 55925 15660
rect 55959 15484 55965 15660
rect 55919 15472 55965 15484
rect 56037 15660 56083 15672
rect 56037 15484 56043 15660
rect 56077 15484 56083 15660
rect 56037 15472 56083 15484
rect 56155 15660 56201 15672
rect 56155 15484 56161 15660
rect 56195 15484 56201 15660
rect 56155 15472 56201 15484
rect 56273 15660 56319 15672
rect 56273 15484 56279 15660
rect 56313 15484 56319 15660
rect 56273 15472 56319 15484
rect 56391 15660 56437 15672
rect 56391 15484 56397 15660
rect 56431 15484 56437 15660
rect 56391 15472 56437 15484
rect 56509 15660 56555 15672
rect 56509 15484 56515 15660
rect 56549 15484 56555 15660
rect 56509 15472 56555 15484
rect 56627 15660 56673 15672
rect 56627 15484 56633 15660
rect 56667 15484 56673 15660
rect 56627 15472 56673 15484
rect 56745 15660 56791 15672
rect 56745 15484 56751 15660
rect 56785 15484 56791 15660
rect 56745 15472 56791 15484
rect 56863 15660 56909 15672
rect 56863 15484 56869 15660
rect 56903 15484 56909 15660
rect 56863 15472 56909 15484
rect 51955 15422 52001 15434
rect 51955 15246 51961 15422
rect 51995 15246 52001 15422
rect 51955 15234 52001 15246
rect 52073 15422 52119 15434
rect 52073 15246 52079 15422
rect 52113 15246 52119 15422
rect 52073 15234 52119 15246
rect 52479 15422 52525 15434
rect 52080 14940 52113 15234
rect 52479 15046 52485 15422
rect 52519 15046 52525 15422
rect 52479 15034 52525 15046
rect 52597 15422 52643 15434
rect 52597 15046 52603 15422
rect 52637 15046 52643 15422
rect 52597 15034 52643 15046
rect 52715 15422 52761 15434
rect 52715 15046 52721 15422
rect 52755 15046 52761 15422
rect 52715 15034 52761 15046
rect 52833 15422 52879 15434
rect 52833 15046 52839 15422
rect 52873 15046 52879 15422
rect 52833 15034 52879 15046
rect 52951 15422 52997 15434
rect 52951 15046 52957 15422
rect 52991 15046 52997 15422
rect 53253 15422 53299 15434
rect 53253 15246 53259 15422
rect 53293 15246 53299 15422
rect 53253 15234 53299 15246
rect 53371 15422 53417 15434
rect 53371 15246 53377 15422
rect 53411 15246 53417 15422
rect 53371 15234 53417 15246
rect 53853 15422 53899 15434
rect 53853 15246 53859 15422
rect 53893 15246 53899 15422
rect 53853 15234 53899 15246
rect 53971 15422 54017 15434
rect 53971 15246 53977 15422
rect 54011 15246 54017 15422
rect 53971 15234 54017 15246
rect 54377 15422 54423 15434
rect 52951 15034 52997 15046
rect 52603 14940 52637 15034
rect 53260 14940 53294 15234
rect 52080 14908 53294 14940
rect 53978 14940 54011 15234
rect 54377 15046 54383 15422
rect 54417 15046 54423 15422
rect 54377 15034 54423 15046
rect 54495 15422 54541 15434
rect 54495 15046 54501 15422
rect 54535 15046 54541 15422
rect 54495 15034 54541 15046
rect 54613 15422 54659 15434
rect 54613 15046 54619 15422
rect 54653 15046 54659 15422
rect 54613 15034 54659 15046
rect 54731 15422 54777 15434
rect 54731 15046 54737 15422
rect 54771 15046 54777 15422
rect 54731 15034 54777 15046
rect 54849 15422 54895 15434
rect 54849 15046 54855 15422
rect 54889 15046 54895 15422
rect 55151 15422 55197 15434
rect 55151 15246 55157 15422
rect 55191 15246 55197 15422
rect 55151 15234 55197 15246
rect 55269 15422 55315 15434
rect 55269 15246 55275 15422
rect 55309 15246 55315 15422
rect 55269 15234 55315 15246
rect 55807 15239 55842 15472
rect 56086 15424 56152 15431
rect 56086 15390 56102 15424
rect 56136 15390 56152 15424
rect 56086 15379 56152 15390
rect 56278 15379 56314 15472
rect 56086 15378 56314 15379
rect 56514 15378 56550 15472
rect 56750 15378 56786 15472
rect 56086 15349 56786 15378
rect 56204 15348 56786 15349
rect 56204 15307 56270 15348
rect 56204 15273 56220 15307
rect 56254 15273 56270 15307
rect 56204 15266 56270 15273
rect 55807 15235 56196 15239
rect 56632 15235 56666 15348
rect 54849 15034 54895 15046
rect 54501 14940 54535 15034
rect 55158 14940 55192 15234
rect 55807 15223 56201 15235
rect 55807 15210 56161 15223
rect 55807 15207 55885 15210
rect 55802 15155 55812 15207
rect 55875 15155 55885 15207
rect 55807 15149 55880 15155
rect 56155 15047 56161 15210
rect 56195 15047 56201 15223
rect 56155 15035 56201 15047
rect 56273 15223 56319 15235
rect 56273 15047 56279 15223
rect 56313 15047 56319 15223
rect 56273 15035 56319 15047
rect 56390 15223 56436 15235
rect 53978 14908 55192 14940
rect 56074 14919 56182 14929
rect 56278 14919 56313 15035
rect 52669 14823 52801 14908
rect 54567 14823 54699 14908
rect 51814 14516 51880 14795
rect 52659 14715 52669 14823
rect 52801 14715 52811 14823
rect 54557 14715 54567 14823
rect 54699 14715 54709 14823
rect 56182 14871 56313 14919
rect 56390 14871 56396 15223
rect 56182 14847 56396 14871
rect 56430 14847 56436 15223
rect 56182 14835 56436 14847
rect 56508 15223 56554 15235
rect 56508 14847 56514 15223
rect 56548 14847 56554 15223
rect 56508 14835 56554 14847
rect 56626 15223 56672 15235
rect 56626 14847 56632 15223
rect 56666 14847 56672 15223
rect 56626 14835 56672 14847
rect 56182 14831 56430 14835
rect 57331 14833 57424 16007
rect 56839 14831 57424 14833
rect 56182 14787 56256 14831
rect 56794 14803 57424 14831
rect 56439 14797 56505 14803
rect 56074 14777 56182 14787
rect 56439 14763 56455 14797
rect 56489 14763 56505 14797
rect 56439 14667 56505 14763
rect 56557 14797 57424 14803
rect 56557 14763 56573 14797
rect 56607 14763 57424 14797
rect 56557 14747 57424 14763
rect 56794 14731 57424 14747
rect 56839 14727 57424 14731
rect 57323 14726 57424 14727
rect 58109 15752 58265 15758
rect 58109 15654 58121 15752
rect 58253 15654 58265 15752
rect 56794 14678 56894 14689
rect 56794 14667 56808 14678
rect 56439 14619 56808 14667
rect 56440 14516 56506 14619
rect 56794 14589 56808 14619
rect 56798 14572 56808 14589
rect 56920 14572 56930 14678
rect 51814 14436 56508 14516
rect 58109 13981 58265 15654
rect 58326 14798 58393 16181
rect 58474 15610 58508 16393
rect 59177 16331 59211 16393
rect 58880 16293 59622 16331
rect 58880 16169 58914 16293
rect 59116 16169 59150 16293
rect 59352 16169 59386 16293
rect 59588 16169 59622 16293
rect 58874 16157 58920 16169
rect 58874 15781 58880 16157
rect 58914 15781 58920 16157
rect 58874 15769 58920 15781
rect 58992 16157 59038 16169
rect 58992 15781 58998 16157
rect 59032 15781 59038 16157
rect 58992 15769 59038 15781
rect 59110 16157 59156 16169
rect 59110 15781 59116 16157
rect 59150 15781 59156 16157
rect 59110 15769 59156 15781
rect 59228 16157 59274 16169
rect 59228 15781 59234 16157
rect 59268 15781 59274 16157
rect 59228 15769 59274 15781
rect 59346 16157 59392 16169
rect 59346 15781 59352 16157
rect 59386 15781 59392 16157
rect 59346 15769 59392 15781
rect 59464 16157 59510 16169
rect 59464 15781 59470 16157
rect 59504 15781 59510 16157
rect 59464 15769 59510 15781
rect 59582 16157 59628 16169
rect 59582 15781 59588 16157
rect 59622 15781 59628 16157
rect 59582 15769 59628 15781
rect 58474 15609 58781 15610
rect 58827 15609 58896 15610
rect 59890 15609 59924 16393
rect 58474 15605 58896 15609
rect 58474 15594 58963 15605
rect 59608 15604 59924 15609
rect 58474 15566 58912 15594
rect 58474 15565 58781 15566
rect 58474 15437 58508 15565
rect 58896 15560 58912 15566
rect 58946 15560 58963 15594
rect 58896 15554 58963 15560
rect 59541 15593 59924 15604
rect 59541 15559 59558 15593
rect 59592 15566 59924 15593
rect 59592 15559 59608 15566
rect 59541 15553 59608 15559
rect 58614 15525 58670 15537
rect 59727 15526 59783 15538
rect 59727 15525 59743 15526
rect 58614 15491 58620 15525
rect 58654 15510 59224 15525
rect 58654 15491 59174 15510
rect 58614 15476 59174 15491
rect 59208 15476 59224 15510
rect 58614 15475 58670 15476
rect 59157 15466 59224 15476
rect 59276 15509 59743 15525
rect 59276 15475 59292 15509
rect 59326 15492 59743 15509
rect 59777 15492 59783 15526
rect 59326 15476 59783 15492
rect 59326 15475 59342 15476
rect 59276 15468 59342 15475
rect 59890 15437 59924 15566
rect 60372 15610 60406 16393
rect 61075 16331 61109 16393
rect 60778 16293 61520 16331
rect 60439 16186 60449 16252
rect 60512 16186 60522 16252
rect 60778 16169 60812 16293
rect 61014 16169 61048 16293
rect 61250 16169 61284 16293
rect 61486 16169 61520 16293
rect 60772 16157 60818 16169
rect 60772 15781 60778 16157
rect 60812 15781 60818 16157
rect 60772 15769 60818 15781
rect 60890 16157 60936 16169
rect 60890 15781 60896 16157
rect 60930 15781 60936 16157
rect 60890 15769 60936 15781
rect 61008 16157 61054 16169
rect 61008 15781 61014 16157
rect 61048 15781 61054 16157
rect 61008 15769 61054 15781
rect 61126 16157 61172 16169
rect 61126 15781 61132 16157
rect 61166 15781 61172 16157
rect 61126 15769 61172 15781
rect 61244 16157 61290 16169
rect 61244 15781 61250 16157
rect 61284 15781 61290 16157
rect 61244 15769 61290 15781
rect 61362 16157 61408 16169
rect 61362 15781 61368 16157
rect 61402 15781 61408 16157
rect 61362 15769 61408 15781
rect 61480 16157 61526 16169
rect 61480 15781 61486 16157
rect 61520 15781 61526 16157
rect 61480 15769 61526 15781
rect 60372 15609 60679 15610
rect 61788 15609 61822 16393
rect 62582 16384 62690 16394
rect 62947 16370 62963 16404
rect 62997 16370 63013 16404
rect 62947 16274 63013 16370
rect 63065 16404 63317 16410
rect 63065 16370 63081 16404
rect 63115 16370 63317 16404
rect 63065 16354 63317 16370
rect 63302 16352 63317 16354
rect 63435 16352 63445 16470
rect 63302 16338 63402 16352
rect 63302 16295 63402 16296
rect 63676 16295 63781 17472
rect 63302 16274 63781 16295
rect 62947 16226 63781 16274
rect 63302 16197 63781 16226
rect 63302 16196 63402 16197
rect 63676 16195 63781 16197
rect 63844 16089 63937 17983
rect 64653 16624 64780 22931
rect 68599 22315 71306 22316
rect 68599 22300 71403 22315
rect 68599 22235 68618 22300
rect 68701 22235 71403 22300
rect 68599 22222 71403 22235
rect 71319 22204 71403 22222
rect 71319 22147 71327 22204
rect 71395 22147 71403 22204
rect 71319 22145 71403 22147
rect 71487 22204 71571 22225
rect 71487 22147 71495 22204
rect 71563 22147 71571 22204
rect 71487 22145 71571 22147
rect 71327 22137 71395 22145
rect 71495 22137 71563 22145
rect 70713 22062 70913 22067
rect 70713 22061 71723 22062
rect 70713 22027 70725 22061
rect 70901 22027 71723 22061
rect 70713 22021 70913 22027
rect 70713 21943 70913 21949
rect 70713 21909 70725 21943
rect 70901 21909 70913 21943
rect 70713 21903 70913 21909
rect 70713 21825 70913 21831
rect 70713 21791 70725 21825
rect 70901 21791 70913 21825
rect 70713 21785 70913 21791
rect 70713 21707 70913 21713
rect 70713 21673 70725 21707
rect 70901 21673 70913 21707
rect 70713 21626 70913 21673
rect 70513 21620 70913 21626
rect 70369 21586 70525 21620
rect 70901 21586 70913 21620
rect 64272 16622 64780 16624
rect 64061 16468 64780 16622
rect 65902 21342 66076 21353
rect 65902 21264 65917 21342
rect 66062 21264 66076 21342
rect 64061 16460 64349 16468
rect 64061 16458 64101 16460
rect 64061 16447 64095 16458
rect 64060 16352 64095 16447
rect 64213 16354 64349 16460
rect 64207 16352 64349 16354
rect 64060 16343 64349 16352
rect 64061 16342 64349 16343
rect 64093 16341 64349 16342
rect 63835 16010 63845 16089
rect 63938 16010 63948 16089
rect 62799 15961 63019 15981
rect 62799 15853 62843 15961
rect 62975 15853 63019 15961
rect 62799 15811 63019 15853
rect 62438 15781 63415 15811
rect 62438 15675 62472 15781
rect 62675 15675 62707 15781
rect 62911 15675 62943 15781
rect 63147 15675 63179 15781
rect 63383 15675 63415 15781
rect 60372 15604 60792 15609
rect 61506 15604 61822 15609
rect 60372 15593 60859 15604
rect 60372 15566 60808 15593
rect 60372 15565 60679 15566
rect 60372 15437 60406 15565
rect 60792 15559 60808 15566
rect 60842 15559 60859 15593
rect 60792 15553 60859 15559
rect 61439 15593 61822 15604
rect 61439 15559 61456 15593
rect 61490 15566 61822 15593
rect 61490 15559 61506 15566
rect 61439 15553 61506 15559
rect 60512 15525 60568 15537
rect 61625 15526 61681 15538
rect 61625 15525 61641 15526
rect 60512 15491 60518 15525
rect 60552 15510 61122 15525
rect 60552 15491 61072 15510
rect 60512 15476 61072 15491
rect 61106 15476 61122 15510
rect 60512 15475 60568 15476
rect 61055 15466 61122 15476
rect 61174 15509 61641 15525
rect 61174 15475 61190 15509
rect 61224 15492 61641 15509
rect 61675 15492 61681 15526
rect 61224 15476 61681 15492
rect 61224 15475 61240 15476
rect 61174 15468 61240 15475
rect 61788 15437 61822 15566
rect 62314 15663 62360 15675
rect 62314 15487 62320 15663
rect 62354 15487 62360 15663
rect 62314 15475 62360 15487
rect 62432 15663 62478 15675
rect 62432 15487 62438 15663
rect 62472 15487 62478 15663
rect 62432 15475 62478 15487
rect 62550 15663 62596 15675
rect 62550 15487 62556 15663
rect 62590 15487 62596 15663
rect 62550 15475 62596 15487
rect 62668 15663 62714 15675
rect 62668 15487 62674 15663
rect 62708 15487 62714 15663
rect 62668 15475 62714 15487
rect 62786 15663 62832 15675
rect 62786 15487 62792 15663
rect 62826 15487 62832 15663
rect 62786 15475 62832 15487
rect 62904 15663 62950 15675
rect 62904 15487 62910 15663
rect 62944 15487 62950 15663
rect 62904 15475 62950 15487
rect 63022 15663 63068 15675
rect 63022 15487 63028 15663
rect 63062 15487 63068 15663
rect 63022 15475 63068 15487
rect 63140 15663 63186 15675
rect 63140 15487 63146 15663
rect 63180 15487 63186 15663
rect 63140 15475 63186 15487
rect 63258 15663 63304 15675
rect 63258 15487 63264 15663
rect 63298 15487 63304 15663
rect 63258 15475 63304 15487
rect 63376 15663 63422 15675
rect 63376 15487 63382 15663
rect 63416 15487 63422 15663
rect 63376 15475 63422 15487
rect 58468 15425 58514 15437
rect 58468 15249 58474 15425
rect 58508 15249 58514 15425
rect 58468 15237 58514 15249
rect 58586 15425 58632 15437
rect 58586 15249 58592 15425
rect 58626 15249 58632 15425
rect 58586 15237 58632 15249
rect 58992 15425 59038 15437
rect 58593 14943 58626 15237
rect 58992 15049 58998 15425
rect 59032 15049 59038 15425
rect 58992 15037 59038 15049
rect 59110 15425 59156 15437
rect 59110 15049 59116 15425
rect 59150 15049 59156 15425
rect 59110 15037 59156 15049
rect 59228 15425 59274 15437
rect 59228 15049 59234 15425
rect 59268 15049 59274 15425
rect 59228 15037 59274 15049
rect 59346 15425 59392 15437
rect 59346 15049 59352 15425
rect 59386 15049 59392 15425
rect 59346 15037 59392 15049
rect 59464 15425 59510 15437
rect 59464 15049 59470 15425
rect 59504 15049 59510 15425
rect 59766 15425 59812 15437
rect 59766 15249 59772 15425
rect 59806 15249 59812 15425
rect 59766 15237 59812 15249
rect 59884 15425 59930 15437
rect 59884 15249 59890 15425
rect 59924 15249 59930 15425
rect 59884 15237 59930 15249
rect 60366 15425 60412 15437
rect 60366 15249 60372 15425
rect 60406 15249 60412 15425
rect 60366 15237 60412 15249
rect 60484 15425 60530 15437
rect 60484 15249 60490 15425
rect 60524 15249 60530 15425
rect 60484 15237 60530 15249
rect 60890 15425 60936 15437
rect 59464 15037 59510 15049
rect 59116 14943 59150 15037
rect 59773 14943 59807 15237
rect 58593 14911 59807 14943
rect 60491 14943 60524 15237
rect 60890 15049 60896 15425
rect 60930 15049 60936 15425
rect 60890 15037 60936 15049
rect 61008 15425 61054 15437
rect 61008 15049 61014 15425
rect 61048 15049 61054 15425
rect 61008 15037 61054 15049
rect 61126 15425 61172 15437
rect 61126 15049 61132 15425
rect 61166 15049 61172 15425
rect 61126 15037 61172 15049
rect 61244 15425 61290 15437
rect 61244 15049 61250 15425
rect 61284 15049 61290 15425
rect 61244 15037 61290 15049
rect 61362 15425 61408 15437
rect 61362 15049 61368 15425
rect 61402 15049 61408 15425
rect 61664 15425 61710 15437
rect 61664 15249 61670 15425
rect 61704 15249 61710 15425
rect 61664 15237 61710 15249
rect 61782 15425 61828 15437
rect 61782 15249 61788 15425
rect 61822 15249 61828 15425
rect 61782 15237 61828 15249
rect 62320 15242 62355 15475
rect 62599 15427 62665 15434
rect 62599 15393 62615 15427
rect 62649 15393 62665 15427
rect 62599 15382 62665 15393
rect 62791 15382 62827 15475
rect 62599 15381 62827 15382
rect 63027 15381 63063 15475
rect 63263 15381 63299 15475
rect 62599 15352 63299 15381
rect 62717 15351 63299 15352
rect 62717 15310 62783 15351
rect 62717 15276 62733 15310
rect 62767 15276 62783 15310
rect 62717 15269 62783 15276
rect 62320 15238 62709 15242
rect 63145 15238 63179 15351
rect 61362 15037 61408 15049
rect 61014 14943 61048 15037
rect 61671 14943 61705 15237
rect 62320 15226 62714 15238
rect 62320 15213 62674 15226
rect 62320 15210 62398 15213
rect 62315 15158 62325 15210
rect 62388 15158 62398 15210
rect 62320 15152 62393 15158
rect 62668 15050 62674 15213
rect 62708 15050 62714 15226
rect 62668 15038 62714 15050
rect 62786 15226 62832 15238
rect 62786 15050 62792 15226
rect 62826 15050 62832 15226
rect 62786 15038 62832 15050
rect 62903 15226 62949 15238
rect 60491 14911 61705 14943
rect 62587 14922 62695 14932
rect 62791 14922 62826 15038
rect 59182 14826 59314 14911
rect 61080 14826 61212 14911
rect 58327 14519 58393 14798
rect 59172 14718 59182 14826
rect 59314 14718 59324 14826
rect 61070 14718 61080 14826
rect 61212 14718 61222 14826
rect 62695 14874 62826 14922
rect 62903 14874 62909 15226
rect 62695 14850 62909 14874
rect 62943 14850 62949 15226
rect 62695 14838 62949 14850
rect 63021 15226 63067 15238
rect 63021 14850 63027 15226
rect 63061 14850 63067 15226
rect 63021 14838 63067 14850
rect 63139 15226 63185 15238
rect 63139 14850 63145 15226
rect 63179 14850 63185 15226
rect 63139 14838 63185 14850
rect 62695 14834 62943 14838
rect 63844 14836 63937 16010
rect 65902 15575 66076 21264
rect 70369 20823 70426 21586
rect 70513 21580 70913 21586
rect 70513 21502 70913 21508
rect 70513 21468 70525 21502
rect 70901 21468 70913 21502
rect 70513 21462 70913 21468
rect 70513 21384 70913 21390
rect 70513 21350 70525 21384
rect 70901 21350 70913 21384
rect 70513 21344 70913 21350
rect 70513 21266 70913 21272
rect 70513 21232 70525 21266
rect 70901 21232 70913 21266
rect 70513 21226 70913 21232
rect 70513 21153 70913 21159
rect 70513 21119 70525 21153
rect 70901 21119 71039 21153
rect 70513 21113 70913 21119
rect 70513 21035 70913 21041
rect 70513 21001 70525 21035
rect 70901 21001 70913 21035
rect 70513 20995 70913 21001
rect 70513 20917 70913 20923
rect 70513 20883 70525 20917
rect 70901 20883 70913 20917
rect 70513 20877 70913 20883
rect 70269 20813 70426 20823
rect 70329 20733 70426 20813
rect 70513 20799 70913 20805
rect 70513 20765 70525 20799
rect 70901 20765 70913 20799
rect 70513 20759 70913 20765
rect 70269 20723 70426 20733
rect 70369 20445 70426 20723
rect 70513 20681 70913 20687
rect 70513 20647 70525 20681
rect 70901 20647 70913 20681
rect 70513 20641 70913 20647
rect 70513 20563 70913 20569
rect 70513 20529 70525 20563
rect 70901 20529 70913 20563
rect 70513 20523 70913 20529
rect 70513 20445 70913 20451
rect 70369 20411 70525 20445
rect 70901 20411 70913 20445
rect 66419 19962 66589 19976
rect 66419 19890 66434 19962
rect 66569 19890 66589 19962
rect 66419 19882 66589 19890
rect 66419 16045 66587 19882
rect 70369 19854 70426 20411
rect 70513 20405 70913 20411
rect 70513 20326 70913 20332
rect 70513 20292 70525 20326
rect 70901 20292 70913 20326
rect 70513 20286 70913 20292
rect 70513 20208 70913 20214
rect 70513 20174 70525 20208
rect 70901 20174 70913 20208
rect 70513 20168 70913 20174
rect 70513 20090 70913 20096
rect 70513 20056 70525 20090
rect 70901 20056 70913 20090
rect 70513 20050 70913 20056
rect 70513 19972 70913 19978
rect 70997 19972 71039 21119
rect 71099 20975 71166 22027
rect 71199 21960 71284 21972
rect 71199 21889 71212 21960
rect 71275 21889 71284 21960
rect 71199 21880 71284 21889
rect 71676 21228 71723 22027
rect 71846 21228 72046 21233
rect 71676 21227 72046 21228
rect 71676 21194 71858 21227
rect 71099 20941 71116 20975
rect 71150 20941 71166 20975
rect 71099 20925 71166 20941
rect 71487 20993 71572 21005
rect 71487 20925 71495 20993
rect 71560 20925 71572 20993
rect 71487 20913 71572 20925
rect 71202 20875 71287 20887
rect 71202 20805 71212 20875
rect 71274 20805 71287 20875
rect 71202 20795 71287 20805
rect 71676 20756 71723 21194
rect 71846 21193 71858 21194
rect 72034 21193 72046 21227
rect 71846 21187 72046 21193
rect 71846 21109 72046 21115
rect 71846 21075 71858 21109
rect 72034 21075 72465 21109
rect 71846 21041 72046 21075
rect 71846 21035 72246 21041
rect 71846 21001 71858 21035
rect 72234 21001 72246 21035
rect 71846 20995 72246 21001
rect 71846 20917 72246 20923
rect 71846 20883 71858 20917
rect 72234 20883 72246 20917
rect 71846 20877 72246 20883
rect 71846 20799 72246 20805
rect 72319 20799 72385 20814
rect 71846 20765 71858 20799
rect 72234 20798 72385 20799
rect 72234 20765 72335 20798
rect 71846 20759 72246 20765
rect 72319 20764 72335 20765
rect 72369 20764 72385 20798
rect 71676 20740 71786 20756
rect 72319 20748 72385 20764
rect 72413 20811 72465 21075
rect 72413 20799 72543 20811
rect 71676 20706 71736 20740
rect 71770 20706 71786 20740
rect 71676 20690 71786 20706
rect 72413 20733 72487 20799
rect 72539 20733 72543 20799
rect 72413 20719 72543 20733
rect 71846 20681 72246 20687
rect 71846 20647 71858 20681
rect 72234 20647 72246 20681
rect 71846 20641 72246 20647
rect 71326 20634 71398 20640
rect 71326 20575 71332 20634
rect 71392 20575 71398 20634
rect 71329 20571 71396 20575
rect 71332 20565 71392 20571
rect 71846 20563 72246 20569
rect 71846 20529 71858 20563
rect 72234 20529 72246 20563
rect 71846 20523 72246 20529
rect 71846 20485 72046 20523
rect 72413 20485 72465 20719
rect 71846 20451 71858 20485
rect 72034 20451 72465 20485
rect 71846 20445 72046 20451
rect 71675 20367 71722 20368
rect 71846 20367 72046 20373
rect 71675 20333 71858 20367
rect 72034 20333 72046 20367
rect 70513 19938 70525 19972
rect 70901 19938 71125 19972
rect 70513 19932 70913 19938
rect 70713 19854 70913 19859
rect 70369 19853 70913 19854
rect 69651 19830 69776 19831
rect 67059 19829 69776 19830
rect 66988 19812 69776 19829
rect 70369 19819 70725 19853
rect 70901 19819 70913 19853
rect 70369 19817 70913 19819
rect 70713 19813 70913 19817
rect 66988 19722 67002 19812
rect 67132 19722 69776 19812
rect 66988 19703 69776 19722
rect 67059 19701 69776 19703
rect 69651 19170 69776 19701
rect 70713 19735 70913 19741
rect 70713 19701 70725 19735
rect 70901 19701 70913 19735
rect 70713 19695 70913 19701
rect 71059 19665 71125 19938
rect 71059 19631 71075 19665
rect 71109 19631 71125 19665
rect 70713 19617 70913 19623
rect 70713 19583 70725 19617
rect 70901 19583 70913 19617
rect 71059 19615 71125 19631
rect 70713 19577 70913 19583
rect 70713 19499 70913 19505
rect 71675 19499 71722 20333
rect 71846 20327 72046 20333
rect 70713 19465 70725 19499
rect 70901 19467 71722 19499
rect 70901 19466 71802 19467
rect 72926 19466 74819 19467
rect 70901 19465 74819 19466
rect 70713 19464 74819 19465
rect 70713 19459 70913 19464
rect 71267 19318 74819 19464
rect 71363 19316 74819 19318
rect 72926 19315 74819 19316
rect 68254 19159 68315 19161
rect 68238 19076 68248 19159
rect 68316 19076 68326 19159
rect 69651 19083 71403 19170
rect 68254 19074 68315 19076
rect 71319 19060 71403 19083
rect 71319 19003 71327 19060
rect 71395 19003 71403 19060
rect 71319 19001 71403 19003
rect 71487 19060 71571 19082
rect 71487 19003 71495 19060
rect 71563 19003 71571 19060
rect 71487 19001 71571 19003
rect 71327 18993 71395 19001
rect 71495 18993 71563 19001
rect 70713 18918 70913 18923
rect 70713 18917 71723 18918
rect 70713 18883 70725 18917
rect 70901 18883 71723 18917
rect 70713 18877 70913 18883
rect 70713 18799 70913 18805
rect 70713 18765 70725 18799
rect 70901 18765 70913 18799
rect 70713 18759 70913 18765
rect 70713 18681 70913 18687
rect 70713 18647 70725 18681
rect 70901 18647 70913 18681
rect 70713 18641 70913 18647
rect 70713 18563 70913 18569
rect 70713 18529 70725 18563
rect 70901 18529 70913 18563
rect 70713 18482 70913 18529
rect 70513 18476 70913 18482
rect 70369 18442 70525 18476
rect 70901 18442 70913 18476
rect 70369 17679 70426 18442
rect 70513 18436 70913 18442
rect 70513 18358 70913 18364
rect 70513 18324 70525 18358
rect 70901 18324 70913 18358
rect 70513 18318 70913 18324
rect 70513 18240 70913 18246
rect 70513 18206 70525 18240
rect 70901 18206 70913 18240
rect 70513 18200 70913 18206
rect 70513 18122 70913 18128
rect 70513 18088 70525 18122
rect 70901 18088 70913 18122
rect 70513 18082 70913 18088
rect 70513 18009 70913 18015
rect 70513 17975 70525 18009
rect 70901 17975 71039 18009
rect 70513 17969 70913 17975
rect 70513 17891 70913 17897
rect 70513 17857 70525 17891
rect 70901 17857 70913 17891
rect 70513 17851 70913 17857
rect 70513 17773 70913 17779
rect 70513 17739 70525 17773
rect 70901 17739 70913 17773
rect 70513 17733 70913 17739
rect 70269 17669 70426 17679
rect 70329 17589 70426 17669
rect 70513 17655 70913 17661
rect 70513 17621 70525 17655
rect 70901 17621 70913 17655
rect 70513 17615 70913 17621
rect 70269 17579 70426 17589
rect 70369 17301 70426 17579
rect 70513 17537 70913 17543
rect 70513 17503 70525 17537
rect 70901 17503 70913 17537
rect 70513 17497 70913 17503
rect 70513 17419 70913 17425
rect 70513 17385 70525 17419
rect 70901 17385 70913 17419
rect 70513 17379 70913 17385
rect 70513 17301 70913 17307
rect 70369 17267 70525 17301
rect 70901 17267 70913 17301
rect 70369 16710 70426 17267
rect 70513 17261 70913 17267
rect 70513 17182 70913 17188
rect 70513 17148 70525 17182
rect 70901 17148 70913 17182
rect 70513 17142 70913 17148
rect 70513 17064 70913 17070
rect 70513 17030 70525 17064
rect 70901 17030 70913 17064
rect 70513 17024 70913 17030
rect 70513 16946 70913 16952
rect 70513 16912 70525 16946
rect 70901 16912 70913 16946
rect 70513 16906 70913 16912
rect 70513 16828 70913 16834
rect 70997 16828 71039 17975
rect 71099 17831 71166 18883
rect 71199 18816 71284 18828
rect 71199 18745 71212 18816
rect 71275 18745 71284 18816
rect 71199 18736 71284 18745
rect 71676 18084 71723 18883
rect 71846 18084 72046 18089
rect 71676 18083 72046 18084
rect 71676 18050 71858 18083
rect 71099 17797 71116 17831
rect 71150 17797 71166 17831
rect 71099 17781 71166 17797
rect 71487 17849 71572 17861
rect 71487 17781 71495 17849
rect 71560 17781 71572 17849
rect 71487 17769 71572 17781
rect 71202 17731 71287 17743
rect 71202 17661 71212 17731
rect 71274 17661 71287 17731
rect 71202 17651 71287 17661
rect 71676 17612 71723 18050
rect 71846 18049 71858 18050
rect 72034 18049 72046 18083
rect 71846 18043 72046 18049
rect 71846 17965 72046 17971
rect 71846 17931 71858 17965
rect 72034 17931 72465 17965
rect 71846 17897 72046 17931
rect 71846 17891 72246 17897
rect 71846 17857 71858 17891
rect 72234 17857 72246 17891
rect 71846 17851 72246 17857
rect 71846 17773 72246 17779
rect 71846 17739 71858 17773
rect 72234 17739 72246 17773
rect 71846 17733 72246 17739
rect 71846 17655 72246 17661
rect 72319 17655 72385 17670
rect 71846 17621 71858 17655
rect 72234 17654 72385 17655
rect 72234 17621 72335 17654
rect 71846 17615 72246 17621
rect 72319 17620 72335 17621
rect 72369 17620 72385 17654
rect 71676 17596 71786 17612
rect 72319 17604 72385 17620
rect 72413 17667 72465 17931
rect 72413 17655 72543 17667
rect 71676 17562 71736 17596
rect 71770 17562 71786 17596
rect 71676 17546 71786 17562
rect 72413 17589 72487 17655
rect 72539 17589 72543 17655
rect 72413 17575 72543 17589
rect 71846 17537 72246 17543
rect 71846 17503 71858 17537
rect 72234 17503 72246 17537
rect 71846 17497 72246 17503
rect 71326 17490 71398 17496
rect 71326 17431 71332 17490
rect 71392 17431 71398 17490
rect 71329 17427 71396 17431
rect 71332 17421 71392 17427
rect 71846 17419 72246 17425
rect 71846 17385 71858 17419
rect 72234 17385 72246 17419
rect 71846 17379 72246 17385
rect 71846 17341 72046 17379
rect 72413 17341 72465 17575
rect 71846 17307 71858 17341
rect 72034 17307 72465 17341
rect 71846 17301 72046 17307
rect 71675 17223 71722 17224
rect 71846 17223 72046 17229
rect 71675 17189 71858 17223
rect 72034 17189 72046 17223
rect 70513 16794 70525 16828
rect 70901 16794 71125 16828
rect 70513 16788 70913 16794
rect 70713 16710 70913 16715
rect 70369 16709 70913 16710
rect 70369 16675 70725 16709
rect 70901 16675 70913 16709
rect 70369 16673 70913 16675
rect 70713 16669 70913 16673
rect 70713 16591 70913 16597
rect 70713 16557 70725 16591
rect 70901 16557 70913 16591
rect 70713 16551 70913 16557
rect 71059 16521 71125 16794
rect 71059 16487 71075 16521
rect 71109 16487 71125 16521
rect 70713 16473 70913 16479
rect 70713 16439 70725 16473
rect 70901 16439 70913 16473
rect 71059 16471 71125 16487
rect 70713 16433 70913 16439
rect 70713 16355 70913 16361
rect 71675 16355 71722 17189
rect 71846 17183 72046 17189
rect 70713 16321 70725 16355
rect 70901 16325 71722 16355
rect 72963 16325 73355 16326
rect 74502 16325 74653 16326
rect 70901 16324 71812 16325
rect 72946 16324 74653 16325
rect 70901 16321 74653 16324
rect 70713 16320 74653 16321
rect 70713 16315 70913 16320
rect 71267 16175 74653 16320
rect 71267 16174 71413 16175
rect 71723 16174 74653 16175
rect 72946 16173 74653 16174
rect 66419 15967 71400 16045
rect 66420 15945 71400 15967
rect 66420 15943 67299 15945
rect 71315 15928 71399 15945
rect 71315 15871 71323 15928
rect 71391 15871 71399 15928
rect 71315 15869 71399 15871
rect 71483 15928 71567 15946
rect 71483 15871 71491 15928
rect 71559 15871 71567 15928
rect 71483 15869 71567 15871
rect 71323 15861 71391 15869
rect 71491 15861 71559 15869
rect 70709 15786 70909 15791
rect 70709 15785 71719 15786
rect 70709 15751 70721 15785
rect 70897 15751 71719 15785
rect 70709 15745 70909 15751
rect 70709 15667 70909 15673
rect 70709 15633 70721 15667
rect 70897 15633 70909 15667
rect 70709 15627 70909 15633
rect 65902 15422 69655 15575
rect 70709 15549 70909 15555
rect 70709 15515 70721 15549
rect 70897 15515 70909 15549
rect 70709 15509 70909 15515
rect 66008 15421 69655 15422
rect 63352 14834 63937 14836
rect 62695 14790 62769 14834
rect 63307 14806 63937 14834
rect 62952 14800 63018 14806
rect 62587 14780 62695 14790
rect 62952 14766 62968 14800
rect 63002 14766 63018 14800
rect 62952 14670 63018 14766
rect 63070 14800 63937 14806
rect 63070 14766 63086 14800
rect 63120 14766 63937 14800
rect 63070 14750 63937 14766
rect 63307 14734 63937 14750
rect 63352 14730 63937 14734
rect 63836 14729 63937 14730
rect 63307 14681 63407 14692
rect 63307 14670 63321 14681
rect 62952 14622 63321 14670
rect 62953 14519 63019 14622
rect 63307 14592 63321 14622
rect 63311 14575 63321 14592
rect 63433 14575 63443 14681
rect 58327 14439 63021 14519
rect 58109 13901 69192 13981
rect 68976 13866 69056 13867
rect 51596 13783 69056 13866
rect 45062 13682 68934 13755
rect 38504 13546 68803 13652
rect 38552 13545 68803 13546
rect 66033 13542 68803 13545
rect 64415 13513 64538 13514
rect 64234 13512 64538 13513
rect 33810 13505 64538 13512
rect 33810 13504 64375 13505
rect 33810 13415 64365 13504
rect 33810 13414 64375 13415
rect 64526 13414 64538 13505
rect 33810 13401 64538 13414
rect 64415 13399 64538 13401
rect 68714 13507 68803 13542
rect 33672 13359 56089 13360
rect 33672 13346 58019 13359
rect 33672 13258 57855 13346
rect 58004 13258 58019 13346
rect 33672 13249 58019 13258
rect 54005 13248 58019 13249
rect 57599 13246 58019 13248
rect 33542 13199 51496 13209
rect 33542 13111 51328 13199
rect 51484 13111 51496 13199
rect 33542 13098 51496 13111
rect 57721 13089 57731 13164
rect 57817 13089 57827 13164
rect 33409 13039 44901 13053
rect 33409 12942 44758 13039
rect 44887 12942 44901 13039
rect 51198 12973 51208 13043
rect 51295 12973 51305 13043
rect 33409 12932 44901 12942
rect 36058 12876 68659 12877
rect 33244 12865 68659 12876
rect 33244 12784 68502 12865
rect 68646 12784 68659 12865
rect 33244 12774 68659 12784
rect 33244 12773 65941 12774
rect 44623 12649 44633 12710
rect 44726 12649 44736 12710
rect 62686 12599 68655 12707
rect 62686 12445 62799 12599
rect 68536 12588 68655 12599
rect 62869 12503 68495 12571
rect 55078 12395 55214 12415
rect 41875 12375 42011 12395
rect 41875 12313 41911 12375
rect 41971 12313 42011 12375
rect 41875 12285 42011 12313
rect 48424 12374 48560 12394
rect 48424 12312 48460 12374
rect 48520 12312 48560 12374
rect 41571 12255 42548 12285
rect 48424 12284 48560 12312
rect 55078 12333 55114 12395
rect 55174 12333 55214 12395
rect 55078 12305 55214 12333
rect 41571 12149 41603 12255
rect 41807 12149 41839 12255
rect 42043 12149 42075 12255
rect 42279 12149 42311 12255
rect 42514 12149 42548 12255
rect 48120 12254 49097 12284
rect 41564 12137 41610 12149
rect 41564 11961 41570 12137
rect 41604 11961 41610 12137
rect 41564 11949 41610 11961
rect 41682 12137 41728 12149
rect 41682 11961 41688 12137
rect 41722 11961 41728 12137
rect 41682 11949 41728 11961
rect 41800 12137 41846 12149
rect 41800 11961 41806 12137
rect 41840 11961 41846 12137
rect 41800 11949 41846 11961
rect 41918 12137 41964 12149
rect 41918 11961 41924 12137
rect 41958 11961 41964 12137
rect 41918 11949 41964 11961
rect 42036 12137 42082 12149
rect 42036 11961 42042 12137
rect 42076 11961 42082 12137
rect 42036 11949 42082 11961
rect 42154 12137 42200 12149
rect 42154 11961 42160 12137
rect 42194 11961 42200 12137
rect 42154 11949 42200 11961
rect 42272 12137 42318 12149
rect 42272 11961 42278 12137
rect 42312 11961 42318 12137
rect 42272 11949 42318 11961
rect 42390 12137 42436 12149
rect 42390 11961 42396 12137
rect 42430 11961 42436 12137
rect 42390 11949 42436 11961
rect 42508 12137 42554 12149
rect 42508 11961 42514 12137
rect 42548 11961 42554 12137
rect 42508 11949 42554 11961
rect 42626 12137 42672 12149
rect 48120 12148 48152 12254
rect 48356 12148 48388 12254
rect 48592 12148 48624 12254
rect 48828 12148 48860 12254
rect 49063 12148 49097 12254
rect 54774 12275 55751 12305
rect 54774 12169 54806 12275
rect 55010 12169 55042 12275
rect 55246 12169 55278 12275
rect 55482 12169 55514 12275
rect 55717 12169 55751 12275
rect 54767 12157 54813 12169
rect 42626 11961 42632 12137
rect 42666 11961 42672 12137
rect 42626 11949 42672 11961
rect 48113 12136 48159 12148
rect 48113 11960 48119 12136
rect 48153 11960 48159 12136
rect 41687 11855 41723 11949
rect 41923 11855 41959 11949
rect 42159 11856 42195 11949
rect 42321 11901 42387 11908
rect 42321 11867 42337 11901
rect 42371 11867 42387 11901
rect 42321 11856 42387 11867
rect 42159 11855 42387 11856
rect 41687 11826 42387 11855
rect 41687 11825 42269 11826
rect 41807 11712 41841 11825
rect 42203 11784 42269 11825
rect 42203 11750 42219 11784
rect 42253 11750 42269 11784
rect 42203 11743 42269 11750
rect 42631 11718 42666 11949
rect 48113 11948 48159 11960
rect 48231 12136 48277 12148
rect 48231 11960 48237 12136
rect 48271 11960 48277 12136
rect 48231 11948 48277 11960
rect 48349 12136 48395 12148
rect 48349 11960 48355 12136
rect 48389 11960 48395 12136
rect 48349 11948 48395 11960
rect 48467 12136 48513 12148
rect 48467 11960 48473 12136
rect 48507 11960 48513 12136
rect 48467 11948 48513 11960
rect 48585 12136 48631 12148
rect 48585 11960 48591 12136
rect 48625 11960 48631 12136
rect 48585 11948 48631 11960
rect 48703 12136 48749 12148
rect 48703 11960 48709 12136
rect 48743 11960 48749 12136
rect 48703 11948 48749 11960
rect 48821 12136 48867 12148
rect 48821 11960 48827 12136
rect 48861 11960 48867 12136
rect 48821 11948 48867 11960
rect 48939 12136 48985 12148
rect 48939 11960 48945 12136
rect 48979 11960 48985 12136
rect 48939 11948 48985 11960
rect 49057 12136 49103 12148
rect 49057 11960 49063 12136
rect 49097 11960 49103 12136
rect 49057 11948 49103 11960
rect 49175 12136 49221 12148
rect 49175 11960 49181 12136
rect 49215 11960 49221 12136
rect 54767 11981 54773 12157
rect 54807 11981 54813 12157
rect 54767 11969 54813 11981
rect 54885 12157 54931 12169
rect 54885 11981 54891 12157
rect 54925 11981 54931 12157
rect 54885 11969 54931 11981
rect 55003 12157 55049 12169
rect 55003 11981 55009 12157
rect 55043 11981 55049 12157
rect 55003 11969 55049 11981
rect 55121 12157 55167 12169
rect 55121 11981 55127 12157
rect 55161 11981 55167 12157
rect 55121 11969 55167 11981
rect 55239 12157 55285 12169
rect 55239 11981 55245 12157
rect 55279 11981 55285 12157
rect 55239 11969 55285 11981
rect 55357 12157 55403 12169
rect 55357 11981 55363 12157
rect 55397 11981 55403 12157
rect 55357 11969 55403 11981
rect 55475 12157 55521 12169
rect 55475 11981 55481 12157
rect 55515 11981 55521 12157
rect 55475 11969 55521 11981
rect 55593 12157 55639 12169
rect 55593 11981 55599 12157
rect 55633 11981 55639 12157
rect 55593 11969 55639 11981
rect 55711 12157 55757 12169
rect 55711 11981 55717 12157
rect 55751 11981 55757 12157
rect 55711 11969 55757 11981
rect 55829 12157 55875 12169
rect 55829 11981 55835 12157
rect 55869 11981 55875 12157
rect 55829 11969 55875 11981
rect 49175 11948 49221 11960
rect 48236 11854 48272 11948
rect 48472 11854 48508 11948
rect 48708 11855 48744 11948
rect 48870 11900 48936 11907
rect 48870 11866 48886 11900
rect 48920 11866 48936 11900
rect 48870 11855 48936 11866
rect 48708 11854 48936 11855
rect 48236 11825 48936 11854
rect 48236 11824 48818 11825
rect 42561 11716 43878 11718
rect 42277 11712 43878 11716
rect 41801 11700 41847 11712
rect 41801 11324 41807 11700
rect 41841 11324 41847 11700
rect 41801 11312 41847 11324
rect 41919 11700 41965 11712
rect 41919 11324 41925 11700
rect 41959 11324 41965 11700
rect 41919 11312 41965 11324
rect 42037 11700 42083 11712
rect 42037 11324 42043 11700
rect 42077 11351 42083 11700
rect 42154 11700 42200 11712
rect 42154 11524 42160 11700
rect 42194 11524 42200 11700
rect 42154 11517 42200 11524
rect 42272 11700 43878 11712
rect 48356 11711 48390 11824
rect 48752 11783 48818 11824
rect 48752 11749 48768 11783
rect 48802 11749 48818 11783
rect 48752 11742 48818 11749
rect 49180 11750 49215 11948
rect 54890 11875 54926 11969
rect 55126 11875 55162 11969
rect 55362 11876 55398 11969
rect 55524 11921 55590 11928
rect 55524 11887 55540 11921
rect 55574 11887 55590 11921
rect 55524 11876 55590 11887
rect 55362 11875 55590 11876
rect 54890 11846 55590 11875
rect 54890 11845 55472 11846
rect 49180 11715 49216 11750
rect 55010 11732 55044 11845
rect 55406 11804 55472 11845
rect 55406 11770 55422 11804
rect 55456 11770 55472 11804
rect 55406 11763 55472 11770
rect 55834 11736 55869 11969
rect 55480 11732 57154 11736
rect 55004 11720 55050 11732
rect 48826 11711 50528 11715
rect 42272 11524 42278 11700
rect 42312 11687 43878 11700
rect 42312 11524 42318 11687
rect 42561 11606 43878 11687
rect 42154 11512 42203 11517
rect 42272 11512 42318 11524
rect 42160 11351 42203 11512
rect 42077 11324 42203 11351
rect 42037 11312 42203 11324
rect 42043 11308 42203 11312
rect 41548 11274 41916 11280
rect 41548 11240 41866 11274
rect 41900 11240 41916 11274
rect 41548 11224 41916 11240
rect 41968 11274 42034 11280
rect 41968 11240 41984 11274
rect 42018 11240 42034 11274
rect 33097 11105 33107 11159
rect 33164 11105 33174 11159
rect 33097 9103 33172 11105
rect 41548 11032 41627 11224
rect 41968 11195 42034 11240
rect 33961 11022 41627 11032
rect 33961 10972 33985 11022
rect 34046 10972 41627 11022
rect 33961 10962 41627 10972
rect 41685 11187 42034 11195
rect 41685 11155 42035 11187
rect 42127 11171 42203 11308
rect 41685 10861 41739 11155
rect 42123 11111 42133 11171
rect 42195 11111 42205 11171
rect 41682 10849 41743 10861
rect 33812 10840 33987 10846
rect 33812 10784 33824 10840
rect 33883 10837 33987 10840
rect 33883 10784 33893 10837
rect 33812 10779 33893 10784
rect 33977 10779 33987 10837
rect 41682 10795 41688 10849
rect 41737 10795 41743 10849
rect 41682 10783 41743 10795
rect 33812 10778 33987 10779
rect 35211 10475 35347 10495
rect 34126 10452 34207 10455
rect 34121 10400 34131 10452
rect 34199 10400 34209 10452
rect 35211 10413 35247 10475
rect 35307 10413 35347 10475
rect 34126 10398 34207 10400
rect 35211 10385 35347 10413
rect 40747 10435 40826 10447
rect 38265 10385 38344 10397
rect 34907 10355 35884 10385
rect 34907 10249 34939 10355
rect 35143 10249 35175 10355
rect 35379 10249 35411 10355
rect 35615 10249 35647 10355
rect 35850 10249 35884 10355
rect 38265 10288 38271 10385
rect 38193 10268 38271 10288
rect 38338 10288 38344 10385
rect 40747 10322 40753 10435
rect 40820 10322 40826 10435
rect 41889 10437 41968 10449
rect 41889 10322 41895 10437
rect 41962 10322 41968 10437
rect 38338 10268 38413 10288
rect 34900 10237 34946 10249
rect 34900 10061 34906 10237
rect 34940 10061 34946 10237
rect 34900 10049 34946 10061
rect 35018 10237 35064 10249
rect 35018 10061 35024 10237
rect 35058 10061 35064 10237
rect 35018 10049 35064 10061
rect 35136 10237 35182 10249
rect 35136 10061 35142 10237
rect 35176 10061 35182 10237
rect 35136 10049 35182 10061
rect 35254 10237 35300 10249
rect 35254 10061 35260 10237
rect 35294 10061 35300 10237
rect 35254 10049 35300 10061
rect 35372 10237 35418 10249
rect 35372 10061 35378 10237
rect 35412 10061 35418 10237
rect 35372 10049 35418 10061
rect 35490 10237 35536 10249
rect 35490 10061 35496 10237
rect 35530 10061 35536 10237
rect 35490 10049 35536 10061
rect 35608 10237 35654 10249
rect 35608 10061 35614 10237
rect 35648 10061 35654 10237
rect 35608 10049 35654 10061
rect 35726 10237 35772 10249
rect 35726 10061 35732 10237
rect 35766 10061 35772 10237
rect 35726 10049 35772 10061
rect 35844 10237 35890 10249
rect 35844 10061 35850 10237
rect 35884 10061 35890 10237
rect 35844 10049 35890 10061
rect 35962 10237 36008 10249
rect 35962 10061 35968 10237
rect 36002 10061 36008 10237
rect 38193 10160 38237 10268
rect 38369 10160 38413 10268
rect 39990 10226 40046 10234
rect 38193 10118 38413 10160
rect 39064 10218 40046 10226
rect 39064 10184 40006 10218
rect 40040 10184 40046 10218
rect 40709 10214 40719 10322
rect 40851 10259 40861 10322
rect 40851 10248 40863 10259
rect 40851 10214 40864 10248
rect 41120 10238 41176 10240
rect 39064 10168 40046 10184
rect 40719 10176 40864 10214
rect 39064 10167 40043 10168
rect 35962 10049 36008 10061
rect 37797 10088 38774 10118
rect 35023 9955 35059 10049
rect 35259 9955 35295 10049
rect 35495 9956 35531 10049
rect 35657 10001 35723 10008
rect 35657 9967 35673 10001
rect 35707 9967 35723 10001
rect 35657 9956 35723 9967
rect 35495 9955 35723 9956
rect 35023 9926 35723 9955
rect 35023 9925 35605 9926
rect 35143 9812 35177 9925
rect 35539 9884 35605 9925
rect 35539 9850 35555 9884
rect 35589 9850 35605 9884
rect 35539 9843 35605 9850
rect 35967 9816 36002 10049
rect 37797 9982 37829 10088
rect 38033 9982 38065 10088
rect 38269 9982 38301 10088
rect 38505 9982 38537 10088
rect 38740 9982 38774 10088
rect 35613 9812 36002 9816
rect 35137 9800 35183 9812
rect 33763 9495 35097 9510
rect 33763 9425 33781 9495
rect 33855 9493 35097 9495
rect 33855 9425 34403 9493
rect 33763 9417 34403 9425
rect 34492 9417 35097 9493
rect 33763 9410 35097 9417
rect 35137 9424 35143 9800
rect 35177 9424 35183 9800
rect 35137 9412 35183 9424
rect 35255 9800 35301 9812
rect 35255 9424 35261 9800
rect 35295 9424 35301 9800
rect 35255 9412 35301 9424
rect 35373 9800 35419 9812
rect 35373 9424 35379 9800
rect 35413 9451 35419 9800
rect 35490 9800 35536 9812
rect 35490 9624 35496 9800
rect 35530 9624 35536 9800
rect 35490 9617 35536 9624
rect 35608 9800 36002 9812
rect 35608 9624 35614 9800
rect 35648 9787 36002 9800
rect 35648 9624 35654 9787
rect 35490 9612 35539 9617
rect 35608 9612 35654 9624
rect 35496 9451 35539 9612
rect 35413 9424 35539 9451
rect 35373 9412 35539 9424
rect 35021 9380 35075 9410
rect 35379 9408 35539 9412
rect 35021 9374 35252 9380
rect 35021 9340 35202 9374
rect 35236 9340 35252 9374
rect 33762 9318 34965 9330
rect 35021 9324 35252 9340
rect 35304 9374 35370 9380
rect 35304 9340 35320 9374
rect 35354 9340 35370 9374
rect 33762 9239 33775 9318
rect 33763 9226 33775 9239
rect 33865 9315 34965 9318
rect 33865 9231 33965 9315
rect 34078 9299 34965 9315
rect 34078 9255 34897 9299
rect 34953 9295 34965 9299
rect 35304 9295 35370 9340
rect 34953 9287 35370 9295
rect 34953 9255 35371 9287
rect 35463 9271 35539 9408
rect 34078 9231 34966 9255
rect 33865 9226 34966 9231
rect 33763 9219 34966 9226
rect 35459 9211 35469 9271
rect 35531 9211 35541 9271
rect 35898 9143 36002 9787
rect 37790 9970 37836 9982
rect 37790 9794 37796 9970
rect 37830 9794 37836 9970
rect 37790 9782 37836 9794
rect 37908 9970 37954 9982
rect 37908 9794 37914 9970
rect 37948 9794 37954 9970
rect 37908 9782 37954 9794
rect 38026 9970 38072 9982
rect 38026 9794 38032 9970
rect 38066 9794 38072 9970
rect 38026 9782 38072 9794
rect 38144 9970 38190 9982
rect 38144 9794 38150 9970
rect 38184 9794 38190 9970
rect 38144 9782 38190 9794
rect 38262 9970 38308 9982
rect 38262 9794 38268 9970
rect 38302 9794 38308 9970
rect 38262 9782 38308 9794
rect 38380 9970 38426 9982
rect 38380 9794 38386 9970
rect 38420 9794 38426 9970
rect 38380 9782 38426 9794
rect 38498 9970 38544 9982
rect 38498 9794 38504 9970
rect 38538 9794 38544 9970
rect 38498 9782 38544 9794
rect 38616 9970 38662 9982
rect 38616 9794 38622 9970
rect 38656 9794 38662 9970
rect 38616 9782 38662 9794
rect 38734 9970 38780 9982
rect 38734 9794 38740 9970
rect 38774 9794 38780 9970
rect 38734 9782 38780 9794
rect 38852 9970 38898 9982
rect 38852 9794 38858 9970
rect 38892 9794 38898 9970
rect 38852 9782 38898 9794
rect 37913 9688 37949 9782
rect 38149 9688 38185 9782
rect 38385 9689 38421 9782
rect 38547 9734 38613 9741
rect 38547 9700 38563 9734
rect 38597 9700 38613 9734
rect 38547 9689 38613 9700
rect 38385 9688 38613 9689
rect 37913 9659 38613 9688
rect 37913 9658 38495 9659
rect 38033 9545 38067 9658
rect 38429 9617 38495 9658
rect 38429 9583 38445 9617
rect 38479 9583 38495 9617
rect 38429 9576 38495 9583
rect 38857 9577 38892 9782
rect 39064 9577 39131 10167
rect 40823 10144 40864 10176
rect 41110 10172 41120 10238
rect 41176 10172 41186 10238
rect 41856 10214 41866 10322
rect 41998 10259 42008 10322
rect 41998 10248 42010 10259
rect 41998 10214 42011 10248
rect 41866 10176 42011 10214
rect 41970 10148 42011 10176
rect 40239 10116 40509 10144
rect 39980 10050 39990 10116
rect 40056 10050 40066 10116
rect 40239 10054 40273 10116
rect 40475 10054 40509 10116
rect 40593 10116 40864 10144
rect 41381 10120 41651 10148
rect 40593 10054 40627 10116
rect 40829 10054 40864 10116
rect 41005 10104 41176 10120
rect 41005 10070 41136 10104
rect 41170 10070 41176 10104
rect 41005 10054 41176 10070
rect 41381 10058 41415 10120
rect 41617 10058 41651 10120
rect 41735 10120 42011 10148
rect 41735 10058 41769 10120
rect 41971 10058 42011 10120
rect 40115 10042 40161 10054
rect 40115 9666 40121 10042
rect 40155 9666 40161 10042
rect 40115 9654 40161 9666
rect 40233 10042 40279 10054
rect 40233 9666 40239 10042
rect 40273 9666 40279 10042
rect 40233 9654 40279 9666
rect 40351 10042 40397 10054
rect 40351 9666 40357 10042
rect 40391 9666 40397 10042
rect 40351 9654 40397 9666
rect 40469 10042 40515 10054
rect 40469 9666 40475 10042
rect 40509 9666 40515 10042
rect 40469 9654 40515 9666
rect 40587 10042 40633 10054
rect 40587 9666 40593 10042
rect 40627 9666 40633 10042
rect 40587 9654 40633 9666
rect 40705 10042 40751 10054
rect 40705 9666 40711 10042
rect 40745 9666 40751 10042
rect 40705 9654 40751 9666
rect 40823 10042 40869 10054
rect 40823 9666 40829 10042
rect 40863 9666 40869 10042
rect 40823 9654 40869 9666
rect 38857 9549 39131 9577
rect 38503 9545 39131 9549
rect 38027 9533 38073 9545
rect 38027 9157 38033 9533
rect 38067 9157 38073 9533
rect 38027 9145 38073 9157
rect 38145 9533 38191 9545
rect 38145 9157 38151 9533
rect 38185 9157 38191 9533
rect 38145 9145 38191 9157
rect 38263 9533 38309 9545
rect 38263 9157 38269 9533
rect 38303 9181 38309 9533
rect 38380 9533 38426 9545
rect 38380 9357 38386 9533
rect 38420 9357 38426 9533
rect 38380 9345 38426 9357
rect 38498 9533 39131 9545
rect 38498 9357 38504 9533
rect 38538 9520 39131 9533
rect 40121 9612 40155 9654
rect 40357 9612 40391 9654
rect 40121 9584 40391 9612
rect 40475 9613 40509 9654
rect 40711 9613 40745 9654
rect 40475 9584 40745 9613
rect 40121 9536 40155 9584
rect 38538 9357 38544 9520
rect 40121 9506 40184 9536
rect 38498 9345 38544 9357
rect 40149 9414 40184 9506
rect 40149 9378 40376 9414
rect 40646 9403 40656 9500
rect 40755 9403 40765 9500
rect 40829 9471 40863 9654
rect 40829 9417 40938 9471
rect 38386 9229 38421 9345
rect 40149 9271 40184 9378
rect 40310 9344 40376 9378
rect 40310 9310 40326 9344
rect 40360 9310 40376 9344
rect 40657 9402 40754 9403
rect 40657 9335 40714 9402
rect 40310 9304 40376 9310
rect 40551 9299 40820 9335
rect 40551 9271 40584 9299
rect 40787 9271 40820 9299
rect 40904 9271 40938 9417
rect 40025 9259 40071 9271
rect 38517 9229 38625 9239
rect 38386 9181 38517 9229
rect 38625 9196 38773 9202
rect 38303 9157 38517 9181
rect 38263 9145 38517 9157
rect 35898 9142 36005 9143
rect 35898 9141 36594 9142
rect 38269 9141 38517 9145
rect 35898 9140 37144 9141
rect 35898 9113 37905 9140
rect 35898 9107 38142 9113
rect 33093 9042 33103 9103
rect 33166 9042 33176 9103
rect 35898 9073 38092 9107
rect 38126 9073 38142 9107
rect 35898 9057 38142 9073
rect 38194 9107 38260 9113
rect 38194 9073 38210 9107
rect 38244 9073 38260 9107
rect 38443 9097 38517 9141
rect 38761 9129 38773 9196
rect 38625 9123 38773 9129
rect 38517 9087 38625 9097
rect 33097 7039 33172 9042
rect 35898 9041 37905 9057
rect 35898 9040 37842 9041
rect 35898 9036 37377 9040
rect 35898 9035 37144 9036
rect 35898 9033 36985 9035
rect 36187 8625 37161 8654
rect 36187 8519 37009 8625
rect 37121 8612 37161 8625
rect 37121 8519 37163 8612
rect 36187 8508 37163 8519
rect 36187 8507 37161 8508
rect 35203 7890 35339 7910
rect 35203 7828 35239 7890
rect 35299 7828 35339 7890
rect 35203 7800 35339 7828
rect 34899 7770 35876 7800
rect 34899 7664 34931 7770
rect 35135 7664 35167 7770
rect 35371 7664 35403 7770
rect 35607 7664 35639 7770
rect 35842 7664 35876 7770
rect 34892 7652 34938 7664
rect 34892 7476 34898 7652
rect 34932 7476 34938 7652
rect 34892 7464 34938 7476
rect 35010 7652 35056 7664
rect 35010 7476 35016 7652
rect 35050 7476 35056 7652
rect 35010 7464 35056 7476
rect 35128 7652 35174 7664
rect 35128 7476 35134 7652
rect 35168 7476 35174 7652
rect 35128 7464 35174 7476
rect 35246 7652 35292 7664
rect 35246 7476 35252 7652
rect 35286 7476 35292 7652
rect 35246 7464 35292 7476
rect 35364 7652 35410 7664
rect 35364 7476 35370 7652
rect 35404 7476 35410 7652
rect 35364 7464 35410 7476
rect 35482 7652 35528 7664
rect 35482 7476 35488 7652
rect 35522 7476 35528 7652
rect 35482 7464 35528 7476
rect 35600 7652 35646 7664
rect 35600 7476 35606 7652
rect 35640 7476 35646 7652
rect 35600 7464 35646 7476
rect 35718 7652 35764 7664
rect 35718 7476 35724 7652
rect 35758 7476 35764 7652
rect 35718 7464 35764 7476
rect 35836 7652 35882 7664
rect 35836 7476 35842 7652
rect 35876 7476 35882 7652
rect 35836 7464 35882 7476
rect 35954 7652 36000 7664
rect 35954 7476 35960 7652
rect 35994 7476 36000 7652
rect 35954 7464 36000 7476
rect 35015 7370 35051 7464
rect 35251 7370 35287 7464
rect 35487 7371 35523 7464
rect 35649 7416 35715 7423
rect 35649 7382 35665 7416
rect 35699 7382 35715 7416
rect 35649 7371 35715 7382
rect 35487 7370 35715 7371
rect 35015 7341 35715 7370
rect 35015 7340 35597 7341
rect 35135 7227 35169 7340
rect 35531 7299 35597 7340
rect 35531 7265 35547 7299
rect 35581 7265 35597 7299
rect 35531 7258 35597 7265
rect 35959 7231 35994 7464
rect 36187 7231 36307 8507
rect 36979 7514 37160 7544
rect 36979 7404 37008 7514
rect 37126 7500 37160 7514
rect 37126 7404 37161 7500
rect 36979 7396 37161 7404
rect 36979 7394 37160 7396
rect 35605 7227 36307 7231
rect 35129 7215 35175 7227
rect 33093 6978 33103 7039
rect 33166 6978 33176 7039
rect 33097 4974 33172 6978
rect 35129 6839 35135 7215
rect 35169 6839 35175 7215
rect 35129 6827 35175 6839
rect 35247 7215 35293 7227
rect 35247 6839 35253 7215
rect 35287 6839 35293 7215
rect 35247 6827 35293 6839
rect 35365 7215 35411 7227
rect 35365 6839 35371 7215
rect 35405 6866 35411 7215
rect 35482 7215 35528 7227
rect 35482 7039 35488 7215
rect 35522 7039 35528 7215
rect 35482 7032 35528 7039
rect 35600 7215 36307 7227
rect 35600 7039 35606 7215
rect 35640 7202 36307 7215
rect 35640 7039 35646 7202
rect 35890 7123 36307 7202
rect 37284 7142 37377 9036
rect 37440 8977 37906 8999
rect 38194 8977 38260 9073
rect 40025 9083 40031 9259
rect 40065 9083 40071 9259
rect 40025 9071 40071 9083
rect 40143 9259 40189 9271
rect 40143 9083 40149 9259
rect 40183 9083 40189 9259
rect 40143 9071 40189 9083
rect 40261 9259 40307 9271
rect 40261 9083 40267 9259
rect 40301 9083 40307 9259
rect 40261 9071 40307 9083
rect 40379 9259 40425 9271
rect 40379 9083 40385 9259
rect 40419 9204 40425 9259
rect 40544 9259 40590 9271
rect 40544 9204 40550 9259
rect 40419 9116 40550 9204
rect 40419 9083 40425 9116
rect 40379 9071 40425 9083
rect 40544 9083 40550 9116
rect 40584 9083 40590 9259
rect 40544 9071 40590 9083
rect 40662 9259 40708 9271
rect 40662 9083 40668 9259
rect 40702 9083 40708 9259
rect 40662 9071 40708 9083
rect 40780 9259 40826 9271
rect 40780 9083 40786 9259
rect 40820 9083 40826 9259
rect 40780 9071 40826 9083
rect 40898 9259 40944 9271
rect 40898 9083 40904 9259
rect 40938 9083 40944 9259
rect 40898 9071 40944 9083
rect 40031 9032 40065 9071
rect 40267 9032 40301 9071
rect 40031 8997 40301 9032
rect 40668 9033 40701 9071
rect 40904 9033 40937 9071
rect 40668 8997 40937 9033
rect 37440 8929 38260 8977
rect 40065 8996 40301 8997
rect 37440 8898 37906 8929
rect 40065 8922 40197 8996
rect 37440 8642 37545 8898
rect 40055 8814 40065 8922
rect 40197 8814 40207 8922
rect 38277 8734 38356 8746
rect 37440 8536 37503 8642
rect 37615 8536 37625 8642
rect 38277 8638 38283 8734
rect 38207 8618 38283 8638
rect 38350 8638 38356 8734
rect 40092 8676 40098 8814
rect 40165 8676 40171 8814
rect 40092 8664 40171 8676
rect 38350 8618 38427 8638
rect 37440 8525 37589 8536
rect 37440 7348 37545 8525
rect 38207 8510 38251 8618
rect 38383 8510 38427 8618
rect 38207 8468 38427 8510
rect 41005 8483 41067 10054
rect 41257 10046 41303 10058
rect 41257 9670 41263 10046
rect 41297 9670 41303 10046
rect 41257 9658 41303 9670
rect 41375 10046 41421 10058
rect 41375 9670 41381 10046
rect 41415 9670 41421 10046
rect 41375 9658 41421 9670
rect 41493 10046 41539 10058
rect 41493 9670 41499 10046
rect 41533 9670 41539 10046
rect 41493 9658 41539 9670
rect 41611 10046 41657 10058
rect 41611 9670 41617 10046
rect 41651 9670 41657 10046
rect 41611 9658 41657 9670
rect 41729 10046 41775 10058
rect 41729 9670 41735 10046
rect 41769 9670 41775 10046
rect 41729 9658 41775 9670
rect 41847 10046 41893 10058
rect 41847 9670 41853 10046
rect 41887 9670 41893 10046
rect 41847 9658 41893 9670
rect 41965 10046 42011 10058
rect 41965 9670 41971 10046
rect 42005 9670 42011 10046
rect 41965 9658 42011 9670
rect 41263 9616 41297 9658
rect 41499 9616 41533 9658
rect 41263 9588 41533 9616
rect 41617 9617 41651 9658
rect 41853 9617 41887 9658
rect 41617 9588 41887 9617
rect 41263 9540 41297 9588
rect 41263 9510 41326 9540
rect 41291 9418 41326 9510
rect 41798 9480 41898 9501
rect 41798 9426 41812 9480
rect 41877 9426 41898 9480
rect 41798 9421 41898 9426
rect 41971 9475 42005 9658
rect 41971 9421 42080 9475
rect 43697 9436 43878 11606
rect 48350 11699 48396 11711
rect 48350 11323 48356 11699
rect 48390 11323 48396 11699
rect 48350 11311 48396 11323
rect 48468 11699 48514 11711
rect 48468 11323 48474 11699
rect 48508 11323 48514 11699
rect 48468 11311 48514 11323
rect 48586 11699 48632 11711
rect 48586 11323 48592 11699
rect 48626 11350 48632 11699
rect 48703 11699 48749 11711
rect 48703 11523 48709 11699
rect 48743 11523 48749 11699
rect 48703 11516 48749 11523
rect 48821 11699 50528 11711
rect 48821 11523 48827 11699
rect 48861 11686 50528 11699
rect 48861 11523 48867 11686
rect 49111 11606 50528 11686
rect 49115 11605 50528 11606
rect 48703 11511 48752 11516
rect 48821 11511 48867 11523
rect 48709 11350 48752 11511
rect 48626 11323 48752 11350
rect 48586 11311 48752 11323
rect 48592 11307 48752 11311
rect 48257 11279 48330 11280
rect 48257 11274 48465 11279
rect 48257 11228 48269 11274
rect 48318 11273 48465 11274
rect 48318 11239 48415 11273
rect 48449 11239 48465 11273
rect 48318 11228 48465 11239
rect 48257 11223 48465 11228
rect 48517 11273 48583 11279
rect 48517 11239 48533 11273
rect 48567 11239 48583 11273
rect 48257 11222 48330 11223
rect 48517 11194 48583 11239
rect 48120 11186 48583 11194
rect 48120 11154 48584 11186
rect 48676 11170 48752 11307
rect 48120 10735 48166 11154
rect 48672 11110 48682 11170
rect 48744 11110 48754 11170
rect 48106 10681 48116 10735
rect 48173 10681 48183 10735
rect 50347 10697 50528 11605
rect 55004 11344 55010 11720
rect 55044 11344 55050 11720
rect 55004 11332 55050 11344
rect 55122 11720 55168 11732
rect 55122 11344 55128 11720
rect 55162 11344 55168 11720
rect 55122 11332 55168 11344
rect 55240 11720 55286 11732
rect 55240 11344 55246 11720
rect 55280 11371 55286 11720
rect 55357 11720 55403 11732
rect 55357 11544 55363 11720
rect 55397 11544 55403 11720
rect 55357 11537 55403 11544
rect 55475 11720 57154 11732
rect 55475 11544 55481 11720
rect 55515 11707 57154 11720
rect 55515 11544 55521 11707
rect 55765 11626 57154 11707
rect 55357 11532 55406 11537
rect 55475 11532 55521 11544
rect 55363 11371 55406 11532
rect 55280 11344 55406 11371
rect 55240 11332 55406 11344
rect 55246 11328 55406 11332
rect 54864 11300 54949 11302
rect 54864 11296 55119 11300
rect 54864 11248 54876 11296
rect 54937 11294 55119 11296
rect 54937 11260 55069 11294
rect 55103 11260 55119 11294
rect 54937 11248 55119 11260
rect 54864 11244 55119 11248
rect 55171 11294 55237 11300
rect 55171 11260 55187 11294
rect 55221 11260 55237 11294
rect 54864 11242 54949 11244
rect 55171 11214 55237 11260
rect 54965 11207 55237 11214
rect 54965 11206 55238 11207
rect 54965 11168 54978 11206
rect 55023 11175 55238 11206
rect 55330 11191 55406 11328
rect 55023 11168 55037 11175
rect 54965 11159 55037 11168
rect 55326 11131 55336 11191
rect 55398 11131 55408 11191
rect 56973 10765 57154 11626
rect 47297 10524 47376 10536
rect 44814 10473 44893 10485
rect 44814 10376 44820 10473
rect 44742 10356 44820 10376
rect 44887 10376 44893 10473
rect 47297 10410 47303 10524
rect 47370 10410 47376 10524
rect 48441 10526 48520 10538
rect 48441 10410 48447 10526
rect 48514 10410 48520 10526
rect 44887 10356 44962 10376
rect 44742 10248 44786 10356
rect 44918 10248 44962 10356
rect 46539 10314 46595 10322
rect 44742 10206 44962 10248
rect 45613 10306 46595 10314
rect 45613 10272 46555 10306
rect 46589 10272 46595 10306
rect 47258 10302 47268 10410
rect 47400 10347 47410 10410
rect 47400 10336 47412 10347
rect 47400 10302 47413 10336
rect 47669 10326 47725 10328
rect 45613 10256 46595 10272
rect 47268 10264 47413 10302
rect 45613 10255 46592 10256
rect 44346 10176 45323 10206
rect 44346 10070 44378 10176
rect 44582 10070 44614 10176
rect 44818 10070 44850 10176
rect 45054 10070 45086 10176
rect 45289 10070 45323 10176
rect 44339 10058 44385 10070
rect 44339 9882 44345 10058
rect 44379 9882 44385 10058
rect 44339 9870 44385 9882
rect 44457 10058 44503 10070
rect 44457 9882 44463 10058
rect 44497 9882 44503 10058
rect 44457 9870 44503 9882
rect 44575 10058 44621 10070
rect 44575 9882 44581 10058
rect 44615 9882 44621 10058
rect 44575 9870 44621 9882
rect 44693 10058 44739 10070
rect 44693 9882 44699 10058
rect 44733 9882 44739 10058
rect 44693 9870 44739 9882
rect 44811 10058 44857 10070
rect 44811 9882 44817 10058
rect 44851 9882 44857 10058
rect 44811 9870 44857 9882
rect 44929 10058 44975 10070
rect 44929 9882 44935 10058
rect 44969 9882 44975 10058
rect 44929 9870 44975 9882
rect 45047 10058 45093 10070
rect 45047 9882 45053 10058
rect 45087 9882 45093 10058
rect 45047 9870 45093 9882
rect 45165 10058 45211 10070
rect 45165 9882 45171 10058
rect 45205 9882 45211 10058
rect 45165 9870 45211 9882
rect 45283 10058 45329 10070
rect 45283 9882 45289 10058
rect 45323 9882 45329 10058
rect 45283 9870 45329 9882
rect 45401 10058 45447 10070
rect 45401 9882 45407 10058
rect 45441 9882 45447 10058
rect 45401 9870 45447 9882
rect 44462 9776 44498 9870
rect 44698 9776 44734 9870
rect 44934 9777 44970 9870
rect 45096 9822 45162 9829
rect 45096 9788 45112 9822
rect 45146 9788 45162 9822
rect 45096 9777 45162 9788
rect 44934 9776 45162 9777
rect 44462 9747 45162 9776
rect 44462 9746 45044 9747
rect 44582 9633 44616 9746
rect 44978 9705 45044 9746
rect 44978 9671 44994 9705
rect 45028 9671 45044 9705
rect 44978 9664 45044 9671
rect 45406 9665 45441 9870
rect 45613 9665 45680 10255
rect 47372 10232 47413 10264
rect 47659 10260 47669 10326
rect 47725 10260 47735 10326
rect 48405 10302 48415 10410
rect 48547 10347 48557 10410
rect 48547 10336 48559 10347
rect 48547 10302 48560 10336
rect 48415 10264 48560 10302
rect 48519 10236 48560 10264
rect 46788 10204 47058 10232
rect 46529 10138 46539 10204
rect 46605 10138 46615 10204
rect 46788 10142 46822 10204
rect 47024 10142 47058 10204
rect 47142 10204 47413 10232
rect 47930 10208 48200 10236
rect 47142 10142 47176 10204
rect 47378 10142 47413 10204
rect 47554 10192 47725 10208
rect 47554 10158 47685 10192
rect 47719 10158 47725 10192
rect 47554 10142 47725 10158
rect 47930 10146 47964 10208
rect 48166 10146 48200 10208
rect 48284 10208 48560 10236
rect 48284 10146 48318 10208
rect 48520 10146 48560 10208
rect 46664 10130 46710 10142
rect 46664 9754 46670 10130
rect 46704 9754 46710 10130
rect 46664 9742 46710 9754
rect 46782 10130 46828 10142
rect 46782 9754 46788 10130
rect 46822 9754 46828 10130
rect 46782 9742 46828 9754
rect 46900 10130 46946 10142
rect 46900 9754 46906 10130
rect 46940 9754 46946 10130
rect 46900 9742 46946 9754
rect 47018 10130 47064 10142
rect 47018 9754 47024 10130
rect 47058 9754 47064 10130
rect 47018 9742 47064 9754
rect 47136 10130 47182 10142
rect 47136 9754 47142 10130
rect 47176 9754 47182 10130
rect 47136 9742 47182 9754
rect 47254 10130 47300 10142
rect 47254 9754 47260 10130
rect 47294 9754 47300 10130
rect 47254 9742 47300 9754
rect 47372 10130 47418 10142
rect 47372 9754 47378 10130
rect 47412 9754 47418 10130
rect 47372 9742 47418 9754
rect 45406 9637 45680 9665
rect 45052 9633 45680 9637
rect 41291 9382 41518 9418
rect 41291 9275 41326 9382
rect 41452 9348 41518 9382
rect 41452 9314 41468 9348
rect 41502 9314 41518 9348
rect 41799 9406 41896 9421
rect 41799 9339 41856 9406
rect 41452 9308 41518 9314
rect 41693 9303 41962 9339
rect 41693 9275 41726 9303
rect 41929 9275 41962 9303
rect 42046 9275 42080 9421
rect 41167 9263 41213 9275
rect 41167 9087 41173 9263
rect 41207 9087 41213 9263
rect 41167 9075 41213 9087
rect 41285 9263 41331 9275
rect 41285 9087 41291 9263
rect 41325 9087 41331 9263
rect 41285 9075 41331 9087
rect 41403 9263 41449 9275
rect 41403 9087 41409 9263
rect 41443 9087 41449 9263
rect 41403 9075 41449 9087
rect 41521 9263 41567 9275
rect 41521 9087 41527 9263
rect 41561 9208 41567 9263
rect 41686 9263 41732 9275
rect 41686 9208 41692 9263
rect 41561 9120 41692 9208
rect 41561 9087 41567 9120
rect 41521 9075 41567 9087
rect 41686 9087 41692 9120
rect 41726 9087 41732 9263
rect 41686 9075 41732 9087
rect 41804 9263 41850 9275
rect 41804 9087 41810 9263
rect 41844 9087 41850 9263
rect 41804 9075 41850 9087
rect 41922 9263 41968 9275
rect 41922 9087 41928 9263
rect 41962 9087 41968 9263
rect 41922 9075 41968 9087
rect 42040 9263 42086 9275
rect 42040 9087 42046 9263
rect 42080 9087 42086 9263
rect 43698 9228 43878 9436
rect 44576 9621 44622 9633
rect 44576 9245 44582 9621
rect 44616 9245 44622 9621
rect 44576 9233 44622 9245
rect 44694 9621 44740 9633
rect 44694 9245 44700 9621
rect 44734 9245 44740 9621
rect 44694 9233 44740 9245
rect 44812 9621 44858 9633
rect 44812 9245 44818 9621
rect 44852 9269 44858 9621
rect 44929 9621 44975 9633
rect 44929 9445 44935 9621
rect 44969 9445 44975 9621
rect 44929 9433 44975 9445
rect 45047 9621 45680 9633
rect 45047 9445 45053 9621
rect 45087 9608 45680 9621
rect 46670 9700 46704 9742
rect 46906 9700 46940 9742
rect 46670 9672 46940 9700
rect 47024 9701 47058 9742
rect 47260 9701 47294 9742
rect 47024 9672 47294 9701
rect 46670 9624 46704 9672
rect 45087 9445 45093 9608
rect 46670 9594 46733 9624
rect 45047 9433 45093 9445
rect 46698 9502 46733 9594
rect 46698 9466 46925 9502
rect 47195 9491 47205 9588
rect 47304 9491 47314 9588
rect 47378 9559 47412 9742
rect 47378 9505 47487 9559
rect 44935 9317 44970 9433
rect 46698 9359 46733 9466
rect 46859 9432 46925 9466
rect 46859 9398 46875 9432
rect 46909 9398 46925 9432
rect 47206 9490 47303 9491
rect 47206 9423 47263 9490
rect 46859 9392 46925 9398
rect 47100 9387 47369 9423
rect 47100 9359 47133 9387
rect 47336 9359 47369 9387
rect 47453 9359 47487 9505
rect 46574 9347 46620 9359
rect 45066 9317 45174 9327
rect 44935 9269 45066 9317
rect 45174 9278 45319 9284
rect 44852 9245 45066 9269
rect 44812 9233 45066 9245
rect 44818 9229 45066 9233
rect 43698 9201 44454 9228
rect 43698 9195 44691 9201
rect 43698 9161 44641 9195
rect 44675 9161 44691 9195
rect 43698 9145 44691 9161
rect 44743 9195 44809 9201
rect 44743 9161 44759 9195
rect 44793 9161 44809 9195
rect 44992 9185 45066 9229
rect 45307 9211 45319 9278
rect 45174 9205 45319 9211
rect 45066 9175 45174 9185
rect 43698 9129 44454 9145
rect 43698 9128 44391 9129
rect 43698 9124 43926 9128
rect 42040 9075 42086 9087
rect 41173 9036 41207 9075
rect 41409 9036 41443 9075
rect 41173 9000 41443 9036
rect 41810 9037 41843 9075
rect 42046 9037 42079 9075
rect 41810 9001 42079 9037
rect 41173 8999 41339 9000
rect 41207 8920 41339 8999
rect 41197 8812 41207 8920
rect 41339 8812 41349 8920
rect 41230 8678 41236 8812
rect 41303 8678 41309 8812
rect 41230 8666 41309 8678
rect 43197 8713 43710 8745
rect 43197 8607 43558 8713
rect 43670 8700 43710 8713
rect 43670 8607 43712 8700
rect 43197 8596 43712 8607
rect 43197 8595 43710 8596
rect 37811 8438 38788 8468
rect 41005 8466 41068 8483
rect 40930 8462 41068 8466
rect 37811 8332 37843 8438
rect 38047 8332 38079 8438
rect 38283 8332 38315 8438
rect 38519 8332 38551 8438
rect 38754 8332 38788 8438
rect 39098 8428 41068 8462
rect 39096 8399 41068 8428
rect 39096 8383 39142 8399
rect 40930 8397 41068 8399
rect 37804 8320 37850 8332
rect 37804 8144 37810 8320
rect 37844 8144 37850 8320
rect 37804 8132 37850 8144
rect 37922 8320 37968 8332
rect 37922 8144 37928 8320
rect 37962 8144 37968 8320
rect 37922 8132 37968 8144
rect 38040 8320 38086 8332
rect 38040 8144 38046 8320
rect 38080 8144 38086 8320
rect 38040 8132 38086 8144
rect 38158 8320 38204 8332
rect 38158 8144 38164 8320
rect 38198 8144 38204 8320
rect 38158 8132 38204 8144
rect 38276 8320 38322 8332
rect 38276 8144 38282 8320
rect 38316 8144 38322 8320
rect 38276 8132 38322 8144
rect 38394 8320 38440 8332
rect 38394 8144 38400 8320
rect 38434 8144 38440 8320
rect 38394 8132 38440 8144
rect 38512 8320 38558 8332
rect 38512 8144 38518 8320
rect 38552 8144 38558 8320
rect 38512 8132 38558 8144
rect 38630 8320 38676 8332
rect 38630 8144 38636 8320
rect 38670 8144 38676 8320
rect 38630 8132 38676 8144
rect 38748 8320 38794 8332
rect 38748 8144 38754 8320
rect 38788 8144 38794 8320
rect 38748 8132 38794 8144
rect 38866 8320 38912 8332
rect 38866 8144 38872 8320
rect 38906 8144 38912 8320
rect 38866 8132 38912 8144
rect 37927 8038 37963 8132
rect 38163 8038 38199 8132
rect 38399 8039 38435 8132
rect 38561 8084 38627 8091
rect 38561 8050 38577 8084
rect 38611 8050 38627 8084
rect 38561 8039 38627 8050
rect 38399 8038 38627 8039
rect 37927 8009 38627 8038
rect 37927 8008 38509 8009
rect 38047 7895 38081 8008
rect 38443 7967 38509 8008
rect 38443 7933 38459 7967
rect 38493 7933 38509 7967
rect 38443 7926 38509 7933
rect 38871 7914 38906 8132
rect 39095 7931 39142 8383
rect 41989 8392 42068 8404
rect 41989 8275 41995 8392
rect 42062 8275 42068 8392
rect 40054 8167 40064 8275
rect 40196 8167 40206 8275
rect 41952 8167 41962 8275
rect 42094 8167 42104 8275
rect 40064 8127 40196 8167
rect 41962 8127 42094 8167
rect 40063 8061 40196 8127
rect 41961 8061 42094 8127
rect 39392 8018 40865 8061
rect 39095 7915 39141 7931
rect 39060 7914 39141 7915
rect 38871 7899 39141 7914
rect 38517 7895 39141 7899
rect 38041 7883 38087 7895
rect 37776 7405 37786 7523
rect 37904 7491 37914 7523
rect 38041 7507 38047 7883
rect 38081 7507 38087 7883
rect 38041 7495 38087 7507
rect 38159 7883 38205 7895
rect 38159 7507 38165 7883
rect 38199 7507 38205 7883
rect 38159 7495 38205 7507
rect 38277 7883 38323 7895
rect 38277 7507 38283 7883
rect 38317 7531 38323 7883
rect 38394 7883 38440 7895
rect 38394 7707 38400 7883
rect 38434 7707 38440 7883
rect 38394 7695 38440 7707
rect 38512 7883 39141 7895
rect 38512 7707 38518 7883
rect 38552 7871 39141 7883
rect 38552 7870 38794 7871
rect 38552 7707 38558 7870
rect 39060 7869 39141 7871
rect 39392 7715 39426 8018
rect 39758 7915 39792 8018
rect 39994 7915 40028 8018
rect 40230 7915 40264 8018
rect 40466 7915 40500 8018
rect 39752 7903 39798 7915
rect 38512 7695 38558 7707
rect 39268 7703 39314 7715
rect 38400 7579 38435 7695
rect 38531 7579 38639 7589
rect 38400 7531 38531 7579
rect 38639 7546 38788 7552
rect 38317 7507 38531 7531
rect 38277 7495 38531 7507
rect 38283 7491 38531 7495
rect 37904 7463 37919 7491
rect 37904 7457 38156 7463
rect 37904 7423 38106 7457
rect 38140 7423 38156 7457
rect 37904 7407 38156 7423
rect 38208 7457 38274 7463
rect 38208 7423 38224 7457
rect 38258 7423 38274 7457
rect 38457 7447 38531 7491
rect 38776 7479 38788 7546
rect 39268 7527 39274 7703
rect 39308 7527 39314 7703
rect 39268 7515 39314 7527
rect 39386 7703 39432 7715
rect 39386 7527 39392 7703
rect 39426 7527 39432 7703
rect 39386 7515 39432 7527
rect 39504 7703 39550 7715
rect 39504 7527 39510 7703
rect 39544 7527 39550 7703
rect 39504 7515 39550 7527
rect 39622 7703 39668 7715
rect 39752 7703 39758 7903
rect 39622 7527 39628 7703
rect 39662 7527 39758 7703
rect 39792 7527 39798 7903
rect 39622 7515 39668 7527
rect 39752 7515 39798 7527
rect 39870 7903 39916 7915
rect 39870 7527 39876 7903
rect 39910 7527 39916 7903
rect 39870 7515 39916 7527
rect 39988 7903 40034 7915
rect 39988 7527 39994 7903
rect 40028 7527 40034 7903
rect 39988 7515 40034 7527
rect 40106 7903 40152 7915
rect 40106 7527 40112 7903
rect 40146 7527 40152 7903
rect 40106 7515 40152 7527
rect 40224 7903 40270 7915
rect 40224 7527 40230 7903
rect 40264 7527 40270 7903
rect 40224 7515 40270 7527
rect 40342 7903 40388 7915
rect 40342 7527 40348 7903
rect 40382 7527 40388 7903
rect 40342 7515 40388 7527
rect 40460 7903 40506 7915
rect 40460 7527 40466 7903
rect 40500 7703 40506 7903
rect 40831 7715 40865 8018
rect 41290 8018 42763 8061
rect 41290 7715 41324 8018
rect 41656 7915 41690 8018
rect 41892 7915 41926 8018
rect 42128 7915 42162 8018
rect 42364 7915 42398 8018
rect 41650 7903 41696 7915
rect 40589 7703 40635 7715
rect 40500 7527 40595 7703
rect 40629 7527 40635 7703
rect 40460 7515 40506 7527
rect 40589 7515 40635 7527
rect 40707 7703 40753 7715
rect 40707 7527 40713 7703
rect 40747 7527 40753 7703
rect 40707 7515 40753 7527
rect 40825 7703 40871 7715
rect 40825 7527 40831 7703
rect 40865 7527 40871 7703
rect 40825 7515 40871 7527
rect 40943 7703 40989 7715
rect 40943 7527 40949 7703
rect 40983 7527 40989 7703
rect 40943 7515 40989 7527
rect 41166 7703 41212 7715
rect 41166 7527 41172 7703
rect 41206 7527 41212 7703
rect 41166 7515 41212 7527
rect 41284 7703 41330 7715
rect 41284 7527 41290 7703
rect 41324 7527 41330 7703
rect 41284 7515 41330 7527
rect 41402 7703 41448 7715
rect 41402 7527 41408 7703
rect 41442 7527 41448 7703
rect 41402 7515 41448 7527
rect 41520 7703 41566 7715
rect 41650 7703 41656 7903
rect 41520 7527 41526 7703
rect 41560 7527 41656 7703
rect 41690 7527 41696 7903
rect 41520 7515 41566 7527
rect 41650 7515 41696 7527
rect 41768 7903 41814 7915
rect 41768 7527 41774 7903
rect 41808 7527 41814 7903
rect 41768 7515 41814 7527
rect 41886 7903 41932 7915
rect 41886 7527 41892 7903
rect 41926 7527 41932 7903
rect 41886 7515 41932 7527
rect 42004 7903 42050 7915
rect 42004 7527 42010 7903
rect 42044 7527 42050 7903
rect 42004 7515 42050 7527
rect 42122 7903 42168 7915
rect 42122 7527 42128 7903
rect 42162 7527 42168 7903
rect 42122 7515 42168 7527
rect 42240 7903 42286 7915
rect 42240 7527 42246 7903
rect 42280 7527 42286 7903
rect 42240 7515 42286 7527
rect 42358 7903 42404 7915
rect 42358 7527 42364 7903
rect 42398 7703 42404 7903
rect 42729 7715 42763 8018
rect 42487 7703 42533 7715
rect 42398 7527 42493 7703
rect 42527 7527 42533 7703
rect 42358 7515 42404 7527
rect 42487 7515 42533 7527
rect 42605 7703 42651 7715
rect 42605 7527 42611 7703
rect 42645 7527 42651 7703
rect 42605 7515 42651 7527
rect 42723 7703 42769 7715
rect 42723 7527 42729 7703
rect 42763 7527 42769 7703
rect 42723 7515 42769 7527
rect 42841 7703 42887 7715
rect 42841 7527 42847 7703
rect 42881 7527 42887 7703
rect 42841 7515 42887 7527
rect 38639 7473 38788 7479
rect 39274 7481 39308 7515
rect 39876 7481 39910 7515
rect 40112 7481 40146 7515
rect 38531 7437 38639 7447
rect 39274 7446 39433 7481
rect 39876 7446 40146 7481
rect 40713 7481 40747 7515
rect 40949 7481 40983 7515
rect 40713 7446 40983 7481
rect 41172 7481 41206 7515
rect 41774 7481 41808 7515
rect 42010 7481 42044 7515
rect 41172 7446 41331 7481
rect 41774 7446 42044 7481
rect 42611 7481 42645 7515
rect 42847 7481 42881 7515
rect 42611 7446 42881 7481
rect 37904 7405 37919 7407
rect 37819 7391 37919 7405
rect 37819 7348 37919 7349
rect 37440 7327 37919 7348
rect 38208 7327 38274 7423
rect 37440 7279 38274 7327
rect 37440 7250 37919 7279
rect 37440 7248 37545 7250
rect 37819 7249 37919 7250
rect 37273 7063 37283 7142
rect 37376 7063 37386 7142
rect 38275 7128 38354 7140
rect 35482 7027 35531 7032
rect 35600 7027 35646 7039
rect 35488 6866 35531 7027
rect 35405 6839 35531 6866
rect 35365 6827 35531 6839
rect 35371 6823 35531 6827
rect 34535 6789 35244 6795
rect 34535 6755 35194 6789
rect 35228 6755 35244 6789
rect 34535 6739 35244 6755
rect 35296 6789 35362 6795
rect 35296 6755 35312 6789
rect 35346 6755 35362 6789
rect 33763 6701 34030 6706
rect 33763 6688 33932 6701
rect 33763 6607 33778 6688
rect 33872 6607 33932 6688
rect 33763 6597 33932 6607
rect 34019 6597 34030 6701
rect 33763 6591 34030 6597
rect 33092 4907 33102 4974
rect 33169 4907 33179 4974
rect 30501 -1213 33035 -1147
rect 33097 2900 33172 4907
rect 33097 2846 33108 2900
rect 33164 2846 33174 2900
rect 33097 832 33172 2846
rect 34535 1049 34640 6739
rect 35296 6710 35362 6755
rect 34698 6702 35362 6710
rect 34698 6696 35363 6702
rect 34698 6600 34729 6696
rect 34806 6670 35363 6696
rect 35455 6686 35531 6823
rect 34806 6600 34816 6670
rect 35451 6626 35461 6686
rect 35523 6626 35533 6686
rect 34698 3809 34816 6600
rect 37284 5889 37377 7063
rect 38275 7034 38281 7128
rect 38202 7014 38281 7034
rect 38348 7034 38354 7128
rect 38348 7014 38422 7034
rect 38202 6906 38246 7014
rect 38378 6906 38422 7014
rect 38202 6864 38422 6906
rect 37806 6834 38783 6864
rect 37806 6728 37838 6834
rect 38042 6728 38074 6834
rect 38278 6728 38310 6834
rect 38514 6728 38546 6834
rect 38749 6728 38783 6834
rect 37799 6716 37845 6728
rect 37799 6540 37805 6716
rect 37839 6540 37845 6716
rect 37799 6528 37845 6540
rect 37917 6716 37963 6728
rect 37917 6540 37923 6716
rect 37957 6540 37963 6716
rect 37917 6528 37963 6540
rect 38035 6716 38081 6728
rect 38035 6540 38041 6716
rect 38075 6540 38081 6716
rect 38035 6528 38081 6540
rect 38153 6716 38199 6728
rect 38153 6540 38159 6716
rect 38193 6540 38199 6716
rect 38153 6528 38199 6540
rect 38271 6716 38317 6728
rect 38271 6540 38277 6716
rect 38311 6540 38317 6716
rect 38271 6528 38317 6540
rect 38389 6716 38435 6728
rect 38389 6540 38395 6716
rect 38429 6540 38435 6716
rect 38389 6528 38435 6540
rect 38507 6716 38553 6728
rect 38507 6540 38513 6716
rect 38547 6540 38553 6716
rect 38507 6528 38553 6540
rect 38625 6716 38671 6728
rect 38625 6540 38631 6716
rect 38665 6540 38671 6716
rect 38625 6528 38671 6540
rect 38743 6716 38789 6728
rect 38743 6540 38749 6716
rect 38783 6540 38789 6716
rect 38743 6528 38789 6540
rect 38861 6716 38907 6728
rect 38861 6540 38867 6716
rect 38901 6540 38907 6716
rect 38861 6528 38907 6540
rect 39399 6662 39433 7446
rect 40112 7384 40146 7446
rect 39701 7346 40443 7384
rect 39701 7222 39735 7346
rect 39937 7222 39971 7346
rect 40173 7222 40207 7346
rect 40409 7222 40443 7346
rect 40699 7239 40709 7305
rect 40772 7239 40782 7305
rect 39695 7210 39741 7222
rect 39695 6834 39701 7210
rect 39735 6834 39741 7210
rect 39695 6822 39741 6834
rect 39813 7210 39859 7222
rect 39813 6834 39819 7210
rect 39853 6834 39859 7210
rect 39813 6822 39859 6834
rect 39931 7210 39977 7222
rect 39931 6834 39937 7210
rect 39971 6834 39977 7210
rect 39931 6822 39977 6834
rect 40049 7210 40095 7222
rect 40049 6834 40055 7210
rect 40089 6834 40095 7210
rect 40049 6822 40095 6834
rect 40167 7210 40213 7222
rect 40167 6834 40173 7210
rect 40207 6834 40213 7210
rect 40167 6822 40213 6834
rect 40285 7210 40331 7222
rect 40285 6834 40291 7210
rect 40325 6834 40331 7210
rect 40285 6822 40331 6834
rect 40403 7210 40449 7222
rect 40403 6834 40409 7210
rect 40443 6834 40449 7210
rect 40403 6822 40449 6834
rect 40815 6663 40849 7446
rect 40542 6662 40849 6663
rect 39399 6657 39715 6662
rect 40429 6657 40849 6662
rect 39399 6646 39782 6657
rect 39399 6619 39731 6646
rect 37922 6434 37958 6528
rect 38158 6434 38194 6528
rect 38394 6435 38430 6528
rect 38556 6480 38622 6487
rect 38556 6446 38572 6480
rect 38606 6446 38622 6480
rect 38556 6435 38622 6446
rect 38394 6434 38622 6435
rect 37922 6405 38622 6434
rect 37922 6404 38504 6405
rect 38042 6291 38076 6404
rect 38438 6363 38504 6404
rect 38438 6329 38454 6363
rect 38488 6329 38504 6363
rect 38438 6322 38504 6329
rect 38866 6295 38901 6528
rect 39399 6490 39433 6619
rect 39715 6612 39731 6619
rect 39765 6612 39782 6646
rect 39715 6606 39782 6612
rect 40362 6646 40849 6657
rect 40362 6612 40379 6646
rect 40413 6619 40849 6646
rect 40413 6612 40429 6619
rect 40542 6618 40849 6619
rect 40362 6606 40429 6612
rect 39540 6579 39596 6591
rect 39540 6545 39546 6579
rect 39580 6578 39596 6579
rect 40653 6578 40709 6590
rect 39580 6562 40047 6578
rect 39580 6545 39997 6562
rect 39540 6529 39997 6545
rect 39981 6528 39997 6529
rect 40031 6528 40047 6562
rect 39981 6521 40047 6528
rect 40099 6563 40669 6578
rect 40099 6529 40115 6563
rect 40149 6544 40669 6563
rect 40703 6544 40709 6578
rect 40149 6529 40709 6544
rect 40099 6519 40166 6529
rect 40653 6528 40709 6529
rect 40815 6490 40849 6618
rect 41297 6662 41331 7446
rect 42010 7384 42044 7446
rect 41599 7346 42341 7384
rect 41599 7222 41633 7346
rect 41835 7222 41869 7346
rect 42071 7222 42105 7346
rect 42307 7222 42341 7346
rect 41593 7210 41639 7222
rect 41593 6834 41599 7210
rect 41633 6834 41639 7210
rect 41593 6822 41639 6834
rect 41711 7210 41757 7222
rect 41711 6834 41717 7210
rect 41751 6834 41757 7210
rect 41711 6822 41757 6834
rect 41829 7210 41875 7222
rect 41829 6834 41835 7210
rect 41869 6834 41875 7210
rect 41829 6822 41875 6834
rect 41947 7210 41993 7222
rect 41947 6834 41953 7210
rect 41987 6834 41993 7210
rect 41947 6822 41993 6834
rect 42065 7210 42111 7222
rect 42065 6834 42071 7210
rect 42105 6834 42111 7210
rect 42065 6822 42111 6834
rect 42183 7210 42229 7222
rect 42183 6834 42189 7210
rect 42223 6834 42229 7210
rect 42183 6822 42229 6834
rect 42301 7210 42347 7222
rect 42301 6834 42307 7210
rect 42341 6834 42347 7210
rect 42301 6822 42347 6834
rect 42713 6663 42747 7446
rect 42325 6662 42394 6663
rect 42440 6662 42747 6663
rect 41297 6657 41613 6662
rect 42325 6658 42747 6662
rect 41297 6646 41680 6657
rect 41297 6619 41629 6646
rect 41297 6490 41331 6619
rect 41613 6612 41629 6619
rect 41663 6612 41680 6646
rect 41613 6606 41680 6612
rect 42258 6647 42747 6658
rect 42258 6613 42275 6647
rect 42309 6619 42747 6647
rect 42309 6613 42325 6619
rect 42440 6618 42747 6619
rect 42258 6607 42325 6613
rect 41438 6579 41494 6591
rect 41438 6545 41444 6579
rect 41478 6578 41494 6579
rect 42551 6578 42607 6590
rect 41478 6562 41945 6578
rect 41478 6545 41895 6562
rect 41438 6529 41895 6545
rect 41879 6528 41895 6529
rect 41929 6528 41945 6562
rect 41879 6521 41945 6528
rect 41997 6563 42567 6578
rect 41997 6529 42013 6563
rect 42047 6544 42567 6563
rect 42601 6544 42607 6578
rect 42047 6529 42607 6544
rect 41997 6519 42064 6529
rect 42551 6528 42607 6529
rect 42713 6490 42747 6618
rect 42828 7268 42895 7292
rect 42828 7234 42845 7268
rect 42879 7234 42895 7268
rect 38512 6291 38901 6295
rect 38036 6279 38082 6291
rect 38036 5903 38042 6279
rect 38076 5903 38082 6279
rect 38036 5891 38082 5903
rect 38154 6279 38200 6291
rect 38154 5903 38160 6279
rect 38194 5903 38200 6279
rect 38154 5891 38200 5903
rect 38272 6279 38318 6291
rect 38272 5903 38278 6279
rect 38312 5927 38318 6279
rect 38389 6279 38435 6291
rect 38389 6103 38395 6279
rect 38429 6103 38435 6279
rect 38389 6091 38435 6103
rect 38507 6279 38901 6291
rect 39393 6478 39439 6490
rect 39393 6302 39399 6478
rect 39433 6302 39439 6478
rect 39393 6290 39439 6302
rect 39511 6478 39557 6490
rect 39511 6302 39517 6478
rect 39551 6302 39557 6478
rect 39511 6290 39557 6302
rect 39813 6478 39859 6490
rect 38507 6103 38513 6279
rect 38547 6266 38901 6279
rect 38547 6103 38553 6266
rect 38823 6263 38901 6266
rect 38823 6211 38833 6263
rect 38896 6211 38906 6263
rect 38828 6205 38901 6211
rect 38507 6091 38553 6103
rect 38395 5975 38430 6091
rect 39516 5996 39550 6290
rect 39813 6102 39819 6478
rect 39853 6102 39859 6478
rect 39813 6090 39859 6102
rect 39931 6478 39977 6490
rect 39931 6102 39937 6478
rect 39971 6102 39977 6478
rect 39931 6090 39977 6102
rect 40049 6478 40095 6490
rect 40049 6102 40055 6478
rect 40089 6102 40095 6478
rect 40049 6090 40095 6102
rect 40167 6478 40213 6490
rect 40167 6102 40173 6478
rect 40207 6102 40213 6478
rect 40167 6090 40213 6102
rect 40285 6478 40331 6490
rect 40285 6102 40291 6478
rect 40325 6102 40331 6478
rect 40691 6478 40737 6490
rect 40691 6302 40697 6478
rect 40731 6302 40737 6478
rect 40691 6290 40737 6302
rect 40809 6478 40855 6490
rect 40809 6302 40815 6478
rect 40849 6302 40855 6478
rect 40809 6290 40855 6302
rect 41291 6478 41337 6490
rect 41291 6302 41297 6478
rect 41331 6302 41337 6478
rect 41291 6290 41337 6302
rect 41409 6478 41455 6490
rect 41409 6302 41415 6478
rect 41449 6302 41455 6478
rect 41409 6290 41455 6302
rect 41711 6478 41757 6490
rect 40285 6090 40331 6102
rect 40173 5996 40207 6090
rect 40697 5996 40730 6290
rect 38526 5975 38634 5985
rect 38395 5927 38526 5975
rect 39516 5964 40730 5996
rect 41414 5996 41448 6290
rect 41711 6102 41717 6478
rect 41751 6102 41757 6478
rect 41711 6090 41757 6102
rect 41829 6478 41875 6490
rect 41829 6102 41835 6478
rect 41869 6102 41875 6478
rect 41829 6090 41875 6102
rect 41947 6478 41993 6490
rect 41947 6102 41953 6478
rect 41987 6102 41993 6478
rect 41947 6090 41993 6102
rect 42065 6478 42111 6490
rect 42065 6102 42071 6478
rect 42105 6102 42111 6478
rect 42065 6090 42111 6102
rect 42183 6478 42229 6490
rect 42183 6102 42189 6478
rect 42223 6102 42229 6478
rect 42589 6478 42635 6490
rect 42589 6302 42595 6478
rect 42629 6302 42635 6478
rect 42589 6290 42635 6302
rect 42707 6478 42753 6490
rect 42707 6302 42713 6478
rect 42747 6302 42753 6478
rect 42707 6290 42753 6302
rect 42183 6090 42229 6102
rect 42071 5996 42105 6090
rect 42595 5996 42628 6290
rect 41414 5964 42628 5996
rect 38634 5938 38786 5944
rect 38312 5903 38526 5927
rect 38272 5891 38526 5903
rect 37284 5887 37869 5889
rect 38278 5887 38526 5891
rect 37284 5859 37914 5887
rect 37284 5853 38151 5859
rect 37284 5819 38101 5853
rect 38135 5819 38151 5853
rect 37284 5803 38151 5819
rect 38203 5853 38269 5859
rect 38203 5819 38219 5853
rect 38253 5819 38269 5853
rect 38452 5843 38526 5887
rect 38774 5871 38786 5938
rect 40009 5879 40141 5964
rect 41907 5879 42039 5964
rect 38634 5865 38786 5871
rect 38526 5833 38634 5843
rect 37284 5787 37914 5803
rect 37284 5783 37869 5787
rect 37284 5782 37385 5783
rect 37814 5734 37914 5745
rect 37778 5628 37788 5734
rect 37900 5723 37914 5734
rect 38203 5723 38269 5819
rect 39999 5771 40009 5879
rect 40141 5771 40151 5879
rect 41897 5771 41907 5879
rect 42039 5771 42049 5879
rect 42828 5851 42895 7234
rect 37900 5675 38269 5723
rect 37900 5645 37914 5675
rect 37900 5628 37910 5645
rect 38202 5572 38268 5675
rect 40032 5636 40038 5771
rect 40105 5636 40111 5771
rect 40032 5624 40111 5636
rect 42828 5572 42894 5851
rect 38200 5492 42894 5572
rect 40733 4660 40812 4672
rect 35184 4612 35320 4632
rect 35184 4550 35220 4612
rect 35280 4550 35320 4612
rect 35184 4522 35320 4550
rect 38253 4605 38332 4617
rect 34880 4492 35857 4522
rect 38253 4508 38259 4605
rect 34880 4386 34912 4492
rect 35116 4386 35148 4492
rect 35352 4386 35384 4492
rect 35588 4386 35620 4492
rect 35823 4386 35857 4492
rect 38185 4488 38259 4508
rect 38326 4508 38332 4605
rect 40733 4542 40739 4660
rect 40806 4542 40812 4660
rect 41889 4657 41968 4669
rect 41889 4542 41895 4657
rect 41962 4542 41968 4657
rect 38326 4488 38405 4508
rect 34873 4374 34919 4386
rect 34873 4198 34879 4374
rect 34913 4198 34919 4374
rect 34873 4186 34919 4198
rect 34991 4374 35037 4386
rect 34991 4198 34997 4374
rect 35031 4198 35037 4374
rect 34991 4186 35037 4198
rect 35109 4374 35155 4386
rect 35109 4198 35115 4374
rect 35149 4198 35155 4374
rect 35109 4186 35155 4198
rect 35227 4374 35273 4386
rect 35227 4198 35233 4374
rect 35267 4198 35273 4374
rect 35227 4186 35273 4198
rect 35345 4374 35391 4386
rect 35345 4198 35351 4374
rect 35385 4198 35391 4374
rect 35345 4186 35391 4198
rect 35463 4374 35509 4386
rect 35463 4198 35469 4374
rect 35503 4198 35509 4374
rect 35463 4186 35509 4198
rect 35581 4374 35627 4386
rect 35581 4198 35587 4374
rect 35621 4198 35627 4374
rect 35581 4186 35627 4198
rect 35699 4374 35745 4386
rect 35699 4198 35705 4374
rect 35739 4198 35745 4374
rect 35699 4186 35745 4198
rect 35817 4374 35863 4386
rect 35817 4198 35823 4374
rect 35857 4198 35863 4374
rect 35817 4186 35863 4198
rect 35935 4374 35981 4386
rect 35935 4198 35941 4374
rect 35975 4198 35981 4374
rect 38185 4380 38229 4488
rect 38361 4380 38405 4488
rect 39982 4446 40038 4454
rect 38185 4338 38405 4380
rect 39056 4438 40038 4446
rect 39056 4404 39998 4438
rect 40032 4404 40038 4438
rect 40701 4434 40711 4542
rect 40843 4479 40853 4542
rect 40843 4468 40855 4479
rect 40843 4434 40856 4468
rect 41112 4458 41168 4460
rect 39056 4388 40038 4404
rect 40711 4396 40856 4434
rect 39056 4387 40035 4388
rect 37789 4308 38766 4338
rect 37789 4202 37821 4308
rect 38025 4202 38057 4308
rect 38261 4202 38293 4308
rect 38497 4202 38529 4308
rect 38732 4202 38766 4308
rect 35935 4186 35981 4198
rect 37782 4190 37828 4202
rect 34996 4092 35032 4186
rect 35232 4092 35268 4186
rect 35468 4093 35504 4186
rect 35630 4138 35696 4145
rect 35630 4104 35646 4138
rect 35680 4104 35696 4138
rect 35630 4093 35696 4104
rect 35468 4092 35696 4093
rect 34996 4063 35696 4092
rect 34996 4062 35578 4063
rect 35116 3949 35150 4062
rect 35512 4021 35578 4062
rect 35512 3987 35528 4021
rect 35562 3987 35578 4021
rect 35512 3980 35578 3987
rect 35940 3953 35975 4186
rect 37782 4014 37788 4190
rect 37822 4014 37828 4190
rect 37782 4002 37828 4014
rect 37900 4190 37946 4202
rect 37900 4014 37906 4190
rect 37940 4014 37946 4190
rect 37900 4002 37946 4014
rect 38018 4190 38064 4202
rect 38018 4014 38024 4190
rect 38058 4014 38064 4190
rect 38018 4002 38064 4014
rect 38136 4190 38182 4202
rect 38136 4014 38142 4190
rect 38176 4014 38182 4190
rect 38136 4002 38182 4014
rect 38254 4190 38300 4202
rect 38254 4014 38260 4190
rect 38294 4014 38300 4190
rect 38254 4002 38300 4014
rect 38372 4190 38418 4202
rect 38372 4014 38378 4190
rect 38412 4014 38418 4190
rect 38372 4002 38418 4014
rect 38490 4190 38536 4202
rect 38490 4014 38496 4190
rect 38530 4014 38536 4190
rect 38490 4002 38536 4014
rect 38608 4190 38654 4202
rect 38608 4014 38614 4190
rect 38648 4014 38654 4190
rect 38608 4002 38654 4014
rect 38726 4190 38772 4202
rect 38726 4014 38732 4190
rect 38766 4014 38772 4190
rect 38726 4002 38772 4014
rect 38844 4190 38890 4202
rect 38844 4014 38850 4190
rect 38884 4014 38890 4190
rect 38844 4002 38890 4014
rect 35586 3949 35975 3953
rect 35110 3937 35156 3949
rect 34698 3709 35070 3809
rect 34994 3517 35048 3709
rect 35110 3561 35116 3937
rect 35150 3561 35156 3937
rect 35110 3549 35156 3561
rect 35228 3937 35274 3949
rect 35228 3561 35234 3937
rect 35268 3561 35274 3937
rect 35228 3549 35274 3561
rect 35346 3937 35392 3949
rect 35346 3561 35352 3937
rect 35386 3588 35392 3937
rect 35463 3937 35509 3949
rect 35463 3761 35469 3937
rect 35503 3761 35509 3937
rect 35463 3754 35509 3761
rect 35581 3937 35975 3949
rect 35581 3761 35587 3937
rect 35621 3928 35975 3937
rect 35621 3924 35977 3928
rect 35621 3761 35627 3924
rect 35463 3749 35512 3754
rect 35581 3749 35627 3761
rect 35469 3588 35512 3749
rect 35386 3561 35512 3588
rect 35346 3549 35512 3561
rect 35352 3545 35512 3549
rect 34994 3511 35225 3517
rect 34994 3477 35175 3511
rect 35209 3477 35225 3511
rect 34994 3461 35225 3477
rect 35277 3511 35343 3517
rect 35277 3477 35293 3511
rect 35327 3477 35343 3511
rect 34829 3440 34913 3446
rect 34829 3387 34841 3440
rect 34901 3432 34913 3440
rect 35277 3432 35343 3477
rect 34901 3424 35343 3432
rect 34901 3392 35344 3424
rect 35436 3408 35512 3545
rect 35870 3448 35977 3924
rect 37905 3908 37941 4002
rect 38141 3908 38177 4002
rect 38377 3909 38413 4002
rect 38539 3954 38605 3961
rect 38539 3920 38555 3954
rect 38589 3920 38605 3954
rect 38539 3909 38605 3920
rect 38377 3908 38605 3909
rect 37905 3879 38605 3908
rect 37905 3878 38487 3879
rect 38025 3765 38059 3878
rect 38421 3837 38487 3878
rect 38421 3803 38437 3837
rect 38471 3803 38487 3837
rect 38421 3796 38487 3803
rect 38849 3797 38884 4002
rect 39056 3797 39123 4387
rect 40815 4364 40856 4396
rect 41102 4392 41112 4458
rect 41168 4392 41178 4458
rect 41848 4434 41858 4542
rect 41990 4479 42000 4542
rect 41990 4468 42002 4479
rect 41990 4434 42003 4468
rect 41858 4396 42003 4434
rect 41962 4368 42003 4396
rect 40231 4336 40501 4364
rect 39972 4270 39982 4336
rect 40048 4270 40058 4336
rect 40231 4274 40265 4336
rect 40467 4274 40501 4336
rect 40585 4336 40856 4364
rect 41373 4340 41643 4368
rect 40585 4274 40619 4336
rect 40821 4274 40856 4336
rect 40997 4324 41168 4340
rect 40997 4290 41128 4324
rect 41162 4290 41168 4324
rect 40997 4274 41168 4290
rect 41373 4278 41407 4340
rect 41609 4278 41643 4340
rect 41727 4340 42003 4368
rect 41727 4278 41761 4340
rect 41963 4278 42003 4340
rect 40107 4262 40153 4274
rect 40107 3886 40113 4262
rect 40147 3886 40153 4262
rect 40107 3874 40153 3886
rect 40225 4262 40271 4274
rect 40225 3886 40231 4262
rect 40265 3886 40271 4262
rect 40225 3874 40271 3886
rect 40343 4262 40389 4274
rect 40343 3886 40349 4262
rect 40383 3886 40389 4262
rect 40343 3874 40389 3886
rect 40461 4262 40507 4274
rect 40461 3886 40467 4262
rect 40501 3886 40507 4262
rect 40461 3874 40507 3886
rect 40579 4262 40625 4274
rect 40579 3886 40585 4262
rect 40619 3886 40625 4262
rect 40579 3874 40625 3886
rect 40697 4262 40743 4274
rect 40697 3886 40703 4262
rect 40737 3886 40743 4262
rect 40697 3874 40743 3886
rect 40815 4262 40861 4274
rect 40815 3886 40821 4262
rect 40855 3886 40861 4262
rect 40815 3874 40861 3886
rect 38849 3769 39123 3797
rect 38495 3765 39123 3769
rect 34901 3387 34913 3392
rect 34829 3381 34913 3387
rect 35432 3348 35442 3408
rect 35504 3348 35514 3408
rect 35869 3360 35977 3448
rect 38019 3753 38065 3765
rect 38019 3377 38025 3753
rect 38059 3377 38065 3753
rect 38019 3365 38065 3377
rect 38137 3753 38183 3765
rect 38137 3377 38143 3753
rect 38177 3377 38183 3753
rect 38137 3365 38183 3377
rect 38255 3753 38301 3765
rect 38255 3377 38261 3753
rect 38295 3401 38301 3753
rect 38372 3753 38418 3765
rect 38372 3577 38378 3753
rect 38412 3577 38418 3753
rect 38372 3565 38418 3577
rect 38490 3753 39123 3765
rect 38490 3577 38496 3753
rect 38530 3740 39123 3753
rect 40113 3832 40147 3874
rect 40349 3832 40383 3874
rect 40113 3804 40383 3832
rect 40467 3833 40501 3874
rect 40703 3833 40737 3874
rect 40467 3804 40737 3833
rect 40113 3756 40147 3804
rect 38530 3577 38536 3740
rect 40113 3726 40176 3756
rect 38490 3565 38536 3577
rect 40141 3634 40176 3726
rect 40141 3598 40368 3634
rect 40638 3623 40648 3720
rect 40747 3623 40757 3720
rect 40821 3691 40855 3874
rect 40821 3637 40930 3691
rect 38378 3449 38413 3565
rect 40141 3491 40176 3598
rect 40302 3564 40368 3598
rect 40302 3530 40318 3564
rect 40352 3530 40368 3564
rect 40649 3622 40746 3623
rect 40649 3555 40706 3622
rect 40302 3524 40368 3530
rect 40543 3519 40812 3555
rect 40543 3491 40576 3519
rect 40779 3491 40812 3519
rect 40896 3491 40930 3637
rect 40017 3479 40063 3491
rect 38509 3449 38617 3459
rect 38378 3401 38509 3449
rect 38617 3409 38763 3415
rect 38295 3377 38509 3401
rect 38255 3365 38509 3377
rect 38261 3361 38509 3365
rect 35869 3333 37897 3360
rect 35869 3327 38134 3333
rect 35869 3293 38084 3327
rect 38118 3293 38134 3327
rect 35869 3277 38134 3293
rect 38186 3327 38252 3333
rect 38186 3293 38202 3327
rect 38236 3293 38252 3327
rect 38435 3317 38509 3361
rect 38751 3342 38763 3409
rect 38617 3336 38763 3342
rect 38509 3307 38617 3317
rect 35869 3261 37897 3277
rect 35869 3260 37834 3261
rect 35869 3259 37369 3260
rect 36864 2872 37153 2873
rect 36368 2871 37153 2872
rect 36185 2845 37153 2871
rect 36185 2739 37001 2845
rect 37113 2832 37153 2845
rect 37113 2739 37155 2832
rect 36185 2728 37155 2739
rect 36185 2727 37153 2728
rect 35200 1852 35336 1872
rect 35200 1790 35236 1852
rect 35296 1790 35336 1852
rect 35200 1762 35336 1790
rect 34896 1732 35873 1762
rect 34896 1626 34928 1732
rect 35132 1626 35164 1732
rect 35368 1626 35400 1732
rect 35604 1626 35636 1732
rect 35839 1626 35873 1732
rect 34889 1614 34935 1626
rect 34889 1438 34895 1614
rect 34929 1438 34935 1614
rect 34889 1426 34935 1438
rect 35007 1614 35053 1626
rect 35007 1438 35013 1614
rect 35047 1438 35053 1614
rect 35007 1426 35053 1438
rect 35125 1614 35171 1626
rect 35125 1438 35131 1614
rect 35165 1438 35171 1614
rect 35125 1426 35171 1438
rect 35243 1614 35289 1626
rect 35243 1438 35249 1614
rect 35283 1438 35289 1614
rect 35243 1426 35289 1438
rect 35361 1614 35407 1626
rect 35361 1438 35367 1614
rect 35401 1438 35407 1614
rect 35361 1426 35407 1438
rect 35479 1614 35525 1626
rect 35479 1438 35485 1614
rect 35519 1438 35525 1614
rect 35479 1426 35525 1438
rect 35597 1614 35643 1626
rect 35597 1438 35603 1614
rect 35637 1438 35643 1614
rect 35597 1426 35643 1438
rect 35715 1614 35761 1626
rect 35715 1438 35721 1614
rect 35755 1438 35761 1614
rect 35715 1426 35761 1438
rect 35833 1614 35879 1626
rect 35833 1438 35839 1614
rect 35873 1438 35879 1614
rect 35833 1426 35879 1438
rect 35951 1614 35997 1626
rect 35951 1438 35957 1614
rect 35991 1438 35997 1614
rect 35951 1426 35997 1438
rect 35012 1332 35048 1426
rect 35248 1332 35284 1426
rect 35484 1333 35520 1426
rect 35646 1378 35712 1385
rect 35646 1344 35662 1378
rect 35696 1344 35712 1378
rect 35646 1333 35712 1344
rect 35484 1332 35712 1333
rect 35012 1303 35712 1332
rect 35012 1302 35594 1303
rect 35132 1189 35166 1302
rect 35528 1261 35594 1302
rect 35528 1227 35544 1261
rect 35578 1227 35594 1261
rect 35528 1220 35594 1227
rect 35956 1193 35991 1426
rect 36185 1193 36308 2727
rect 37276 1362 37369 3259
rect 37432 3197 37898 3219
rect 38186 3197 38252 3293
rect 40017 3303 40023 3479
rect 40057 3303 40063 3479
rect 40017 3291 40063 3303
rect 40135 3479 40181 3491
rect 40135 3303 40141 3479
rect 40175 3303 40181 3479
rect 40135 3291 40181 3303
rect 40253 3479 40299 3491
rect 40253 3303 40259 3479
rect 40293 3303 40299 3479
rect 40253 3291 40299 3303
rect 40371 3479 40417 3491
rect 40371 3303 40377 3479
rect 40411 3424 40417 3479
rect 40536 3479 40582 3491
rect 40536 3424 40542 3479
rect 40411 3336 40542 3424
rect 40411 3303 40417 3336
rect 40371 3291 40417 3303
rect 40536 3303 40542 3336
rect 40576 3303 40582 3479
rect 40536 3291 40582 3303
rect 40654 3479 40700 3491
rect 40654 3303 40660 3479
rect 40694 3303 40700 3479
rect 40654 3291 40700 3303
rect 40772 3479 40818 3491
rect 40772 3303 40778 3479
rect 40812 3303 40818 3479
rect 40772 3291 40818 3303
rect 40890 3479 40936 3491
rect 40890 3303 40896 3479
rect 40930 3303 40936 3479
rect 40890 3291 40936 3303
rect 40023 3252 40057 3291
rect 40259 3252 40293 3291
rect 40023 3217 40293 3252
rect 40660 3253 40693 3291
rect 40896 3253 40929 3291
rect 40660 3217 40929 3253
rect 37432 3149 38252 3197
rect 40057 3216 40293 3217
rect 37432 3118 37898 3149
rect 40057 3142 40189 3216
rect 37432 2862 37537 3118
rect 40047 3034 40057 3142
rect 40189 3034 40199 3142
rect 38274 2952 38353 2964
rect 37432 2756 37495 2862
rect 37607 2756 37617 2862
rect 38274 2858 38280 2952
rect 38199 2838 38280 2858
rect 38347 2858 38353 2952
rect 40073 2899 40079 3034
rect 40146 2899 40152 3034
rect 40073 2887 40152 2899
rect 38347 2838 38419 2858
rect 37432 2745 37581 2756
rect 37432 1568 37537 2745
rect 38199 2730 38243 2838
rect 38375 2730 38419 2838
rect 38199 2688 38419 2730
rect 40997 2703 41059 4274
rect 41249 4266 41295 4278
rect 41249 3890 41255 4266
rect 41289 3890 41295 4266
rect 41249 3878 41295 3890
rect 41367 4266 41413 4278
rect 41367 3890 41373 4266
rect 41407 3890 41413 4266
rect 41367 3878 41413 3890
rect 41485 4266 41531 4278
rect 41485 3890 41491 4266
rect 41525 3890 41531 4266
rect 41485 3878 41531 3890
rect 41603 4266 41649 4278
rect 41603 3890 41609 4266
rect 41643 3890 41649 4266
rect 41603 3878 41649 3890
rect 41721 4266 41767 4278
rect 41721 3890 41727 4266
rect 41761 3890 41767 4266
rect 41721 3878 41767 3890
rect 41839 4266 41885 4278
rect 41839 3890 41845 4266
rect 41879 3890 41885 4266
rect 41839 3878 41885 3890
rect 41957 4266 42003 4278
rect 41957 3890 41963 4266
rect 41997 3890 42003 4266
rect 41957 3878 42003 3890
rect 41255 3836 41289 3878
rect 41491 3836 41525 3878
rect 41255 3808 41525 3836
rect 41609 3837 41643 3878
rect 41845 3837 41879 3878
rect 41609 3808 41879 3837
rect 41255 3760 41289 3808
rect 41255 3730 41318 3760
rect 41283 3638 41318 3730
rect 41790 3700 41890 3721
rect 41790 3646 41804 3700
rect 41869 3646 41890 3700
rect 41790 3641 41890 3646
rect 41963 3695 41997 3878
rect 43197 3710 43309 8595
rect 43833 7230 43926 9124
rect 43989 9065 44455 9087
rect 44743 9065 44809 9161
rect 46574 9171 46580 9347
rect 46614 9171 46620 9347
rect 46574 9159 46620 9171
rect 46692 9347 46738 9359
rect 46692 9171 46698 9347
rect 46732 9171 46738 9347
rect 46692 9159 46738 9171
rect 46810 9347 46856 9359
rect 46810 9171 46816 9347
rect 46850 9171 46856 9347
rect 46810 9159 46856 9171
rect 46928 9347 46974 9359
rect 46928 9171 46934 9347
rect 46968 9292 46974 9347
rect 47093 9347 47139 9359
rect 47093 9292 47099 9347
rect 46968 9204 47099 9292
rect 46968 9171 46974 9204
rect 46928 9159 46974 9171
rect 47093 9171 47099 9204
rect 47133 9171 47139 9347
rect 47093 9159 47139 9171
rect 47211 9347 47257 9359
rect 47211 9171 47217 9347
rect 47251 9171 47257 9347
rect 47211 9159 47257 9171
rect 47329 9347 47375 9359
rect 47329 9171 47335 9347
rect 47369 9171 47375 9347
rect 47329 9159 47375 9171
rect 47447 9347 47493 9359
rect 47447 9171 47453 9347
rect 47487 9171 47493 9347
rect 47447 9159 47493 9171
rect 46580 9120 46614 9159
rect 46816 9120 46850 9159
rect 46580 9085 46850 9120
rect 47217 9121 47250 9159
rect 47453 9121 47486 9159
rect 47217 9085 47486 9121
rect 43989 9017 44809 9065
rect 46614 9084 46850 9085
rect 43989 8986 44455 9017
rect 46614 9010 46746 9084
rect 43989 8730 44094 8986
rect 46604 8902 46614 9010
rect 46746 8902 46756 9010
rect 44828 8821 44907 8833
rect 43989 8624 44052 8730
rect 44164 8624 44174 8730
rect 44828 8726 44834 8821
rect 44756 8706 44834 8726
rect 44901 8726 44907 8821
rect 46637 8772 46643 8902
rect 46710 8772 46716 8902
rect 46637 8760 46716 8772
rect 44901 8706 44976 8726
rect 43989 8613 44138 8624
rect 43989 7436 44094 8613
rect 44756 8598 44800 8706
rect 44932 8598 44976 8706
rect 44756 8556 44976 8598
rect 47554 8571 47616 10142
rect 47806 10134 47852 10146
rect 47806 9758 47812 10134
rect 47846 9758 47852 10134
rect 47806 9746 47852 9758
rect 47924 10134 47970 10146
rect 47924 9758 47930 10134
rect 47964 9758 47970 10134
rect 47924 9746 47970 9758
rect 48042 10134 48088 10146
rect 48042 9758 48048 10134
rect 48082 9758 48088 10134
rect 48042 9746 48088 9758
rect 48160 10134 48206 10146
rect 48160 9758 48166 10134
rect 48200 9758 48206 10134
rect 48160 9746 48206 9758
rect 48278 10134 48324 10146
rect 48278 9758 48284 10134
rect 48318 9758 48324 10134
rect 48278 9746 48324 9758
rect 48396 10134 48442 10146
rect 48396 9758 48402 10134
rect 48436 9758 48442 10134
rect 48396 9746 48442 9758
rect 48514 10134 48560 10146
rect 48514 9758 48520 10134
rect 48554 9758 48560 10134
rect 48514 9746 48560 9758
rect 47812 9704 47846 9746
rect 48048 9704 48082 9746
rect 47812 9676 48082 9704
rect 48166 9705 48200 9746
rect 48402 9705 48436 9746
rect 48166 9676 48436 9705
rect 47812 9628 47846 9676
rect 47812 9598 47875 9628
rect 47840 9506 47875 9598
rect 48347 9568 48447 9589
rect 48347 9514 48361 9568
rect 48426 9514 48447 9568
rect 48347 9509 48447 9514
rect 48520 9563 48554 9746
rect 48520 9509 48629 9563
rect 47840 9470 48067 9506
rect 47840 9363 47875 9470
rect 48001 9436 48067 9470
rect 48001 9402 48017 9436
rect 48051 9402 48067 9436
rect 48348 9494 48445 9509
rect 48348 9427 48405 9494
rect 48001 9396 48067 9402
rect 48242 9391 48511 9427
rect 48242 9363 48275 9391
rect 48478 9363 48511 9391
rect 48595 9363 48629 9509
rect 49446 9502 49456 9577
rect 49524 9502 49918 9577
rect 49473 9501 49918 9502
rect 47716 9351 47762 9363
rect 47716 9175 47722 9351
rect 47756 9175 47762 9351
rect 47716 9163 47762 9175
rect 47834 9351 47880 9363
rect 47834 9175 47840 9351
rect 47874 9175 47880 9351
rect 47834 9163 47880 9175
rect 47952 9351 47998 9363
rect 47952 9175 47958 9351
rect 47992 9175 47998 9351
rect 47952 9163 47998 9175
rect 48070 9351 48116 9363
rect 48070 9175 48076 9351
rect 48110 9296 48116 9351
rect 48235 9351 48281 9363
rect 48235 9296 48241 9351
rect 48110 9208 48241 9296
rect 48110 9175 48116 9208
rect 48070 9163 48116 9175
rect 48235 9175 48241 9208
rect 48275 9175 48281 9351
rect 48235 9163 48281 9175
rect 48353 9351 48399 9363
rect 48353 9175 48359 9351
rect 48393 9175 48399 9351
rect 48353 9163 48399 9175
rect 48471 9351 48517 9363
rect 48471 9175 48477 9351
rect 48511 9175 48517 9351
rect 48471 9163 48517 9175
rect 48589 9351 48635 9363
rect 48589 9175 48595 9351
rect 48629 9175 48635 9351
rect 48589 9163 48635 9175
rect 47722 9124 47756 9163
rect 47958 9124 47992 9163
rect 47722 9088 47992 9124
rect 48359 9125 48392 9163
rect 48595 9125 48628 9163
rect 48359 9089 48628 9125
rect 47722 9087 47888 9088
rect 47756 9008 47888 9087
rect 47746 8900 47756 9008
rect 47888 8900 47898 9008
rect 47776 8764 47782 8900
rect 47849 8764 47855 8900
rect 47776 8752 47855 8764
rect 44360 8526 45337 8556
rect 47554 8554 47617 8571
rect 47479 8550 47617 8554
rect 44360 8420 44392 8526
rect 44596 8420 44628 8526
rect 44832 8420 44864 8526
rect 45068 8420 45100 8526
rect 45303 8420 45337 8526
rect 45647 8516 47617 8550
rect 45645 8487 47617 8516
rect 45645 8471 45691 8487
rect 47479 8485 47617 8487
rect 44353 8408 44399 8420
rect 44353 8232 44359 8408
rect 44393 8232 44399 8408
rect 44353 8220 44399 8232
rect 44471 8408 44517 8420
rect 44471 8232 44477 8408
rect 44511 8232 44517 8408
rect 44471 8220 44517 8232
rect 44589 8408 44635 8420
rect 44589 8232 44595 8408
rect 44629 8232 44635 8408
rect 44589 8220 44635 8232
rect 44707 8408 44753 8420
rect 44707 8232 44713 8408
rect 44747 8232 44753 8408
rect 44707 8220 44753 8232
rect 44825 8408 44871 8420
rect 44825 8232 44831 8408
rect 44865 8232 44871 8408
rect 44825 8220 44871 8232
rect 44943 8408 44989 8420
rect 44943 8232 44949 8408
rect 44983 8232 44989 8408
rect 44943 8220 44989 8232
rect 45061 8408 45107 8420
rect 45061 8232 45067 8408
rect 45101 8232 45107 8408
rect 45061 8220 45107 8232
rect 45179 8408 45225 8420
rect 45179 8232 45185 8408
rect 45219 8232 45225 8408
rect 45179 8220 45225 8232
rect 45297 8408 45343 8420
rect 45297 8232 45303 8408
rect 45337 8232 45343 8408
rect 45297 8220 45343 8232
rect 45415 8408 45461 8420
rect 45415 8232 45421 8408
rect 45455 8232 45461 8408
rect 45415 8220 45461 8232
rect 44476 8126 44512 8220
rect 44712 8126 44748 8220
rect 44948 8127 44984 8220
rect 45110 8172 45176 8179
rect 45110 8138 45126 8172
rect 45160 8138 45176 8172
rect 45110 8127 45176 8138
rect 44948 8126 45176 8127
rect 44476 8097 45176 8126
rect 44476 8096 45058 8097
rect 44596 7983 44630 8096
rect 44992 8055 45058 8096
rect 44992 8021 45008 8055
rect 45042 8021 45058 8055
rect 44992 8014 45058 8021
rect 45420 8002 45455 8220
rect 45644 8019 45691 8471
rect 48543 8479 48622 8491
rect 48543 8363 48549 8479
rect 48616 8363 48622 8479
rect 46603 8255 46613 8363
rect 46745 8255 46755 8363
rect 48501 8255 48511 8363
rect 48643 8255 48653 8363
rect 46613 8215 46745 8255
rect 48511 8215 48643 8255
rect 46612 8149 46745 8215
rect 48510 8149 48643 8215
rect 45941 8106 47414 8149
rect 45644 8003 45690 8019
rect 45609 8002 45690 8003
rect 45420 7987 45690 8002
rect 45066 7983 45690 7987
rect 44590 7971 44636 7983
rect 44325 7493 44335 7611
rect 44453 7579 44463 7611
rect 44590 7595 44596 7971
rect 44630 7595 44636 7971
rect 44590 7583 44636 7595
rect 44708 7971 44754 7983
rect 44708 7595 44714 7971
rect 44748 7595 44754 7971
rect 44708 7583 44754 7595
rect 44826 7971 44872 7983
rect 44826 7595 44832 7971
rect 44866 7619 44872 7971
rect 44943 7971 44989 7983
rect 44943 7795 44949 7971
rect 44983 7795 44989 7971
rect 44943 7783 44989 7795
rect 45061 7971 45690 7983
rect 45061 7795 45067 7971
rect 45101 7959 45690 7971
rect 45101 7958 45343 7959
rect 45101 7795 45107 7958
rect 45609 7957 45690 7959
rect 45941 7803 45975 8106
rect 46307 8003 46341 8106
rect 46543 8003 46577 8106
rect 46779 8003 46813 8106
rect 47015 8003 47049 8106
rect 46301 7991 46347 8003
rect 45061 7783 45107 7795
rect 45817 7791 45863 7803
rect 44949 7667 44984 7783
rect 45080 7667 45188 7677
rect 44949 7619 45080 7667
rect 45188 7628 45337 7634
rect 44866 7595 45080 7619
rect 44826 7583 45080 7595
rect 44832 7579 45080 7583
rect 44453 7551 44468 7579
rect 44453 7545 44705 7551
rect 44453 7511 44655 7545
rect 44689 7511 44705 7545
rect 44453 7495 44705 7511
rect 44757 7545 44823 7551
rect 44757 7511 44773 7545
rect 44807 7511 44823 7545
rect 45006 7535 45080 7579
rect 45325 7561 45337 7628
rect 45817 7615 45823 7791
rect 45857 7615 45863 7791
rect 45817 7603 45863 7615
rect 45935 7791 45981 7803
rect 45935 7615 45941 7791
rect 45975 7615 45981 7791
rect 45935 7603 45981 7615
rect 46053 7791 46099 7803
rect 46053 7615 46059 7791
rect 46093 7615 46099 7791
rect 46053 7603 46099 7615
rect 46171 7791 46217 7803
rect 46301 7791 46307 7991
rect 46171 7615 46177 7791
rect 46211 7615 46307 7791
rect 46341 7615 46347 7991
rect 46171 7603 46217 7615
rect 46301 7603 46347 7615
rect 46419 7991 46465 8003
rect 46419 7615 46425 7991
rect 46459 7615 46465 7991
rect 46419 7603 46465 7615
rect 46537 7991 46583 8003
rect 46537 7615 46543 7991
rect 46577 7615 46583 7991
rect 46537 7603 46583 7615
rect 46655 7991 46701 8003
rect 46655 7615 46661 7991
rect 46695 7615 46701 7991
rect 46655 7603 46701 7615
rect 46773 7991 46819 8003
rect 46773 7615 46779 7991
rect 46813 7615 46819 7991
rect 46773 7603 46819 7615
rect 46891 7991 46937 8003
rect 46891 7615 46897 7991
rect 46931 7615 46937 7991
rect 46891 7603 46937 7615
rect 47009 7991 47055 8003
rect 47009 7615 47015 7991
rect 47049 7791 47055 7991
rect 47380 7803 47414 8106
rect 47839 8106 49312 8149
rect 47839 7803 47873 8106
rect 48205 8003 48239 8106
rect 48441 8003 48475 8106
rect 48677 8003 48711 8106
rect 48913 8003 48947 8106
rect 48199 7991 48245 8003
rect 47138 7791 47184 7803
rect 47049 7615 47144 7791
rect 47178 7615 47184 7791
rect 47009 7603 47055 7615
rect 47138 7603 47184 7615
rect 47256 7791 47302 7803
rect 47256 7615 47262 7791
rect 47296 7615 47302 7791
rect 47256 7603 47302 7615
rect 47374 7791 47420 7803
rect 47374 7615 47380 7791
rect 47414 7615 47420 7791
rect 47374 7603 47420 7615
rect 47492 7791 47538 7803
rect 47492 7615 47498 7791
rect 47532 7615 47538 7791
rect 47492 7603 47538 7615
rect 47715 7791 47761 7803
rect 47715 7615 47721 7791
rect 47755 7615 47761 7791
rect 47715 7603 47761 7615
rect 47833 7791 47879 7803
rect 47833 7615 47839 7791
rect 47873 7615 47879 7791
rect 47833 7603 47879 7615
rect 47951 7791 47997 7803
rect 47951 7615 47957 7791
rect 47991 7615 47997 7791
rect 47951 7603 47997 7615
rect 48069 7791 48115 7803
rect 48199 7791 48205 7991
rect 48069 7615 48075 7791
rect 48109 7615 48205 7791
rect 48239 7615 48245 7991
rect 48069 7603 48115 7615
rect 48199 7603 48245 7615
rect 48317 7991 48363 8003
rect 48317 7615 48323 7991
rect 48357 7615 48363 7991
rect 48317 7603 48363 7615
rect 48435 7991 48481 8003
rect 48435 7615 48441 7991
rect 48475 7615 48481 7991
rect 48435 7603 48481 7615
rect 48553 7991 48599 8003
rect 48553 7615 48559 7991
rect 48593 7615 48599 7991
rect 48553 7603 48599 7615
rect 48671 7991 48717 8003
rect 48671 7615 48677 7991
rect 48711 7615 48717 7991
rect 48671 7603 48717 7615
rect 48789 7991 48835 8003
rect 48789 7615 48795 7991
rect 48829 7615 48835 7991
rect 48789 7603 48835 7615
rect 48907 7991 48953 8003
rect 48907 7615 48913 7991
rect 48947 7791 48953 7991
rect 49278 7803 49312 8106
rect 49036 7791 49082 7803
rect 48947 7615 49042 7791
rect 49076 7615 49082 7791
rect 48907 7603 48953 7615
rect 49036 7603 49082 7615
rect 49154 7791 49200 7803
rect 49154 7615 49160 7791
rect 49194 7615 49200 7791
rect 49154 7603 49200 7615
rect 49272 7791 49318 7803
rect 49272 7615 49278 7791
rect 49312 7615 49318 7791
rect 49272 7603 49318 7615
rect 49390 7791 49436 7803
rect 49390 7615 49396 7791
rect 49430 7615 49436 7791
rect 49390 7603 49436 7615
rect 45188 7555 45337 7561
rect 45823 7569 45857 7603
rect 46425 7569 46459 7603
rect 46661 7569 46695 7603
rect 45080 7525 45188 7535
rect 45823 7534 45982 7569
rect 46425 7534 46695 7569
rect 47262 7569 47296 7603
rect 47498 7569 47532 7603
rect 47262 7534 47532 7569
rect 47721 7569 47755 7603
rect 48323 7569 48357 7603
rect 48559 7569 48593 7603
rect 47721 7534 47880 7569
rect 48323 7534 48593 7569
rect 49160 7569 49194 7603
rect 49396 7569 49430 7603
rect 49160 7534 49430 7569
rect 44453 7493 44468 7495
rect 44368 7479 44468 7493
rect 44368 7436 44468 7437
rect 43989 7415 44468 7436
rect 44757 7415 44823 7511
rect 43989 7367 44823 7415
rect 43989 7338 44468 7367
rect 43989 7336 44094 7338
rect 44368 7337 44468 7338
rect 43822 7151 43832 7230
rect 43925 7151 43935 7230
rect 44820 7221 44899 7233
rect 43833 5977 43926 7151
rect 44820 7122 44826 7221
rect 44751 7102 44826 7122
rect 44893 7122 44899 7221
rect 44893 7102 44971 7122
rect 44751 6994 44795 7102
rect 44927 6994 44971 7102
rect 44751 6952 44971 6994
rect 44355 6922 45332 6952
rect 44355 6816 44387 6922
rect 44591 6816 44623 6922
rect 44827 6816 44859 6922
rect 45063 6816 45095 6922
rect 45298 6816 45332 6922
rect 44348 6804 44394 6816
rect 44348 6628 44354 6804
rect 44388 6628 44394 6804
rect 44348 6616 44394 6628
rect 44466 6804 44512 6816
rect 44466 6628 44472 6804
rect 44506 6628 44512 6804
rect 44466 6616 44512 6628
rect 44584 6804 44630 6816
rect 44584 6628 44590 6804
rect 44624 6628 44630 6804
rect 44584 6616 44630 6628
rect 44702 6804 44748 6816
rect 44702 6628 44708 6804
rect 44742 6628 44748 6804
rect 44702 6616 44748 6628
rect 44820 6804 44866 6816
rect 44820 6628 44826 6804
rect 44860 6628 44866 6804
rect 44820 6616 44866 6628
rect 44938 6804 44984 6816
rect 44938 6628 44944 6804
rect 44978 6628 44984 6804
rect 44938 6616 44984 6628
rect 45056 6804 45102 6816
rect 45056 6628 45062 6804
rect 45096 6628 45102 6804
rect 45056 6616 45102 6628
rect 45174 6804 45220 6816
rect 45174 6628 45180 6804
rect 45214 6628 45220 6804
rect 45174 6616 45220 6628
rect 45292 6804 45338 6816
rect 45292 6628 45298 6804
rect 45332 6628 45338 6804
rect 45292 6616 45338 6628
rect 45410 6804 45456 6816
rect 45410 6628 45416 6804
rect 45450 6628 45456 6804
rect 45410 6616 45456 6628
rect 45948 6750 45982 7534
rect 46661 7472 46695 7534
rect 46250 7434 46992 7472
rect 46250 7310 46284 7434
rect 46486 7310 46520 7434
rect 46722 7310 46756 7434
rect 46958 7310 46992 7434
rect 47248 7327 47258 7393
rect 47321 7327 47331 7393
rect 46244 7298 46290 7310
rect 46244 6922 46250 7298
rect 46284 6922 46290 7298
rect 46244 6910 46290 6922
rect 46362 7298 46408 7310
rect 46362 6922 46368 7298
rect 46402 6922 46408 7298
rect 46362 6910 46408 6922
rect 46480 7298 46526 7310
rect 46480 6922 46486 7298
rect 46520 6922 46526 7298
rect 46480 6910 46526 6922
rect 46598 7298 46644 7310
rect 46598 6922 46604 7298
rect 46638 6922 46644 7298
rect 46598 6910 46644 6922
rect 46716 7298 46762 7310
rect 46716 6922 46722 7298
rect 46756 6922 46762 7298
rect 46716 6910 46762 6922
rect 46834 7298 46880 7310
rect 46834 6922 46840 7298
rect 46874 6922 46880 7298
rect 46834 6910 46880 6922
rect 46952 7298 46998 7310
rect 46952 6922 46958 7298
rect 46992 6922 46998 7298
rect 46952 6910 46998 6922
rect 47364 6751 47398 7534
rect 47091 6750 47398 6751
rect 45948 6745 46264 6750
rect 46978 6745 47398 6750
rect 45948 6734 46331 6745
rect 45948 6707 46280 6734
rect 44471 6522 44507 6616
rect 44707 6522 44743 6616
rect 44943 6523 44979 6616
rect 45105 6568 45171 6575
rect 45105 6534 45121 6568
rect 45155 6534 45171 6568
rect 45105 6523 45171 6534
rect 44943 6522 45171 6523
rect 44471 6493 45171 6522
rect 44471 6492 45053 6493
rect 44591 6379 44625 6492
rect 44987 6451 45053 6492
rect 44987 6417 45003 6451
rect 45037 6417 45053 6451
rect 44987 6410 45053 6417
rect 45415 6383 45450 6616
rect 45948 6578 45982 6707
rect 46264 6700 46280 6707
rect 46314 6700 46331 6734
rect 46264 6694 46331 6700
rect 46911 6734 47398 6745
rect 46911 6700 46928 6734
rect 46962 6707 47398 6734
rect 46962 6700 46978 6707
rect 47091 6706 47398 6707
rect 46911 6694 46978 6700
rect 46089 6667 46145 6679
rect 46089 6633 46095 6667
rect 46129 6666 46145 6667
rect 47202 6666 47258 6678
rect 46129 6650 46596 6666
rect 46129 6633 46546 6650
rect 46089 6617 46546 6633
rect 46530 6616 46546 6617
rect 46580 6616 46596 6650
rect 46530 6609 46596 6616
rect 46648 6651 47218 6666
rect 46648 6617 46664 6651
rect 46698 6632 47218 6651
rect 47252 6632 47258 6666
rect 46698 6617 47258 6632
rect 46648 6607 46715 6617
rect 47202 6616 47258 6617
rect 47364 6578 47398 6706
rect 47846 6750 47880 7534
rect 48559 7472 48593 7534
rect 48148 7434 48890 7472
rect 48148 7310 48182 7434
rect 48384 7310 48418 7434
rect 48620 7310 48654 7434
rect 48856 7310 48890 7434
rect 48142 7298 48188 7310
rect 48142 6922 48148 7298
rect 48182 6922 48188 7298
rect 48142 6910 48188 6922
rect 48260 7298 48306 7310
rect 48260 6922 48266 7298
rect 48300 6922 48306 7298
rect 48260 6910 48306 6922
rect 48378 7298 48424 7310
rect 48378 6922 48384 7298
rect 48418 6922 48424 7298
rect 48378 6910 48424 6922
rect 48496 7298 48542 7310
rect 48496 6922 48502 7298
rect 48536 6922 48542 7298
rect 48496 6910 48542 6922
rect 48614 7298 48660 7310
rect 48614 6922 48620 7298
rect 48654 6922 48660 7298
rect 48614 6910 48660 6922
rect 48732 7298 48778 7310
rect 48732 6922 48738 7298
rect 48772 6922 48778 7298
rect 48732 6910 48778 6922
rect 48850 7298 48896 7310
rect 48850 6922 48856 7298
rect 48890 6922 48896 7298
rect 48850 6910 48896 6922
rect 49262 6751 49296 7534
rect 48874 6750 48943 6751
rect 48989 6750 49296 6751
rect 47846 6745 48162 6750
rect 48874 6746 49296 6750
rect 47846 6734 48229 6745
rect 47846 6707 48178 6734
rect 47846 6578 47880 6707
rect 48162 6700 48178 6707
rect 48212 6700 48229 6734
rect 48162 6694 48229 6700
rect 48807 6735 49296 6746
rect 48807 6701 48824 6735
rect 48858 6707 49296 6735
rect 48858 6701 48874 6707
rect 48989 6706 49296 6707
rect 48807 6695 48874 6701
rect 47987 6667 48043 6679
rect 47987 6633 47993 6667
rect 48027 6666 48043 6667
rect 49100 6666 49156 6678
rect 48027 6650 48494 6666
rect 48027 6633 48444 6650
rect 47987 6617 48444 6633
rect 48428 6616 48444 6617
rect 48478 6616 48494 6650
rect 48428 6609 48494 6616
rect 48546 6651 49116 6666
rect 48546 6617 48562 6651
rect 48596 6632 49116 6651
rect 49150 6632 49156 6666
rect 48596 6617 49156 6632
rect 48546 6607 48613 6617
rect 49100 6616 49156 6617
rect 49262 6578 49296 6706
rect 49377 7356 49444 7380
rect 49377 7322 49394 7356
rect 49428 7322 49444 7356
rect 45061 6379 45450 6383
rect 44585 6367 44631 6379
rect 44585 5991 44591 6367
rect 44625 5991 44631 6367
rect 44585 5979 44631 5991
rect 44703 6367 44749 6379
rect 44703 5991 44709 6367
rect 44743 5991 44749 6367
rect 44703 5979 44749 5991
rect 44821 6367 44867 6379
rect 44821 5991 44827 6367
rect 44861 6015 44867 6367
rect 44938 6367 44984 6379
rect 44938 6191 44944 6367
rect 44978 6191 44984 6367
rect 44938 6179 44984 6191
rect 45056 6367 45450 6379
rect 45942 6566 45988 6578
rect 45942 6390 45948 6566
rect 45982 6390 45988 6566
rect 45942 6378 45988 6390
rect 46060 6566 46106 6578
rect 46060 6390 46066 6566
rect 46100 6390 46106 6566
rect 46060 6378 46106 6390
rect 46362 6566 46408 6578
rect 45056 6191 45062 6367
rect 45096 6354 45450 6367
rect 45096 6191 45102 6354
rect 45372 6351 45450 6354
rect 45372 6299 45382 6351
rect 45445 6299 45455 6351
rect 45377 6293 45450 6299
rect 45056 6179 45102 6191
rect 44944 6063 44979 6179
rect 46065 6084 46099 6378
rect 46362 6190 46368 6566
rect 46402 6190 46408 6566
rect 46362 6178 46408 6190
rect 46480 6566 46526 6578
rect 46480 6190 46486 6566
rect 46520 6190 46526 6566
rect 46480 6178 46526 6190
rect 46598 6566 46644 6578
rect 46598 6190 46604 6566
rect 46638 6190 46644 6566
rect 46598 6178 46644 6190
rect 46716 6566 46762 6578
rect 46716 6190 46722 6566
rect 46756 6190 46762 6566
rect 46716 6178 46762 6190
rect 46834 6566 46880 6578
rect 46834 6190 46840 6566
rect 46874 6190 46880 6566
rect 47240 6566 47286 6578
rect 47240 6390 47246 6566
rect 47280 6390 47286 6566
rect 47240 6378 47286 6390
rect 47358 6566 47404 6578
rect 47358 6390 47364 6566
rect 47398 6390 47404 6566
rect 47358 6378 47404 6390
rect 47840 6566 47886 6578
rect 47840 6390 47846 6566
rect 47880 6390 47886 6566
rect 47840 6378 47886 6390
rect 47958 6566 48004 6578
rect 47958 6390 47964 6566
rect 47998 6390 48004 6566
rect 47958 6378 48004 6390
rect 48260 6566 48306 6578
rect 46834 6178 46880 6190
rect 46722 6084 46756 6178
rect 47246 6084 47279 6378
rect 45075 6063 45183 6073
rect 44944 6015 45075 6063
rect 46065 6052 47279 6084
rect 47963 6084 47997 6378
rect 48260 6190 48266 6566
rect 48300 6190 48306 6566
rect 48260 6178 48306 6190
rect 48378 6566 48424 6578
rect 48378 6190 48384 6566
rect 48418 6190 48424 6566
rect 48378 6178 48424 6190
rect 48496 6566 48542 6578
rect 48496 6190 48502 6566
rect 48536 6190 48542 6566
rect 48496 6178 48542 6190
rect 48614 6566 48660 6578
rect 48614 6190 48620 6566
rect 48654 6190 48660 6566
rect 48614 6178 48660 6190
rect 48732 6566 48778 6578
rect 48732 6190 48738 6566
rect 48772 6190 48778 6566
rect 49138 6566 49184 6578
rect 49138 6390 49144 6566
rect 49178 6390 49184 6566
rect 49138 6378 49184 6390
rect 49256 6566 49302 6578
rect 49256 6390 49262 6566
rect 49296 6390 49302 6566
rect 49256 6378 49302 6390
rect 48732 6178 48778 6190
rect 48620 6084 48654 6178
rect 49144 6084 49177 6378
rect 47963 6052 49177 6084
rect 45183 6027 45334 6033
rect 44861 5991 45075 6015
rect 44821 5979 45075 5991
rect 43833 5975 44418 5977
rect 44827 5975 45075 5979
rect 43833 5947 44463 5975
rect 43833 5941 44700 5947
rect 43833 5907 44650 5941
rect 44684 5907 44700 5941
rect 43833 5891 44700 5907
rect 44752 5941 44818 5947
rect 44752 5907 44768 5941
rect 44802 5907 44818 5941
rect 45001 5931 45075 5975
rect 45322 5960 45334 6027
rect 46558 5967 46690 6052
rect 48456 5967 48588 6052
rect 45183 5954 45334 5960
rect 45075 5921 45183 5931
rect 43833 5875 44463 5891
rect 43833 5871 44418 5875
rect 43833 5870 43934 5871
rect 44363 5822 44463 5833
rect 44327 5716 44337 5822
rect 44449 5811 44463 5822
rect 44752 5811 44818 5907
rect 46548 5859 46558 5967
rect 46690 5859 46700 5967
rect 48446 5859 48456 5967
rect 48588 5859 48598 5967
rect 49377 5939 49444 7322
rect 49505 6893 49661 6899
rect 49505 6795 49517 6893
rect 49649 6795 49661 6893
rect 49505 6789 49661 6795
rect 44449 5763 44818 5811
rect 44449 5733 44463 5763
rect 44449 5716 44459 5733
rect 44751 5660 44817 5763
rect 46581 5721 46587 5859
rect 46654 5721 46660 5859
rect 46581 5709 46660 5721
rect 49377 5660 49443 5939
rect 44749 5580 49443 5660
rect 47289 4656 47368 4668
rect 44808 4603 44887 4615
rect 44808 4506 44814 4603
rect 44736 4486 44814 4506
rect 44881 4506 44887 4603
rect 47289 4540 47295 4656
rect 47362 4540 47368 4656
rect 48437 4656 48516 4668
rect 48437 4540 48443 4656
rect 48510 4540 48516 4656
rect 44881 4486 44956 4506
rect 44736 4378 44780 4486
rect 44912 4378 44956 4486
rect 46533 4444 46589 4452
rect 44736 4336 44956 4378
rect 45607 4436 46589 4444
rect 45607 4402 46549 4436
rect 46583 4402 46589 4436
rect 47252 4432 47262 4540
rect 47394 4477 47404 4540
rect 47394 4466 47406 4477
rect 47394 4432 47407 4466
rect 47663 4456 47719 4458
rect 45607 4386 46589 4402
rect 47262 4394 47407 4432
rect 45607 4385 46586 4386
rect 44340 4306 45317 4336
rect 44340 4200 44372 4306
rect 44576 4200 44608 4306
rect 44812 4200 44844 4306
rect 45048 4200 45080 4306
rect 45283 4200 45317 4306
rect 44333 4188 44379 4200
rect 44333 4012 44339 4188
rect 44373 4012 44379 4188
rect 44333 4000 44379 4012
rect 44451 4188 44497 4200
rect 44451 4012 44457 4188
rect 44491 4012 44497 4188
rect 44451 4000 44497 4012
rect 44569 4188 44615 4200
rect 44569 4012 44575 4188
rect 44609 4012 44615 4188
rect 44569 4000 44615 4012
rect 44687 4188 44733 4200
rect 44687 4012 44693 4188
rect 44727 4012 44733 4188
rect 44687 4000 44733 4012
rect 44805 4188 44851 4200
rect 44805 4012 44811 4188
rect 44845 4012 44851 4188
rect 44805 4000 44851 4012
rect 44923 4188 44969 4200
rect 44923 4012 44929 4188
rect 44963 4012 44969 4188
rect 44923 4000 44969 4012
rect 45041 4188 45087 4200
rect 45041 4012 45047 4188
rect 45081 4012 45087 4188
rect 45041 4000 45087 4012
rect 45159 4188 45205 4200
rect 45159 4012 45165 4188
rect 45199 4012 45205 4188
rect 45159 4000 45205 4012
rect 45277 4188 45323 4200
rect 45277 4012 45283 4188
rect 45317 4012 45323 4188
rect 45277 4000 45323 4012
rect 45395 4188 45441 4200
rect 45395 4012 45401 4188
rect 45435 4012 45441 4188
rect 45395 4000 45441 4012
rect 44456 3906 44492 4000
rect 44692 3906 44728 4000
rect 44928 3907 44964 4000
rect 45090 3952 45156 3959
rect 45090 3918 45106 3952
rect 45140 3918 45156 3952
rect 45090 3907 45156 3918
rect 44928 3906 45156 3907
rect 44456 3877 45156 3906
rect 44456 3876 45038 3877
rect 44576 3763 44610 3876
rect 44972 3835 45038 3876
rect 44972 3801 44988 3835
rect 45022 3801 45038 3835
rect 44972 3794 45038 3801
rect 45400 3795 45435 4000
rect 45607 3795 45674 4385
rect 47366 4362 47407 4394
rect 47653 4390 47663 4456
rect 47719 4390 47729 4456
rect 48399 4432 48409 4540
rect 48541 4477 48551 4540
rect 48541 4466 48553 4477
rect 48541 4432 48554 4466
rect 48409 4394 48554 4432
rect 48513 4366 48554 4394
rect 46782 4334 47052 4362
rect 46523 4268 46533 4334
rect 46599 4268 46609 4334
rect 46782 4272 46816 4334
rect 47018 4272 47052 4334
rect 47136 4334 47407 4362
rect 47924 4338 48194 4366
rect 47136 4272 47170 4334
rect 47372 4272 47407 4334
rect 47548 4322 47719 4338
rect 47548 4288 47679 4322
rect 47713 4288 47719 4322
rect 47548 4272 47719 4288
rect 47924 4276 47958 4338
rect 48160 4276 48194 4338
rect 48278 4338 48554 4366
rect 48278 4276 48312 4338
rect 48514 4276 48554 4338
rect 46658 4260 46704 4272
rect 46658 3884 46664 4260
rect 46698 3884 46704 4260
rect 46658 3872 46704 3884
rect 46776 4260 46822 4272
rect 46776 3884 46782 4260
rect 46816 3884 46822 4260
rect 46776 3872 46822 3884
rect 46894 4260 46940 4272
rect 46894 3884 46900 4260
rect 46934 3884 46940 4260
rect 46894 3872 46940 3884
rect 47012 4260 47058 4272
rect 47012 3884 47018 4260
rect 47052 3884 47058 4260
rect 47012 3872 47058 3884
rect 47130 4260 47176 4272
rect 47130 3884 47136 4260
rect 47170 3884 47176 4260
rect 47130 3872 47176 3884
rect 47248 4260 47294 4272
rect 47248 3884 47254 4260
rect 47288 3884 47294 4260
rect 47248 3872 47294 3884
rect 47366 4260 47412 4272
rect 47366 3884 47372 4260
rect 47406 3884 47412 4260
rect 47366 3872 47412 3884
rect 45400 3767 45674 3795
rect 45046 3763 45674 3767
rect 42954 3709 43309 3710
rect 41963 3641 42072 3695
rect 41283 3602 41510 3638
rect 41283 3495 41318 3602
rect 41444 3568 41510 3602
rect 41444 3534 41460 3568
rect 41494 3534 41510 3568
rect 41791 3626 41888 3641
rect 41791 3559 41848 3626
rect 41444 3528 41510 3534
rect 41685 3523 41954 3559
rect 41685 3495 41718 3523
rect 41921 3495 41954 3523
rect 42038 3495 42072 3641
rect 42889 3634 42899 3709
rect 42967 3634 43309 3709
rect 42916 3633 43309 3634
rect 42954 3632 43309 3633
rect 44570 3751 44616 3763
rect 41159 3483 41205 3495
rect 41159 3307 41165 3483
rect 41199 3307 41205 3483
rect 41159 3295 41205 3307
rect 41277 3483 41323 3495
rect 41277 3307 41283 3483
rect 41317 3307 41323 3483
rect 41277 3295 41323 3307
rect 41395 3483 41441 3495
rect 41395 3307 41401 3483
rect 41435 3307 41441 3483
rect 41395 3295 41441 3307
rect 41513 3483 41559 3495
rect 41513 3307 41519 3483
rect 41553 3428 41559 3483
rect 41678 3483 41724 3495
rect 41678 3428 41684 3483
rect 41553 3340 41684 3428
rect 41553 3307 41559 3340
rect 41513 3295 41559 3307
rect 41678 3307 41684 3340
rect 41718 3307 41724 3483
rect 41678 3295 41724 3307
rect 41796 3483 41842 3495
rect 41796 3307 41802 3483
rect 41836 3307 41842 3483
rect 41796 3295 41842 3307
rect 41914 3483 41960 3495
rect 41914 3307 41920 3483
rect 41954 3307 41960 3483
rect 41914 3295 41960 3307
rect 42032 3483 42078 3495
rect 42032 3307 42038 3483
rect 42072 3307 42078 3483
rect 44570 3375 44576 3751
rect 44610 3375 44616 3751
rect 44570 3363 44616 3375
rect 44688 3751 44734 3763
rect 44688 3375 44694 3751
rect 44728 3375 44734 3751
rect 44688 3363 44734 3375
rect 44806 3751 44852 3763
rect 44806 3375 44812 3751
rect 44846 3399 44852 3751
rect 44923 3751 44969 3763
rect 44923 3575 44929 3751
rect 44963 3575 44969 3751
rect 44923 3563 44969 3575
rect 45041 3751 45674 3763
rect 45041 3575 45047 3751
rect 45081 3738 45674 3751
rect 46664 3830 46698 3872
rect 46900 3830 46934 3872
rect 46664 3802 46934 3830
rect 47018 3831 47052 3872
rect 47254 3831 47288 3872
rect 47018 3802 47288 3831
rect 46664 3754 46698 3802
rect 45081 3575 45087 3738
rect 46664 3724 46727 3754
rect 45041 3563 45087 3575
rect 46692 3632 46727 3724
rect 46692 3596 46919 3632
rect 47189 3621 47199 3718
rect 47298 3621 47308 3718
rect 47372 3689 47406 3872
rect 47372 3635 47481 3689
rect 44929 3447 44964 3563
rect 46692 3489 46727 3596
rect 46853 3562 46919 3596
rect 46853 3528 46869 3562
rect 46903 3528 46919 3562
rect 47200 3620 47297 3621
rect 47200 3553 47257 3620
rect 46853 3522 46919 3528
rect 47094 3517 47363 3553
rect 47094 3489 47127 3517
rect 47330 3489 47363 3517
rect 47447 3489 47481 3635
rect 46568 3477 46614 3489
rect 45060 3447 45168 3457
rect 44929 3399 45060 3447
rect 45168 3403 45313 3409
rect 44846 3375 45060 3399
rect 44806 3363 45060 3375
rect 44812 3359 45060 3363
rect 42032 3295 42078 3307
rect 42948 3331 44448 3358
rect 42948 3325 44685 3331
rect 41165 3256 41199 3295
rect 41401 3256 41435 3295
rect 41165 3220 41435 3256
rect 41802 3257 41835 3295
rect 42038 3257 42071 3295
rect 41802 3221 42071 3257
rect 42948 3291 44635 3325
rect 44669 3291 44685 3325
rect 42948 3275 44685 3291
rect 44737 3325 44803 3331
rect 44737 3291 44753 3325
rect 44787 3291 44803 3325
rect 44986 3315 45060 3359
rect 45301 3336 45313 3403
rect 45168 3330 45313 3336
rect 45060 3305 45168 3315
rect 42948 3259 44448 3275
rect 42948 3258 44385 3259
rect 42948 3252 43920 3258
rect 41165 3219 41331 3220
rect 41199 3140 41331 3219
rect 41189 3032 41199 3140
rect 41331 3032 41341 3140
rect 41226 2894 41232 3032
rect 41299 2894 41305 3032
rect 41226 2882 41305 2894
rect 37803 2658 38780 2688
rect 40997 2686 41060 2703
rect 40922 2682 41060 2686
rect 37803 2552 37835 2658
rect 38039 2552 38071 2658
rect 38275 2552 38307 2658
rect 38511 2552 38543 2658
rect 38746 2552 38780 2658
rect 39090 2648 41060 2682
rect 39088 2619 41060 2648
rect 39088 2603 39134 2619
rect 40922 2617 41060 2619
rect 37796 2540 37842 2552
rect 37796 2364 37802 2540
rect 37836 2364 37842 2540
rect 37796 2352 37842 2364
rect 37914 2540 37960 2552
rect 37914 2364 37920 2540
rect 37954 2364 37960 2540
rect 37914 2352 37960 2364
rect 38032 2540 38078 2552
rect 38032 2364 38038 2540
rect 38072 2364 38078 2540
rect 38032 2352 38078 2364
rect 38150 2540 38196 2552
rect 38150 2364 38156 2540
rect 38190 2364 38196 2540
rect 38150 2352 38196 2364
rect 38268 2540 38314 2552
rect 38268 2364 38274 2540
rect 38308 2364 38314 2540
rect 38268 2352 38314 2364
rect 38386 2540 38432 2552
rect 38386 2364 38392 2540
rect 38426 2364 38432 2540
rect 38386 2352 38432 2364
rect 38504 2540 38550 2552
rect 38504 2364 38510 2540
rect 38544 2364 38550 2540
rect 38504 2352 38550 2364
rect 38622 2540 38668 2552
rect 38622 2364 38628 2540
rect 38662 2364 38668 2540
rect 38622 2352 38668 2364
rect 38740 2540 38786 2552
rect 38740 2364 38746 2540
rect 38780 2364 38786 2540
rect 38740 2352 38786 2364
rect 38858 2540 38904 2552
rect 38858 2364 38864 2540
rect 38898 2364 38904 2540
rect 38858 2352 38904 2364
rect 37919 2258 37955 2352
rect 38155 2258 38191 2352
rect 38391 2259 38427 2352
rect 38553 2304 38619 2311
rect 38553 2270 38569 2304
rect 38603 2270 38619 2304
rect 38553 2259 38619 2270
rect 38391 2258 38619 2259
rect 37919 2229 38619 2258
rect 37919 2228 38501 2229
rect 38039 2115 38073 2228
rect 38435 2187 38501 2228
rect 38435 2153 38451 2187
rect 38485 2153 38501 2187
rect 38435 2146 38501 2153
rect 38863 2134 38898 2352
rect 39087 2151 39134 2603
rect 41980 2611 42059 2623
rect 41980 2495 41986 2611
rect 42053 2495 42059 2611
rect 40046 2387 40056 2495
rect 40188 2387 40198 2495
rect 41944 2387 41954 2495
rect 42086 2387 42096 2495
rect 40056 2347 40188 2387
rect 41954 2347 42086 2387
rect 40055 2281 40188 2347
rect 41953 2281 42086 2347
rect 39384 2238 40857 2281
rect 39087 2135 39133 2151
rect 39052 2134 39133 2135
rect 38863 2119 39133 2134
rect 38509 2115 39133 2119
rect 38033 2103 38079 2115
rect 37768 1625 37778 1743
rect 37896 1711 37906 1743
rect 38033 1727 38039 2103
rect 38073 1727 38079 2103
rect 38033 1715 38079 1727
rect 38151 2103 38197 2115
rect 38151 1727 38157 2103
rect 38191 1727 38197 2103
rect 38151 1715 38197 1727
rect 38269 2103 38315 2115
rect 38269 1727 38275 2103
rect 38309 1751 38315 2103
rect 38386 2103 38432 2115
rect 38386 1927 38392 2103
rect 38426 1927 38432 2103
rect 38386 1915 38432 1927
rect 38504 2103 39133 2115
rect 38504 1927 38510 2103
rect 38544 2091 39133 2103
rect 38544 2090 38786 2091
rect 38544 1927 38550 2090
rect 39052 2089 39133 2091
rect 39384 1935 39418 2238
rect 39750 2135 39784 2238
rect 39986 2135 40020 2238
rect 40222 2135 40256 2238
rect 40458 2135 40492 2238
rect 39744 2123 39790 2135
rect 38504 1915 38550 1927
rect 39260 1923 39306 1935
rect 38392 1799 38427 1915
rect 38523 1799 38631 1809
rect 38392 1751 38523 1799
rect 38631 1759 38771 1765
rect 38309 1727 38523 1751
rect 38269 1715 38523 1727
rect 38275 1711 38523 1715
rect 37896 1683 37911 1711
rect 37896 1677 38148 1683
rect 37896 1643 38098 1677
rect 38132 1643 38148 1677
rect 37896 1627 38148 1643
rect 38200 1677 38266 1683
rect 38200 1643 38216 1677
rect 38250 1643 38266 1677
rect 38449 1667 38523 1711
rect 38759 1692 38771 1759
rect 39260 1747 39266 1923
rect 39300 1747 39306 1923
rect 39260 1735 39306 1747
rect 39378 1923 39424 1935
rect 39378 1747 39384 1923
rect 39418 1747 39424 1923
rect 39378 1735 39424 1747
rect 39496 1923 39542 1935
rect 39496 1747 39502 1923
rect 39536 1747 39542 1923
rect 39496 1735 39542 1747
rect 39614 1923 39660 1935
rect 39744 1923 39750 2123
rect 39614 1747 39620 1923
rect 39654 1747 39750 1923
rect 39784 1747 39790 2123
rect 39614 1735 39660 1747
rect 39744 1735 39790 1747
rect 39862 2123 39908 2135
rect 39862 1747 39868 2123
rect 39902 1747 39908 2123
rect 39862 1735 39908 1747
rect 39980 2123 40026 2135
rect 39980 1747 39986 2123
rect 40020 1747 40026 2123
rect 39980 1735 40026 1747
rect 40098 2123 40144 2135
rect 40098 1747 40104 2123
rect 40138 1747 40144 2123
rect 40098 1735 40144 1747
rect 40216 2123 40262 2135
rect 40216 1747 40222 2123
rect 40256 1747 40262 2123
rect 40216 1735 40262 1747
rect 40334 2123 40380 2135
rect 40334 1747 40340 2123
rect 40374 1747 40380 2123
rect 40334 1735 40380 1747
rect 40452 2123 40498 2135
rect 40452 1747 40458 2123
rect 40492 1923 40498 2123
rect 40823 1935 40857 2238
rect 41282 2238 42755 2281
rect 41282 1935 41316 2238
rect 41648 2135 41682 2238
rect 41884 2135 41918 2238
rect 42120 2135 42154 2238
rect 42356 2135 42390 2238
rect 41642 2123 41688 2135
rect 40581 1923 40627 1935
rect 40492 1747 40587 1923
rect 40621 1747 40627 1923
rect 40452 1735 40498 1747
rect 40581 1735 40627 1747
rect 40699 1923 40745 1935
rect 40699 1747 40705 1923
rect 40739 1747 40745 1923
rect 40699 1735 40745 1747
rect 40817 1923 40863 1935
rect 40817 1747 40823 1923
rect 40857 1747 40863 1923
rect 40817 1735 40863 1747
rect 40935 1923 40981 1935
rect 40935 1747 40941 1923
rect 40975 1747 40981 1923
rect 40935 1735 40981 1747
rect 41158 1923 41204 1935
rect 41158 1747 41164 1923
rect 41198 1747 41204 1923
rect 41158 1735 41204 1747
rect 41276 1923 41322 1935
rect 41276 1747 41282 1923
rect 41316 1747 41322 1923
rect 41276 1735 41322 1747
rect 41394 1923 41440 1935
rect 41394 1747 41400 1923
rect 41434 1747 41440 1923
rect 41394 1735 41440 1747
rect 41512 1923 41558 1935
rect 41642 1923 41648 2123
rect 41512 1747 41518 1923
rect 41552 1747 41648 1923
rect 41682 1747 41688 2123
rect 41512 1735 41558 1747
rect 41642 1735 41688 1747
rect 41760 2123 41806 2135
rect 41760 1747 41766 2123
rect 41800 1747 41806 2123
rect 41760 1735 41806 1747
rect 41878 2123 41924 2135
rect 41878 1747 41884 2123
rect 41918 1747 41924 2123
rect 41878 1735 41924 1747
rect 41996 2123 42042 2135
rect 41996 1747 42002 2123
rect 42036 1747 42042 2123
rect 41996 1735 42042 1747
rect 42114 2123 42160 2135
rect 42114 1747 42120 2123
rect 42154 1747 42160 2123
rect 42114 1735 42160 1747
rect 42232 2123 42278 2135
rect 42232 1747 42238 2123
rect 42272 1747 42278 2123
rect 42232 1735 42278 1747
rect 42350 2123 42396 2135
rect 42350 1747 42356 2123
rect 42390 1923 42396 2123
rect 42721 1935 42755 2238
rect 42479 1923 42525 1935
rect 42390 1747 42485 1923
rect 42519 1747 42525 1923
rect 42350 1735 42396 1747
rect 42479 1735 42525 1747
rect 42597 1923 42643 1935
rect 42597 1747 42603 1923
rect 42637 1747 42643 1923
rect 42597 1735 42643 1747
rect 42715 1923 42761 1935
rect 42715 1747 42721 1923
rect 42755 1747 42761 1923
rect 42715 1735 42761 1747
rect 42833 1923 42879 1935
rect 42833 1747 42839 1923
rect 42873 1747 42879 1923
rect 42833 1735 42879 1747
rect 38631 1686 38771 1692
rect 39266 1701 39300 1735
rect 39868 1701 39902 1735
rect 40104 1701 40138 1735
rect 38523 1657 38631 1667
rect 39266 1666 39425 1701
rect 39868 1666 40138 1701
rect 40705 1701 40739 1735
rect 40941 1701 40975 1735
rect 40705 1666 40975 1701
rect 41164 1701 41198 1735
rect 41766 1701 41800 1735
rect 42002 1701 42036 1735
rect 41164 1666 41323 1701
rect 41766 1666 42036 1701
rect 42603 1701 42637 1735
rect 42839 1701 42873 1735
rect 42603 1666 42873 1701
rect 37896 1625 37911 1627
rect 37811 1611 37911 1625
rect 37811 1568 37911 1569
rect 37432 1547 37911 1568
rect 38200 1547 38266 1643
rect 37432 1499 38266 1547
rect 37432 1470 37911 1499
rect 37432 1468 37537 1470
rect 37811 1469 37911 1470
rect 37265 1283 37275 1362
rect 37368 1283 37378 1362
rect 38263 1353 38342 1365
rect 35602 1189 36308 1193
rect 35126 1177 35172 1189
rect 33763 1038 35086 1049
rect 33763 957 33774 1038
rect 33861 1032 35086 1038
rect 33861 969 34127 1032
rect 34208 969 35086 1032
rect 33861 957 35086 969
rect 33763 951 35086 957
rect 35010 949 35086 951
rect 33766 921 34910 922
rect 33766 914 34974 921
rect 33766 832 33779 914
rect 33861 913 34974 914
rect 33861 832 34257 913
rect 34359 832 34974 913
rect 33097 778 33108 832
rect 33164 778 33174 832
rect 33766 821 34974 832
rect 30150 -1311 30350 -1305
rect 30150 -1345 30162 -1311
rect 30338 -1345 30419 -1311
rect 30150 -1351 30350 -1345
rect 30150 -1429 30350 -1423
rect 29804 -1463 30162 -1429
rect 30338 -1463 30350 -1429
rect 29804 -1795 29847 -1463
rect 30150 -1469 30350 -1463
rect 30384 -1436 30419 -1345
rect 30501 -1315 30568 -1213
rect 33097 -1230 33172 778
rect 33097 -1284 33108 -1230
rect 33164 -1284 33174 -1230
rect 33097 -1296 33172 -1284
rect 30501 -1330 30567 -1315
rect 30691 -1318 30763 -1300
rect 30688 -1383 30697 -1318
rect 30757 -1383 30767 -1318
rect 30691 -1384 30697 -1383
rect 30757 -1384 30763 -1383
rect 30691 -1396 30763 -1384
rect 30501 -1406 30567 -1396
rect 31375 -1436 31575 -1430
rect 30384 -1470 31387 -1436
rect 31563 -1470 31575 -1436
rect 30150 -1547 30350 -1541
rect 30150 -1581 30162 -1547
rect 30338 -1581 30350 -1547
rect 30150 -1587 30350 -1581
rect 30150 -1665 30350 -1659
rect 30150 -1699 30162 -1665
rect 30338 -1699 30350 -1665
rect 30150 -1705 30350 -1699
rect 30162 -1789 30338 -1705
rect 30643 -1738 31043 -1732
rect 30481 -1772 30655 -1738
rect 31031 -1772 31043 -1738
rect 31203 -1752 31246 -1470
rect 31375 -1476 31575 -1470
rect 31375 -1553 31575 -1548
rect 31375 -1554 31901 -1553
rect 31274 -1583 31336 -1577
rect 31274 -1617 31286 -1583
rect 31320 -1617 31336 -1583
rect 31375 -1588 31387 -1554
rect 31563 -1587 31901 -1554
rect 31563 -1588 31575 -1587
rect 31375 -1594 31575 -1588
rect 31274 -1633 31336 -1617
rect 29950 -1795 30350 -1789
rect 29804 -1829 29962 -1795
rect 30338 -1829 30350 -1795
rect 29804 -2031 29847 -1829
rect 29950 -1835 30350 -1829
rect 29950 -1913 30350 -1907
rect 29950 -1947 29962 -1913
rect 30338 -1947 30419 -1913
rect 29950 -1953 30350 -1947
rect 29950 -2031 30350 -2025
rect 29804 -2065 29962 -2031
rect 30338 -2065 30350 -2031
rect 29804 -2100 29847 -2065
rect 29950 -2071 30350 -2065
rect 29721 -2128 29847 -2100
rect 29699 -2138 29847 -2128
rect 29753 -2192 29847 -2138
rect 29950 -2149 30350 -2143
rect 30384 -2149 30419 -1947
rect 30481 -1974 30519 -1772
rect 30643 -1778 31043 -1772
rect 31208 -1768 31259 -1752
rect 31208 -1802 31219 -1768
rect 31253 -1802 31259 -1768
rect 31208 -1819 31259 -1802
rect 30643 -1856 31043 -1850
rect 30643 -1890 30655 -1856
rect 31031 -1890 31043 -1856
rect 30643 -1896 31043 -1890
rect 30643 -1974 31043 -1968
rect 30481 -2008 30655 -1974
rect 31031 -2008 31043 -1974
rect 30481 -2149 30519 -2008
rect 30643 -2014 31043 -2008
rect 31287 -2018 31336 -1633
rect 31375 -1856 31775 -1850
rect 31375 -1890 31387 -1856
rect 31763 -1890 31775 -1856
rect 31375 -1896 31775 -1890
rect 31375 -1974 31775 -1968
rect 31375 -2008 31387 -1974
rect 31763 -2008 31775 -1974
rect 31375 -2014 31775 -2008
rect 31287 -2034 31344 -2018
rect 31287 -2068 31303 -2034
rect 31337 -2068 31344 -2034
rect 31287 -2084 31344 -2068
rect 31869 -2046 31901 -1587
rect 31869 -2080 31986 -2046
rect 30643 -2092 31043 -2086
rect 30643 -2126 30655 -2092
rect 31031 -2126 31043 -2092
rect 30643 -2132 31043 -2126
rect 31375 -2092 31775 -2086
rect 31375 -2126 31387 -2092
rect 31763 -2126 31775 -2092
rect 31375 -2132 31775 -2126
rect 29950 -2183 29962 -2149
rect 30338 -2183 30519 -2149
rect 29950 -2189 30350 -2183
rect 29699 -2202 29847 -2192
rect 29721 -2234 29847 -2202
rect 29804 -2267 29847 -2234
rect 30481 -2210 30519 -2183
rect 31287 -2152 31346 -2136
rect 31287 -2186 31302 -2152
rect 31336 -2186 31346 -2152
rect 31287 -2203 31346 -2186
rect 31869 -2142 31923 -2080
rect 31981 -2142 31986 -2080
rect 31869 -2178 31986 -2142
rect 34530 -2059 34648 821
rect 34896 672 34950 821
rect 35010 757 35064 949
rect 35126 801 35132 1177
rect 35166 801 35172 1177
rect 35126 789 35172 801
rect 35244 1177 35290 1189
rect 35244 801 35250 1177
rect 35284 801 35290 1177
rect 35244 789 35290 801
rect 35362 1177 35408 1189
rect 35362 801 35368 1177
rect 35402 828 35408 1177
rect 35479 1177 35525 1189
rect 35479 1001 35485 1177
rect 35519 1001 35525 1177
rect 35479 994 35525 1001
rect 35597 1177 36308 1189
rect 35597 1001 35603 1177
rect 35637 1164 36308 1177
rect 35637 1001 35643 1164
rect 35887 1085 36308 1164
rect 35887 1084 35991 1085
rect 35479 989 35528 994
rect 35597 989 35643 1001
rect 35485 828 35528 989
rect 35402 801 35528 828
rect 35362 789 35528 801
rect 35368 785 35528 789
rect 35010 751 35241 757
rect 35010 717 35191 751
rect 35225 717 35241 751
rect 35010 701 35241 717
rect 35293 751 35359 757
rect 35293 717 35309 751
rect 35343 717 35359 751
rect 35293 672 35359 717
rect 34896 664 35359 672
rect 34896 632 35360 664
rect 35452 648 35528 785
rect 35448 588 35458 648
rect 35520 588 35530 648
rect 37276 109 37369 1283
rect 38263 1254 38269 1353
rect 38194 1234 38269 1254
rect 38336 1254 38342 1353
rect 38336 1234 38414 1254
rect 38194 1126 38238 1234
rect 38370 1126 38414 1234
rect 38194 1084 38414 1126
rect 37798 1054 38775 1084
rect 37798 948 37830 1054
rect 38034 948 38066 1054
rect 38270 948 38302 1054
rect 38506 948 38538 1054
rect 38741 948 38775 1054
rect 37791 936 37837 948
rect 37791 760 37797 936
rect 37831 760 37837 936
rect 37791 748 37837 760
rect 37909 936 37955 948
rect 37909 760 37915 936
rect 37949 760 37955 936
rect 37909 748 37955 760
rect 38027 936 38073 948
rect 38027 760 38033 936
rect 38067 760 38073 936
rect 38027 748 38073 760
rect 38145 936 38191 948
rect 38145 760 38151 936
rect 38185 760 38191 936
rect 38145 748 38191 760
rect 38263 936 38309 948
rect 38263 760 38269 936
rect 38303 760 38309 936
rect 38263 748 38309 760
rect 38381 936 38427 948
rect 38381 760 38387 936
rect 38421 760 38427 936
rect 38381 748 38427 760
rect 38499 936 38545 948
rect 38499 760 38505 936
rect 38539 760 38545 936
rect 38499 748 38545 760
rect 38617 936 38663 948
rect 38617 760 38623 936
rect 38657 760 38663 936
rect 38617 748 38663 760
rect 38735 936 38781 948
rect 38735 760 38741 936
rect 38775 760 38781 936
rect 38735 748 38781 760
rect 38853 936 38899 948
rect 38853 760 38859 936
rect 38893 760 38899 936
rect 38853 748 38899 760
rect 39391 882 39425 1666
rect 40104 1604 40138 1666
rect 39693 1566 40435 1604
rect 39693 1442 39727 1566
rect 39929 1442 39963 1566
rect 40165 1442 40199 1566
rect 40401 1442 40435 1566
rect 40691 1459 40701 1525
rect 40764 1459 40774 1525
rect 39687 1430 39733 1442
rect 39687 1054 39693 1430
rect 39727 1054 39733 1430
rect 39687 1042 39733 1054
rect 39805 1430 39851 1442
rect 39805 1054 39811 1430
rect 39845 1054 39851 1430
rect 39805 1042 39851 1054
rect 39923 1430 39969 1442
rect 39923 1054 39929 1430
rect 39963 1054 39969 1430
rect 39923 1042 39969 1054
rect 40041 1430 40087 1442
rect 40041 1054 40047 1430
rect 40081 1054 40087 1430
rect 40041 1042 40087 1054
rect 40159 1430 40205 1442
rect 40159 1054 40165 1430
rect 40199 1054 40205 1430
rect 40159 1042 40205 1054
rect 40277 1430 40323 1442
rect 40277 1054 40283 1430
rect 40317 1054 40323 1430
rect 40277 1042 40323 1054
rect 40395 1430 40441 1442
rect 40395 1054 40401 1430
rect 40435 1054 40441 1430
rect 40395 1042 40441 1054
rect 40807 883 40841 1666
rect 40534 882 40841 883
rect 39391 877 39707 882
rect 40421 877 40841 882
rect 39391 866 39774 877
rect 39391 839 39723 866
rect 37914 654 37950 748
rect 38150 654 38186 748
rect 38386 655 38422 748
rect 38548 700 38614 707
rect 38548 666 38564 700
rect 38598 666 38614 700
rect 38548 655 38614 666
rect 38386 654 38614 655
rect 37914 625 38614 654
rect 37914 624 38496 625
rect 38034 511 38068 624
rect 38430 583 38496 624
rect 38430 549 38446 583
rect 38480 549 38496 583
rect 38430 542 38496 549
rect 38858 515 38893 748
rect 39391 710 39425 839
rect 39707 832 39723 839
rect 39757 832 39774 866
rect 39707 826 39774 832
rect 40354 866 40841 877
rect 40354 832 40371 866
rect 40405 839 40841 866
rect 40405 832 40421 839
rect 40534 838 40841 839
rect 40354 826 40421 832
rect 39532 799 39588 811
rect 39532 765 39538 799
rect 39572 798 39588 799
rect 40645 798 40701 810
rect 39572 782 40039 798
rect 39572 765 39989 782
rect 39532 749 39989 765
rect 39973 748 39989 749
rect 40023 748 40039 782
rect 39973 741 40039 748
rect 40091 783 40661 798
rect 40091 749 40107 783
rect 40141 764 40661 783
rect 40695 764 40701 798
rect 40141 749 40701 764
rect 40091 739 40158 749
rect 40645 748 40701 749
rect 40807 710 40841 838
rect 41289 882 41323 1666
rect 42002 1604 42036 1666
rect 41591 1566 42333 1604
rect 41591 1442 41625 1566
rect 41827 1442 41861 1566
rect 42063 1442 42097 1566
rect 42299 1442 42333 1566
rect 41585 1430 41631 1442
rect 41585 1054 41591 1430
rect 41625 1054 41631 1430
rect 41585 1042 41631 1054
rect 41703 1430 41749 1442
rect 41703 1054 41709 1430
rect 41743 1054 41749 1430
rect 41703 1042 41749 1054
rect 41821 1430 41867 1442
rect 41821 1054 41827 1430
rect 41861 1054 41867 1430
rect 41821 1042 41867 1054
rect 41939 1430 41985 1442
rect 41939 1054 41945 1430
rect 41979 1054 41985 1430
rect 41939 1042 41985 1054
rect 42057 1430 42103 1442
rect 42057 1054 42063 1430
rect 42097 1054 42103 1430
rect 42057 1042 42103 1054
rect 42175 1430 42221 1442
rect 42175 1054 42181 1430
rect 42215 1054 42221 1430
rect 42175 1042 42221 1054
rect 42293 1430 42339 1442
rect 42293 1054 42299 1430
rect 42333 1054 42339 1430
rect 42293 1042 42339 1054
rect 42705 883 42739 1666
rect 42317 882 42386 883
rect 42432 882 42739 883
rect 41289 877 41605 882
rect 42317 878 42739 882
rect 41289 866 41672 877
rect 41289 839 41621 866
rect 41289 710 41323 839
rect 41605 832 41621 839
rect 41655 832 41672 866
rect 41605 826 41672 832
rect 42250 867 42739 878
rect 42250 833 42267 867
rect 42301 839 42739 867
rect 42301 833 42317 839
rect 42432 838 42739 839
rect 42250 827 42317 833
rect 41430 799 41486 811
rect 41430 765 41436 799
rect 41470 798 41486 799
rect 42543 798 42599 810
rect 41470 782 41937 798
rect 41470 765 41887 782
rect 41430 749 41887 765
rect 41871 748 41887 749
rect 41921 748 41937 782
rect 41871 741 41937 748
rect 41989 783 42559 798
rect 41989 749 42005 783
rect 42039 764 42559 783
rect 42593 764 42599 798
rect 42039 749 42599 764
rect 41989 739 42056 749
rect 42543 748 42599 749
rect 42705 710 42739 838
rect 42820 1488 42887 1512
rect 42820 1454 42837 1488
rect 42871 1454 42887 1488
rect 38504 511 38893 515
rect 38028 499 38074 511
rect 38028 123 38034 499
rect 38068 123 38074 499
rect 38028 111 38074 123
rect 38146 499 38192 511
rect 38146 123 38152 499
rect 38186 123 38192 499
rect 38146 111 38192 123
rect 38264 499 38310 511
rect 38264 123 38270 499
rect 38304 147 38310 499
rect 38381 499 38427 511
rect 38381 323 38387 499
rect 38421 323 38427 499
rect 38381 311 38427 323
rect 38499 499 38893 511
rect 39385 698 39431 710
rect 39385 522 39391 698
rect 39425 522 39431 698
rect 39385 510 39431 522
rect 39503 698 39549 710
rect 39503 522 39509 698
rect 39543 522 39549 698
rect 39503 510 39549 522
rect 39805 698 39851 710
rect 38499 323 38505 499
rect 38539 486 38893 499
rect 38539 323 38545 486
rect 38815 483 38893 486
rect 38815 431 38825 483
rect 38888 431 38898 483
rect 38820 425 38893 431
rect 38499 311 38545 323
rect 38387 195 38422 311
rect 39508 216 39542 510
rect 39805 322 39811 698
rect 39845 322 39851 698
rect 39805 310 39851 322
rect 39923 698 39969 710
rect 39923 322 39929 698
rect 39963 322 39969 698
rect 39923 310 39969 322
rect 40041 698 40087 710
rect 40041 322 40047 698
rect 40081 322 40087 698
rect 40041 310 40087 322
rect 40159 698 40205 710
rect 40159 322 40165 698
rect 40199 322 40205 698
rect 40159 310 40205 322
rect 40277 698 40323 710
rect 40277 322 40283 698
rect 40317 322 40323 698
rect 40683 698 40729 710
rect 40683 522 40689 698
rect 40723 522 40729 698
rect 40683 510 40729 522
rect 40801 698 40847 710
rect 40801 522 40807 698
rect 40841 522 40847 698
rect 40801 510 40847 522
rect 41283 698 41329 710
rect 41283 522 41289 698
rect 41323 522 41329 698
rect 41283 510 41329 522
rect 41401 698 41447 710
rect 41401 522 41407 698
rect 41441 522 41447 698
rect 41401 510 41447 522
rect 41703 698 41749 710
rect 40277 310 40323 322
rect 40165 216 40199 310
rect 40689 216 40722 510
rect 38518 195 38626 205
rect 38387 147 38518 195
rect 39508 184 40722 216
rect 41406 216 41440 510
rect 41703 322 41709 698
rect 41743 322 41749 698
rect 41703 310 41749 322
rect 41821 698 41867 710
rect 41821 322 41827 698
rect 41861 322 41867 698
rect 41821 310 41867 322
rect 41939 698 41985 710
rect 41939 322 41945 698
rect 41979 322 41985 698
rect 41939 310 41985 322
rect 42057 698 42103 710
rect 42057 322 42063 698
rect 42097 322 42103 698
rect 42057 310 42103 322
rect 42175 698 42221 710
rect 42175 322 42181 698
rect 42215 322 42221 698
rect 42581 698 42627 710
rect 42581 522 42587 698
rect 42621 522 42627 698
rect 42581 510 42627 522
rect 42699 698 42745 710
rect 42699 522 42705 698
rect 42739 522 42745 698
rect 42699 510 42745 522
rect 42175 310 42221 322
rect 42063 216 42097 310
rect 42587 216 42620 510
rect 41406 184 42620 216
rect 38626 167 38771 173
rect 38304 123 38518 147
rect 38264 111 38518 123
rect 37276 107 37861 109
rect 38270 107 38518 111
rect 37276 79 37906 107
rect 37276 73 38143 79
rect 37276 39 38093 73
rect 38127 39 38143 73
rect 37276 23 38143 39
rect 38195 73 38261 79
rect 38195 39 38211 73
rect 38245 39 38261 73
rect 38444 63 38518 107
rect 38759 100 38771 167
rect 38626 94 38771 100
rect 40001 99 40133 184
rect 41899 99 42031 184
rect 38518 53 38626 63
rect 37276 7 37906 23
rect 37276 3 37861 7
rect 37276 2 37377 3
rect 37806 -46 37906 -35
rect 37770 -152 37780 -46
rect 37892 -57 37906 -46
rect 38195 -57 38261 39
rect 39991 -9 40001 99
rect 40133 -9 40143 99
rect 41889 -9 41899 99
rect 42031 -9 42041 99
rect 42820 71 42887 1454
rect 42948 1025 43106 3252
rect 42948 927 42960 1025
rect 43092 950 43106 1025
rect 43190 2843 43704 2867
rect 43190 2737 43552 2843
rect 43664 2830 43704 2843
rect 43664 2737 43706 2830
rect 43190 2726 43706 2737
rect 43190 2725 43704 2726
rect 43092 927 43104 950
rect 42948 921 43104 927
rect 37892 -105 38261 -57
rect 37892 -135 37906 -105
rect 37892 -152 37902 -135
rect 38194 -208 38260 -105
rect 40025 -150 40031 -9
rect 40098 -150 40104 -9
rect 40025 -162 40104 -150
rect 42820 -208 42886 71
rect 38192 -288 42886 -208
rect 41606 -793 42070 -761
rect 42158 -777 42168 -717
rect 42230 -777 42240 -717
rect 41606 -801 42069 -793
rect 41606 -950 41660 -801
rect 41221 -956 41660 -950
rect 41219 -1042 41229 -956
rect 41305 -1042 41660 -956
rect 41221 -1050 41660 -1042
rect 41720 -846 41951 -830
rect 41720 -880 41901 -846
rect 41935 -880 41951 -846
rect 41720 -886 41951 -880
rect 42003 -846 42069 -801
rect 42003 -880 42019 -846
rect 42053 -880 42069 -846
rect 42003 -886 42069 -880
rect 41720 -1078 41774 -886
rect 42162 -914 42238 -777
rect 42078 -918 42238 -914
rect 41456 -1083 41774 -1078
rect 41450 -1174 41460 -1083
rect 41589 -1174 41774 -1083
rect 41456 -1178 41774 -1174
rect 41836 -930 41882 -918
rect 41836 -1306 41842 -930
rect 41876 -1306 41882 -930
rect 41836 -1318 41882 -1306
rect 41954 -930 42000 -918
rect 41954 -1306 41960 -930
rect 41994 -1306 42000 -930
rect 41954 -1318 42000 -1306
rect 42072 -930 42238 -918
rect 42072 -1306 42078 -930
rect 42112 -957 42238 -930
rect 42112 -1306 42118 -957
rect 42195 -1118 42238 -957
rect 42072 -1318 42118 -1306
rect 42189 -1123 42238 -1118
rect 42189 -1130 42235 -1123
rect 42189 -1306 42195 -1130
rect 42229 -1306 42235 -1130
rect 42189 -1318 42235 -1306
rect 42307 -1130 42353 -1118
rect 42307 -1306 42313 -1130
rect 42347 -1293 42353 -1130
rect 43190 -1213 43326 2725
rect 43827 1360 43920 3252
rect 43983 3195 44449 3217
rect 44737 3195 44803 3291
rect 46568 3301 46574 3477
rect 46608 3301 46614 3477
rect 46568 3289 46614 3301
rect 46686 3477 46732 3489
rect 46686 3301 46692 3477
rect 46726 3301 46732 3477
rect 46686 3289 46732 3301
rect 46804 3477 46850 3489
rect 46804 3301 46810 3477
rect 46844 3301 46850 3477
rect 46804 3289 46850 3301
rect 46922 3477 46968 3489
rect 46922 3301 46928 3477
rect 46962 3422 46968 3477
rect 47087 3477 47133 3489
rect 47087 3422 47093 3477
rect 46962 3334 47093 3422
rect 46962 3301 46968 3334
rect 46922 3289 46968 3301
rect 47087 3301 47093 3334
rect 47127 3301 47133 3477
rect 47087 3289 47133 3301
rect 47205 3477 47251 3489
rect 47205 3301 47211 3477
rect 47245 3301 47251 3477
rect 47205 3289 47251 3301
rect 47323 3477 47369 3489
rect 47323 3301 47329 3477
rect 47363 3301 47369 3477
rect 47323 3289 47369 3301
rect 47441 3477 47487 3489
rect 47441 3301 47447 3477
rect 47481 3301 47487 3477
rect 47441 3289 47487 3301
rect 46574 3250 46608 3289
rect 46810 3250 46844 3289
rect 46574 3215 46844 3250
rect 47211 3251 47244 3289
rect 47447 3251 47480 3289
rect 47211 3215 47480 3251
rect 43983 3147 44803 3195
rect 46608 3214 46844 3215
rect 43983 3116 44449 3147
rect 46608 3140 46740 3214
rect 43983 2860 44088 3116
rect 46598 3032 46608 3140
rect 46740 3032 46750 3140
rect 44819 2959 44898 2971
rect 43983 2754 44046 2860
rect 44158 2754 44168 2860
rect 44819 2856 44825 2959
rect 44750 2836 44825 2856
rect 44892 2856 44898 2959
rect 46631 2896 46637 3032
rect 46704 2896 46710 3032
rect 46631 2884 46710 2896
rect 44892 2836 44970 2856
rect 43983 2743 44132 2754
rect 43983 1566 44088 2743
rect 44750 2728 44794 2836
rect 44926 2728 44970 2836
rect 44750 2686 44970 2728
rect 47548 2701 47610 4272
rect 47800 4264 47846 4276
rect 47800 3888 47806 4264
rect 47840 3888 47846 4264
rect 47800 3876 47846 3888
rect 47918 4264 47964 4276
rect 47918 3888 47924 4264
rect 47958 3888 47964 4264
rect 47918 3876 47964 3888
rect 48036 4264 48082 4276
rect 48036 3888 48042 4264
rect 48076 3888 48082 4264
rect 48036 3876 48082 3888
rect 48154 4264 48200 4276
rect 48154 3888 48160 4264
rect 48194 3888 48200 4264
rect 48154 3876 48200 3888
rect 48272 4264 48318 4276
rect 48272 3888 48278 4264
rect 48312 3888 48318 4264
rect 48272 3876 48318 3888
rect 48390 4264 48436 4276
rect 48390 3888 48396 4264
rect 48430 3888 48436 4264
rect 48390 3876 48436 3888
rect 48508 4264 48554 4276
rect 48508 3888 48514 4264
rect 48548 3888 48554 4264
rect 48508 3876 48554 3888
rect 47806 3834 47840 3876
rect 48042 3834 48076 3876
rect 47806 3806 48076 3834
rect 48160 3835 48194 3876
rect 48396 3835 48430 3876
rect 48160 3806 48430 3835
rect 47806 3758 47840 3806
rect 47806 3728 47869 3758
rect 47834 3636 47869 3728
rect 48341 3698 48441 3719
rect 48341 3644 48355 3698
rect 48420 3644 48441 3698
rect 48341 3639 48441 3644
rect 48514 3693 48548 3876
rect 48514 3639 48623 3693
rect 47834 3600 48061 3636
rect 47834 3493 47869 3600
rect 47995 3566 48061 3600
rect 47995 3532 48011 3566
rect 48045 3532 48061 3566
rect 48342 3624 48439 3639
rect 48342 3557 48399 3624
rect 47995 3526 48061 3532
rect 48236 3521 48505 3557
rect 48236 3493 48269 3521
rect 48472 3493 48505 3521
rect 48589 3493 48623 3639
rect 47710 3481 47756 3493
rect 47710 3305 47716 3481
rect 47750 3305 47756 3481
rect 47710 3293 47756 3305
rect 47828 3481 47874 3493
rect 47828 3305 47834 3481
rect 47868 3305 47874 3481
rect 47828 3293 47874 3305
rect 47946 3481 47992 3493
rect 47946 3305 47952 3481
rect 47986 3305 47992 3481
rect 47946 3293 47992 3305
rect 48064 3481 48110 3493
rect 48064 3305 48070 3481
rect 48104 3426 48110 3481
rect 48229 3481 48275 3493
rect 48229 3426 48235 3481
rect 48104 3338 48235 3426
rect 48104 3305 48110 3338
rect 48064 3293 48110 3305
rect 48229 3305 48235 3338
rect 48269 3305 48275 3481
rect 48229 3293 48275 3305
rect 48347 3481 48393 3493
rect 48347 3305 48353 3481
rect 48387 3305 48393 3481
rect 48347 3293 48393 3305
rect 48465 3481 48511 3493
rect 48465 3305 48471 3481
rect 48505 3305 48511 3481
rect 48465 3293 48511 3305
rect 48583 3481 48629 3493
rect 48583 3305 48589 3481
rect 48623 3305 48629 3481
rect 48583 3293 48629 3305
rect 49778 3360 49918 9501
rect 50347 9209 50529 10697
rect 53948 10459 54027 10471
rect 51467 10403 51546 10415
rect 51467 10308 51473 10403
rect 51396 10288 51473 10308
rect 51540 10308 51546 10403
rect 53948 10342 53954 10459
rect 54021 10342 54027 10459
rect 55095 10458 55174 10470
rect 55095 10342 55101 10458
rect 55168 10342 55174 10458
rect 51540 10288 51616 10308
rect 51396 10180 51440 10288
rect 51572 10180 51616 10288
rect 53193 10246 53249 10254
rect 51396 10138 51616 10180
rect 52267 10238 53249 10246
rect 52267 10204 53209 10238
rect 53243 10204 53249 10238
rect 53912 10234 53922 10342
rect 54054 10279 54064 10342
rect 54054 10268 54066 10279
rect 54054 10234 54067 10268
rect 54323 10258 54379 10260
rect 52267 10188 53249 10204
rect 53922 10196 54067 10234
rect 52267 10187 53246 10188
rect 51000 10108 51977 10138
rect 51000 10002 51032 10108
rect 51236 10002 51268 10108
rect 51472 10002 51504 10108
rect 51708 10002 51740 10108
rect 51943 10002 51977 10108
rect 50993 9990 51039 10002
rect 50993 9814 50999 9990
rect 51033 9814 51039 9990
rect 50993 9802 51039 9814
rect 51111 9990 51157 10002
rect 51111 9814 51117 9990
rect 51151 9814 51157 9990
rect 51111 9802 51157 9814
rect 51229 9990 51275 10002
rect 51229 9814 51235 9990
rect 51269 9814 51275 9990
rect 51229 9802 51275 9814
rect 51347 9990 51393 10002
rect 51347 9814 51353 9990
rect 51387 9814 51393 9990
rect 51347 9802 51393 9814
rect 51465 9990 51511 10002
rect 51465 9814 51471 9990
rect 51505 9814 51511 9990
rect 51465 9802 51511 9814
rect 51583 9990 51629 10002
rect 51583 9814 51589 9990
rect 51623 9814 51629 9990
rect 51583 9802 51629 9814
rect 51701 9990 51747 10002
rect 51701 9814 51707 9990
rect 51741 9814 51747 9990
rect 51701 9802 51747 9814
rect 51819 9990 51865 10002
rect 51819 9814 51825 9990
rect 51859 9814 51865 9990
rect 51819 9802 51865 9814
rect 51937 9990 51983 10002
rect 51937 9814 51943 9990
rect 51977 9814 51983 9990
rect 51937 9802 51983 9814
rect 52055 9990 52101 10002
rect 52055 9814 52061 9990
rect 52095 9814 52101 9990
rect 52055 9802 52101 9814
rect 51116 9708 51152 9802
rect 51352 9708 51388 9802
rect 51588 9709 51624 9802
rect 51750 9754 51816 9761
rect 51750 9720 51766 9754
rect 51800 9720 51816 9754
rect 51750 9709 51816 9720
rect 51588 9708 51816 9709
rect 51116 9679 51816 9708
rect 51116 9678 51698 9679
rect 51236 9565 51270 9678
rect 51632 9637 51698 9678
rect 51632 9603 51648 9637
rect 51682 9603 51698 9637
rect 51632 9596 51698 9603
rect 52060 9597 52095 9802
rect 52267 9597 52334 10187
rect 54026 10164 54067 10196
rect 54313 10192 54323 10258
rect 54379 10192 54389 10258
rect 55059 10234 55069 10342
rect 55201 10279 55211 10342
rect 55201 10268 55213 10279
rect 55201 10234 55214 10268
rect 55069 10196 55214 10234
rect 55173 10168 55214 10196
rect 53442 10136 53712 10164
rect 53183 10070 53193 10136
rect 53259 10070 53269 10136
rect 53442 10074 53476 10136
rect 53678 10074 53712 10136
rect 53796 10136 54067 10164
rect 54584 10140 54854 10168
rect 53796 10074 53830 10136
rect 54032 10074 54067 10136
rect 54208 10124 54379 10140
rect 54208 10090 54339 10124
rect 54373 10090 54379 10124
rect 54208 10074 54379 10090
rect 54584 10078 54618 10140
rect 54820 10078 54854 10140
rect 54938 10140 55214 10168
rect 54938 10078 54972 10140
rect 55174 10078 55214 10140
rect 53318 10062 53364 10074
rect 53318 9686 53324 10062
rect 53358 9686 53364 10062
rect 53318 9674 53364 9686
rect 53436 10062 53482 10074
rect 53436 9686 53442 10062
rect 53476 9686 53482 10062
rect 53436 9674 53482 9686
rect 53554 10062 53600 10074
rect 53554 9686 53560 10062
rect 53594 9686 53600 10062
rect 53554 9674 53600 9686
rect 53672 10062 53718 10074
rect 53672 9686 53678 10062
rect 53712 9686 53718 10062
rect 53672 9674 53718 9686
rect 53790 10062 53836 10074
rect 53790 9686 53796 10062
rect 53830 9686 53836 10062
rect 53790 9674 53836 9686
rect 53908 10062 53954 10074
rect 53908 9686 53914 10062
rect 53948 9686 53954 10062
rect 53908 9674 53954 9686
rect 54026 10062 54072 10074
rect 54026 9686 54032 10062
rect 54066 9686 54072 10062
rect 54026 9674 54072 9686
rect 52060 9569 52334 9597
rect 51706 9565 52334 9569
rect 50346 9160 50529 9209
rect 51230 9553 51276 9565
rect 51230 9177 51236 9553
rect 51270 9177 51276 9553
rect 51230 9165 51276 9177
rect 51348 9553 51394 9565
rect 51348 9177 51354 9553
rect 51388 9177 51394 9553
rect 51348 9165 51394 9177
rect 51466 9553 51512 9565
rect 51466 9177 51472 9553
rect 51506 9201 51512 9553
rect 51583 9553 51629 9565
rect 51583 9377 51589 9553
rect 51623 9377 51629 9553
rect 51583 9365 51629 9377
rect 51701 9553 52334 9565
rect 51701 9377 51707 9553
rect 51741 9540 52334 9553
rect 53324 9632 53358 9674
rect 53560 9632 53594 9674
rect 53324 9604 53594 9632
rect 53678 9633 53712 9674
rect 53914 9633 53948 9674
rect 53678 9604 53948 9633
rect 53324 9556 53358 9604
rect 51741 9377 51747 9540
rect 53324 9526 53387 9556
rect 51701 9365 51747 9377
rect 53352 9434 53387 9526
rect 53352 9398 53579 9434
rect 53849 9423 53859 9520
rect 53958 9423 53968 9520
rect 54032 9491 54066 9674
rect 54032 9437 54141 9491
rect 51589 9249 51624 9365
rect 53352 9291 53387 9398
rect 53513 9364 53579 9398
rect 53513 9330 53529 9364
rect 53563 9330 53579 9364
rect 53860 9422 53957 9423
rect 53860 9355 53917 9422
rect 53513 9324 53579 9330
rect 53754 9319 54023 9355
rect 53754 9291 53787 9319
rect 53990 9291 54023 9319
rect 54107 9291 54141 9437
rect 53228 9279 53274 9291
rect 51720 9249 51828 9259
rect 51589 9201 51720 9249
rect 51828 9212 51969 9218
rect 51506 9177 51720 9201
rect 51466 9165 51720 9177
rect 51472 9161 51720 9165
rect 50346 9133 51108 9160
rect 50346 9127 51345 9133
rect 50346 9093 51295 9127
rect 51329 9093 51345 9127
rect 50346 9077 51345 9093
rect 51397 9127 51463 9133
rect 51397 9093 51413 9127
rect 51447 9093 51463 9127
rect 51646 9117 51720 9161
rect 51957 9145 51969 9212
rect 51828 9139 51969 9145
rect 51720 9107 51828 9117
rect 50346 9061 51108 9077
rect 50346 9060 51045 9061
rect 50346 9056 50580 9060
rect 50198 7543 50363 7563
rect 50198 7426 50210 7543
rect 50349 7520 50363 7543
rect 50349 7426 50364 7520
rect 50198 7425 50217 7426
rect 50329 7425 50364 7426
rect 50198 7416 50364 7425
rect 50198 7415 50363 7416
rect 50198 7414 50331 7415
rect 50487 7162 50580 9056
rect 50643 8997 51109 9019
rect 51397 8997 51463 9093
rect 53228 9103 53234 9279
rect 53268 9103 53274 9279
rect 53228 9091 53274 9103
rect 53346 9279 53392 9291
rect 53346 9103 53352 9279
rect 53386 9103 53392 9279
rect 53346 9091 53392 9103
rect 53464 9279 53510 9291
rect 53464 9103 53470 9279
rect 53504 9103 53510 9279
rect 53464 9091 53510 9103
rect 53582 9279 53628 9291
rect 53582 9103 53588 9279
rect 53622 9224 53628 9279
rect 53747 9279 53793 9291
rect 53747 9224 53753 9279
rect 53622 9136 53753 9224
rect 53622 9103 53628 9136
rect 53582 9091 53628 9103
rect 53747 9103 53753 9136
rect 53787 9103 53793 9279
rect 53747 9091 53793 9103
rect 53865 9279 53911 9291
rect 53865 9103 53871 9279
rect 53905 9103 53911 9279
rect 53865 9091 53911 9103
rect 53983 9279 54029 9291
rect 53983 9103 53989 9279
rect 54023 9103 54029 9279
rect 53983 9091 54029 9103
rect 54101 9279 54147 9291
rect 54101 9103 54107 9279
rect 54141 9103 54147 9279
rect 54101 9091 54147 9103
rect 53234 9052 53268 9091
rect 53470 9052 53504 9091
rect 53234 9017 53504 9052
rect 53871 9053 53904 9091
rect 54107 9053 54140 9091
rect 53871 9017 54140 9053
rect 50643 8949 51463 8997
rect 53268 9016 53504 9017
rect 50643 8918 51109 8949
rect 53268 8942 53400 9016
rect 50643 8662 50748 8918
rect 53258 8834 53268 8942
rect 53400 8834 53410 8942
rect 51482 8755 51561 8767
rect 50643 8556 50706 8662
rect 50818 8556 50828 8662
rect 51482 8658 51488 8755
rect 51410 8638 51488 8658
rect 51555 8658 51561 8755
rect 53290 8700 53296 8834
rect 53363 8700 53369 8834
rect 53290 8688 53369 8700
rect 51555 8638 51630 8658
rect 50643 8545 50792 8556
rect 50643 7368 50748 8545
rect 51410 8530 51454 8638
rect 51586 8530 51630 8638
rect 51410 8488 51630 8530
rect 54208 8503 54270 10074
rect 54460 10066 54506 10078
rect 54460 9690 54466 10066
rect 54500 9690 54506 10066
rect 54460 9678 54506 9690
rect 54578 10066 54624 10078
rect 54578 9690 54584 10066
rect 54618 9690 54624 10066
rect 54578 9678 54624 9690
rect 54696 10066 54742 10078
rect 54696 9690 54702 10066
rect 54736 9690 54742 10066
rect 54696 9678 54742 9690
rect 54814 10066 54860 10078
rect 54814 9690 54820 10066
rect 54854 9690 54860 10066
rect 54814 9678 54860 9690
rect 54932 10066 54978 10078
rect 54932 9690 54938 10066
rect 54972 9690 54978 10066
rect 54932 9678 54978 9690
rect 55050 10066 55096 10078
rect 55050 9690 55056 10066
rect 55090 9690 55096 10066
rect 55050 9678 55096 9690
rect 55168 10066 55214 10078
rect 55168 9690 55174 10066
rect 55208 9690 55214 10066
rect 55168 9678 55214 9690
rect 54466 9636 54500 9678
rect 54702 9636 54736 9678
rect 54466 9608 54736 9636
rect 54820 9637 54854 9678
rect 55056 9637 55090 9678
rect 54820 9608 55090 9637
rect 54466 9560 54500 9608
rect 54466 9530 54529 9560
rect 54494 9438 54529 9530
rect 55001 9500 55101 9521
rect 55001 9446 55015 9500
rect 55080 9446 55101 9500
rect 55001 9441 55101 9446
rect 55174 9495 55208 9678
rect 55174 9441 55283 9495
rect 54494 9402 54721 9438
rect 54494 9295 54529 9402
rect 54655 9368 54721 9402
rect 54655 9334 54671 9368
rect 54705 9334 54721 9368
rect 55002 9426 55099 9441
rect 55002 9359 55059 9426
rect 54655 9328 54721 9334
rect 54896 9323 55165 9359
rect 54896 9295 54929 9323
rect 55132 9295 55165 9323
rect 55249 9295 55283 9441
rect 54370 9283 54416 9295
rect 54370 9107 54376 9283
rect 54410 9107 54416 9283
rect 54370 9095 54416 9107
rect 54488 9283 54534 9295
rect 54488 9107 54494 9283
rect 54528 9107 54534 9283
rect 54488 9095 54534 9107
rect 54606 9283 54652 9295
rect 54606 9107 54612 9283
rect 54646 9107 54652 9283
rect 54606 9095 54652 9107
rect 54724 9283 54770 9295
rect 54724 9107 54730 9283
rect 54764 9228 54770 9283
rect 54889 9283 54935 9295
rect 54889 9228 54895 9283
rect 54764 9140 54895 9228
rect 54764 9107 54770 9140
rect 54724 9095 54770 9107
rect 54889 9107 54895 9140
rect 54929 9107 54935 9283
rect 54889 9095 54935 9107
rect 55007 9283 55053 9295
rect 55007 9107 55013 9283
rect 55047 9107 55053 9283
rect 55007 9095 55053 9107
rect 55125 9283 55171 9295
rect 55125 9107 55131 9283
rect 55165 9107 55171 9283
rect 55125 9095 55171 9107
rect 55243 9283 55289 9295
rect 55243 9107 55249 9283
rect 55283 9107 55289 9283
rect 56973 9228 57155 10765
rect 60571 10524 60650 10536
rect 58087 10472 58166 10484
rect 58087 10376 58093 10472
rect 58021 10356 58093 10376
rect 58160 10376 58166 10472
rect 60571 10410 60577 10524
rect 60644 10410 60650 10524
rect 61720 10530 61799 10542
rect 61720 10410 61726 10530
rect 61793 10410 61799 10530
rect 58160 10356 58241 10376
rect 58021 10248 58065 10356
rect 58197 10248 58241 10356
rect 59818 10314 59874 10322
rect 58021 10206 58241 10248
rect 58892 10306 59874 10314
rect 58892 10272 59834 10306
rect 59868 10272 59874 10306
rect 60537 10302 60547 10410
rect 60679 10347 60689 10410
rect 60679 10336 60691 10347
rect 60679 10302 60692 10336
rect 60948 10326 61004 10328
rect 58892 10256 59874 10272
rect 60547 10264 60692 10302
rect 58892 10255 59871 10256
rect 57625 10176 58602 10206
rect 57625 10070 57657 10176
rect 57861 10070 57893 10176
rect 58097 10070 58129 10176
rect 58333 10070 58365 10176
rect 58568 10070 58602 10176
rect 57618 10058 57664 10070
rect 57618 9882 57624 10058
rect 57658 9882 57664 10058
rect 57618 9870 57664 9882
rect 57736 10058 57782 10070
rect 57736 9882 57742 10058
rect 57776 9882 57782 10058
rect 57736 9870 57782 9882
rect 57854 10058 57900 10070
rect 57854 9882 57860 10058
rect 57894 9882 57900 10058
rect 57854 9870 57900 9882
rect 57972 10058 58018 10070
rect 57972 9882 57978 10058
rect 58012 9882 58018 10058
rect 57972 9870 58018 9882
rect 58090 10058 58136 10070
rect 58090 9882 58096 10058
rect 58130 9882 58136 10058
rect 58090 9870 58136 9882
rect 58208 10058 58254 10070
rect 58208 9882 58214 10058
rect 58248 9882 58254 10058
rect 58208 9870 58254 9882
rect 58326 10058 58372 10070
rect 58326 9882 58332 10058
rect 58366 9882 58372 10058
rect 58326 9870 58372 9882
rect 58444 10058 58490 10070
rect 58444 9882 58450 10058
rect 58484 9882 58490 10058
rect 58444 9870 58490 9882
rect 58562 10058 58608 10070
rect 58562 9882 58568 10058
rect 58602 9882 58608 10058
rect 58562 9870 58608 9882
rect 58680 10058 58726 10070
rect 58680 9882 58686 10058
rect 58720 9882 58726 10058
rect 58680 9870 58726 9882
rect 57741 9776 57777 9870
rect 57977 9776 58013 9870
rect 58213 9777 58249 9870
rect 58375 9822 58441 9829
rect 58375 9788 58391 9822
rect 58425 9788 58441 9822
rect 58375 9777 58441 9788
rect 58213 9776 58441 9777
rect 57741 9747 58441 9776
rect 57741 9746 58323 9747
rect 57861 9633 57895 9746
rect 58257 9705 58323 9746
rect 58257 9671 58273 9705
rect 58307 9671 58323 9705
rect 58257 9664 58323 9671
rect 58685 9665 58720 9870
rect 58892 9665 58959 10255
rect 60651 10232 60692 10264
rect 60938 10260 60948 10326
rect 61004 10260 61014 10326
rect 61684 10302 61694 10410
rect 61826 10347 61836 10410
rect 61826 10336 61838 10347
rect 61826 10302 61839 10336
rect 61694 10264 61839 10302
rect 61798 10236 61839 10264
rect 60067 10204 60337 10232
rect 59808 10138 59818 10204
rect 59884 10138 59894 10204
rect 60067 10142 60101 10204
rect 60303 10142 60337 10204
rect 60421 10204 60692 10232
rect 61209 10208 61479 10236
rect 60421 10142 60455 10204
rect 60657 10142 60692 10204
rect 60833 10192 61004 10208
rect 60833 10158 60964 10192
rect 60998 10158 61004 10192
rect 60833 10142 61004 10158
rect 61209 10146 61243 10208
rect 61445 10146 61479 10208
rect 61563 10208 61839 10236
rect 61563 10146 61597 10208
rect 61799 10146 61839 10208
rect 59943 10130 59989 10142
rect 59943 9754 59949 10130
rect 59983 9754 59989 10130
rect 59943 9742 59989 9754
rect 60061 10130 60107 10142
rect 60061 9754 60067 10130
rect 60101 9754 60107 10130
rect 60061 9742 60107 9754
rect 60179 10130 60225 10142
rect 60179 9754 60185 10130
rect 60219 9754 60225 10130
rect 60179 9742 60225 9754
rect 60297 10130 60343 10142
rect 60297 9754 60303 10130
rect 60337 9754 60343 10130
rect 60297 9742 60343 9754
rect 60415 10130 60461 10142
rect 60415 9754 60421 10130
rect 60455 9754 60461 10130
rect 60415 9742 60461 9754
rect 60533 10130 60579 10142
rect 60533 9754 60539 10130
rect 60573 9754 60579 10130
rect 60533 9742 60579 9754
rect 60651 10130 60697 10142
rect 60651 9754 60657 10130
rect 60691 9754 60697 10130
rect 60651 9742 60697 9754
rect 58685 9637 58959 9665
rect 58331 9633 58959 9637
rect 57855 9621 57901 9633
rect 57855 9245 57861 9621
rect 57895 9245 57901 9621
rect 57855 9233 57901 9245
rect 57973 9621 58019 9633
rect 57973 9245 57979 9621
rect 58013 9245 58019 9621
rect 57973 9233 58019 9245
rect 58091 9621 58137 9633
rect 58091 9245 58097 9621
rect 58131 9269 58137 9621
rect 58208 9621 58254 9633
rect 58208 9445 58214 9621
rect 58248 9445 58254 9621
rect 58208 9433 58254 9445
rect 58326 9621 58959 9633
rect 58326 9445 58332 9621
rect 58366 9608 58959 9621
rect 59949 9700 59983 9742
rect 60185 9700 60219 9742
rect 59949 9672 60219 9700
rect 60303 9701 60337 9742
rect 60539 9701 60573 9742
rect 60303 9672 60573 9701
rect 59949 9624 59983 9672
rect 58366 9445 58372 9608
rect 59949 9594 60012 9624
rect 58326 9433 58372 9445
rect 59977 9502 60012 9594
rect 59977 9466 60204 9502
rect 60474 9491 60484 9588
rect 60583 9491 60593 9588
rect 60657 9559 60691 9742
rect 60657 9505 60766 9559
rect 58214 9317 58249 9433
rect 59977 9359 60012 9466
rect 60138 9432 60204 9466
rect 60138 9398 60154 9432
rect 60188 9398 60204 9432
rect 60485 9490 60582 9491
rect 60485 9423 60542 9490
rect 60138 9392 60204 9398
rect 60379 9387 60648 9423
rect 60379 9359 60412 9387
rect 60615 9359 60648 9387
rect 60732 9359 60766 9505
rect 59853 9347 59899 9359
rect 58345 9317 58453 9327
rect 58214 9269 58345 9317
rect 58453 9288 58601 9294
rect 58131 9245 58345 9269
rect 58091 9233 58345 9245
rect 58097 9229 58345 9233
rect 56973 9201 57733 9228
rect 56973 9195 57970 9201
rect 56973 9161 57920 9195
rect 57954 9161 57970 9195
rect 56973 9145 57970 9161
rect 58022 9195 58088 9201
rect 58022 9161 58038 9195
rect 58072 9161 58088 9195
rect 58271 9185 58345 9229
rect 58589 9221 58601 9288
rect 58453 9215 58601 9221
rect 58345 9175 58453 9185
rect 56973 9129 57733 9145
rect 56973 9128 57670 9129
rect 56973 9124 57205 9128
rect 55243 9095 55289 9107
rect 54376 9056 54410 9095
rect 54612 9056 54646 9095
rect 54376 9020 54646 9056
rect 55013 9057 55046 9095
rect 55249 9057 55282 9095
rect 55013 9021 55282 9057
rect 54376 9019 54542 9020
rect 54410 8940 54542 9019
rect 54400 8832 54410 8940
rect 54542 8832 54552 8940
rect 54436 8703 54442 8832
rect 54509 8703 54515 8832
rect 54436 8691 54515 8703
rect 56385 8713 56989 8741
rect 56385 8607 56837 8713
rect 56949 8700 56989 8713
rect 56949 8607 56991 8700
rect 56385 8596 56991 8607
rect 51014 8458 51991 8488
rect 54208 8486 54271 8503
rect 54133 8482 54271 8486
rect 51014 8352 51046 8458
rect 51250 8352 51282 8458
rect 51486 8352 51518 8458
rect 51722 8352 51754 8458
rect 51957 8352 51991 8458
rect 52301 8448 54271 8482
rect 52299 8419 54271 8448
rect 52299 8403 52345 8419
rect 54133 8417 54271 8419
rect 51007 8340 51053 8352
rect 51007 8164 51013 8340
rect 51047 8164 51053 8340
rect 51007 8152 51053 8164
rect 51125 8340 51171 8352
rect 51125 8164 51131 8340
rect 51165 8164 51171 8340
rect 51125 8152 51171 8164
rect 51243 8340 51289 8352
rect 51243 8164 51249 8340
rect 51283 8164 51289 8340
rect 51243 8152 51289 8164
rect 51361 8340 51407 8352
rect 51361 8164 51367 8340
rect 51401 8164 51407 8340
rect 51361 8152 51407 8164
rect 51479 8340 51525 8352
rect 51479 8164 51485 8340
rect 51519 8164 51525 8340
rect 51479 8152 51525 8164
rect 51597 8340 51643 8352
rect 51597 8164 51603 8340
rect 51637 8164 51643 8340
rect 51597 8152 51643 8164
rect 51715 8340 51761 8352
rect 51715 8164 51721 8340
rect 51755 8164 51761 8340
rect 51715 8152 51761 8164
rect 51833 8340 51879 8352
rect 51833 8164 51839 8340
rect 51873 8164 51879 8340
rect 51833 8152 51879 8164
rect 51951 8340 51997 8352
rect 51951 8164 51957 8340
rect 51991 8164 51997 8340
rect 51951 8152 51997 8164
rect 52069 8340 52115 8352
rect 52069 8164 52075 8340
rect 52109 8164 52115 8340
rect 52069 8152 52115 8164
rect 51130 8058 51166 8152
rect 51366 8058 51402 8152
rect 51602 8059 51638 8152
rect 51764 8104 51830 8111
rect 51764 8070 51780 8104
rect 51814 8070 51830 8104
rect 51764 8059 51830 8070
rect 51602 8058 51830 8059
rect 51130 8029 51830 8058
rect 51130 8028 51712 8029
rect 51250 7915 51284 8028
rect 51646 7987 51712 8028
rect 51646 7953 51662 7987
rect 51696 7953 51712 7987
rect 51646 7946 51712 7953
rect 52074 7934 52109 8152
rect 52298 7951 52345 8403
rect 55189 8407 55268 8419
rect 55189 8295 55195 8407
rect 55262 8295 55268 8407
rect 53257 8187 53267 8295
rect 53399 8187 53409 8295
rect 55155 8187 55165 8295
rect 55297 8187 55307 8295
rect 53267 8147 53399 8187
rect 55165 8147 55297 8187
rect 53266 8081 53399 8147
rect 55164 8081 55297 8147
rect 56385 8096 56535 8596
rect 56596 8595 56989 8596
rect 52595 8038 54068 8081
rect 52298 7935 52344 7951
rect 52263 7934 52344 7935
rect 52074 7919 52344 7934
rect 51720 7915 52344 7919
rect 51244 7903 51290 7915
rect 50979 7425 50989 7543
rect 51107 7511 51117 7543
rect 51244 7527 51250 7903
rect 51284 7527 51290 7903
rect 51244 7515 51290 7527
rect 51362 7903 51408 7915
rect 51362 7527 51368 7903
rect 51402 7527 51408 7903
rect 51362 7515 51408 7527
rect 51480 7903 51526 7915
rect 51480 7527 51486 7903
rect 51520 7551 51526 7903
rect 51597 7903 51643 7915
rect 51597 7727 51603 7903
rect 51637 7727 51643 7903
rect 51597 7715 51643 7727
rect 51715 7903 52344 7915
rect 51715 7727 51721 7903
rect 51755 7891 52344 7903
rect 51755 7890 51997 7891
rect 51755 7727 51761 7890
rect 52263 7889 52344 7891
rect 52595 7735 52629 8038
rect 52961 7935 52995 8038
rect 53197 7935 53231 8038
rect 53433 7935 53467 8038
rect 53669 7935 53703 8038
rect 52955 7923 53001 7935
rect 51715 7715 51761 7727
rect 52471 7723 52517 7735
rect 51603 7599 51638 7715
rect 51734 7599 51842 7609
rect 51603 7551 51734 7599
rect 51842 7561 51986 7567
rect 51520 7527 51734 7551
rect 51480 7515 51734 7527
rect 51486 7511 51734 7515
rect 51107 7483 51122 7511
rect 51107 7477 51359 7483
rect 51107 7443 51309 7477
rect 51343 7443 51359 7477
rect 51107 7427 51359 7443
rect 51411 7477 51477 7483
rect 51411 7443 51427 7477
rect 51461 7443 51477 7477
rect 51660 7467 51734 7511
rect 51974 7494 51986 7561
rect 52471 7547 52477 7723
rect 52511 7547 52517 7723
rect 52471 7535 52517 7547
rect 52589 7723 52635 7735
rect 52589 7547 52595 7723
rect 52629 7547 52635 7723
rect 52589 7535 52635 7547
rect 52707 7723 52753 7735
rect 52707 7547 52713 7723
rect 52747 7547 52753 7723
rect 52707 7535 52753 7547
rect 52825 7723 52871 7735
rect 52955 7723 52961 7923
rect 52825 7547 52831 7723
rect 52865 7547 52961 7723
rect 52995 7547 53001 7923
rect 52825 7535 52871 7547
rect 52955 7535 53001 7547
rect 53073 7923 53119 7935
rect 53073 7547 53079 7923
rect 53113 7547 53119 7923
rect 53073 7535 53119 7547
rect 53191 7923 53237 7935
rect 53191 7547 53197 7923
rect 53231 7547 53237 7923
rect 53191 7535 53237 7547
rect 53309 7923 53355 7935
rect 53309 7547 53315 7923
rect 53349 7547 53355 7923
rect 53309 7535 53355 7547
rect 53427 7923 53473 7935
rect 53427 7547 53433 7923
rect 53467 7547 53473 7923
rect 53427 7535 53473 7547
rect 53545 7923 53591 7935
rect 53545 7547 53551 7923
rect 53585 7547 53591 7923
rect 53545 7535 53591 7547
rect 53663 7923 53709 7935
rect 53663 7547 53669 7923
rect 53703 7723 53709 7923
rect 54034 7735 54068 8038
rect 54493 8038 55966 8081
rect 54493 7735 54527 8038
rect 54859 7935 54893 8038
rect 55095 7935 55129 8038
rect 55331 7935 55365 8038
rect 55567 7935 55601 8038
rect 54853 7923 54899 7935
rect 53792 7723 53838 7735
rect 53703 7547 53798 7723
rect 53832 7547 53838 7723
rect 53663 7535 53709 7547
rect 53792 7535 53838 7547
rect 53910 7723 53956 7735
rect 53910 7547 53916 7723
rect 53950 7547 53956 7723
rect 53910 7535 53956 7547
rect 54028 7723 54074 7735
rect 54028 7547 54034 7723
rect 54068 7547 54074 7723
rect 54028 7535 54074 7547
rect 54146 7723 54192 7735
rect 54146 7547 54152 7723
rect 54186 7547 54192 7723
rect 54146 7535 54192 7547
rect 54369 7723 54415 7735
rect 54369 7547 54375 7723
rect 54409 7547 54415 7723
rect 54369 7535 54415 7547
rect 54487 7723 54533 7735
rect 54487 7547 54493 7723
rect 54527 7547 54533 7723
rect 54487 7535 54533 7547
rect 54605 7723 54651 7735
rect 54605 7547 54611 7723
rect 54645 7547 54651 7723
rect 54605 7535 54651 7547
rect 54723 7723 54769 7735
rect 54853 7723 54859 7923
rect 54723 7547 54729 7723
rect 54763 7547 54859 7723
rect 54893 7547 54899 7923
rect 54723 7535 54769 7547
rect 54853 7535 54899 7547
rect 54971 7923 55017 7935
rect 54971 7547 54977 7923
rect 55011 7547 55017 7923
rect 54971 7535 55017 7547
rect 55089 7923 55135 7935
rect 55089 7547 55095 7923
rect 55129 7547 55135 7923
rect 55089 7535 55135 7547
rect 55207 7923 55253 7935
rect 55207 7547 55213 7923
rect 55247 7547 55253 7923
rect 55207 7535 55253 7547
rect 55325 7923 55371 7935
rect 55325 7547 55331 7923
rect 55365 7547 55371 7923
rect 55325 7535 55371 7547
rect 55443 7923 55489 7935
rect 55443 7547 55449 7923
rect 55483 7547 55489 7923
rect 55443 7535 55489 7547
rect 55561 7923 55607 7935
rect 55561 7547 55567 7923
rect 55601 7723 55607 7923
rect 55932 7735 55966 8038
rect 56384 8030 56535 8096
rect 55690 7723 55736 7735
rect 55601 7547 55696 7723
rect 55730 7547 55736 7723
rect 55561 7535 55607 7547
rect 55690 7535 55736 7547
rect 55808 7723 55854 7735
rect 55808 7547 55814 7723
rect 55848 7547 55854 7723
rect 55808 7535 55854 7547
rect 55926 7723 55972 7735
rect 55926 7547 55932 7723
rect 55966 7547 55972 7723
rect 55926 7535 55972 7547
rect 56044 7723 56090 7735
rect 56044 7547 56050 7723
rect 56084 7547 56090 7723
rect 56044 7535 56090 7547
rect 51842 7488 51986 7494
rect 52477 7501 52511 7535
rect 53079 7501 53113 7535
rect 53315 7501 53349 7535
rect 51734 7457 51842 7467
rect 52477 7466 52636 7501
rect 53079 7466 53349 7501
rect 53916 7501 53950 7535
rect 54152 7501 54186 7535
rect 53916 7466 54186 7501
rect 54375 7501 54409 7535
rect 54977 7501 55011 7535
rect 55213 7501 55247 7535
rect 54375 7466 54534 7501
rect 54977 7466 55247 7501
rect 55814 7501 55848 7535
rect 56050 7501 56084 7535
rect 55814 7466 56084 7501
rect 51107 7425 51122 7427
rect 51022 7411 51122 7425
rect 51022 7368 51122 7369
rect 50643 7347 51122 7368
rect 51411 7347 51477 7443
rect 50643 7299 51477 7347
rect 50643 7270 51122 7299
rect 50643 7268 50748 7270
rect 51022 7269 51122 7270
rect 50476 7083 50486 7162
rect 50579 7083 50589 7162
rect 51477 7152 51556 7164
rect 50487 5909 50580 7083
rect 51477 7054 51483 7152
rect 51405 7034 51483 7054
rect 51550 7054 51556 7152
rect 51550 7034 51625 7054
rect 51405 6926 51449 7034
rect 51581 6926 51625 7034
rect 51405 6884 51625 6926
rect 51009 6854 51986 6884
rect 51009 6748 51041 6854
rect 51245 6748 51277 6854
rect 51481 6748 51513 6854
rect 51717 6748 51749 6854
rect 51952 6748 51986 6854
rect 51002 6736 51048 6748
rect 51002 6560 51008 6736
rect 51042 6560 51048 6736
rect 51002 6548 51048 6560
rect 51120 6736 51166 6748
rect 51120 6560 51126 6736
rect 51160 6560 51166 6736
rect 51120 6548 51166 6560
rect 51238 6736 51284 6748
rect 51238 6560 51244 6736
rect 51278 6560 51284 6736
rect 51238 6548 51284 6560
rect 51356 6736 51402 6748
rect 51356 6560 51362 6736
rect 51396 6560 51402 6736
rect 51356 6548 51402 6560
rect 51474 6736 51520 6748
rect 51474 6560 51480 6736
rect 51514 6560 51520 6736
rect 51474 6548 51520 6560
rect 51592 6736 51638 6748
rect 51592 6560 51598 6736
rect 51632 6560 51638 6736
rect 51592 6548 51638 6560
rect 51710 6736 51756 6748
rect 51710 6560 51716 6736
rect 51750 6560 51756 6736
rect 51710 6548 51756 6560
rect 51828 6736 51874 6748
rect 51828 6560 51834 6736
rect 51868 6560 51874 6736
rect 51828 6548 51874 6560
rect 51946 6736 51992 6748
rect 51946 6560 51952 6736
rect 51986 6560 51992 6736
rect 51946 6548 51992 6560
rect 52064 6736 52110 6748
rect 52064 6560 52070 6736
rect 52104 6560 52110 6736
rect 52064 6548 52110 6560
rect 52602 6682 52636 7466
rect 53315 7404 53349 7466
rect 52904 7366 53646 7404
rect 52904 7242 52938 7366
rect 53140 7242 53174 7366
rect 53376 7242 53410 7366
rect 53612 7242 53646 7366
rect 53902 7259 53912 7325
rect 53975 7259 53985 7325
rect 52898 7230 52944 7242
rect 52898 6854 52904 7230
rect 52938 6854 52944 7230
rect 52898 6842 52944 6854
rect 53016 7230 53062 7242
rect 53016 6854 53022 7230
rect 53056 6854 53062 7230
rect 53016 6842 53062 6854
rect 53134 7230 53180 7242
rect 53134 6854 53140 7230
rect 53174 6854 53180 7230
rect 53134 6842 53180 6854
rect 53252 7230 53298 7242
rect 53252 6854 53258 7230
rect 53292 6854 53298 7230
rect 53252 6842 53298 6854
rect 53370 7230 53416 7242
rect 53370 6854 53376 7230
rect 53410 6854 53416 7230
rect 53370 6842 53416 6854
rect 53488 7230 53534 7242
rect 53488 6854 53494 7230
rect 53528 6854 53534 7230
rect 53488 6842 53534 6854
rect 53606 7230 53652 7242
rect 53606 6854 53612 7230
rect 53646 6854 53652 7230
rect 53606 6842 53652 6854
rect 54018 6683 54052 7466
rect 53745 6682 54052 6683
rect 52602 6677 52918 6682
rect 53632 6677 54052 6682
rect 52602 6666 52985 6677
rect 52602 6639 52934 6666
rect 51125 6454 51161 6548
rect 51361 6454 51397 6548
rect 51597 6455 51633 6548
rect 51759 6500 51825 6507
rect 51759 6466 51775 6500
rect 51809 6466 51825 6500
rect 51759 6455 51825 6466
rect 51597 6454 51825 6455
rect 51125 6425 51825 6454
rect 51125 6424 51707 6425
rect 51245 6311 51279 6424
rect 51641 6383 51707 6424
rect 51641 6349 51657 6383
rect 51691 6349 51707 6383
rect 51641 6342 51707 6349
rect 52069 6315 52104 6548
rect 52602 6510 52636 6639
rect 52918 6632 52934 6639
rect 52968 6632 52985 6666
rect 52918 6626 52985 6632
rect 53565 6666 54052 6677
rect 53565 6632 53582 6666
rect 53616 6639 54052 6666
rect 53616 6632 53632 6639
rect 53745 6638 54052 6639
rect 53565 6626 53632 6632
rect 52743 6599 52799 6611
rect 52743 6565 52749 6599
rect 52783 6598 52799 6599
rect 53856 6598 53912 6610
rect 52783 6582 53250 6598
rect 52783 6565 53200 6582
rect 52743 6549 53200 6565
rect 53184 6548 53200 6549
rect 53234 6548 53250 6582
rect 53184 6541 53250 6548
rect 53302 6583 53872 6598
rect 53302 6549 53318 6583
rect 53352 6564 53872 6583
rect 53906 6564 53912 6598
rect 53352 6549 53912 6564
rect 53302 6539 53369 6549
rect 53856 6548 53912 6549
rect 54018 6510 54052 6638
rect 54500 6682 54534 7466
rect 55213 7404 55247 7466
rect 54802 7366 55544 7404
rect 54802 7242 54836 7366
rect 55038 7242 55072 7366
rect 55274 7242 55308 7366
rect 55510 7242 55544 7366
rect 54796 7230 54842 7242
rect 54796 6854 54802 7230
rect 54836 6854 54842 7230
rect 54796 6842 54842 6854
rect 54914 7230 54960 7242
rect 54914 6854 54920 7230
rect 54954 6854 54960 7230
rect 54914 6842 54960 6854
rect 55032 7230 55078 7242
rect 55032 6854 55038 7230
rect 55072 6854 55078 7230
rect 55032 6842 55078 6854
rect 55150 7230 55196 7242
rect 55150 6854 55156 7230
rect 55190 6854 55196 7230
rect 55150 6842 55196 6854
rect 55268 7230 55314 7242
rect 55268 6854 55274 7230
rect 55308 6854 55314 7230
rect 55268 6842 55314 6854
rect 55386 7230 55432 7242
rect 55386 6854 55392 7230
rect 55426 6854 55432 7230
rect 55386 6842 55432 6854
rect 55504 7230 55550 7242
rect 55504 6854 55510 7230
rect 55544 6854 55550 7230
rect 55504 6842 55550 6854
rect 55916 6683 55950 7466
rect 55528 6682 55597 6683
rect 55643 6682 55950 6683
rect 54500 6677 54816 6682
rect 55528 6678 55950 6682
rect 54500 6666 54883 6677
rect 54500 6639 54832 6666
rect 54500 6510 54534 6639
rect 54816 6632 54832 6639
rect 54866 6632 54883 6666
rect 54816 6626 54883 6632
rect 55461 6667 55950 6678
rect 55461 6633 55478 6667
rect 55512 6639 55950 6667
rect 55512 6633 55528 6639
rect 55643 6638 55950 6639
rect 55461 6627 55528 6633
rect 54641 6599 54697 6611
rect 54641 6565 54647 6599
rect 54681 6598 54697 6599
rect 55754 6598 55810 6610
rect 54681 6582 55148 6598
rect 54681 6565 55098 6582
rect 54641 6549 55098 6565
rect 55082 6548 55098 6549
rect 55132 6548 55148 6582
rect 55082 6541 55148 6548
rect 55200 6583 55770 6598
rect 55200 6549 55216 6583
rect 55250 6564 55770 6583
rect 55804 6564 55810 6598
rect 55250 6549 55810 6564
rect 55200 6539 55267 6549
rect 55754 6548 55810 6549
rect 55916 6510 55950 6638
rect 56031 7288 56098 7312
rect 56031 7254 56048 7288
rect 56082 7254 56098 7288
rect 51715 6311 52104 6315
rect 51239 6299 51285 6311
rect 51239 5923 51245 6299
rect 51279 5923 51285 6299
rect 51239 5911 51285 5923
rect 51357 6299 51403 6311
rect 51357 5923 51363 6299
rect 51397 5923 51403 6299
rect 51357 5911 51403 5923
rect 51475 6299 51521 6311
rect 51475 5923 51481 6299
rect 51515 5947 51521 6299
rect 51592 6299 51638 6311
rect 51592 6123 51598 6299
rect 51632 6123 51638 6299
rect 51592 6111 51638 6123
rect 51710 6299 52104 6311
rect 52596 6498 52642 6510
rect 52596 6322 52602 6498
rect 52636 6322 52642 6498
rect 52596 6310 52642 6322
rect 52714 6498 52760 6510
rect 52714 6322 52720 6498
rect 52754 6322 52760 6498
rect 52714 6310 52760 6322
rect 53016 6498 53062 6510
rect 51710 6123 51716 6299
rect 51750 6286 52104 6299
rect 51750 6123 51756 6286
rect 52026 6283 52104 6286
rect 52026 6231 52036 6283
rect 52099 6231 52109 6283
rect 52031 6225 52104 6231
rect 51710 6111 51756 6123
rect 51598 5995 51633 6111
rect 52719 6016 52753 6310
rect 53016 6122 53022 6498
rect 53056 6122 53062 6498
rect 53016 6110 53062 6122
rect 53134 6498 53180 6510
rect 53134 6122 53140 6498
rect 53174 6122 53180 6498
rect 53134 6110 53180 6122
rect 53252 6498 53298 6510
rect 53252 6122 53258 6498
rect 53292 6122 53298 6498
rect 53252 6110 53298 6122
rect 53370 6498 53416 6510
rect 53370 6122 53376 6498
rect 53410 6122 53416 6498
rect 53370 6110 53416 6122
rect 53488 6498 53534 6510
rect 53488 6122 53494 6498
rect 53528 6122 53534 6498
rect 53894 6498 53940 6510
rect 53894 6322 53900 6498
rect 53934 6322 53940 6498
rect 53894 6310 53940 6322
rect 54012 6498 54058 6510
rect 54012 6322 54018 6498
rect 54052 6322 54058 6498
rect 54012 6310 54058 6322
rect 54494 6498 54540 6510
rect 54494 6322 54500 6498
rect 54534 6322 54540 6498
rect 54494 6310 54540 6322
rect 54612 6498 54658 6510
rect 54612 6322 54618 6498
rect 54652 6322 54658 6498
rect 54612 6310 54658 6322
rect 54914 6498 54960 6510
rect 53488 6110 53534 6122
rect 53376 6016 53410 6110
rect 53900 6016 53933 6310
rect 51729 5995 51837 6005
rect 51598 5947 51729 5995
rect 52719 5984 53933 6016
rect 54617 6016 54651 6310
rect 54914 6122 54920 6498
rect 54954 6122 54960 6498
rect 54914 6110 54960 6122
rect 55032 6498 55078 6510
rect 55032 6122 55038 6498
rect 55072 6122 55078 6498
rect 55032 6110 55078 6122
rect 55150 6498 55196 6510
rect 55150 6122 55156 6498
rect 55190 6122 55196 6498
rect 55150 6110 55196 6122
rect 55268 6498 55314 6510
rect 55268 6122 55274 6498
rect 55308 6122 55314 6498
rect 55268 6110 55314 6122
rect 55386 6498 55432 6510
rect 55386 6122 55392 6498
rect 55426 6122 55432 6498
rect 55792 6498 55838 6510
rect 55792 6322 55798 6498
rect 55832 6322 55838 6498
rect 55792 6310 55838 6322
rect 55910 6498 55956 6510
rect 55910 6322 55916 6498
rect 55950 6322 55956 6498
rect 55910 6310 55956 6322
rect 55386 6110 55432 6122
rect 55274 6016 55308 6110
rect 55798 6016 55831 6310
rect 54617 5984 55831 6016
rect 51837 5956 51988 5962
rect 51515 5923 51729 5947
rect 51475 5911 51729 5923
rect 50487 5907 51072 5909
rect 51481 5907 51729 5911
rect 50487 5879 51117 5907
rect 50487 5873 51354 5879
rect 50487 5839 51304 5873
rect 51338 5839 51354 5873
rect 50487 5823 51354 5839
rect 51406 5873 51472 5879
rect 51406 5839 51422 5873
rect 51456 5839 51472 5873
rect 51655 5863 51729 5907
rect 51976 5889 51988 5956
rect 53212 5899 53344 5984
rect 55110 5899 55242 5984
rect 51837 5883 51988 5889
rect 51729 5853 51837 5863
rect 50487 5807 51117 5823
rect 50487 5803 51072 5807
rect 50487 5802 50588 5803
rect 51017 5754 51117 5765
rect 50981 5648 50991 5754
rect 51103 5743 51117 5754
rect 51406 5743 51472 5839
rect 53202 5791 53212 5899
rect 53344 5791 53354 5899
rect 55100 5791 55110 5899
rect 55242 5791 55252 5899
rect 56031 5871 56098 7254
rect 51103 5695 51472 5743
rect 51103 5665 51117 5695
rect 51103 5648 51113 5665
rect 51405 5592 51471 5695
rect 53230 5655 53236 5791
rect 53303 5655 53309 5791
rect 53230 5643 53309 5655
rect 56031 5592 56097 5871
rect 51403 5512 56097 5592
rect 50145 5478 50308 5492
rect 50145 5410 50189 5478
rect 50259 5410 50308 5478
rect 50145 4691 50308 5410
rect 56153 5398 56163 5512
rect 56286 5398 56296 5512
rect 50145 4661 50309 4691
rect 50145 4593 50188 4661
rect 50258 4593 50309 4661
rect 53944 4660 54023 4672
rect 50145 4579 50309 4593
rect 51459 4600 51538 4612
rect 51459 4507 51465 4600
rect 51391 4487 51465 4507
rect 51532 4507 51538 4600
rect 53944 4541 53950 4660
rect 54017 4541 54023 4660
rect 55093 4657 55172 4669
rect 55093 4541 55099 4657
rect 55166 4541 55172 4657
rect 51532 4487 51611 4507
rect 51391 4379 51435 4487
rect 51567 4379 51611 4487
rect 53188 4445 53244 4453
rect 51391 4337 51611 4379
rect 52262 4437 53244 4445
rect 52262 4403 53204 4437
rect 53238 4403 53244 4437
rect 53907 4433 53917 4541
rect 54049 4478 54059 4541
rect 54049 4467 54061 4478
rect 54049 4433 54062 4467
rect 54318 4457 54374 4459
rect 52262 4387 53244 4403
rect 53917 4395 54062 4433
rect 52262 4386 53241 4387
rect 50995 4307 51972 4337
rect 50995 4201 51027 4307
rect 51231 4201 51263 4307
rect 51467 4201 51499 4307
rect 51703 4201 51735 4307
rect 51938 4201 51972 4307
rect 50988 4189 51034 4201
rect 50988 4013 50994 4189
rect 51028 4013 51034 4189
rect 50988 4001 51034 4013
rect 51106 4189 51152 4201
rect 51106 4013 51112 4189
rect 51146 4013 51152 4189
rect 51106 4001 51152 4013
rect 51224 4189 51270 4201
rect 51224 4013 51230 4189
rect 51264 4013 51270 4189
rect 51224 4001 51270 4013
rect 51342 4189 51388 4201
rect 51342 4013 51348 4189
rect 51382 4013 51388 4189
rect 51342 4001 51388 4013
rect 51460 4189 51506 4201
rect 51460 4013 51466 4189
rect 51500 4013 51506 4189
rect 51460 4001 51506 4013
rect 51578 4189 51624 4201
rect 51578 4013 51584 4189
rect 51618 4013 51624 4189
rect 51578 4001 51624 4013
rect 51696 4189 51742 4201
rect 51696 4013 51702 4189
rect 51736 4013 51742 4189
rect 51696 4001 51742 4013
rect 51814 4189 51860 4201
rect 51814 4013 51820 4189
rect 51854 4013 51860 4189
rect 51814 4001 51860 4013
rect 51932 4189 51978 4201
rect 51932 4013 51938 4189
rect 51972 4013 51978 4189
rect 51932 4001 51978 4013
rect 52050 4189 52096 4201
rect 52050 4013 52056 4189
rect 52090 4013 52096 4189
rect 52050 4001 52096 4013
rect 51111 3907 51147 4001
rect 51347 3907 51383 4001
rect 51583 3908 51619 4001
rect 51745 3953 51811 3960
rect 51745 3919 51761 3953
rect 51795 3919 51811 3953
rect 51745 3908 51811 3919
rect 51583 3907 51811 3908
rect 51111 3878 51811 3907
rect 51111 3877 51693 3878
rect 51231 3764 51265 3877
rect 51627 3836 51693 3877
rect 51627 3802 51643 3836
rect 51677 3802 51693 3836
rect 51627 3795 51693 3802
rect 52055 3796 52090 4001
rect 52262 3796 52329 4386
rect 54021 4363 54062 4395
rect 54308 4391 54318 4457
rect 54374 4391 54384 4457
rect 55054 4433 55064 4541
rect 55196 4478 55206 4541
rect 55196 4467 55208 4478
rect 55196 4433 55209 4467
rect 55064 4395 55209 4433
rect 55168 4367 55209 4395
rect 53437 4335 53707 4363
rect 53178 4269 53188 4335
rect 53254 4269 53264 4335
rect 53437 4273 53471 4335
rect 53673 4273 53707 4335
rect 53791 4335 54062 4363
rect 54579 4339 54849 4367
rect 53791 4273 53825 4335
rect 54027 4273 54062 4335
rect 54203 4323 54374 4339
rect 54203 4289 54334 4323
rect 54368 4289 54374 4323
rect 54203 4273 54374 4289
rect 54579 4277 54613 4339
rect 54815 4277 54849 4339
rect 54933 4339 55209 4367
rect 54933 4277 54967 4339
rect 55169 4277 55209 4339
rect 53313 4261 53359 4273
rect 53313 3885 53319 4261
rect 53353 3885 53359 4261
rect 53313 3873 53359 3885
rect 53431 4261 53477 4273
rect 53431 3885 53437 4261
rect 53471 3885 53477 4261
rect 53431 3873 53477 3885
rect 53549 4261 53595 4273
rect 53549 3885 53555 4261
rect 53589 3885 53595 4261
rect 53549 3873 53595 3885
rect 53667 4261 53713 4273
rect 53667 3885 53673 4261
rect 53707 3885 53713 4261
rect 53667 3873 53713 3885
rect 53785 4261 53831 4273
rect 53785 3885 53791 4261
rect 53825 3885 53831 4261
rect 53785 3873 53831 3885
rect 53903 4261 53949 4273
rect 53903 3885 53909 4261
rect 53943 3885 53949 4261
rect 53903 3873 53949 3885
rect 54021 4261 54067 4273
rect 54021 3885 54027 4261
rect 54061 3885 54067 4261
rect 54021 3873 54067 3885
rect 52055 3768 52329 3796
rect 51701 3764 52329 3768
rect 51225 3752 51271 3764
rect 51225 3376 51231 3752
rect 51265 3376 51271 3752
rect 51225 3364 51271 3376
rect 51343 3752 51389 3764
rect 51343 3376 51349 3752
rect 51383 3376 51389 3752
rect 51343 3364 51389 3376
rect 51461 3752 51507 3764
rect 51461 3376 51467 3752
rect 51501 3400 51507 3752
rect 51578 3752 51624 3764
rect 51578 3576 51584 3752
rect 51618 3576 51624 3752
rect 51578 3564 51624 3576
rect 51696 3752 52329 3764
rect 51696 3576 51702 3752
rect 51736 3739 52329 3752
rect 53319 3831 53353 3873
rect 53555 3831 53589 3873
rect 53319 3803 53589 3831
rect 53673 3832 53707 3873
rect 53909 3832 53943 3873
rect 53673 3803 53943 3832
rect 53319 3755 53353 3803
rect 51736 3576 51742 3739
rect 53319 3725 53382 3755
rect 51696 3564 51742 3576
rect 53347 3633 53382 3725
rect 53347 3597 53574 3633
rect 53844 3622 53854 3719
rect 53953 3622 53963 3719
rect 54027 3690 54061 3873
rect 54027 3636 54136 3690
rect 51584 3448 51619 3564
rect 53347 3490 53382 3597
rect 53508 3563 53574 3597
rect 53508 3529 53524 3563
rect 53558 3529 53574 3563
rect 53855 3621 53952 3622
rect 53855 3554 53912 3621
rect 53508 3523 53574 3529
rect 53749 3518 54018 3554
rect 53749 3490 53782 3518
rect 53985 3490 54018 3518
rect 54102 3490 54136 3636
rect 53223 3478 53269 3490
rect 51715 3448 51823 3458
rect 51584 3400 51715 3448
rect 51823 3412 51974 3418
rect 51501 3376 51715 3400
rect 51461 3364 51715 3376
rect 51467 3360 51715 3364
rect 49778 3359 50401 3360
rect 49778 3332 51103 3359
rect 49778 3326 51340 3332
rect 47716 3254 47750 3293
rect 47952 3254 47986 3293
rect 47716 3218 47986 3254
rect 48353 3255 48386 3293
rect 48589 3255 48622 3293
rect 48353 3219 48622 3255
rect 49778 3292 51290 3326
rect 51324 3292 51340 3326
rect 49778 3276 51340 3292
rect 51392 3326 51458 3332
rect 51392 3292 51408 3326
rect 51442 3292 51458 3326
rect 51641 3316 51715 3360
rect 51962 3345 51974 3412
rect 51823 3339 51974 3345
rect 51715 3306 51823 3316
rect 49778 3260 51103 3276
rect 49778 3259 51040 3260
rect 49778 3255 50575 3259
rect 49778 3254 50401 3255
rect 47716 3217 47882 3218
rect 47750 3138 47882 3217
rect 47740 3030 47750 3138
rect 47882 3030 47892 3138
rect 47772 2885 47778 3030
rect 47845 2885 47851 3030
rect 47772 2873 47851 2885
rect 49779 2867 50360 2875
rect 49778 2849 50360 2867
rect 49778 2736 50140 2849
rect 50344 2831 50360 2849
rect 49778 2735 50292 2736
rect 50344 2735 50361 2831
rect 49778 2725 50361 2735
rect 44354 2656 45331 2686
rect 47548 2684 47611 2701
rect 47473 2680 47611 2684
rect 44354 2550 44386 2656
rect 44590 2550 44622 2656
rect 44826 2550 44858 2656
rect 45062 2550 45094 2656
rect 45297 2550 45331 2656
rect 45641 2646 47611 2680
rect 45639 2617 47611 2646
rect 45639 2601 45685 2617
rect 47473 2615 47611 2617
rect 44347 2538 44393 2550
rect 44347 2362 44353 2538
rect 44387 2362 44393 2538
rect 44347 2350 44393 2362
rect 44465 2538 44511 2550
rect 44465 2362 44471 2538
rect 44505 2362 44511 2538
rect 44465 2350 44511 2362
rect 44583 2538 44629 2550
rect 44583 2362 44589 2538
rect 44623 2362 44629 2538
rect 44583 2350 44629 2362
rect 44701 2538 44747 2550
rect 44701 2362 44707 2538
rect 44741 2362 44747 2538
rect 44701 2350 44747 2362
rect 44819 2538 44865 2550
rect 44819 2362 44825 2538
rect 44859 2362 44865 2538
rect 44819 2350 44865 2362
rect 44937 2538 44983 2550
rect 44937 2362 44943 2538
rect 44977 2362 44983 2538
rect 44937 2350 44983 2362
rect 45055 2538 45101 2550
rect 45055 2362 45061 2538
rect 45095 2362 45101 2538
rect 45055 2350 45101 2362
rect 45173 2538 45219 2550
rect 45173 2362 45179 2538
rect 45213 2362 45219 2538
rect 45173 2350 45219 2362
rect 45291 2538 45337 2550
rect 45291 2362 45297 2538
rect 45331 2362 45337 2538
rect 45291 2350 45337 2362
rect 45409 2538 45455 2550
rect 45409 2362 45415 2538
rect 45449 2362 45455 2538
rect 45409 2350 45455 2362
rect 44470 2256 44506 2350
rect 44706 2256 44742 2350
rect 44942 2257 44978 2350
rect 45104 2302 45170 2309
rect 45104 2268 45120 2302
rect 45154 2268 45170 2302
rect 45104 2257 45170 2268
rect 44942 2256 45170 2257
rect 44470 2227 45170 2256
rect 44470 2226 45052 2227
rect 44590 2113 44624 2226
rect 44986 2185 45052 2226
rect 44986 2151 45002 2185
rect 45036 2151 45052 2185
rect 44986 2144 45052 2151
rect 45414 2132 45449 2350
rect 45638 2149 45685 2601
rect 48536 2610 48615 2622
rect 48536 2493 48542 2610
rect 48609 2493 48615 2610
rect 46597 2385 46607 2493
rect 46739 2385 46749 2493
rect 48495 2385 48505 2493
rect 48637 2385 48647 2493
rect 46607 2345 46739 2385
rect 48505 2345 48637 2385
rect 46606 2279 46739 2345
rect 48504 2279 48637 2345
rect 45935 2236 47408 2279
rect 45638 2133 45684 2149
rect 45603 2132 45684 2133
rect 45414 2117 45684 2132
rect 45060 2113 45684 2117
rect 44584 2101 44630 2113
rect 44319 1623 44329 1741
rect 44447 1709 44457 1741
rect 44584 1725 44590 2101
rect 44624 1725 44630 2101
rect 44584 1713 44630 1725
rect 44702 2101 44748 2113
rect 44702 1725 44708 2101
rect 44742 1725 44748 2101
rect 44702 1713 44748 1725
rect 44820 2101 44866 2113
rect 44820 1725 44826 2101
rect 44860 1749 44866 2101
rect 44937 2101 44983 2113
rect 44937 1925 44943 2101
rect 44977 1925 44983 2101
rect 44937 1913 44983 1925
rect 45055 2101 45684 2113
rect 45055 1925 45061 2101
rect 45095 2089 45684 2101
rect 45095 2088 45337 2089
rect 45095 1925 45101 2088
rect 45603 2087 45684 2089
rect 45935 1933 45969 2236
rect 46301 2133 46335 2236
rect 46537 2133 46571 2236
rect 46773 2133 46807 2236
rect 47009 2133 47043 2236
rect 46295 2121 46341 2133
rect 45055 1913 45101 1925
rect 45811 1921 45857 1933
rect 44943 1797 44978 1913
rect 45074 1797 45182 1807
rect 44943 1749 45074 1797
rect 45182 1758 45329 1764
rect 44860 1725 45074 1749
rect 44820 1713 45074 1725
rect 44826 1709 45074 1713
rect 44447 1681 44462 1709
rect 44447 1675 44699 1681
rect 44447 1641 44649 1675
rect 44683 1641 44699 1675
rect 44447 1625 44699 1641
rect 44751 1675 44817 1681
rect 44751 1641 44767 1675
rect 44801 1641 44817 1675
rect 45000 1665 45074 1709
rect 45317 1691 45329 1758
rect 45811 1745 45817 1921
rect 45851 1745 45857 1921
rect 45811 1733 45857 1745
rect 45929 1921 45975 1933
rect 45929 1745 45935 1921
rect 45969 1745 45975 1921
rect 45929 1733 45975 1745
rect 46047 1921 46093 1933
rect 46047 1745 46053 1921
rect 46087 1745 46093 1921
rect 46047 1733 46093 1745
rect 46165 1921 46211 1933
rect 46295 1921 46301 2121
rect 46165 1745 46171 1921
rect 46205 1745 46301 1921
rect 46335 1745 46341 2121
rect 46165 1733 46211 1745
rect 46295 1733 46341 1745
rect 46413 2121 46459 2133
rect 46413 1745 46419 2121
rect 46453 1745 46459 2121
rect 46413 1733 46459 1745
rect 46531 2121 46577 2133
rect 46531 1745 46537 2121
rect 46571 1745 46577 2121
rect 46531 1733 46577 1745
rect 46649 2121 46695 2133
rect 46649 1745 46655 2121
rect 46689 1745 46695 2121
rect 46649 1733 46695 1745
rect 46767 2121 46813 2133
rect 46767 1745 46773 2121
rect 46807 1745 46813 2121
rect 46767 1733 46813 1745
rect 46885 2121 46931 2133
rect 46885 1745 46891 2121
rect 46925 1745 46931 2121
rect 46885 1733 46931 1745
rect 47003 2121 47049 2133
rect 47003 1745 47009 2121
rect 47043 1921 47049 2121
rect 47374 1933 47408 2236
rect 47833 2236 49306 2279
rect 47833 1933 47867 2236
rect 48199 2133 48233 2236
rect 48435 2133 48469 2236
rect 48671 2133 48705 2236
rect 48907 2133 48941 2236
rect 48193 2121 48239 2133
rect 47132 1921 47178 1933
rect 47043 1745 47138 1921
rect 47172 1745 47178 1921
rect 47003 1733 47049 1745
rect 47132 1733 47178 1745
rect 47250 1921 47296 1933
rect 47250 1745 47256 1921
rect 47290 1745 47296 1921
rect 47250 1733 47296 1745
rect 47368 1921 47414 1933
rect 47368 1745 47374 1921
rect 47408 1745 47414 1921
rect 47368 1733 47414 1745
rect 47486 1921 47532 1933
rect 47486 1745 47492 1921
rect 47526 1745 47532 1921
rect 47486 1733 47532 1745
rect 47709 1921 47755 1933
rect 47709 1745 47715 1921
rect 47749 1745 47755 1921
rect 47709 1733 47755 1745
rect 47827 1921 47873 1933
rect 47827 1745 47833 1921
rect 47867 1745 47873 1921
rect 47827 1733 47873 1745
rect 47945 1921 47991 1933
rect 47945 1745 47951 1921
rect 47985 1745 47991 1921
rect 47945 1733 47991 1745
rect 48063 1921 48109 1933
rect 48193 1921 48199 2121
rect 48063 1745 48069 1921
rect 48103 1745 48199 1921
rect 48233 1745 48239 2121
rect 48063 1733 48109 1745
rect 48193 1733 48239 1745
rect 48311 2121 48357 2133
rect 48311 1745 48317 2121
rect 48351 1745 48357 2121
rect 48311 1733 48357 1745
rect 48429 2121 48475 2133
rect 48429 1745 48435 2121
rect 48469 1745 48475 2121
rect 48429 1733 48475 1745
rect 48547 2121 48593 2133
rect 48547 1745 48553 2121
rect 48587 1745 48593 2121
rect 48547 1733 48593 1745
rect 48665 2121 48711 2133
rect 48665 1745 48671 2121
rect 48705 1745 48711 2121
rect 48665 1733 48711 1745
rect 48783 2121 48829 2133
rect 48783 1745 48789 2121
rect 48823 1745 48829 2121
rect 48783 1733 48829 1745
rect 48901 2121 48947 2133
rect 48901 1745 48907 2121
rect 48941 1921 48947 2121
rect 49272 1933 49306 2236
rect 49030 1921 49076 1933
rect 48941 1745 49036 1921
rect 49070 1745 49076 1921
rect 48901 1733 48947 1745
rect 49030 1733 49076 1745
rect 49148 1921 49194 1933
rect 49148 1745 49154 1921
rect 49188 1745 49194 1921
rect 49148 1733 49194 1745
rect 49266 1921 49312 1933
rect 49266 1745 49272 1921
rect 49306 1745 49312 1921
rect 49266 1733 49312 1745
rect 49384 1921 49430 1933
rect 49384 1745 49390 1921
rect 49424 1745 49430 1921
rect 49384 1733 49430 1745
rect 45182 1685 45329 1691
rect 45817 1699 45851 1733
rect 46419 1699 46453 1733
rect 46655 1699 46689 1733
rect 45074 1655 45182 1665
rect 45817 1664 45976 1699
rect 46419 1664 46689 1699
rect 47256 1699 47290 1733
rect 47492 1699 47526 1733
rect 47256 1664 47526 1699
rect 47715 1699 47749 1733
rect 48317 1699 48351 1733
rect 48553 1699 48587 1733
rect 47715 1664 47874 1699
rect 48317 1664 48587 1699
rect 49154 1699 49188 1733
rect 49390 1699 49424 1733
rect 49154 1664 49424 1699
rect 44447 1623 44462 1625
rect 44362 1609 44462 1623
rect 44362 1566 44462 1567
rect 43983 1545 44462 1566
rect 44751 1545 44817 1641
rect 43983 1497 44817 1545
rect 43983 1468 44462 1497
rect 43983 1466 44088 1468
rect 44362 1467 44462 1468
rect 43816 1281 43826 1360
rect 43919 1281 43929 1360
rect 44819 1348 44898 1360
rect 43827 107 43920 1281
rect 44819 1252 44825 1348
rect 44745 1232 44825 1252
rect 44892 1252 44898 1348
rect 44892 1232 44965 1252
rect 44745 1124 44789 1232
rect 44921 1124 44965 1232
rect 44745 1082 44965 1124
rect 44349 1052 45326 1082
rect 44349 946 44381 1052
rect 44585 946 44617 1052
rect 44821 946 44853 1052
rect 45057 946 45089 1052
rect 45292 946 45326 1052
rect 44342 934 44388 946
rect 44342 758 44348 934
rect 44382 758 44388 934
rect 44342 746 44388 758
rect 44460 934 44506 946
rect 44460 758 44466 934
rect 44500 758 44506 934
rect 44460 746 44506 758
rect 44578 934 44624 946
rect 44578 758 44584 934
rect 44618 758 44624 934
rect 44578 746 44624 758
rect 44696 934 44742 946
rect 44696 758 44702 934
rect 44736 758 44742 934
rect 44696 746 44742 758
rect 44814 934 44860 946
rect 44814 758 44820 934
rect 44854 758 44860 934
rect 44814 746 44860 758
rect 44932 934 44978 946
rect 44932 758 44938 934
rect 44972 758 44978 934
rect 44932 746 44978 758
rect 45050 934 45096 946
rect 45050 758 45056 934
rect 45090 758 45096 934
rect 45050 746 45096 758
rect 45168 934 45214 946
rect 45168 758 45174 934
rect 45208 758 45214 934
rect 45168 746 45214 758
rect 45286 934 45332 946
rect 45286 758 45292 934
rect 45326 758 45332 934
rect 45286 746 45332 758
rect 45404 934 45450 946
rect 45404 758 45410 934
rect 45444 758 45450 934
rect 45404 746 45450 758
rect 45942 880 45976 1664
rect 46655 1602 46689 1664
rect 46244 1564 46986 1602
rect 46244 1440 46278 1564
rect 46480 1440 46514 1564
rect 46716 1440 46750 1564
rect 46952 1440 46986 1564
rect 47242 1457 47252 1523
rect 47315 1457 47325 1523
rect 46238 1428 46284 1440
rect 46238 1052 46244 1428
rect 46278 1052 46284 1428
rect 46238 1040 46284 1052
rect 46356 1428 46402 1440
rect 46356 1052 46362 1428
rect 46396 1052 46402 1428
rect 46356 1040 46402 1052
rect 46474 1428 46520 1440
rect 46474 1052 46480 1428
rect 46514 1052 46520 1428
rect 46474 1040 46520 1052
rect 46592 1428 46638 1440
rect 46592 1052 46598 1428
rect 46632 1052 46638 1428
rect 46592 1040 46638 1052
rect 46710 1428 46756 1440
rect 46710 1052 46716 1428
rect 46750 1052 46756 1428
rect 46710 1040 46756 1052
rect 46828 1428 46874 1440
rect 46828 1052 46834 1428
rect 46868 1052 46874 1428
rect 46828 1040 46874 1052
rect 46946 1428 46992 1440
rect 46946 1052 46952 1428
rect 46986 1052 46992 1428
rect 46946 1040 46992 1052
rect 47358 881 47392 1664
rect 47085 880 47392 881
rect 45942 875 46258 880
rect 46972 875 47392 880
rect 45942 864 46325 875
rect 45942 837 46274 864
rect 44465 652 44501 746
rect 44701 652 44737 746
rect 44937 653 44973 746
rect 45099 698 45165 705
rect 45099 664 45115 698
rect 45149 664 45165 698
rect 45099 653 45165 664
rect 44937 652 45165 653
rect 44465 623 45165 652
rect 44465 622 45047 623
rect 44585 509 44619 622
rect 44981 581 45047 622
rect 44981 547 44997 581
rect 45031 547 45047 581
rect 44981 540 45047 547
rect 45409 513 45444 746
rect 45942 708 45976 837
rect 46258 830 46274 837
rect 46308 830 46325 864
rect 46258 824 46325 830
rect 46905 864 47392 875
rect 46905 830 46922 864
rect 46956 837 47392 864
rect 46956 830 46972 837
rect 47085 836 47392 837
rect 46905 824 46972 830
rect 46083 797 46139 809
rect 46083 763 46089 797
rect 46123 796 46139 797
rect 47196 796 47252 808
rect 46123 780 46590 796
rect 46123 763 46540 780
rect 46083 747 46540 763
rect 46524 746 46540 747
rect 46574 746 46590 780
rect 46524 739 46590 746
rect 46642 781 47212 796
rect 46642 747 46658 781
rect 46692 762 47212 781
rect 47246 762 47252 796
rect 46692 747 47252 762
rect 46642 737 46709 747
rect 47196 746 47252 747
rect 47358 708 47392 836
rect 47840 880 47874 1664
rect 48553 1602 48587 1664
rect 48142 1564 48884 1602
rect 48142 1440 48176 1564
rect 48378 1440 48412 1564
rect 48614 1440 48648 1564
rect 48850 1440 48884 1564
rect 48136 1428 48182 1440
rect 48136 1052 48142 1428
rect 48176 1052 48182 1428
rect 48136 1040 48182 1052
rect 48254 1428 48300 1440
rect 48254 1052 48260 1428
rect 48294 1052 48300 1428
rect 48254 1040 48300 1052
rect 48372 1428 48418 1440
rect 48372 1052 48378 1428
rect 48412 1052 48418 1428
rect 48372 1040 48418 1052
rect 48490 1428 48536 1440
rect 48490 1052 48496 1428
rect 48530 1052 48536 1428
rect 48490 1040 48536 1052
rect 48608 1428 48654 1440
rect 48608 1052 48614 1428
rect 48648 1052 48654 1428
rect 48608 1040 48654 1052
rect 48726 1428 48772 1440
rect 48726 1052 48732 1428
rect 48766 1052 48772 1428
rect 48726 1040 48772 1052
rect 48844 1428 48890 1440
rect 48844 1052 48850 1428
rect 48884 1052 48890 1428
rect 48844 1040 48890 1052
rect 49256 881 49290 1664
rect 48868 880 48937 881
rect 48983 880 49290 881
rect 47840 875 48156 880
rect 48868 876 49290 880
rect 47840 864 48223 875
rect 47840 837 48172 864
rect 47840 708 47874 837
rect 48156 830 48172 837
rect 48206 830 48223 864
rect 48156 824 48223 830
rect 48801 865 49290 876
rect 48801 831 48818 865
rect 48852 837 49290 865
rect 48852 831 48868 837
rect 48983 836 49290 837
rect 48801 825 48868 831
rect 47981 797 48037 809
rect 47981 763 47987 797
rect 48021 796 48037 797
rect 49094 796 49150 808
rect 48021 780 48488 796
rect 48021 763 48438 780
rect 47981 747 48438 763
rect 48422 746 48438 747
rect 48472 746 48488 780
rect 48422 739 48488 746
rect 48540 781 49110 796
rect 48540 747 48556 781
rect 48590 762 49110 781
rect 49144 762 49150 796
rect 48590 747 49150 762
rect 48540 737 48607 747
rect 49094 746 49150 747
rect 49256 708 49290 836
rect 49371 1486 49438 1510
rect 49371 1452 49388 1486
rect 49422 1452 49438 1486
rect 45055 509 45444 513
rect 44579 497 44625 509
rect 44579 121 44585 497
rect 44619 121 44625 497
rect 44579 109 44625 121
rect 44697 497 44743 509
rect 44697 121 44703 497
rect 44737 121 44743 497
rect 44697 109 44743 121
rect 44815 497 44861 509
rect 44815 121 44821 497
rect 44855 145 44861 497
rect 44932 497 44978 509
rect 44932 321 44938 497
rect 44972 321 44978 497
rect 44932 309 44978 321
rect 45050 497 45444 509
rect 45936 696 45982 708
rect 45936 520 45942 696
rect 45976 520 45982 696
rect 45936 508 45982 520
rect 46054 696 46100 708
rect 46054 520 46060 696
rect 46094 520 46100 696
rect 46054 508 46100 520
rect 46356 696 46402 708
rect 45050 321 45056 497
rect 45090 484 45444 497
rect 45090 321 45096 484
rect 45366 481 45444 484
rect 45366 429 45376 481
rect 45439 429 45449 481
rect 45371 423 45444 429
rect 45050 309 45096 321
rect 44938 193 44973 309
rect 46059 214 46093 508
rect 46356 320 46362 696
rect 46396 320 46402 696
rect 46356 308 46402 320
rect 46474 696 46520 708
rect 46474 320 46480 696
rect 46514 320 46520 696
rect 46474 308 46520 320
rect 46592 696 46638 708
rect 46592 320 46598 696
rect 46632 320 46638 696
rect 46592 308 46638 320
rect 46710 696 46756 708
rect 46710 320 46716 696
rect 46750 320 46756 696
rect 46710 308 46756 320
rect 46828 696 46874 708
rect 46828 320 46834 696
rect 46868 320 46874 696
rect 47234 696 47280 708
rect 47234 520 47240 696
rect 47274 520 47280 696
rect 47234 508 47280 520
rect 47352 696 47398 708
rect 47352 520 47358 696
rect 47392 520 47398 696
rect 47352 508 47398 520
rect 47834 696 47880 708
rect 47834 520 47840 696
rect 47874 520 47880 696
rect 47834 508 47880 520
rect 47952 696 47998 708
rect 47952 520 47958 696
rect 47992 520 47998 696
rect 47952 508 47998 520
rect 48254 696 48300 708
rect 46828 308 46874 320
rect 46716 214 46750 308
rect 47240 214 47273 508
rect 45069 193 45177 203
rect 44938 145 45069 193
rect 46059 182 47273 214
rect 47957 214 47991 508
rect 48254 320 48260 696
rect 48294 320 48300 696
rect 48254 308 48300 320
rect 48372 696 48418 708
rect 48372 320 48378 696
rect 48412 320 48418 696
rect 48372 308 48418 320
rect 48490 696 48536 708
rect 48490 320 48496 696
rect 48530 320 48536 696
rect 48490 308 48536 320
rect 48608 696 48654 708
rect 48608 320 48614 696
rect 48648 320 48654 696
rect 48608 308 48654 320
rect 48726 696 48772 708
rect 48726 320 48732 696
rect 48766 320 48772 696
rect 49132 696 49178 708
rect 49132 520 49138 696
rect 49172 520 49178 696
rect 49132 508 49178 520
rect 49250 696 49296 708
rect 49250 520 49256 696
rect 49290 520 49296 696
rect 49250 508 49296 520
rect 48726 308 48772 320
rect 48614 214 48648 308
rect 49138 214 49171 508
rect 47957 182 49171 214
rect 45177 158 45318 164
rect 44855 121 45069 145
rect 44815 109 45069 121
rect 43827 105 44412 107
rect 44821 105 45069 109
rect 43827 77 44457 105
rect 43827 71 44694 77
rect 43827 37 44644 71
rect 44678 37 44694 71
rect 43827 21 44694 37
rect 44746 71 44812 77
rect 44746 37 44762 71
rect 44796 37 44812 71
rect 44995 61 45069 105
rect 45306 91 45318 158
rect 46552 97 46684 182
rect 48450 97 48582 182
rect 45177 85 45318 91
rect 45069 51 45177 61
rect 43827 5 44457 21
rect 43827 1 44412 5
rect 43827 0 43928 1
rect 44357 -48 44457 -37
rect 44321 -154 44331 -48
rect 44443 -59 44457 -48
rect 44746 -59 44812 37
rect 46542 -11 46552 97
rect 46684 -11 46694 97
rect 48440 -11 48450 97
rect 48582 -11 48592 97
rect 49371 69 49438 1452
rect 44443 -107 44812 -59
rect 44443 -137 44457 -107
rect 44443 -154 44453 -137
rect 44745 -210 44811 -107
rect 46573 -151 46579 -11
rect 46646 -151 46652 -11
rect 46573 -163 46652 -151
rect 49371 -210 49437 69
rect 44743 -290 49437 -210
rect 48160 -788 48624 -756
rect 48712 -772 48722 -712
rect 48784 -772 48794 -712
rect 48160 -796 48623 -788
rect 48160 -945 48214 -796
rect 42597 -1293 43326 -1213
rect 42347 -1306 43326 -1293
rect 42307 -1318 43326 -1306
rect 41842 -1431 41876 -1318
rect 42312 -1322 43326 -1318
rect 47840 -1045 48214 -945
rect 48274 -841 48505 -825
rect 48274 -875 48455 -841
rect 48489 -875 48505 -841
rect 48274 -881 48505 -875
rect 48557 -841 48623 -796
rect 48557 -875 48573 -841
rect 48607 -875 48623 -841
rect 48557 -881 48623 -875
rect 42238 -1356 42304 -1349
rect 42238 -1390 42254 -1356
rect 42288 -1390 42304 -1356
rect 42238 -1431 42304 -1390
rect 41722 -1432 42304 -1431
rect 41722 -1461 42422 -1432
rect 41722 -1555 41758 -1461
rect 41958 -1555 41994 -1461
rect 42194 -1462 42422 -1461
rect 42194 -1555 42230 -1462
rect 42356 -1473 42422 -1462
rect 42356 -1507 42372 -1473
rect 42406 -1507 42422 -1473
rect 42356 -1514 42422 -1507
rect 42666 -1555 42701 -1322
rect 41599 -1567 41645 -1555
rect 41599 -1743 41605 -1567
rect 41639 -1743 41645 -1567
rect 41599 -1755 41645 -1743
rect 41717 -1567 41763 -1555
rect 41717 -1743 41723 -1567
rect 41757 -1743 41763 -1567
rect 41717 -1755 41763 -1743
rect 41835 -1567 41881 -1555
rect 41835 -1743 41841 -1567
rect 41875 -1743 41881 -1567
rect 41835 -1755 41881 -1743
rect 41953 -1567 41999 -1555
rect 41953 -1743 41959 -1567
rect 41993 -1743 41999 -1567
rect 41953 -1755 41999 -1743
rect 42071 -1567 42117 -1555
rect 42071 -1743 42077 -1567
rect 42111 -1743 42117 -1567
rect 42071 -1755 42117 -1743
rect 42189 -1567 42235 -1555
rect 42189 -1743 42195 -1567
rect 42229 -1743 42235 -1567
rect 42189 -1755 42235 -1743
rect 42307 -1567 42353 -1555
rect 42307 -1743 42313 -1567
rect 42347 -1743 42353 -1567
rect 42307 -1755 42353 -1743
rect 42425 -1567 42471 -1555
rect 42425 -1743 42431 -1567
rect 42465 -1743 42471 -1567
rect 42425 -1755 42471 -1743
rect 42543 -1567 42589 -1555
rect 42543 -1743 42549 -1567
rect 42583 -1743 42589 -1567
rect 42543 -1755 42589 -1743
rect 42661 -1567 42707 -1555
rect 42661 -1743 42667 -1567
rect 42701 -1743 42707 -1567
rect 42661 -1755 42707 -1743
rect 41606 -1861 41638 -1755
rect 41842 -1861 41874 -1755
rect 42078 -1861 42110 -1755
rect 42314 -1861 42346 -1755
rect 42549 -1861 42583 -1755
rect 41606 -1891 42583 -1861
rect 41910 -1919 42046 -1891
rect 41910 -1981 41946 -1919
rect 42006 -1981 42046 -1919
rect 41910 -2001 42046 -1981
rect 34530 -2060 35303 -2059
rect 47840 -2060 47963 -1045
rect 48274 -1074 48328 -881
rect 48716 -909 48792 -772
rect 48632 -913 48792 -909
rect 34530 -2159 47963 -2060
rect 48001 -1173 48328 -1074
rect 48390 -925 48436 -913
rect 34629 -2160 47564 -2159
rect 30643 -2210 31043 -2204
rect 30481 -2244 30655 -2210
rect 31031 -2244 31043 -2210
rect 29950 -2267 30350 -2261
rect 29804 -2301 29962 -2267
rect 30338 -2301 30350 -2267
rect 29804 -2503 29847 -2301
rect 29950 -2307 30350 -2301
rect 29950 -2385 30350 -2379
rect 29950 -2419 29962 -2385
rect 30338 -2419 30350 -2385
rect 29950 -2425 30350 -2419
rect 30481 -2446 30519 -2244
rect 30643 -2250 31043 -2244
rect 30643 -2328 31043 -2322
rect 30643 -2362 30655 -2328
rect 31031 -2362 31043 -2328
rect 30643 -2368 31043 -2362
rect 31208 -2416 31259 -2399
rect 30643 -2446 31043 -2440
rect 30481 -2480 30655 -2446
rect 31031 -2480 31043 -2446
rect 31208 -2450 31219 -2416
rect 31253 -2450 31259 -2416
rect 31208 -2466 31259 -2450
rect 30643 -2486 31043 -2480
rect 29950 -2503 30350 -2497
rect 29804 -2537 29962 -2503
rect 30338 -2537 30350 -2503
rect 29804 -2868 29847 -2537
rect 29950 -2543 30350 -2537
rect 30162 -2626 30338 -2543
rect 31203 -2579 31246 -2466
rect 30150 -2632 30350 -2626
rect 30150 -2666 30162 -2632
rect 30338 -2666 30350 -2632
rect 30150 -2672 30350 -2666
rect 30501 -2718 30567 -2706
rect 30150 -2750 30350 -2744
rect 30150 -2784 30162 -2750
rect 30338 -2784 30419 -2750
rect 30501 -2772 30507 -2718
rect 30561 -2772 30567 -2718
rect 30501 -2784 30567 -2772
rect 30150 -2790 30350 -2784
rect 30384 -2852 30419 -2784
rect 31202 -2852 31247 -2579
rect 31287 -2690 31336 -2203
rect 31375 -2210 31775 -2204
rect 31869 -2210 31901 -2178
rect 33763 -2184 33888 -2178
rect 31375 -2244 31387 -2210
rect 31763 -2244 31901 -2210
rect 31375 -2250 31775 -2244
rect 31375 -2328 31775 -2322
rect 31375 -2362 31387 -2328
rect 31763 -2362 31775 -2328
rect 31375 -2368 31775 -2362
rect 31275 -2706 31337 -2690
rect 31275 -2740 31287 -2706
rect 31321 -2740 31337 -2706
rect 31275 -2746 31337 -2740
rect 31375 -2734 31575 -2728
rect 31869 -2734 31901 -2244
rect 33761 -2189 33888 -2184
rect 48001 -2189 48106 -1173
rect 48390 -1301 48396 -925
rect 48430 -1301 48436 -925
rect 48390 -1313 48436 -1301
rect 48508 -925 48554 -913
rect 48508 -1301 48514 -925
rect 48548 -1301 48554 -925
rect 48508 -1313 48554 -1301
rect 48626 -925 48792 -913
rect 48626 -1301 48632 -925
rect 48666 -952 48792 -925
rect 48666 -1301 48672 -952
rect 48749 -1113 48792 -952
rect 48626 -1313 48672 -1301
rect 48743 -1118 48792 -1113
rect 48743 -1125 48789 -1118
rect 48743 -1301 48749 -1125
rect 48783 -1301 48789 -1125
rect 48743 -1313 48789 -1301
rect 48861 -1125 48907 -1113
rect 48861 -1301 48867 -1125
rect 48901 -1288 48907 -1125
rect 49778 -1208 49914 2725
rect 50482 1361 50575 3255
rect 50638 3196 51104 3218
rect 51392 3196 51458 3292
rect 53223 3302 53229 3478
rect 53263 3302 53269 3478
rect 53223 3290 53269 3302
rect 53341 3478 53387 3490
rect 53341 3302 53347 3478
rect 53381 3302 53387 3478
rect 53341 3290 53387 3302
rect 53459 3478 53505 3490
rect 53459 3302 53465 3478
rect 53499 3302 53505 3478
rect 53459 3290 53505 3302
rect 53577 3478 53623 3490
rect 53577 3302 53583 3478
rect 53617 3423 53623 3478
rect 53742 3478 53788 3490
rect 53742 3423 53748 3478
rect 53617 3335 53748 3423
rect 53617 3302 53623 3335
rect 53577 3290 53623 3302
rect 53742 3302 53748 3335
rect 53782 3302 53788 3478
rect 53742 3290 53788 3302
rect 53860 3478 53906 3490
rect 53860 3302 53866 3478
rect 53900 3302 53906 3478
rect 53860 3290 53906 3302
rect 53978 3478 54024 3490
rect 53978 3302 53984 3478
rect 54018 3302 54024 3478
rect 53978 3290 54024 3302
rect 54096 3478 54142 3490
rect 54096 3302 54102 3478
rect 54136 3302 54142 3478
rect 54096 3290 54142 3302
rect 53229 3251 53263 3290
rect 53465 3251 53499 3290
rect 53229 3216 53499 3251
rect 53866 3252 53899 3290
rect 54102 3252 54135 3290
rect 53866 3216 54135 3252
rect 50638 3148 51458 3196
rect 53263 3215 53499 3216
rect 50638 3117 51104 3148
rect 53263 3141 53395 3215
rect 50638 2861 50743 3117
rect 53253 3033 53263 3141
rect 53395 3033 53405 3141
rect 51479 2954 51558 2966
rect 50638 2755 50701 2861
rect 50813 2755 50823 2861
rect 51479 2857 51485 2954
rect 51405 2837 51485 2857
rect 51552 2857 51558 2954
rect 53283 2900 53289 3033
rect 53356 2900 53362 3033
rect 53283 2888 53362 2900
rect 51552 2837 51625 2857
rect 50638 2744 50787 2755
rect 50638 1567 50743 2744
rect 51405 2729 51449 2837
rect 51581 2729 51625 2837
rect 51405 2687 51625 2729
rect 54203 2702 54265 4273
rect 54455 4265 54501 4277
rect 54455 3889 54461 4265
rect 54495 3889 54501 4265
rect 54455 3877 54501 3889
rect 54573 4265 54619 4277
rect 54573 3889 54579 4265
rect 54613 3889 54619 4265
rect 54573 3877 54619 3889
rect 54691 4265 54737 4277
rect 54691 3889 54697 4265
rect 54731 3889 54737 4265
rect 54691 3877 54737 3889
rect 54809 4265 54855 4277
rect 54809 3889 54815 4265
rect 54849 3889 54855 4265
rect 54809 3877 54855 3889
rect 54927 4265 54973 4277
rect 54927 3889 54933 4265
rect 54967 3889 54973 4265
rect 54927 3877 54973 3889
rect 55045 4265 55091 4277
rect 55045 3889 55051 4265
rect 55085 3889 55091 4265
rect 55045 3877 55091 3889
rect 55163 4265 55209 4277
rect 55163 3889 55169 4265
rect 55203 3889 55209 4265
rect 55163 3877 55209 3889
rect 54461 3835 54495 3877
rect 54697 3835 54731 3877
rect 54461 3807 54731 3835
rect 54815 3836 54849 3877
rect 55051 3836 55085 3877
rect 54815 3807 55085 3836
rect 54461 3759 54495 3807
rect 54461 3729 54524 3759
rect 54489 3637 54524 3729
rect 54996 3699 55096 3720
rect 54996 3645 55010 3699
rect 55075 3645 55096 3699
rect 54996 3640 55096 3645
rect 55169 3694 55203 3877
rect 56384 3846 56536 8030
rect 57112 7230 57205 9124
rect 57268 9065 57734 9087
rect 58022 9065 58088 9161
rect 59853 9171 59859 9347
rect 59893 9171 59899 9347
rect 59853 9159 59899 9171
rect 59971 9347 60017 9359
rect 59971 9171 59977 9347
rect 60011 9171 60017 9347
rect 59971 9159 60017 9171
rect 60089 9347 60135 9359
rect 60089 9171 60095 9347
rect 60129 9171 60135 9347
rect 60089 9159 60135 9171
rect 60207 9347 60253 9359
rect 60207 9171 60213 9347
rect 60247 9292 60253 9347
rect 60372 9347 60418 9359
rect 60372 9292 60378 9347
rect 60247 9204 60378 9292
rect 60247 9171 60253 9204
rect 60207 9159 60253 9171
rect 60372 9171 60378 9204
rect 60412 9171 60418 9347
rect 60372 9159 60418 9171
rect 60490 9347 60536 9359
rect 60490 9171 60496 9347
rect 60530 9171 60536 9347
rect 60490 9159 60536 9171
rect 60608 9347 60654 9359
rect 60608 9171 60614 9347
rect 60648 9171 60654 9347
rect 60608 9159 60654 9171
rect 60726 9347 60772 9359
rect 60726 9171 60732 9347
rect 60766 9171 60772 9347
rect 60726 9159 60772 9171
rect 59859 9120 59893 9159
rect 60095 9120 60129 9159
rect 59859 9085 60129 9120
rect 60496 9121 60529 9159
rect 60732 9121 60765 9159
rect 60496 9085 60765 9121
rect 57268 9017 58088 9065
rect 59893 9084 60129 9085
rect 57268 8986 57734 9017
rect 59893 9010 60025 9084
rect 57268 8730 57373 8986
rect 59883 8902 59893 9010
rect 60025 8902 60035 9010
rect 58110 8821 58189 8833
rect 57268 8624 57331 8730
rect 57443 8624 57453 8730
rect 58110 8726 58116 8821
rect 58035 8706 58116 8726
rect 58183 8726 58189 8821
rect 59911 8759 59917 8902
rect 59984 8759 59990 8902
rect 59911 8747 59990 8759
rect 58183 8706 58255 8726
rect 57268 8613 57417 8624
rect 57268 7436 57373 8613
rect 58035 8598 58079 8706
rect 58211 8598 58255 8706
rect 58035 8556 58255 8598
rect 60833 8571 60895 10142
rect 61085 10134 61131 10146
rect 61085 9758 61091 10134
rect 61125 9758 61131 10134
rect 61085 9746 61131 9758
rect 61203 10134 61249 10146
rect 61203 9758 61209 10134
rect 61243 9758 61249 10134
rect 61203 9746 61249 9758
rect 61321 10134 61367 10146
rect 61321 9758 61327 10134
rect 61361 9758 61367 10134
rect 61321 9746 61367 9758
rect 61439 10134 61485 10146
rect 61439 9758 61445 10134
rect 61479 9758 61485 10134
rect 61439 9746 61485 9758
rect 61557 10134 61603 10146
rect 61557 9758 61563 10134
rect 61597 9758 61603 10134
rect 61557 9746 61603 9758
rect 61675 10134 61721 10146
rect 61675 9758 61681 10134
rect 61715 9758 61721 10134
rect 61675 9746 61721 9758
rect 61793 10134 61839 10146
rect 61793 9758 61799 10134
rect 61833 9758 61839 10134
rect 61793 9746 61839 9758
rect 61091 9704 61125 9746
rect 61327 9704 61361 9746
rect 61091 9676 61361 9704
rect 61445 9705 61479 9746
rect 61681 9705 61715 9746
rect 61445 9676 61715 9705
rect 61091 9628 61125 9676
rect 61091 9598 61154 9628
rect 61119 9506 61154 9598
rect 61626 9568 61726 9589
rect 61626 9514 61640 9568
rect 61705 9514 61726 9568
rect 61626 9509 61726 9514
rect 61799 9563 61833 9746
rect 61799 9509 61908 9563
rect 61119 9470 61346 9506
rect 61119 9363 61154 9470
rect 61280 9436 61346 9470
rect 61280 9402 61296 9436
rect 61330 9402 61346 9436
rect 61627 9494 61724 9509
rect 61627 9427 61684 9494
rect 61280 9396 61346 9402
rect 61521 9391 61790 9427
rect 61521 9363 61554 9391
rect 61757 9363 61790 9391
rect 61874 9363 61908 9509
rect 62608 9502 62618 9577
rect 62686 9502 62798 12445
rect 62635 9501 62798 9502
rect 62687 9491 62798 9501
rect 60995 9351 61041 9363
rect 60995 9175 61001 9351
rect 61035 9175 61041 9351
rect 60995 9163 61041 9175
rect 61113 9351 61159 9363
rect 61113 9175 61119 9351
rect 61153 9175 61159 9351
rect 61113 9163 61159 9175
rect 61231 9351 61277 9363
rect 61231 9175 61237 9351
rect 61271 9175 61277 9351
rect 61231 9163 61277 9175
rect 61349 9351 61395 9363
rect 61349 9175 61355 9351
rect 61389 9296 61395 9351
rect 61514 9351 61560 9363
rect 61514 9296 61520 9351
rect 61389 9208 61520 9296
rect 61389 9175 61395 9208
rect 61349 9163 61395 9175
rect 61514 9175 61520 9208
rect 61554 9175 61560 9351
rect 61514 9163 61560 9175
rect 61632 9351 61678 9363
rect 61632 9175 61638 9351
rect 61672 9175 61678 9351
rect 61632 9163 61678 9175
rect 61750 9351 61796 9363
rect 61750 9175 61756 9351
rect 61790 9175 61796 9351
rect 61750 9163 61796 9175
rect 61868 9351 61914 9363
rect 61868 9175 61874 9351
rect 61908 9175 61914 9351
rect 61868 9163 61914 9175
rect 61001 9124 61035 9163
rect 61237 9124 61271 9163
rect 61001 9088 61271 9124
rect 61638 9125 61671 9163
rect 61874 9125 61907 9163
rect 61638 9089 61907 9125
rect 61001 9087 61167 9088
rect 61035 9008 61167 9087
rect 61025 8900 61035 9008
rect 61167 8900 61177 9008
rect 61054 8761 61060 8900
rect 61127 8761 61133 8900
rect 61054 8749 61133 8761
rect 57639 8526 58616 8556
rect 60833 8554 60896 8571
rect 60758 8550 60896 8554
rect 57639 8420 57671 8526
rect 57875 8420 57907 8526
rect 58111 8420 58143 8526
rect 58347 8420 58379 8526
rect 58582 8420 58616 8526
rect 58926 8516 60896 8550
rect 58924 8487 60896 8516
rect 58924 8471 58970 8487
rect 60758 8485 60896 8487
rect 57632 8408 57678 8420
rect 57632 8232 57638 8408
rect 57672 8232 57678 8408
rect 57632 8220 57678 8232
rect 57750 8408 57796 8420
rect 57750 8232 57756 8408
rect 57790 8232 57796 8408
rect 57750 8220 57796 8232
rect 57868 8408 57914 8420
rect 57868 8232 57874 8408
rect 57908 8232 57914 8408
rect 57868 8220 57914 8232
rect 57986 8408 58032 8420
rect 57986 8232 57992 8408
rect 58026 8232 58032 8408
rect 57986 8220 58032 8232
rect 58104 8408 58150 8420
rect 58104 8232 58110 8408
rect 58144 8232 58150 8408
rect 58104 8220 58150 8232
rect 58222 8408 58268 8420
rect 58222 8232 58228 8408
rect 58262 8232 58268 8408
rect 58222 8220 58268 8232
rect 58340 8408 58386 8420
rect 58340 8232 58346 8408
rect 58380 8232 58386 8408
rect 58340 8220 58386 8232
rect 58458 8408 58504 8420
rect 58458 8232 58464 8408
rect 58498 8232 58504 8408
rect 58458 8220 58504 8232
rect 58576 8408 58622 8420
rect 58576 8232 58582 8408
rect 58616 8232 58622 8408
rect 58576 8220 58622 8232
rect 58694 8408 58740 8420
rect 58694 8232 58700 8408
rect 58734 8232 58740 8408
rect 58694 8220 58740 8232
rect 57755 8126 57791 8220
rect 57991 8126 58027 8220
rect 58227 8127 58263 8220
rect 58389 8172 58455 8179
rect 58389 8138 58405 8172
rect 58439 8138 58455 8172
rect 58389 8127 58455 8138
rect 58227 8126 58455 8127
rect 57755 8097 58455 8126
rect 57755 8096 58337 8097
rect 57875 7983 57909 8096
rect 58271 8055 58337 8096
rect 58271 8021 58287 8055
rect 58321 8021 58337 8055
rect 58271 8014 58337 8021
rect 58699 8002 58734 8220
rect 58923 8019 58970 8471
rect 61817 8476 61896 8488
rect 61817 8363 61823 8476
rect 61890 8363 61896 8476
rect 59882 8255 59892 8363
rect 60024 8255 60034 8363
rect 61780 8255 61790 8363
rect 61922 8255 61932 8363
rect 59892 8215 60024 8255
rect 61790 8215 61922 8255
rect 59891 8149 60024 8215
rect 61789 8149 61922 8215
rect 59220 8106 60693 8149
rect 58923 8003 58969 8019
rect 58888 8002 58969 8003
rect 58699 7987 58969 8002
rect 58345 7983 58969 7987
rect 57869 7971 57915 7983
rect 57604 7493 57614 7611
rect 57732 7579 57742 7611
rect 57869 7595 57875 7971
rect 57909 7595 57915 7971
rect 57869 7583 57915 7595
rect 57987 7971 58033 7983
rect 57987 7595 57993 7971
rect 58027 7595 58033 7971
rect 57987 7583 58033 7595
rect 58105 7971 58151 7983
rect 58105 7595 58111 7971
rect 58145 7619 58151 7971
rect 58222 7971 58268 7983
rect 58222 7795 58228 7971
rect 58262 7795 58268 7971
rect 58222 7783 58268 7795
rect 58340 7971 58969 7983
rect 58340 7795 58346 7971
rect 58380 7959 58969 7971
rect 58380 7958 58622 7959
rect 58380 7795 58386 7958
rect 58888 7957 58969 7959
rect 59220 7803 59254 8106
rect 59586 8003 59620 8106
rect 59822 8003 59856 8106
rect 60058 8003 60092 8106
rect 60294 8003 60328 8106
rect 59580 7991 59626 8003
rect 58340 7783 58386 7795
rect 59096 7791 59142 7803
rect 58228 7667 58263 7783
rect 58359 7667 58467 7677
rect 58228 7619 58359 7667
rect 58467 7627 58606 7633
rect 58145 7595 58359 7619
rect 58105 7583 58359 7595
rect 58111 7579 58359 7583
rect 57732 7551 57747 7579
rect 57732 7545 57984 7551
rect 57732 7511 57934 7545
rect 57968 7511 57984 7545
rect 57732 7495 57984 7511
rect 58036 7545 58102 7551
rect 58036 7511 58052 7545
rect 58086 7511 58102 7545
rect 58285 7535 58359 7579
rect 58594 7560 58606 7627
rect 59096 7615 59102 7791
rect 59136 7615 59142 7791
rect 59096 7603 59142 7615
rect 59214 7791 59260 7803
rect 59214 7615 59220 7791
rect 59254 7615 59260 7791
rect 59214 7603 59260 7615
rect 59332 7791 59378 7803
rect 59332 7615 59338 7791
rect 59372 7615 59378 7791
rect 59332 7603 59378 7615
rect 59450 7791 59496 7803
rect 59580 7791 59586 7991
rect 59450 7615 59456 7791
rect 59490 7615 59586 7791
rect 59620 7615 59626 7991
rect 59450 7603 59496 7615
rect 59580 7603 59626 7615
rect 59698 7991 59744 8003
rect 59698 7615 59704 7991
rect 59738 7615 59744 7991
rect 59698 7603 59744 7615
rect 59816 7991 59862 8003
rect 59816 7615 59822 7991
rect 59856 7615 59862 7991
rect 59816 7603 59862 7615
rect 59934 7991 59980 8003
rect 59934 7615 59940 7991
rect 59974 7615 59980 7991
rect 59934 7603 59980 7615
rect 60052 7991 60098 8003
rect 60052 7615 60058 7991
rect 60092 7615 60098 7991
rect 60052 7603 60098 7615
rect 60170 7991 60216 8003
rect 60170 7615 60176 7991
rect 60210 7615 60216 7991
rect 60170 7603 60216 7615
rect 60288 7991 60334 8003
rect 60288 7615 60294 7991
rect 60328 7791 60334 7991
rect 60659 7803 60693 8106
rect 61118 8106 62591 8149
rect 61118 7803 61152 8106
rect 61484 8003 61518 8106
rect 61720 8003 61754 8106
rect 61956 8003 61990 8106
rect 62192 8003 62226 8106
rect 61478 7991 61524 8003
rect 60417 7791 60463 7803
rect 60328 7615 60423 7791
rect 60457 7615 60463 7791
rect 60288 7603 60334 7615
rect 60417 7603 60463 7615
rect 60535 7791 60581 7803
rect 60535 7615 60541 7791
rect 60575 7615 60581 7791
rect 60535 7603 60581 7615
rect 60653 7791 60699 7803
rect 60653 7615 60659 7791
rect 60693 7615 60699 7791
rect 60653 7603 60699 7615
rect 60771 7791 60817 7803
rect 60771 7615 60777 7791
rect 60811 7615 60817 7791
rect 60771 7603 60817 7615
rect 60994 7791 61040 7803
rect 60994 7615 61000 7791
rect 61034 7615 61040 7791
rect 60994 7603 61040 7615
rect 61112 7791 61158 7803
rect 61112 7615 61118 7791
rect 61152 7615 61158 7791
rect 61112 7603 61158 7615
rect 61230 7791 61276 7803
rect 61230 7615 61236 7791
rect 61270 7615 61276 7791
rect 61230 7603 61276 7615
rect 61348 7791 61394 7803
rect 61478 7791 61484 7991
rect 61348 7615 61354 7791
rect 61388 7615 61484 7791
rect 61518 7615 61524 7991
rect 61348 7603 61394 7615
rect 61478 7603 61524 7615
rect 61596 7991 61642 8003
rect 61596 7615 61602 7991
rect 61636 7615 61642 7991
rect 61596 7603 61642 7615
rect 61714 7991 61760 8003
rect 61714 7615 61720 7991
rect 61754 7615 61760 7991
rect 61714 7603 61760 7615
rect 61832 7991 61878 8003
rect 61832 7615 61838 7991
rect 61872 7615 61878 7991
rect 61832 7603 61878 7615
rect 61950 7991 61996 8003
rect 61950 7615 61956 7991
rect 61990 7615 61996 7991
rect 61950 7603 61996 7615
rect 62068 7991 62114 8003
rect 62068 7615 62074 7991
rect 62108 7615 62114 7991
rect 62068 7603 62114 7615
rect 62186 7991 62232 8003
rect 62186 7615 62192 7991
rect 62226 7791 62232 7991
rect 62557 7803 62591 8106
rect 62315 7791 62361 7803
rect 62226 7615 62321 7791
rect 62355 7615 62361 7791
rect 62186 7603 62232 7615
rect 62315 7603 62361 7615
rect 62433 7791 62479 7803
rect 62433 7615 62439 7791
rect 62473 7615 62479 7791
rect 62433 7603 62479 7615
rect 62551 7791 62597 7803
rect 62551 7615 62557 7791
rect 62591 7615 62597 7791
rect 62551 7603 62597 7615
rect 62669 7791 62715 7803
rect 62669 7615 62675 7791
rect 62709 7615 62715 7791
rect 62669 7603 62715 7615
rect 58467 7554 58606 7560
rect 59102 7569 59136 7603
rect 59704 7569 59738 7603
rect 59940 7569 59974 7603
rect 58359 7525 58467 7535
rect 59102 7534 59261 7569
rect 59704 7534 59974 7569
rect 60541 7569 60575 7603
rect 60777 7569 60811 7603
rect 60541 7534 60811 7569
rect 61000 7569 61034 7603
rect 61602 7569 61636 7603
rect 61838 7569 61872 7603
rect 61000 7534 61159 7569
rect 61602 7534 61872 7569
rect 62439 7569 62473 7603
rect 62675 7569 62709 7603
rect 62439 7534 62709 7569
rect 57732 7493 57747 7495
rect 57647 7479 57747 7493
rect 57647 7436 57747 7437
rect 57268 7415 57747 7436
rect 58036 7415 58102 7511
rect 57268 7367 58102 7415
rect 57268 7338 57747 7367
rect 57268 7336 57373 7338
rect 57647 7337 57747 7338
rect 57101 7151 57111 7230
rect 57204 7151 57214 7230
rect 58102 7213 58181 7225
rect 56626 6824 56734 6836
rect 56622 6724 56632 6824
rect 56728 6724 56738 6824
rect 56626 6712 56734 6724
rect 57112 5977 57205 7151
rect 58102 7122 58108 7213
rect 58030 7102 58108 7122
rect 58175 7122 58181 7213
rect 58175 7102 58250 7122
rect 58030 6994 58074 7102
rect 58206 6994 58250 7102
rect 58030 6952 58250 6994
rect 57634 6922 58611 6952
rect 57634 6816 57666 6922
rect 57870 6816 57902 6922
rect 58106 6816 58138 6922
rect 58342 6816 58374 6922
rect 58577 6816 58611 6922
rect 57627 6804 57673 6816
rect 57627 6628 57633 6804
rect 57667 6628 57673 6804
rect 57627 6616 57673 6628
rect 57745 6804 57791 6816
rect 57745 6628 57751 6804
rect 57785 6628 57791 6804
rect 57745 6616 57791 6628
rect 57863 6804 57909 6816
rect 57863 6628 57869 6804
rect 57903 6628 57909 6804
rect 57863 6616 57909 6628
rect 57981 6804 58027 6816
rect 57981 6628 57987 6804
rect 58021 6628 58027 6804
rect 57981 6616 58027 6628
rect 58099 6804 58145 6816
rect 58099 6628 58105 6804
rect 58139 6628 58145 6804
rect 58099 6616 58145 6628
rect 58217 6804 58263 6816
rect 58217 6628 58223 6804
rect 58257 6628 58263 6804
rect 58217 6616 58263 6628
rect 58335 6804 58381 6816
rect 58335 6628 58341 6804
rect 58375 6628 58381 6804
rect 58335 6616 58381 6628
rect 58453 6804 58499 6816
rect 58453 6628 58459 6804
rect 58493 6628 58499 6804
rect 58453 6616 58499 6628
rect 58571 6804 58617 6816
rect 58571 6628 58577 6804
rect 58611 6628 58617 6804
rect 58571 6616 58617 6628
rect 58689 6804 58735 6816
rect 58689 6628 58695 6804
rect 58729 6628 58735 6804
rect 58689 6616 58735 6628
rect 59227 6750 59261 7534
rect 59940 7472 59974 7534
rect 59529 7434 60271 7472
rect 59529 7310 59563 7434
rect 59765 7310 59799 7434
rect 60001 7310 60035 7434
rect 60237 7310 60271 7434
rect 60527 7327 60537 7393
rect 60600 7327 60610 7393
rect 59523 7298 59569 7310
rect 59523 6922 59529 7298
rect 59563 6922 59569 7298
rect 59523 6910 59569 6922
rect 59641 7298 59687 7310
rect 59641 6922 59647 7298
rect 59681 6922 59687 7298
rect 59641 6910 59687 6922
rect 59759 7298 59805 7310
rect 59759 6922 59765 7298
rect 59799 6922 59805 7298
rect 59759 6910 59805 6922
rect 59877 7298 59923 7310
rect 59877 6922 59883 7298
rect 59917 6922 59923 7298
rect 59877 6910 59923 6922
rect 59995 7298 60041 7310
rect 59995 6922 60001 7298
rect 60035 6922 60041 7298
rect 59995 6910 60041 6922
rect 60113 7298 60159 7310
rect 60113 6922 60119 7298
rect 60153 6922 60159 7298
rect 60113 6910 60159 6922
rect 60231 7298 60277 7310
rect 60231 6922 60237 7298
rect 60271 6922 60277 7298
rect 60231 6910 60277 6922
rect 60643 6751 60677 7534
rect 60370 6750 60677 6751
rect 59227 6745 59543 6750
rect 60257 6745 60677 6750
rect 59227 6734 59610 6745
rect 59227 6707 59559 6734
rect 57750 6522 57786 6616
rect 57986 6522 58022 6616
rect 58222 6523 58258 6616
rect 58384 6568 58450 6575
rect 58384 6534 58400 6568
rect 58434 6534 58450 6568
rect 58384 6523 58450 6534
rect 58222 6522 58450 6523
rect 57750 6493 58450 6522
rect 57750 6492 58332 6493
rect 57870 6379 57904 6492
rect 58266 6451 58332 6492
rect 58266 6417 58282 6451
rect 58316 6417 58332 6451
rect 58266 6410 58332 6417
rect 58694 6383 58729 6616
rect 59227 6578 59261 6707
rect 59543 6700 59559 6707
rect 59593 6700 59610 6734
rect 59543 6694 59610 6700
rect 60190 6734 60677 6745
rect 60190 6700 60207 6734
rect 60241 6707 60677 6734
rect 60241 6700 60257 6707
rect 60370 6706 60677 6707
rect 60190 6694 60257 6700
rect 59368 6667 59424 6679
rect 59368 6633 59374 6667
rect 59408 6666 59424 6667
rect 60481 6666 60537 6678
rect 59408 6650 59875 6666
rect 59408 6633 59825 6650
rect 59368 6617 59825 6633
rect 59809 6616 59825 6617
rect 59859 6616 59875 6650
rect 59809 6609 59875 6616
rect 59927 6651 60497 6666
rect 59927 6617 59943 6651
rect 59977 6632 60497 6651
rect 60531 6632 60537 6666
rect 59977 6617 60537 6632
rect 59927 6607 59994 6617
rect 60481 6616 60537 6617
rect 60643 6578 60677 6706
rect 61125 6750 61159 7534
rect 61838 7472 61872 7534
rect 61427 7434 62169 7472
rect 61427 7310 61461 7434
rect 61663 7310 61697 7434
rect 61899 7310 61933 7434
rect 62135 7310 62169 7434
rect 61421 7298 61467 7310
rect 61421 6922 61427 7298
rect 61461 6922 61467 7298
rect 61421 6910 61467 6922
rect 61539 7298 61585 7310
rect 61539 6922 61545 7298
rect 61579 6922 61585 7298
rect 61539 6910 61585 6922
rect 61657 7298 61703 7310
rect 61657 6922 61663 7298
rect 61697 6922 61703 7298
rect 61657 6910 61703 6922
rect 61775 7298 61821 7310
rect 61775 6922 61781 7298
rect 61815 6922 61821 7298
rect 61775 6910 61821 6922
rect 61893 7298 61939 7310
rect 61893 6922 61899 7298
rect 61933 6922 61939 7298
rect 61893 6910 61939 6922
rect 62011 7298 62057 7310
rect 62011 6922 62017 7298
rect 62051 6922 62057 7298
rect 62011 6910 62057 6922
rect 62129 7298 62175 7310
rect 62129 6922 62135 7298
rect 62169 6922 62175 7298
rect 62129 6910 62175 6922
rect 62541 6751 62575 7534
rect 62153 6750 62222 6751
rect 62268 6750 62575 6751
rect 61125 6745 61441 6750
rect 62153 6746 62575 6750
rect 61125 6734 61508 6745
rect 61125 6707 61457 6734
rect 61125 6578 61159 6707
rect 61441 6700 61457 6707
rect 61491 6700 61508 6734
rect 61441 6694 61508 6700
rect 62086 6735 62575 6746
rect 62086 6701 62103 6735
rect 62137 6707 62575 6735
rect 62137 6701 62153 6707
rect 62268 6706 62575 6707
rect 62086 6695 62153 6701
rect 61266 6667 61322 6679
rect 61266 6633 61272 6667
rect 61306 6666 61322 6667
rect 62379 6666 62435 6678
rect 61306 6650 61773 6666
rect 61306 6633 61723 6650
rect 61266 6617 61723 6633
rect 61707 6616 61723 6617
rect 61757 6616 61773 6650
rect 61707 6609 61773 6616
rect 61825 6651 62395 6666
rect 61825 6617 61841 6651
rect 61875 6632 62395 6651
rect 62429 6632 62435 6666
rect 61875 6617 62435 6632
rect 61825 6607 61892 6617
rect 62379 6616 62435 6617
rect 62541 6578 62575 6706
rect 62656 7356 62723 7380
rect 62656 7322 62673 7356
rect 62707 7322 62723 7356
rect 58340 6379 58729 6383
rect 57864 6367 57910 6379
rect 57864 5991 57870 6367
rect 57904 5991 57910 6367
rect 57864 5979 57910 5991
rect 57982 6367 58028 6379
rect 57982 5991 57988 6367
rect 58022 5991 58028 6367
rect 57982 5979 58028 5991
rect 58100 6367 58146 6379
rect 58100 5991 58106 6367
rect 58140 6015 58146 6367
rect 58217 6367 58263 6379
rect 58217 6191 58223 6367
rect 58257 6191 58263 6367
rect 58217 6179 58263 6191
rect 58335 6367 58729 6379
rect 59221 6566 59267 6578
rect 59221 6390 59227 6566
rect 59261 6390 59267 6566
rect 59221 6378 59267 6390
rect 59339 6566 59385 6578
rect 59339 6390 59345 6566
rect 59379 6390 59385 6566
rect 59339 6378 59385 6390
rect 59641 6566 59687 6578
rect 58335 6191 58341 6367
rect 58375 6354 58729 6367
rect 58375 6191 58381 6354
rect 58651 6351 58729 6354
rect 58651 6299 58661 6351
rect 58724 6299 58734 6351
rect 58656 6293 58729 6299
rect 58335 6179 58381 6191
rect 58223 6063 58258 6179
rect 59344 6084 59378 6378
rect 59641 6190 59647 6566
rect 59681 6190 59687 6566
rect 59641 6178 59687 6190
rect 59759 6566 59805 6578
rect 59759 6190 59765 6566
rect 59799 6190 59805 6566
rect 59759 6178 59805 6190
rect 59877 6566 59923 6578
rect 59877 6190 59883 6566
rect 59917 6190 59923 6566
rect 59877 6178 59923 6190
rect 59995 6566 60041 6578
rect 59995 6190 60001 6566
rect 60035 6190 60041 6566
rect 59995 6178 60041 6190
rect 60113 6566 60159 6578
rect 60113 6190 60119 6566
rect 60153 6190 60159 6566
rect 60519 6566 60565 6578
rect 60519 6390 60525 6566
rect 60559 6390 60565 6566
rect 60519 6378 60565 6390
rect 60637 6566 60683 6578
rect 60637 6390 60643 6566
rect 60677 6390 60683 6566
rect 60637 6378 60683 6390
rect 61119 6566 61165 6578
rect 61119 6390 61125 6566
rect 61159 6390 61165 6566
rect 61119 6378 61165 6390
rect 61237 6566 61283 6578
rect 61237 6390 61243 6566
rect 61277 6390 61283 6566
rect 61237 6378 61283 6390
rect 61539 6566 61585 6578
rect 60113 6178 60159 6190
rect 60001 6084 60035 6178
rect 60525 6084 60558 6378
rect 58354 6063 58462 6073
rect 58223 6015 58354 6063
rect 59344 6052 60558 6084
rect 61242 6084 61276 6378
rect 61539 6190 61545 6566
rect 61579 6190 61585 6566
rect 61539 6178 61585 6190
rect 61657 6566 61703 6578
rect 61657 6190 61663 6566
rect 61697 6190 61703 6566
rect 61657 6178 61703 6190
rect 61775 6566 61821 6578
rect 61775 6190 61781 6566
rect 61815 6190 61821 6566
rect 61775 6178 61821 6190
rect 61893 6566 61939 6578
rect 61893 6190 61899 6566
rect 61933 6190 61939 6566
rect 61893 6178 61939 6190
rect 62011 6566 62057 6578
rect 62011 6190 62017 6566
rect 62051 6190 62057 6566
rect 62417 6566 62463 6578
rect 62417 6390 62423 6566
rect 62457 6390 62463 6566
rect 62417 6378 62463 6390
rect 62535 6566 62581 6578
rect 62535 6390 62541 6566
rect 62575 6390 62581 6566
rect 62535 6378 62581 6390
rect 62011 6178 62057 6190
rect 61899 6084 61933 6178
rect 62423 6084 62456 6378
rect 61242 6052 62456 6084
rect 58462 6022 58612 6028
rect 58140 5991 58354 6015
rect 58100 5979 58354 5991
rect 57112 5975 57697 5977
rect 58106 5975 58354 5979
rect 57112 5947 57742 5975
rect 57112 5941 57979 5947
rect 57112 5907 57929 5941
rect 57963 5907 57979 5941
rect 57112 5891 57979 5907
rect 58031 5941 58097 5947
rect 58031 5907 58047 5941
rect 58081 5907 58097 5941
rect 58280 5931 58354 5975
rect 58600 5955 58612 6022
rect 59837 5967 59969 6052
rect 61735 5967 61867 6052
rect 58462 5949 58612 5955
rect 58354 5921 58462 5931
rect 57112 5875 57742 5891
rect 57112 5871 57697 5875
rect 57112 5870 57213 5871
rect 57642 5822 57742 5833
rect 57606 5716 57616 5822
rect 57728 5811 57742 5822
rect 58031 5811 58097 5907
rect 59827 5859 59837 5967
rect 59969 5859 59979 5967
rect 61725 5859 61735 5967
rect 61867 5859 61877 5967
rect 62656 5939 62723 7322
rect 62869 6899 62969 12503
rect 64603 12371 64698 12374
rect 64598 12365 64700 12371
rect 64598 12293 64610 12365
rect 64688 12293 64700 12365
rect 64598 12287 64700 12293
rect 65856 12323 66301 12329
rect 63731 12228 63867 12248
rect 63731 12166 63767 12228
rect 63827 12166 63867 12228
rect 63731 12138 63867 12166
rect 63427 12108 64404 12138
rect 63427 12002 63459 12108
rect 63663 12002 63695 12108
rect 63899 12002 63931 12108
rect 64135 12002 64167 12108
rect 64370 12002 64404 12108
rect 63420 11990 63466 12002
rect 63420 11814 63426 11990
rect 63460 11814 63466 11990
rect 63420 11802 63466 11814
rect 63538 11990 63584 12002
rect 63538 11814 63544 11990
rect 63578 11814 63584 11990
rect 63538 11802 63584 11814
rect 63656 11990 63702 12002
rect 63656 11814 63662 11990
rect 63696 11814 63702 11990
rect 63656 11802 63702 11814
rect 63774 11990 63820 12002
rect 63774 11814 63780 11990
rect 63814 11814 63820 11990
rect 63774 11802 63820 11814
rect 63892 11990 63938 12002
rect 63892 11814 63898 11990
rect 63932 11814 63938 11990
rect 63892 11802 63938 11814
rect 64010 11990 64056 12002
rect 64010 11814 64016 11990
rect 64050 11814 64056 11990
rect 64010 11802 64056 11814
rect 64128 11990 64174 12002
rect 64128 11814 64134 11990
rect 64168 11814 64174 11990
rect 64128 11802 64174 11814
rect 64246 11990 64292 12002
rect 64246 11814 64252 11990
rect 64286 11814 64292 11990
rect 64246 11802 64292 11814
rect 64364 11990 64410 12002
rect 64364 11814 64370 11990
rect 64404 11814 64410 11990
rect 64364 11802 64410 11814
rect 64482 11990 64528 12002
rect 64482 11814 64488 11990
rect 64522 11814 64528 11990
rect 64482 11802 64528 11814
rect 63543 11708 63579 11802
rect 63779 11708 63815 11802
rect 64015 11709 64051 11802
rect 64177 11754 64243 11761
rect 64177 11720 64193 11754
rect 64227 11720 64243 11754
rect 64177 11709 64243 11720
rect 64015 11708 64243 11709
rect 63543 11679 64243 11708
rect 63543 11678 64125 11679
rect 63663 11565 63697 11678
rect 64059 11637 64125 11678
rect 64059 11603 64075 11637
rect 64109 11603 64125 11637
rect 64059 11596 64125 11603
rect 64487 11570 64522 11802
rect 64603 11570 64698 12287
rect 65856 12123 65868 12323
rect 66289 12123 66301 12323
rect 65856 12117 66024 12123
rect 66014 12049 66024 12117
rect 66156 12117 66301 12123
rect 66156 12049 66166 12117
rect 66024 12009 66156 12049
rect 66023 11943 66156 12009
rect 65352 11900 66825 11943
rect 65352 11597 65386 11900
rect 65718 11797 65752 11900
rect 65954 11797 65988 11900
rect 66190 11797 66224 11900
rect 66426 11797 66460 11900
rect 65712 11785 65758 11797
rect 64432 11569 64698 11570
rect 64133 11565 64698 11569
rect 63657 11553 63703 11565
rect 63657 11177 63663 11553
rect 63697 11177 63703 11553
rect 63657 11165 63703 11177
rect 63775 11553 63821 11565
rect 63775 11177 63781 11553
rect 63815 11177 63821 11553
rect 63775 11165 63821 11177
rect 63893 11553 63939 11565
rect 63893 11177 63899 11553
rect 63933 11204 63939 11553
rect 64010 11553 64056 11565
rect 64010 11377 64016 11553
rect 64050 11377 64056 11553
rect 64010 11370 64056 11377
rect 64128 11553 64698 11565
rect 64128 11377 64134 11553
rect 64168 11540 64698 11553
rect 64168 11377 64174 11540
rect 64418 11460 64698 11540
rect 64432 11459 64698 11460
rect 65228 11585 65274 11597
rect 65228 11409 65234 11585
rect 65268 11409 65274 11585
rect 65228 11397 65274 11409
rect 65346 11585 65392 11597
rect 65346 11409 65352 11585
rect 65386 11409 65392 11585
rect 65346 11397 65392 11409
rect 65464 11585 65510 11597
rect 65464 11409 65470 11585
rect 65504 11409 65510 11585
rect 65464 11397 65510 11409
rect 65582 11585 65628 11597
rect 65712 11585 65718 11785
rect 65582 11409 65588 11585
rect 65622 11409 65718 11585
rect 65752 11409 65758 11785
rect 65582 11397 65628 11409
rect 65712 11397 65758 11409
rect 65830 11785 65876 11797
rect 65830 11409 65836 11785
rect 65870 11409 65876 11785
rect 65830 11397 65876 11409
rect 65948 11785 65994 11797
rect 65948 11409 65954 11785
rect 65988 11409 65994 11785
rect 65948 11397 65994 11409
rect 66066 11785 66112 11797
rect 66066 11409 66072 11785
rect 66106 11409 66112 11785
rect 66066 11397 66112 11409
rect 66184 11785 66230 11797
rect 66184 11409 66190 11785
rect 66224 11409 66230 11785
rect 66184 11397 66230 11409
rect 66302 11785 66348 11797
rect 66302 11409 66308 11785
rect 66342 11409 66348 11785
rect 66302 11397 66348 11409
rect 66420 11785 66466 11797
rect 66420 11409 66426 11785
rect 66460 11585 66466 11785
rect 66791 11597 66825 11900
rect 67332 11820 67468 11840
rect 67332 11758 67368 11820
rect 67428 11758 67468 11820
rect 67332 11730 67468 11758
rect 67028 11700 68005 11730
rect 66549 11585 66595 11597
rect 66460 11409 66555 11585
rect 66589 11409 66595 11585
rect 66420 11397 66466 11409
rect 66549 11397 66595 11409
rect 66667 11585 66713 11597
rect 66667 11409 66673 11585
rect 66707 11409 66713 11585
rect 66667 11397 66713 11409
rect 66785 11585 66831 11597
rect 66785 11409 66791 11585
rect 66825 11409 66831 11585
rect 66785 11397 66831 11409
rect 66903 11585 66949 11597
rect 67028 11594 67060 11700
rect 67264 11594 67296 11700
rect 67500 11594 67532 11700
rect 67736 11594 67768 11700
rect 67971 11594 68005 11700
rect 66903 11409 66909 11585
rect 66943 11409 66949 11585
rect 66903 11397 66949 11409
rect 67021 11582 67067 11594
rect 67021 11406 67027 11582
rect 67061 11406 67067 11582
rect 64010 11365 64059 11370
rect 64128 11365 64174 11377
rect 64016 11204 64059 11365
rect 65234 11363 65268 11397
rect 65836 11363 65870 11397
rect 66072 11363 66106 11397
rect 65234 11328 65393 11363
rect 65836 11328 66106 11363
rect 66673 11363 66707 11397
rect 66909 11363 66943 11397
rect 67021 11394 67067 11406
rect 67139 11582 67185 11594
rect 67139 11406 67145 11582
rect 67179 11406 67185 11582
rect 67139 11394 67185 11406
rect 67257 11582 67303 11594
rect 67257 11406 67263 11582
rect 67297 11406 67303 11582
rect 67257 11394 67303 11406
rect 67375 11582 67421 11594
rect 67375 11406 67381 11582
rect 67415 11406 67421 11582
rect 67375 11394 67421 11406
rect 67493 11582 67539 11594
rect 67493 11406 67499 11582
rect 67533 11406 67539 11582
rect 67493 11394 67539 11406
rect 67611 11582 67657 11594
rect 67611 11406 67617 11582
rect 67651 11406 67657 11582
rect 67611 11394 67657 11406
rect 67729 11582 67775 11594
rect 67729 11406 67735 11582
rect 67769 11406 67775 11582
rect 67729 11394 67775 11406
rect 67847 11582 67893 11594
rect 67847 11406 67853 11582
rect 67887 11406 67893 11582
rect 67847 11394 67893 11406
rect 67965 11582 68011 11594
rect 67965 11406 67971 11582
rect 68005 11406 68011 11582
rect 67965 11394 68011 11406
rect 68083 11582 68129 11594
rect 68083 11406 68089 11582
rect 68123 11406 68129 11582
rect 68083 11394 68129 11406
rect 66673 11328 66943 11363
rect 65170 11246 65299 11247
rect 63933 11177 64059 11204
rect 63893 11165 64059 11177
rect 63899 11161 64059 11165
rect 63107 11159 63194 11160
rect 63107 11155 63490 11159
rect 63102 11081 63112 11155
rect 63191 11134 63490 11155
rect 63191 11133 63624 11134
rect 63191 11127 63772 11133
rect 63191 11093 63722 11127
rect 63756 11093 63772 11127
rect 63191 11081 63772 11093
rect 62784 6893 62969 6899
rect 62784 6795 62796 6893
rect 62928 6795 62969 6893
rect 62784 6789 62969 6795
rect 62869 6788 62969 6789
rect 63107 11077 63772 11081
rect 63824 11127 63890 11133
rect 63824 11093 63840 11127
rect 63874 11093 63890 11127
rect 57728 5763 58097 5811
rect 57728 5733 57742 5763
rect 57728 5716 57738 5733
rect 58030 5660 58096 5763
rect 59861 5721 59867 5859
rect 59934 5721 59940 5859
rect 59861 5709 59940 5721
rect 62656 5660 62722 5939
rect 58028 5580 62722 5660
rect 63107 5693 63197 11077
rect 63824 11048 63890 11093
rect 63257 11041 63890 11048
rect 63254 10945 63264 11041
rect 63345 11040 63890 11041
rect 63345 11008 63891 11040
rect 63983 11024 64059 11161
rect 64769 11243 65299 11246
rect 64769 11180 65221 11243
rect 65288 11180 65299 11243
rect 64769 11177 65299 11180
rect 63345 10945 63490 11008
rect 63979 10964 63989 11024
rect 64051 10964 64061 11024
rect 64769 10957 64911 11177
rect 65201 11121 65305 11127
rect 65201 11053 65213 11121
rect 65293 11053 65305 11121
rect 65201 11047 65305 11053
rect 63257 8854 63351 10945
rect 63726 9657 63862 9677
rect 63726 9595 63762 9657
rect 63822 9595 63862 9657
rect 63726 9567 63862 9595
rect 63422 9537 64399 9567
rect 63422 9431 63454 9537
rect 63658 9431 63690 9537
rect 63894 9431 63926 9537
rect 64130 9431 64162 9537
rect 64365 9431 64399 9537
rect 63415 9419 63461 9431
rect 63415 9243 63421 9419
rect 63455 9243 63461 9419
rect 63415 9231 63461 9243
rect 63533 9419 63579 9431
rect 63533 9243 63539 9419
rect 63573 9243 63579 9419
rect 63533 9231 63579 9243
rect 63651 9419 63697 9431
rect 63651 9243 63657 9419
rect 63691 9243 63697 9419
rect 63651 9231 63697 9243
rect 63769 9419 63815 9431
rect 63769 9243 63775 9419
rect 63809 9243 63815 9419
rect 63769 9231 63815 9243
rect 63887 9419 63933 9431
rect 63887 9243 63893 9419
rect 63927 9243 63933 9419
rect 63887 9231 63933 9243
rect 64005 9419 64051 9431
rect 64005 9243 64011 9419
rect 64045 9243 64051 9419
rect 64005 9231 64051 9243
rect 64123 9419 64169 9431
rect 64123 9243 64129 9419
rect 64163 9243 64169 9419
rect 64123 9231 64169 9243
rect 64241 9419 64287 9431
rect 64241 9243 64247 9419
rect 64281 9243 64287 9419
rect 64241 9231 64287 9243
rect 64359 9419 64405 9431
rect 64359 9243 64365 9419
rect 64399 9243 64405 9419
rect 64359 9231 64405 9243
rect 64477 9419 64523 9431
rect 64477 9243 64483 9419
rect 64517 9243 64523 9419
rect 64477 9231 64523 9243
rect 63538 9137 63574 9231
rect 63774 9137 63810 9231
rect 64010 9138 64046 9231
rect 64172 9183 64238 9190
rect 64172 9149 64188 9183
rect 64222 9149 64238 9183
rect 64172 9138 64238 9149
rect 64010 9137 64238 9138
rect 63538 9108 64238 9137
rect 63538 9107 64120 9108
rect 63658 8994 63692 9107
rect 64054 9066 64120 9107
rect 64054 9032 64070 9066
rect 64104 9032 64120 9066
rect 64054 9025 64120 9032
rect 64482 8998 64517 9231
rect 64769 8998 64910 10957
rect 65359 10544 65393 11328
rect 66072 11266 66106 11328
rect 65661 11228 66403 11266
rect 65471 11057 65481 11125
rect 65536 11057 65546 11125
rect 65661 11104 65695 11228
rect 65897 11104 65931 11228
rect 66133 11104 66167 11228
rect 66369 11104 66403 11228
rect 65655 11092 65701 11104
rect 65655 10716 65661 11092
rect 65695 10716 65701 11092
rect 65655 10704 65701 10716
rect 65773 11092 65819 11104
rect 65773 10716 65779 11092
rect 65813 10716 65819 11092
rect 65773 10704 65819 10716
rect 65891 11092 65937 11104
rect 65891 10716 65897 11092
rect 65931 10716 65937 11092
rect 65891 10704 65937 10716
rect 66009 11092 66055 11104
rect 66009 10716 66015 11092
rect 66049 10716 66055 11092
rect 66009 10704 66055 10716
rect 66127 11092 66173 11104
rect 66127 10716 66133 11092
rect 66167 10716 66173 11092
rect 66127 10704 66173 10716
rect 66245 11092 66291 11104
rect 66245 10716 66251 11092
rect 66285 10716 66291 11092
rect 66245 10704 66291 10716
rect 66363 11092 66409 11104
rect 66363 10716 66369 11092
rect 66403 10716 66409 11092
rect 66529 10887 66603 10899
rect 66525 10796 66535 10887
rect 66597 10796 66607 10887
rect 66529 10784 66603 10796
rect 66363 10704 66409 10716
rect 66775 10545 66809 11328
rect 67144 11300 67180 11394
rect 67380 11300 67416 11394
rect 67616 11301 67652 11394
rect 67778 11346 67844 11353
rect 67778 11312 67794 11346
rect 67828 11312 67844 11346
rect 67778 11301 67844 11312
rect 67616 11300 67844 11301
rect 67144 11271 67844 11300
rect 67144 11270 67726 11271
rect 66870 11238 66946 11243
rect 66867 11182 66877 11238
rect 66930 11237 66946 11238
rect 66930 11182 67196 11237
rect 66870 11177 67196 11182
rect 66991 11135 67082 11140
rect 66991 11046 67001 11135
rect 67074 11046 67082 11135
rect 66991 11034 67082 11046
rect 67028 10640 67082 11034
rect 67142 10725 67196 11177
rect 67264 11157 67298 11270
rect 67660 11229 67726 11270
rect 67660 11195 67676 11229
rect 67710 11195 67726 11229
rect 67660 11188 67726 11195
rect 68088 11161 68123 11394
rect 67734 11157 68123 11161
rect 67258 11145 67304 11157
rect 67258 10769 67264 11145
rect 67298 10769 67304 11145
rect 67258 10757 67304 10769
rect 67376 11145 67422 11157
rect 67376 10769 67382 11145
rect 67416 10769 67422 11145
rect 67376 10757 67422 10769
rect 67494 11145 67540 11157
rect 67494 10769 67500 11145
rect 67534 10796 67540 11145
rect 67611 11145 67657 11157
rect 67611 10969 67617 11145
rect 67651 10969 67657 11145
rect 67611 10962 67657 10969
rect 67729 11145 68123 11157
rect 67729 10969 67735 11145
rect 67769 11132 68123 11145
rect 67769 10969 67775 11132
rect 67948 11130 68123 11132
rect 67948 11072 67990 11130
rect 68102 11072 68123 11130
rect 67948 11043 68123 11072
rect 67611 10957 67660 10962
rect 67729 10957 67775 10969
rect 67617 10796 67660 10957
rect 67534 10769 67660 10796
rect 67758 10897 68086 10898
rect 67758 10890 68152 10897
rect 67758 10882 68012 10890
rect 67758 10801 67774 10882
rect 67882 10801 68012 10882
rect 67758 10796 68012 10801
rect 68135 10796 68152 10890
rect 67758 10784 68152 10796
rect 68002 10783 68152 10784
rect 67494 10757 67660 10769
rect 67500 10753 67660 10757
rect 67142 10719 67373 10725
rect 67142 10685 67323 10719
rect 67357 10685 67373 10719
rect 67142 10669 67373 10685
rect 67425 10719 67491 10725
rect 67425 10685 67441 10719
rect 67475 10685 67491 10719
rect 67425 10640 67491 10685
rect 67028 10632 67491 10640
rect 67028 10600 67492 10632
rect 67584 10616 67660 10753
rect 67580 10556 67590 10616
rect 67652 10556 67662 10616
rect 66502 10544 66809 10545
rect 65359 10539 65675 10544
rect 66389 10539 66809 10544
rect 65359 10528 65742 10539
rect 65359 10501 65691 10528
rect 65359 10372 65393 10501
rect 65675 10494 65691 10501
rect 65725 10494 65742 10528
rect 65675 10488 65742 10494
rect 66322 10528 66809 10539
rect 67588 10530 67658 10556
rect 66322 10494 66339 10528
rect 66373 10501 66809 10528
rect 66373 10494 66389 10501
rect 66502 10500 66809 10501
rect 66322 10488 66389 10494
rect 65500 10461 65556 10473
rect 65500 10427 65506 10461
rect 65540 10460 65556 10461
rect 66613 10460 66669 10472
rect 65540 10444 66007 10460
rect 65540 10427 65957 10444
rect 65500 10411 65957 10427
rect 65941 10410 65957 10411
rect 65991 10410 66007 10444
rect 65941 10403 66007 10410
rect 66059 10445 66629 10460
rect 66059 10411 66075 10445
rect 66109 10426 66629 10445
rect 66663 10426 66669 10460
rect 66109 10411 66669 10426
rect 66059 10401 66126 10411
rect 66613 10410 66669 10411
rect 66775 10372 66809 10500
rect 65353 10360 65399 10372
rect 65353 10184 65359 10360
rect 65393 10184 65399 10360
rect 65353 10172 65399 10184
rect 65471 10360 65517 10372
rect 65471 10184 65477 10360
rect 65511 10184 65517 10360
rect 65471 10172 65517 10184
rect 65773 10360 65819 10372
rect 65476 9878 65510 10172
rect 65773 9984 65779 10360
rect 65813 9984 65819 10360
rect 65773 9972 65819 9984
rect 65891 10360 65937 10372
rect 65891 9984 65897 10360
rect 65931 9984 65937 10360
rect 65891 9972 65937 9984
rect 66009 10360 66055 10372
rect 66009 9984 66015 10360
rect 66049 9984 66055 10360
rect 66009 9972 66055 9984
rect 66127 10360 66173 10372
rect 66127 9984 66133 10360
rect 66167 9984 66173 10360
rect 66127 9972 66173 9984
rect 66245 10360 66291 10372
rect 66245 9984 66251 10360
rect 66285 9984 66291 10360
rect 66651 10360 66697 10372
rect 66651 10184 66657 10360
rect 66691 10184 66697 10360
rect 66651 10172 66697 10184
rect 66769 10360 66815 10372
rect 66769 10184 66775 10360
rect 66809 10184 66815 10360
rect 66769 10172 66815 10184
rect 66245 9972 66291 9984
rect 66133 9878 66167 9972
rect 66657 9878 66690 10172
rect 65476 9846 66690 9878
rect 65842 9822 66248 9846
rect 65842 9699 65954 9822
rect 66128 9699 66248 9822
rect 65842 9655 66248 9699
rect 64128 8994 64910 8998
rect 63652 8982 63698 8994
rect 63257 8757 63590 8854
rect 63400 8714 63500 8726
rect 63400 8633 63411 8714
rect 63493 8633 63503 8714
rect 63400 8626 63500 8633
rect 63422 8477 63476 8626
rect 63536 8562 63590 8757
rect 63652 8606 63658 8982
rect 63692 8606 63698 8982
rect 63652 8594 63698 8606
rect 63770 8982 63816 8994
rect 63770 8606 63776 8982
rect 63810 8606 63816 8982
rect 63770 8594 63816 8606
rect 63888 8982 63934 8994
rect 63888 8606 63894 8982
rect 63928 8633 63934 8982
rect 64005 8982 64051 8994
rect 64005 8806 64011 8982
rect 64045 8806 64051 8982
rect 64005 8799 64051 8806
rect 64123 8982 64910 8994
rect 64123 8806 64129 8982
rect 64163 8969 64910 8982
rect 64163 8806 64169 8969
rect 64413 8887 64910 8969
rect 64005 8794 64054 8799
rect 64123 8794 64169 8806
rect 64011 8633 64054 8794
rect 63928 8606 64054 8633
rect 63888 8594 64054 8606
rect 63894 8590 64054 8594
rect 63536 8556 63767 8562
rect 63536 8522 63717 8556
rect 63751 8522 63767 8556
rect 63536 8506 63767 8522
rect 63819 8556 63885 8562
rect 63819 8522 63835 8556
rect 63869 8522 63885 8556
rect 63819 8477 63885 8522
rect 63422 8469 63885 8477
rect 63422 8437 63886 8469
rect 63978 8453 64054 8590
rect 63974 8393 63984 8453
rect 64046 8393 64056 8453
rect 65858 8232 66303 8238
rect 65858 8032 65870 8232
rect 66291 8032 66303 8232
rect 65858 8026 66026 8032
rect 66016 7958 66026 8026
rect 66158 8026 66303 8032
rect 66158 7958 66168 8026
rect 66026 7918 66158 7958
rect 66025 7852 66158 7918
rect 65354 7809 66827 7852
rect 65354 7506 65388 7809
rect 65720 7706 65754 7809
rect 65956 7706 65990 7809
rect 66192 7706 66226 7809
rect 66428 7706 66462 7809
rect 65714 7694 65760 7706
rect 65230 7494 65276 7506
rect 65230 7318 65236 7494
rect 65270 7318 65276 7494
rect 65230 7306 65276 7318
rect 65348 7494 65394 7506
rect 65348 7318 65354 7494
rect 65388 7318 65394 7494
rect 65348 7306 65394 7318
rect 65466 7494 65512 7506
rect 65466 7318 65472 7494
rect 65506 7318 65512 7494
rect 65466 7306 65512 7318
rect 65584 7494 65630 7506
rect 65714 7494 65720 7694
rect 65584 7318 65590 7494
rect 65624 7318 65720 7494
rect 65754 7318 65760 7694
rect 65584 7306 65630 7318
rect 65714 7306 65760 7318
rect 65832 7694 65878 7706
rect 65832 7318 65838 7694
rect 65872 7318 65878 7694
rect 65832 7306 65878 7318
rect 65950 7694 65996 7706
rect 65950 7318 65956 7694
rect 65990 7318 65996 7694
rect 65950 7306 65996 7318
rect 66068 7694 66114 7706
rect 66068 7318 66074 7694
rect 66108 7318 66114 7694
rect 66068 7306 66114 7318
rect 66186 7694 66232 7706
rect 66186 7318 66192 7694
rect 66226 7318 66232 7694
rect 66186 7306 66232 7318
rect 66304 7694 66350 7706
rect 66304 7318 66310 7694
rect 66344 7318 66350 7694
rect 66304 7306 66350 7318
rect 66422 7694 66468 7706
rect 66422 7318 66428 7694
rect 66462 7494 66468 7694
rect 66793 7506 66827 7809
rect 67334 7729 67470 7749
rect 67334 7667 67370 7729
rect 67430 7667 67470 7729
rect 67334 7639 67470 7667
rect 67030 7609 68007 7639
rect 66551 7494 66597 7506
rect 66462 7318 66557 7494
rect 66591 7318 66597 7494
rect 66422 7306 66468 7318
rect 66551 7306 66597 7318
rect 66669 7494 66715 7506
rect 66669 7318 66675 7494
rect 66709 7318 66715 7494
rect 66669 7306 66715 7318
rect 66787 7494 66833 7506
rect 66787 7318 66793 7494
rect 66827 7318 66833 7494
rect 66787 7306 66833 7318
rect 66905 7494 66951 7506
rect 67030 7503 67062 7609
rect 67266 7503 67298 7609
rect 67502 7503 67534 7609
rect 67738 7503 67770 7609
rect 67973 7503 68007 7609
rect 66905 7318 66911 7494
rect 66945 7318 66951 7494
rect 66905 7306 66951 7318
rect 67023 7491 67069 7503
rect 67023 7315 67029 7491
rect 67063 7315 67069 7491
rect 65236 7272 65270 7306
rect 65838 7272 65872 7306
rect 66074 7272 66108 7306
rect 65236 7237 65395 7272
rect 65838 7237 66108 7272
rect 66675 7272 66709 7306
rect 66911 7272 66945 7306
rect 67023 7303 67069 7315
rect 67141 7491 67187 7503
rect 67141 7315 67147 7491
rect 67181 7315 67187 7491
rect 67141 7303 67187 7315
rect 67259 7491 67305 7503
rect 67259 7315 67265 7491
rect 67299 7315 67305 7491
rect 67259 7303 67305 7315
rect 67377 7491 67423 7503
rect 67377 7315 67383 7491
rect 67417 7315 67423 7491
rect 67377 7303 67423 7315
rect 67495 7491 67541 7503
rect 67495 7315 67501 7491
rect 67535 7315 67541 7491
rect 67495 7303 67541 7315
rect 67613 7491 67659 7503
rect 67613 7315 67619 7491
rect 67653 7315 67659 7491
rect 67613 7303 67659 7315
rect 67731 7491 67777 7503
rect 67731 7315 67737 7491
rect 67771 7315 67777 7491
rect 67731 7303 67777 7315
rect 67849 7491 67895 7503
rect 67849 7315 67855 7491
rect 67889 7315 67895 7491
rect 67849 7303 67895 7315
rect 67967 7491 68013 7503
rect 67967 7315 67973 7491
rect 68007 7315 68013 7491
rect 67967 7303 68013 7315
rect 68085 7491 68131 7503
rect 68085 7315 68091 7491
rect 68125 7315 68131 7491
rect 68085 7303 68131 7315
rect 66675 7237 66945 7272
rect 64605 7089 65223 7152
rect 65290 7089 65300 7152
rect 64605 7088 65259 7089
rect 63726 6624 63862 6644
rect 63726 6562 63762 6624
rect 63822 6562 63862 6624
rect 63726 6534 63862 6562
rect 63422 6504 64399 6534
rect 63422 6398 63454 6504
rect 63658 6398 63690 6504
rect 63894 6398 63926 6504
rect 64130 6398 64162 6504
rect 64365 6398 64399 6504
rect 63415 6386 63461 6398
rect 63415 6210 63421 6386
rect 63455 6210 63461 6386
rect 63415 6198 63461 6210
rect 63533 6386 63579 6398
rect 63533 6210 63539 6386
rect 63573 6210 63579 6386
rect 63533 6198 63579 6210
rect 63651 6386 63697 6398
rect 63651 6210 63657 6386
rect 63691 6210 63697 6386
rect 63651 6198 63697 6210
rect 63769 6386 63815 6398
rect 63769 6210 63775 6386
rect 63809 6210 63815 6386
rect 63769 6198 63815 6210
rect 63887 6386 63933 6398
rect 63887 6210 63893 6386
rect 63927 6210 63933 6386
rect 63887 6198 63933 6210
rect 64005 6386 64051 6398
rect 64005 6210 64011 6386
rect 64045 6210 64051 6386
rect 64005 6198 64051 6210
rect 64123 6386 64169 6398
rect 64123 6210 64129 6386
rect 64163 6210 64169 6386
rect 64123 6198 64169 6210
rect 64241 6386 64287 6398
rect 64241 6210 64247 6386
rect 64281 6210 64287 6386
rect 64241 6198 64287 6210
rect 64359 6386 64405 6398
rect 64359 6210 64365 6386
rect 64399 6210 64405 6386
rect 64359 6198 64405 6210
rect 64477 6386 64523 6398
rect 64477 6210 64483 6386
rect 64517 6210 64523 6386
rect 64477 6198 64523 6210
rect 63538 6104 63574 6198
rect 63774 6104 63810 6198
rect 64010 6105 64046 6198
rect 64172 6150 64238 6157
rect 64172 6116 64188 6150
rect 64222 6116 64238 6150
rect 64172 6105 64238 6116
rect 64010 6104 64238 6105
rect 63538 6075 64238 6104
rect 63538 6074 64120 6075
rect 63658 5961 63692 6074
rect 64054 6033 64120 6074
rect 64054 5999 64070 6033
rect 64104 5999 64120 6033
rect 64054 5992 64120 5999
rect 64482 5965 64517 6198
rect 64605 5965 64696 7088
rect 64128 5961 64696 5965
rect 63652 5949 63698 5961
rect 63512 5813 63612 5821
rect 63506 5726 63516 5813
rect 63605 5726 63615 5813
rect 63512 5721 63612 5726
rect 63107 5593 63476 5693
rect 57262 5398 57272 5512
rect 57395 5398 57405 5512
rect 63422 5444 63476 5593
rect 63536 5529 63590 5721
rect 63652 5573 63658 5949
rect 63692 5573 63698 5949
rect 63652 5561 63698 5573
rect 63770 5949 63816 5961
rect 63770 5573 63776 5949
rect 63810 5573 63816 5949
rect 63770 5561 63816 5573
rect 63888 5949 63934 5961
rect 63888 5573 63894 5949
rect 63928 5600 63934 5949
rect 64005 5949 64051 5961
rect 64005 5773 64011 5949
rect 64045 5773 64051 5949
rect 64005 5766 64051 5773
rect 64123 5949 64696 5961
rect 64123 5773 64129 5949
rect 64163 5936 64696 5949
rect 64163 5773 64169 5936
rect 64413 5856 64696 5936
rect 64785 6963 65223 7026
rect 65290 6963 65300 7026
rect 64005 5761 64054 5766
rect 64123 5761 64169 5773
rect 64011 5600 64054 5761
rect 63928 5573 64054 5600
rect 63888 5561 64054 5573
rect 63894 5557 64054 5561
rect 63536 5523 63767 5529
rect 63536 5489 63717 5523
rect 63751 5489 63767 5523
rect 63536 5473 63767 5489
rect 63819 5523 63885 5529
rect 63819 5489 63835 5523
rect 63869 5489 63885 5523
rect 63819 5444 63885 5489
rect 63422 5436 63885 5444
rect 63422 5404 63886 5436
rect 63978 5420 64054 5557
rect 63974 5360 63984 5420
rect 64046 5360 64056 5420
rect 63797 4704 63933 4724
rect 60562 4653 60641 4665
rect 58083 4605 58162 4617
rect 58083 4508 58089 4605
rect 58013 4488 58089 4508
rect 58156 4508 58162 4605
rect 60562 4542 60568 4653
rect 60635 4542 60641 4653
rect 61710 4659 61789 4671
rect 61710 4542 61716 4659
rect 61783 4542 61789 4659
rect 63797 4642 63833 4704
rect 63893 4642 63933 4704
rect 63797 4614 63933 4642
rect 63493 4584 64470 4614
rect 58156 4488 58233 4508
rect 58013 4380 58057 4488
rect 58189 4380 58233 4488
rect 59810 4446 59866 4454
rect 58013 4338 58233 4380
rect 58884 4438 59866 4446
rect 58884 4404 59826 4438
rect 59860 4404 59866 4438
rect 60529 4434 60539 4542
rect 60671 4479 60681 4542
rect 60671 4468 60683 4479
rect 60671 4434 60684 4468
rect 60940 4458 60996 4460
rect 58884 4388 59866 4404
rect 60539 4396 60684 4434
rect 58884 4387 59863 4388
rect 57617 4308 58594 4338
rect 57617 4202 57649 4308
rect 57853 4202 57885 4308
rect 58089 4202 58121 4308
rect 58325 4202 58357 4308
rect 58560 4202 58594 4308
rect 57610 4190 57656 4202
rect 57610 4014 57616 4190
rect 57650 4014 57656 4190
rect 57610 4002 57656 4014
rect 57728 4190 57774 4202
rect 57728 4014 57734 4190
rect 57768 4014 57774 4190
rect 57728 4002 57774 4014
rect 57846 4190 57892 4202
rect 57846 4014 57852 4190
rect 57886 4014 57892 4190
rect 57846 4002 57892 4014
rect 57964 4190 58010 4202
rect 57964 4014 57970 4190
rect 58004 4014 58010 4190
rect 57964 4002 58010 4014
rect 58082 4190 58128 4202
rect 58082 4014 58088 4190
rect 58122 4014 58128 4190
rect 58082 4002 58128 4014
rect 58200 4190 58246 4202
rect 58200 4014 58206 4190
rect 58240 4014 58246 4190
rect 58200 4002 58246 4014
rect 58318 4190 58364 4202
rect 58318 4014 58324 4190
rect 58358 4014 58364 4190
rect 58318 4002 58364 4014
rect 58436 4190 58482 4202
rect 58436 4014 58442 4190
rect 58476 4014 58482 4190
rect 58436 4002 58482 4014
rect 58554 4190 58600 4202
rect 58554 4014 58560 4190
rect 58594 4014 58600 4190
rect 58554 4002 58600 4014
rect 58672 4190 58718 4202
rect 58672 4014 58678 4190
rect 58712 4014 58718 4190
rect 58672 4002 58718 4014
rect 57733 3908 57769 4002
rect 57969 3908 58005 4002
rect 58205 3909 58241 4002
rect 58367 3954 58433 3961
rect 58367 3920 58383 3954
rect 58417 3920 58433 3954
rect 58367 3909 58433 3920
rect 58205 3908 58433 3909
rect 57733 3879 58433 3908
rect 57733 3878 58315 3879
rect 56384 3708 56537 3846
rect 57853 3765 57887 3878
rect 58249 3837 58315 3878
rect 58249 3803 58265 3837
rect 58299 3803 58315 3837
rect 58249 3796 58315 3803
rect 58677 3797 58712 4002
rect 58884 3797 58951 4387
rect 60643 4364 60684 4396
rect 60930 4392 60940 4458
rect 60996 4392 61006 4458
rect 61676 4434 61686 4542
rect 61818 4479 61828 4542
rect 61818 4468 61830 4479
rect 63493 4478 63525 4584
rect 63729 4478 63761 4584
rect 63965 4478 63997 4584
rect 64201 4478 64233 4584
rect 64436 4478 64470 4584
rect 61818 4434 61831 4468
rect 61686 4396 61831 4434
rect 61790 4368 61831 4396
rect 60059 4336 60329 4364
rect 59800 4270 59810 4336
rect 59876 4270 59886 4336
rect 60059 4274 60093 4336
rect 60295 4274 60329 4336
rect 60413 4336 60684 4364
rect 61201 4340 61471 4368
rect 60413 4274 60447 4336
rect 60649 4274 60684 4336
rect 60825 4324 60996 4340
rect 60825 4290 60956 4324
rect 60990 4290 60996 4324
rect 60825 4274 60996 4290
rect 61201 4278 61235 4340
rect 61437 4278 61471 4340
rect 61555 4340 61831 4368
rect 61555 4278 61589 4340
rect 61791 4278 61831 4340
rect 63486 4466 63532 4478
rect 63486 4290 63492 4466
rect 63526 4290 63532 4466
rect 63486 4278 63532 4290
rect 63604 4466 63650 4478
rect 63604 4290 63610 4466
rect 63644 4290 63650 4466
rect 63604 4278 63650 4290
rect 63722 4466 63768 4478
rect 63722 4290 63728 4466
rect 63762 4290 63768 4466
rect 63722 4278 63768 4290
rect 63840 4466 63886 4478
rect 63840 4290 63846 4466
rect 63880 4290 63886 4466
rect 63840 4278 63886 4290
rect 63958 4466 64004 4478
rect 63958 4290 63964 4466
rect 63998 4290 64004 4466
rect 63958 4278 64004 4290
rect 64076 4466 64122 4478
rect 64076 4290 64082 4466
rect 64116 4290 64122 4466
rect 64076 4278 64122 4290
rect 64194 4466 64240 4478
rect 64194 4290 64200 4466
rect 64234 4290 64240 4466
rect 64194 4278 64240 4290
rect 64312 4466 64358 4478
rect 64312 4290 64318 4466
rect 64352 4290 64358 4466
rect 64312 4278 64358 4290
rect 64430 4466 64476 4478
rect 64430 4290 64436 4466
rect 64470 4290 64476 4466
rect 64430 4278 64476 4290
rect 64548 4466 64594 4478
rect 64548 4290 64554 4466
rect 64588 4290 64594 4466
rect 64548 4278 64594 4290
rect 59935 4262 59981 4274
rect 59935 3886 59941 4262
rect 59975 3886 59981 4262
rect 59935 3874 59981 3886
rect 60053 4262 60099 4274
rect 60053 3886 60059 4262
rect 60093 3886 60099 4262
rect 60053 3874 60099 3886
rect 60171 4262 60217 4274
rect 60171 3886 60177 4262
rect 60211 3886 60217 4262
rect 60171 3874 60217 3886
rect 60289 4262 60335 4274
rect 60289 3886 60295 4262
rect 60329 3886 60335 4262
rect 60289 3874 60335 3886
rect 60407 4262 60453 4274
rect 60407 3886 60413 4262
rect 60447 3886 60453 4262
rect 60407 3874 60453 3886
rect 60525 4262 60571 4274
rect 60525 3886 60531 4262
rect 60565 3886 60571 4262
rect 60525 3874 60571 3886
rect 60643 4262 60689 4274
rect 60643 3886 60649 4262
rect 60683 3886 60689 4262
rect 60643 3874 60689 3886
rect 58677 3769 58951 3797
rect 58323 3765 58951 3769
rect 55169 3640 55278 3694
rect 54489 3601 54716 3637
rect 54489 3494 54524 3601
rect 54650 3567 54716 3601
rect 54650 3533 54666 3567
rect 54700 3533 54716 3567
rect 54997 3625 55094 3640
rect 54997 3558 55054 3625
rect 54650 3527 54716 3533
rect 54891 3522 55160 3558
rect 54891 3494 54924 3522
rect 55127 3494 55160 3522
rect 55244 3494 55278 3640
rect 56095 3633 56105 3708
rect 56173 3633 56537 3708
rect 56122 3632 56537 3633
rect 57847 3753 57893 3765
rect 54365 3482 54411 3494
rect 54365 3306 54371 3482
rect 54405 3306 54411 3482
rect 54365 3294 54411 3306
rect 54483 3482 54529 3494
rect 54483 3306 54489 3482
rect 54523 3306 54529 3482
rect 54483 3294 54529 3306
rect 54601 3482 54647 3494
rect 54601 3306 54607 3482
rect 54641 3306 54647 3482
rect 54601 3294 54647 3306
rect 54719 3482 54765 3494
rect 54719 3306 54725 3482
rect 54759 3427 54765 3482
rect 54884 3482 54930 3494
rect 54884 3427 54890 3482
rect 54759 3339 54890 3427
rect 54759 3306 54765 3339
rect 54719 3294 54765 3306
rect 54884 3306 54890 3339
rect 54924 3306 54930 3482
rect 54884 3294 54930 3306
rect 55002 3482 55048 3494
rect 55002 3306 55008 3482
rect 55042 3306 55048 3482
rect 55002 3294 55048 3306
rect 55120 3482 55166 3494
rect 55120 3306 55126 3482
rect 55160 3306 55166 3482
rect 55120 3294 55166 3306
rect 55238 3482 55284 3494
rect 55238 3306 55244 3482
rect 55278 3306 55284 3482
rect 57847 3377 57853 3753
rect 57887 3377 57893 3753
rect 57847 3365 57893 3377
rect 57965 3753 58011 3765
rect 57965 3377 57971 3753
rect 58005 3377 58011 3753
rect 57965 3365 58011 3377
rect 58083 3753 58129 3765
rect 58083 3377 58089 3753
rect 58123 3401 58129 3753
rect 58200 3753 58246 3765
rect 58200 3577 58206 3753
rect 58240 3577 58246 3753
rect 58200 3565 58246 3577
rect 58318 3753 58951 3765
rect 58318 3577 58324 3753
rect 58358 3740 58951 3753
rect 59941 3832 59975 3874
rect 60177 3832 60211 3874
rect 59941 3804 60211 3832
rect 60295 3833 60329 3874
rect 60531 3833 60565 3874
rect 60295 3804 60565 3833
rect 59941 3756 59975 3804
rect 58358 3577 58364 3740
rect 59941 3726 60004 3756
rect 58318 3565 58364 3577
rect 59969 3634 60004 3726
rect 59969 3598 60196 3634
rect 60466 3623 60476 3720
rect 60575 3623 60585 3720
rect 60649 3691 60683 3874
rect 60649 3637 60758 3691
rect 58206 3449 58241 3565
rect 59969 3491 60004 3598
rect 60130 3564 60196 3598
rect 60130 3530 60146 3564
rect 60180 3530 60196 3564
rect 60477 3622 60574 3623
rect 60477 3555 60534 3622
rect 60130 3524 60196 3530
rect 60371 3519 60640 3555
rect 60371 3491 60404 3519
rect 60607 3491 60640 3519
rect 60724 3491 60758 3637
rect 59845 3479 59891 3491
rect 58337 3449 58445 3459
rect 58206 3401 58337 3449
rect 58445 3417 58590 3423
rect 58123 3377 58337 3401
rect 58083 3365 58337 3377
rect 58089 3361 58337 3365
rect 55238 3294 55284 3306
rect 56154 3360 57000 3361
rect 56154 3333 57725 3360
rect 56154 3327 57962 3333
rect 54371 3255 54405 3294
rect 54607 3255 54641 3294
rect 54371 3219 54641 3255
rect 55008 3256 55041 3294
rect 55244 3256 55277 3294
rect 55008 3220 55277 3256
rect 56154 3293 57912 3327
rect 57946 3293 57962 3327
rect 56154 3277 57962 3293
rect 58014 3327 58080 3333
rect 58014 3293 58030 3327
rect 58064 3293 58080 3327
rect 58263 3317 58337 3361
rect 58578 3350 58590 3417
rect 58445 3344 58590 3350
rect 58337 3307 58445 3317
rect 56154 3261 57725 3277
rect 56154 3260 57662 3261
rect 56154 3257 57197 3260
rect 54371 3218 54537 3219
rect 54405 3139 54537 3218
rect 54395 3031 54405 3139
rect 54537 3031 54547 3139
rect 54429 2903 54435 3031
rect 54502 2903 54508 3031
rect 54429 2891 54508 2903
rect 51009 2657 51986 2687
rect 54203 2685 54266 2702
rect 54128 2681 54266 2685
rect 51009 2551 51041 2657
rect 51245 2551 51277 2657
rect 51481 2551 51513 2657
rect 51717 2551 51749 2657
rect 51952 2551 51986 2657
rect 52296 2647 54266 2681
rect 52294 2618 54266 2647
rect 52294 2602 52340 2618
rect 54128 2616 54266 2618
rect 51002 2539 51048 2551
rect 51002 2363 51008 2539
rect 51042 2363 51048 2539
rect 51002 2351 51048 2363
rect 51120 2539 51166 2551
rect 51120 2363 51126 2539
rect 51160 2363 51166 2539
rect 51120 2351 51166 2363
rect 51238 2539 51284 2551
rect 51238 2363 51244 2539
rect 51278 2363 51284 2539
rect 51238 2351 51284 2363
rect 51356 2539 51402 2551
rect 51356 2363 51362 2539
rect 51396 2363 51402 2539
rect 51356 2351 51402 2363
rect 51474 2539 51520 2551
rect 51474 2363 51480 2539
rect 51514 2363 51520 2539
rect 51474 2351 51520 2363
rect 51592 2539 51638 2551
rect 51592 2363 51598 2539
rect 51632 2363 51638 2539
rect 51592 2351 51638 2363
rect 51710 2539 51756 2551
rect 51710 2363 51716 2539
rect 51750 2363 51756 2539
rect 51710 2351 51756 2363
rect 51828 2539 51874 2551
rect 51828 2363 51834 2539
rect 51868 2363 51874 2539
rect 51828 2351 51874 2363
rect 51946 2539 51992 2551
rect 51946 2363 51952 2539
rect 51986 2363 51992 2539
rect 51946 2351 51992 2363
rect 52064 2539 52110 2551
rect 52064 2363 52070 2539
rect 52104 2363 52110 2539
rect 52064 2351 52110 2363
rect 51125 2257 51161 2351
rect 51361 2257 51397 2351
rect 51597 2258 51633 2351
rect 51759 2303 51825 2310
rect 51759 2269 51775 2303
rect 51809 2269 51825 2303
rect 51759 2258 51825 2269
rect 51597 2257 51825 2258
rect 51125 2228 51825 2257
rect 51125 2227 51707 2228
rect 51245 2114 51279 2227
rect 51641 2186 51707 2227
rect 51641 2152 51657 2186
rect 51691 2152 51707 2186
rect 51641 2145 51707 2152
rect 52069 2133 52104 2351
rect 52293 2150 52340 2602
rect 55190 2612 55269 2624
rect 55190 2494 55196 2612
rect 55263 2494 55269 2612
rect 53252 2386 53262 2494
rect 53394 2386 53404 2494
rect 55150 2386 55160 2494
rect 55292 2386 55302 2494
rect 53262 2346 53394 2386
rect 55160 2346 55292 2386
rect 53261 2280 53394 2346
rect 55159 2280 55292 2346
rect 52590 2237 54063 2280
rect 52293 2134 52339 2150
rect 52258 2133 52339 2134
rect 52069 2118 52339 2133
rect 51715 2114 52339 2118
rect 51239 2102 51285 2114
rect 50974 1624 50984 1742
rect 51102 1710 51112 1742
rect 51239 1726 51245 2102
rect 51279 1726 51285 2102
rect 51239 1714 51285 1726
rect 51357 2102 51403 2114
rect 51357 1726 51363 2102
rect 51397 1726 51403 2102
rect 51357 1714 51403 1726
rect 51475 2102 51521 2114
rect 51475 1726 51481 2102
rect 51515 1750 51521 2102
rect 51592 2102 51638 2114
rect 51592 1926 51598 2102
rect 51632 1926 51638 2102
rect 51592 1914 51638 1926
rect 51710 2102 52339 2114
rect 51710 1926 51716 2102
rect 51750 2090 52339 2102
rect 51750 2089 51992 2090
rect 51750 1926 51756 2089
rect 52258 2088 52339 2090
rect 52590 1934 52624 2237
rect 52956 2134 52990 2237
rect 53192 2134 53226 2237
rect 53428 2134 53462 2237
rect 53664 2134 53698 2237
rect 52950 2122 52996 2134
rect 51710 1914 51756 1926
rect 52466 1922 52512 1934
rect 51598 1798 51633 1914
rect 51729 1798 51837 1808
rect 51598 1750 51729 1798
rect 51837 1761 51985 1767
rect 51515 1726 51729 1750
rect 51475 1714 51729 1726
rect 51481 1710 51729 1714
rect 51102 1682 51117 1710
rect 51102 1676 51354 1682
rect 51102 1642 51304 1676
rect 51338 1642 51354 1676
rect 51102 1626 51354 1642
rect 51406 1676 51472 1682
rect 51406 1642 51422 1676
rect 51456 1642 51472 1676
rect 51655 1666 51729 1710
rect 51973 1694 51985 1761
rect 52466 1746 52472 1922
rect 52506 1746 52512 1922
rect 52466 1734 52512 1746
rect 52584 1922 52630 1934
rect 52584 1746 52590 1922
rect 52624 1746 52630 1922
rect 52584 1734 52630 1746
rect 52702 1922 52748 1934
rect 52702 1746 52708 1922
rect 52742 1746 52748 1922
rect 52702 1734 52748 1746
rect 52820 1922 52866 1934
rect 52950 1922 52956 2122
rect 52820 1746 52826 1922
rect 52860 1746 52956 1922
rect 52990 1746 52996 2122
rect 52820 1734 52866 1746
rect 52950 1734 52996 1746
rect 53068 2122 53114 2134
rect 53068 1746 53074 2122
rect 53108 1746 53114 2122
rect 53068 1734 53114 1746
rect 53186 2122 53232 2134
rect 53186 1746 53192 2122
rect 53226 1746 53232 2122
rect 53186 1734 53232 1746
rect 53304 2122 53350 2134
rect 53304 1746 53310 2122
rect 53344 1746 53350 2122
rect 53304 1734 53350 1746
rect 53422 2122 53468 2134
rect 53422 1746 53428 2122
rect 53462 1746 53468 2122
rect 53422 1734 53468 1746
rect 53540 2122 53586 2134
rect 53540 1746 53546 2122
rect 53580 1746 53586 2122
rect 53540 1734 53586 1746
rect 53658 2122 53704 2134
rect 53658 1746 53664 2122
rect 53698 1922 53704 2122
rect 54029 1934 54063 2237
rect 54488 2237 55961 2280
rect 54488 1934 54522 2237
rect 54854 2134 54888 2237
rect 55090 2134 55124 2237
rect 55326 2134 55360 2237
rect 55562 2134 55596 2237
rect 54848 2122 54894 2134
rect 53787 1922 53833 1934
rect 53698 1746 53793 1922
rect 53827 1746 53833 1922
rect 53658 1734 53704 1746
rect 53787 1734 53833 1746
rect 53905 1922 53951 1934
rect 53905 1746 53911 1922
rect 53945 1746 53951 1922
rect 53905 1734 53951 1746
rect 54023 1922 54069 1934
rect 54023 1746 54029 1922
rect 54063 1746 54069 1922
rect 54023 1734 54069 1746
rect 54141 1922 54187 1934
rect 54141 1746 54147 1922
rect 54181 1746 54187 1922
rect 54141 1734 54187 1746
rect 54364 1922 54410 1934
rect 54364 1746 54370 1922
rect 54404 1746 54410 1922
rect 54364 1734 54410 1746
rect 54482 1922 54528 1934
rect 54482 1746 54488 1922
rect 54522 1746 54528 1922
rect 54482 1734 54528 1746
rect 54600 1922 54646 1934
rect 54600 1746 54606 1922
rect 54640 1746 54646 1922
rect 54600 1734 54646 1746
rect 54718 1922 54764 1934
rect 54848 1922 54854 2122
rect 54718 1746 54724 1922
rect 54758 1746 54854 1922
rect 54888 1746 54894 2122
rect 54718 1734 54764 1746
rect 54848 1734 54894 1746
rect 54966 2122 55012 2134
rect 54966 1746 54972 2122
rect 55006 1746 55012 2122
rect 54966 1734 55012 1746
rect 55084 2122 55130 2134
rect 55084 1746 55090 2122
rect 55124 1746 55130 2122
rect 55084 1734 55130 1746
rect 55202 2122 55248 2134
rect 55202 1746 55208 2122
rect 55242 1746 55248 2122
rect 55202 1734 55248 1746
rect 55320 2122 55366 2134
rect 55320 1746 55326 2122
rect 55360 1746 55366 2122
rect 55320 1734 55366 1746
rect 55438 2122 55484 2134
rect 55438 1746 55444 2122
rect 55478 1746 55484 2122
rect 55438 1734 55484 1746
rect 55556 2122 55602 2134
rect 55556 1746 55562 2122
rect 55596 1922 55602 2122
rect 55927 1934 55961 2237
rect 55685 1922 55731 1934
rect 55596 1746 55691 1922
rect 55725 1746 55731 1922
rect 55556 1734 55602 1746
rect 55685 1734 55731 1746
rect 55803 1922 55849 1934
rect 55803 1746 55809 1922
rect 55843 1746 55849 1922
rect 55803 1734 55849 1746
rect 55921 1922 55967 1934
rect 55921 1746 55927 1922
rect 55961 1746 55967 1922
rect 55921 1734 55967 1746
rect 56039 1922 56085 1934
rect 56039 1746 56045 1922
rect 56079 1746 56085 1922
rect 56039 1734 56085 1746
rect 51837 1688 51985 1694
rect 52472 1700 52506 1734
rect 53074 1700 53108 1734
rect 53310 1700 53344 1734
rect 51729 1656 51837 1666
rect 52472 1665 52631 1700
rect 53074 1665 53344 1700
rect 53911 1700 53945 1734
rect 54147 1700 54181 1734
rect 53911 1665 54181 1700
rect 54370 1700 54404 1734
rect 54972 1700 55006 1734
rect 55208 1700 55242 1734
rect 54370 1665 54529 1700
rect 54972 1665 55242 1700
rect 55809 1700 55843 1734
rect 56045 1700 56079 1734
rect 55809 1665 56079 1700
rect 51102 1624 51117 1626
rect 51017 1610 51117 1624
rect 51017 1567 51117 1568
rect 50638 1546 51117 1567
rect 51406 1546 51472 1642
rect 50638 1498 51472 1546
rect 50638 1469 51117 1498
rect 50638 1467 50743 1469
rect 51017 1468 51117 1469
rect 50471 1282 50481 1361
rect 50574 1282 50584 1361
rect 51474 1346 51553 1358
rect 50482 108 50575 1282
rect 51474 1253 51480 1346
rect 51400 1233 51480 1253
rect 51547 1253 51553 1346
rect 51547 1233 51620 1253
rect 51400 1125 51444 1233
rect 51576 1125 51620 1233
rect 51400 1083 51620 1125
rect 51004 1053 51981 1083
rect 51004 947 51036 1053
rect 51240 947 51272 1053
rect 51476 947 51508 1053
rect 51712 947 51744 1053
rect 51947 947 51981 1053
rect 50997 935 51043 947
rect 50997 759 51003 935
rect 51037 759 51043 935
rect 50997 747 51043 759
rect 51115 935 51161 947
rect 51115 759 51121 935
rect 51155 759 51161 935
rect 51115 747 51161 759
rect 51233 935 51279 947
rect 51233 759 51239 935
rect 51273 759 51279 935
rect 51233 747 51279 759
rect 51351 935 51397 947
rect 51351 759 51357 935
rect 51391 759 51397 935
rect 51351 747 51397 759
rect 51469 935 51515 947
rect 51469 759 51475 935
rect 51509 759 51515 935
rect 51469 747 51515 759
rect 51587 935 51633 947
rect 51587 759 51593 935
rect 51627 759 51633 935
rect 51587 747 51633 759
rect 51705 935 51751 947
rect 51705 759 51711 935
rect 51745 759 51751 935
rect 51705 747 51751 759
rect 51823 935 51869 947
rect 51823 759 51829 935
rect 51863 759 51869 935
rect 51823 747 51869 759
rect 51941 935 51987 947
rect 51941 759 51947 935
rect 51981 759 51987 935
rect 51941 747 51987 759
rect 52059 935 52105 947
rect 52059 759 52065 935
rect 52099 759 52105 935
rect 52059 747 52105 759
rect 52597 881 52631 1665
rect 53310 1603 53344 1665
rect 52899 1565 53641 1603
rect 52899 1441 52933 1565
rect 53135 1441 53169 1565
rect 53371 1441 53405 1565
rect 53607 1441 53641 1565
rect 53897 1458 53907 1524
rect 53970 1458 53980 1524
rect 52893 1429 52939 1441
rect 52893 1053 52899 1429
rect 52933 1053 52939 1429
rect 52893 1041 52939 1053
rect 53011 1429 53057 1441
rect 53011 1053 53017 1429
rect 53051 1053 53057 1429
rect 53011 1041 53057 1053
rect 53129 1429 53175 1441
rect 53129 1053 53135 1429
rect 53169 1053 53175 1429
rect 53129 1041 53175 1053
rect 53247 1429 53293 1441
rect 53247 1053 53253 1429
rect 53287 1053 53293 1429
rect 53247 1041 53293 1053
rect 53365 1429 53411 1441
rect 53365 1053 53371 1429
rect 53405 1053 53411 1429
rect 53365 1041 53411 1053
rect 53483 1429 53529 1441
rect 53483 1053 53489 1429
rect 53523 1053 53529 1429
rect 53483 1041 53529 1053
rect 53601 1429 53647 1441
rect 53601 1053 53607 1429
rect 53641 1053 53647 1429
rect 53601 1041 53647 1053
rect 54013 882 54047 1665
rect 53740 881 54047 882
rect 52597 876 52913 881
rect 53627 876 54047 881
rect 52597 865 52980 876
rect 52597 838 52929 865
rect 51120 653 51156 747
rect 51356 653 51392 747
rect 51592 654 51628 747
rect 51754 699 51820 706
rect 51754 665 51770 699
rect 51804 665 51820 699
rect 51754 654 51820 665
rect 51592 653 51820 654
rect 51120 624 51820 653
rect 51120 623 51702 624
rect 51240 510 51274 623
rect 51636 582 51702 623
rect 51636 548 51652 582
rect 51686 548 51702 582
rect 51636 541 51702 548
rect 52064 514 52099 747
rect 52597 709 52631 838
rect 52913 831 52929 838
rect 52963 831 52980 865
rect 52913 825 52980 831
rect 53560 865 54047 876
rect 53560 831 53577 865
rect 53611 838 54047 865
rect 53611 831 53627 838
rect 53740 837 54047 838
rect 53560 825 53627 831
rect 52738 798 52794 810
rect 52738 764 52744 798
rect 52778 797 52794 798
rect 53851 797 53907 809
rect 52778 781 53245 797
rect 52778 764 53195 781
rect 52738 748 53195 764
rect 53179 747 53195 748
rect 53229 747 53245 781
rect 53179 740 53245 747
rect 53297 782 53867 797
rect 53297 748 53313 782
rect 53347 763 53867 782
rect 53901 763 53907 797
rect 53347 748 53907 763
rect 53297 738 53364 748
rect 53851 747 53907 748
rect 54013 709 54047 837
rect 54495 881 54529 1665
rect 55208 1603 55242 1665
rect 54797 1565 55539 1603
rect 54797 1441 54831 1565
rect 55033 1441 55067 1565
rect 55269 1441 55303 1565
rect 55505 1441 55539 1565
rect 54791 1429 54837 1441
rect 54791 1053 54797 1429
rect 54831 1053 54837 1429
rect 54791 1041 54837 1053
rect 54909 1429 54955 1441
rect 54909 1053 54915 1429
rect 54949 1053 54955 1429
rect 54909 1041 54955 1053
rect 55027 1429 55073 1441
rect 55027 1053 55033 1429
rect 55067 1053 55073 1429
rect 55027 1041 55073 1053
rect 55145 1429 55191 1441
rect 55145 1053 55151 1429
rect 55185 1053 55191 1429
rect 55145 1041 55191 1053
rect 55263 1429 55309 1441
rect 55263 1053 55269 1429
rect 55303 1053 55309 1429
rect 55263 1041 55309 1053
rect 55381 1429 55427 1441
rect 55381 1053 55387 1429
rect 55421 1053 55427 1429
rect 55381 1041 55427 1053
rect 55499 1429 55545 1441
rect 55499 1053 55505 1429
rect 55539 1053 55545 1429
rect 55499 1041 55545 1053
rect 55911 882 55945 1665
rect 55523 881 55592 882
rect 55638 881 55945 882
rect 54495 876 54811 881
rect 55523 877 55945 881
rect 54495 865 54878 876
rect 54495 838 54827 865
rect 54495 709 54529 838
rect 54811 831 54827 838
rect 54861 831 54878 865
rect 54811 825 54878 831
rect 55456 866 55945 877
rect 55456 832 55473 866
rect 55507 838 55945 866
rect 55507 832 55523 838
rect 55638 837 55945 838
rect 55456 826 55523 832
rect 54636 798 54692 810
rect 54636 764 54642 798
rect 54676 797 54692 798
rect 55749 797 55805 809
rect 54676 781 55143 797
rect 54676 764 55093 781
rect 54636 748 55093 764
rect 55077 747 55093 748
rect 55127 747 55143 781
rect 55077 740 55143 747
rect 55195 782 55765 797
rect 55195 748 55211 782
rect 55245 763 55765 782
rect 55799 763 55805 797
rect 55245 748 55805 763
rect 55195 738 55262 748
rect 55749 747 55805 748
rect 55911 709 55945 837
rect 56026 1487 56093 1511
rect 56026 1453 56043 1487
rect 56077 1453 56093 1487
rect 51710 510 52099 514
rect 51234 498 51280 510
rect 51234 122 51240 498
rect 51274 122 51280 498
rect 51234 110 51280 122
rect 51352 498 51398 510
rect 51352 122 51358 498
rect 51392 122 51398 498
rect 51352 110 51398 122
rect 51470 498 51516 510
rect 51470 122 51476 498
rect 51510 146 51516 498
rect 51587 498 51633 510
rect 51587 322 51593 498
rect 51627 322 51633 498
rect 51587 310 51633 322
rect 51705 498 52099 510
rect 52591 697 52637 709
rect 52591 521 52597 697
rect 52631 521 52637 697
rect 52591 509 52637 521
rect 52709 697 52755 709
rect 52709 521 52715 697
rect 52749 521 52755 697
rect 52709 509 52755 521
rect 53011 697 53057 709
rect 51705 322 51711 498
rect 51745 485 52099 498
rect 51745 322 51751 485
rect 52021 482 52099 485
rect 52021 430 52031 482
rect 52094 430 52104 482
rect 52026 424 52099 430
rect 51705 310 51751 322
rect 51593 194 51628 310
rect 52714 215 52748 509
rect 53011 321 53017 697
rect 53051 321 53057 697
rect 53011 309 53057 321
rect 53129 697 53175 709
rect 53129 321 53135 697
rect 53169 321 53175 697
rect 53129 309 53175 321
rect 53247 697 53293 709
rect 53247 321 53253 697
rect 53287 321 53293 697
rect 53247 309 53293 321
rect 53365 697 53411 709
rect 53365 321 53371 697
rect 53405 321 53411 697
rect 53365 309 53411 321
rect 53483 697 53529 709
rect 53483 321 53489 697
rect 53523 321 53529 697
rect 53889 697 53935 709
rect 53889 521 53895 697
rect 53929 521 53935 697
rect 53889 509 53935 521
rect 54007 697 54053 709
rect 54007 521 54013 697
rect 54047 521 54053 697
rect 54007 509 54053 521
rect 54489 697 54535 709
rect 54489 521 54495 697
rect 54529 521 54535 697
rect 54489 509 54535 521
rect 54607 697 54653 709
rect 54607 521 54613 697
rect 54647 521 54653 697
rect 54607 509 54653 521
rect 54909 697 54955 709
rect 53483 309 53529 321
rect 53371 215 53405 309
rect 53895 215 53928 509
rect 51724 194 51832 204
rect 51593 146 51724 194
rect 52714 183 53928 215
rect 54612 215 54646 509
rect 54909 321 54915 697
rect 54949 321 54955 697
rect 54909 309 54955 321
rect 55027 697 55073 709
rect 55027 321 55033 697
rect 55067 321 55073 697
rect 55027 309 55073 321
rect 55145 697 55191 709
rect 55145 321 55151 697
rect 55185 321 55191 697
rect 55145 309 55191 321
rect 55263 697 55309 709
rect 55263 321 55269 697
rect 55303 321 55309 697
rect 55263 309 55309 321
rect 55381 697 55427 709
rect 55381 321 55387 697
rect 55421 321 55427 697
rect 55787 697 55833 709
rect 55787 521 55793 697
rect 55827 521 55833 697
rect 55787 509 55833 521
rect 55905 697 55951 709
rect 55905 521 55911 697
rect 55945 521 55951 697
rect 55905 509 55951 521
rect 55381 309 55427 321
rect 55269 215 55303 309
rect 55793 215 55826 509
rect 54612 183 55826 215
rect 51832 152 51988 158
rect 51510 122 51724 146
rect 51470 110 51724 122
rect 50482 106 51067 108
rect 51476 106 51724 110
rect 50482 78 51112 106
rect 50482 72 51349 78
rect 50482 38 51299 72
rect 51333 38 51349 72
rect 50482 22 51349 38
rect 51401 72 51467 78
rect 51401 38 51417 72
rect 51451 38 51467 72
rect 51650 62 51724 106
rect 51976 85 51988 152
rect 53207 98 53339 183
rect 55105 98 55237 183
rect 51832 79 51988 85
rect 51724 52 51832 62
rect 50482 6 51112 22
rect 50482 2 51067 6
rect 50482 1 50583 2
rect 51012 -47 51112 -36
rect 50142 -85 50310 -66
rect 50142 -172 50169 -85
rect 50271 -172 50310 -85
rect 50976 -153 50986 -47
rect 51098 -58 51112 -47
rect 51401 -58 51467 38
rect 53197 -10 53207 98
rect 53339 -10 53349 98
rect 55095 -10 55105 98
rect 55237 -10 55247 98
rect 56026 70 56093 1453
rect 56154 1024 56310 3257
rect 56995 3256 57197 3257
rect 56154 926 56166 1024
rect 56298 926 56310 1024
rect 56154 920 56310 926
rect 56437 2845 56981 2872
rect 56437 2739 56829 2845
rect 56941 2832 56981 2845
rect 56941 2739 56983 2832
rect 56437 2728 56983 2739
rect 56437 2727 56981 2728
rect 51098 -106 51467 -58
rect 51098 -136 51112 -106
rect 51098 -153 51108 -136
rect 50142 -178 50310 -172
rect 51400 -209 51466 -106
rect 53223 -150 53229 -10
rect 53296 -150 53302 -10
rect 53223 -162 53302 -150
rect 56026 -209 56092 70
rect 51398 -289 56092 -209
rect 54809 -800 55273 -768
rect 55361 -784 55371 -724
rect 55433 -784 55443 -724
rect 54809 -808 55272 -800
rect 54809 -956 54863 -808
rect 49151 -1288 49914 -1208
rect 48901 -1301 49914 -1288
rect 48861 -1313 49914 -1301
rect 48396 -1426 48430 -1313
rect 48866 -1317 49914 -1313
rect 49216 -1318 49914 -1317
rect 54498 -1057 54863 -956
rect 54923 -853 55154 -837
rect 54923 -887 55104 -853
rect 55138 -887 55154 -853
rect 54923 -893 55154 -887
rect 55206 -853 55272 -808
rect 55206 -887 55222 -853
rect 55256 -887 55272 -853
rect 55206 -893 55272 -887
rect 48792 -1351 48858 -1344
rect 48792 -1385 48808 -1351
rect 48842 -1385 48858 -1351
rect 48792 -1426 48858 -1385
rect 48276 -1427 48858 -1426
rect 48276 -1456 48976 -1427
rect 48276 -1550 48312 -1456
rect 48512 -1550 48548 -1456
rect 48748 -1457 48976 -1456
rect 48748 -1550 48784 -1457
rect 48910 -1468 48976 -1457
rect 48910 -1502 48926 -1468
rect 48960 -1502 48976 -1468
rect 48910 -1509 48976 -1502
rect 49220 -1550 49255 -1318
rect 48153 -1562 48199 -1550
rect 48153 -1738 48159 -1562
rect 48193 -1738 48199 -1562
rect 48153 -1750 48199 -1738
rect 48271 -1562 48317 -1550
rect 48271 -1738 48277 -1562
rect 48311 -1738 48317 -1562
rect 48271 -1750 48317 -1738
rect 48389 -1562 48435 -1550
rect 48389 -1738 48395 -1562
rect 48429 -1738 48435 -1562
rect 48389 -1750 48435 -1738
rect 48507 -1562 48553 -1550
rect 48507 -1738 48513 -1562
rect 48547 -1738 48553 -1562
rect 48507 -1750 48553 -1738
rect 48625 -1562 48671 -1550
rect 48625 -1738 48631 -1562
rect 48665 -1738 48671 -1562
rect 48625 -1750 48671 -1738
rect 48743 -1562 48789 -1550
rect 48743 -1738 48749 -1562
rect 48783 -1738 48789 -1562
rect 48743 -1750 48789 -1738
rect 48861 -1562 48907 -1550
rect 48861 -1738 48867 -1562
rect 48901 -1738 48907 -1562
rect 48861 -1750 48907 -1738
rect 48979 -1562 49025 -1550
rect 48979 -1738 48985 -1562
rect 49019 -1738 49025 -1562
rect 48979 -1750 49025 -1738
rect 49097 -1562 49143 -1550
rect 49097 -1738 49103 -1562
rect 49137 -1738 49143 -1562
rect 49097 -1750 49143 -1738
rect 49215 -1562 49261 -1550
rect 49215 -1738 49221 -1562
rect 49255 -1738 49261 -1562
rect 49215 -1750 49261 -1738
rect 48160 -1856 48192 -1750
rect 48396 -1856 48428 -1750
rect 48632 -1856 48664 -1750
rect 48868 -1856 48900 -1750
rect 49103 -1856 49137 -1750
rect 48160 -1886 49137 -1856
rect 48464 -1914 48600 -1886
rect 48464 -1976 48500 -1914
rect 48560 -1976 48600 -1914
rect 48464 -1996 48600 -1976
rect 54498 -2086 54584 -1057
rect 54923 -1085 54977 -893
rect 55365 -921 55441 -784
rect 55281 -925 55441 -921
rect 54652 -1092 54977 -1085
rect 54647 -1181 54657 -1092
rect 54726 -1181 54977 -1092
rect 54652 -1185 54977 -1181
rect 55039 -937 55085 -925
rect 55039 -1313 55045 -937
rect 55079 -1313 55085 -937
rect 55039 -1325 55085 -1313
rect 55157 -937 55203 -925
rect 55157 -1313 55163 -937
rect 55197 -1313 55203 -937
rect 55157 -1325 55203 -1313
rect 55275 -937 55441 -925
rect 55275 -1313 55281 -937
rect 55315 -964 55441 -937
rect 55315 -1313 55321 -964
rect 55398 -1125 55441 -964
rect 55275 -1325 55321 -1313
rect 55392 -1130 55441 -1125
rect 55392 -1137 55438 -1130
rect 55392 -1313 55398 -1137
rect 55432 -1313 55438 -1137
rect 55392 -1325 55438 -1313
rect 55510 -1137 55556 -1125
rect 55510 -1313 55516 -1137
rect 55550 -1300 55556 -1137
rect 56437 -1220 56593 2727
rect 56693 1733 56980 1762
rect 56693 1627 56828 1733
rect 56940 1731 56980 1733
rect 56946 1720 56980 1731
rect 56693 1625 56834 1627
rect 56946 1625 56981 1720
rect 56693 1616 56981 1625
rect 56693 1615 56980 1616
rect 56693 1614 56948 1615
rect 56696 -723 56848 1614
rect 57104 1362 57197 3256
rect 57260 3197 57726 3219
rect 58014 3197 58080 3293
rect 59845 3303 59851 3479
rect 59885 3303 59891 3479
rect 59845 3291 59891 3303
rect 59963 3479 60009 3491
rect 59963 3303 59969 3479
rect 60003 3303 60009 3479
rect 59963 3291 60009 3303
rect 60081 3479 60127 3491
rect 60081 3303 60087 3479
rect 60121 3303 60127 3479
rect 60081 3291 60127 3303
rect 60199 3479 60245 3491
rect 60199 3303 60205 3479
rect 60239 3424 60245 3479
rect 60364 3479 60410 3491
rect 60364 3424 60370 3479
rect 60239 3336 60370 3424
rect 60239 3303 60245 3336
rect 60199 3291 60245 3303
rect 60364 3303 60370 3336
rect 60404 3303 60410 3479
rect 60364 3291 60410 3303
rect 60482 3479 60528 3491
rect 60482 3303 60488 3479
rect 60522 3303 60528 3479
rect 60482 3291 60528 3303
rect 60600 3479 60646 3491
rect 60600 3303 60606 3479
rect 60640 3303 60646 3479
rect 60600 3291 60646 3303
rect 60718 3479 60764 3491
rect 60718 3303 60724 3479
rect 60758 3303 60764 3479
rect 60718 3291 60764 3303
rect 59851 3252 59885 3291
rect 60087 3252 60121 3291
rect 59851 3217 60121 3252
rect 60488 3253 60521 3291
rect 60724 3253 60757 3291
rect 60488 3217 60757 3253
rect 57260 3149 58080 3197
rect 59885 3216 60121 3217
rect 57260 3118 57726 3149
rect 59885 3142 60017 3216
rect 57260 2862 57365 3118
rect 59875 3034 59885 3142
rect 60017 3034 60027 3142
rect 58098 2955 58177 2967
rect 57260 2756 57323 2862
rect 57435 2756 57445 2862
rect 58098 2858 58104 2955
rect 58027 2838 58104 2858
rect 58171 2858 58177 2955
rect 59914 2904 59920 3034
rect 59987 2904 59993 3034
rect 59914 2892 59993 2904
rect 58171 2838 58247 2858
rect 57260 2745 57409 2756
rect 57260 1568 57365 2745
rect 58027 2730 58071 2838
rect 58203 2730 58247 2838
rect 58027 2688 58247 2730
rect 60825 2703 60887 4274
rect 61077 4266 61123 4278
rect 61077 3890 61083 4266
rect 61117 3890 61123 4266
rect 61077 3878 61123 3890
rect 61195 4266 61241 4278
rect 61195 3890 61201 4266
rect 61235 3890 61241 4266
rect 61195 3878 61241 3890
rect 61313 4266 61359 4278
rect 61313 3890 61319 4266
rect 61353 3890 61359 4266
rect 61313 3878 61359 3890
rect 61431 4266 61477 4278
rect 61431 3890 61437 4266
rect 61471 3890 61477 4266
rect 61431 3878 61477 3890
rect 61549 4266 61595 4278
rect 61549 3890 61555 4266
rect 61589 3890 61595 4266
rect 61549 3878 61595 3890
rect 61667 4266 61713 4278
rect 61667 3890 61673 4266
rect 61707 3890 61713 4266
rect 61667 3878 61713 3890
rect 61785 4266 61831 4278
rect 61785 3890 61791 4266
rect 61825 3890 61831 4266
rect 63609 4184 63645 4278
rect 63845 4184 63881 4278
rect 64081 4185 64117 4278
rect 64243 4230 64309 4237
rect 64243 4196 64259 4230
rect 64293 4196 64309 4230
rect 64243 4185 64309 4196
rect 64081 4184 64309 4185
rect 63609 4155 64309 4184
rect 63609 4154 64191 4155
rect 63729 4041 63763 4154
rect 64125 4113 64191 4154
rect 64125 4079 64141 4113
rect 64175 4079 64191 4113
rect 64125 4072 64191 4079
rect 64553 4045 64588 4278
rect 64199 4044 64588 4045
rect 64785 4044 64876 6963
rect 65361 6453 65395 7237
rect 66074 7175 66108 7237
rect 65663 7137 66405 7175
rect 65473 6966 65483 7034
rect 65538 6966 65548 7034
rect 65663 7013 65697 7137
rect 65899 7013 65933 7137
rect 66135 7013 66169 7137
rect 66371 7013 66405 7137
rect 65657 7001 65703 7013
rect 65657 6625 65663 7001
rect 65697 6625 65703 7001
rect 65657 6613 65703 6625
rect 65775 7001 65821 7013
rect 65775 6625 65781 7001
rect 65815 6625 65821 7001
rect 65775 6613 65821 6625
rect 65893 7001 65939 7013
rect 65893 6625 65899 7001
rect 65933 6625 65939 7001
rect 65893 6613 65939 6625
rect 66011 7001 66057 7013
rect 66011 6625 66017 7001
rect 66051 6625 66057 7001
rect 66011 6613 66057 6625
rect 66129 7001 66175 7013
rect 66129 6625 66135 7001
rect 66169 6625 66175 7001
rect 66129 6613 66175 6625
rect 66247 7001 66293 7013
rect 66247 6625 66253 7001
rect 66287 6625 66293 7001
rect 66247 6613 66293 6625
rect 66365 7001 66411 7013
rect 66365 6625 66371 7001
rect 66405 6625 66411 7001
rect 66531 6796 66605 6808
rect 66527 6705 66537 6796
rect 66599 6705 66609 6796
rect 66531 6693 66605 6705
rect 66365 6613 66411 6625
rect 66777 6454 66811 7237
rect 67146 7209 67182 7303
rect 67382 7209 67418 7303
rect 67618 7210 67654 7303
rect 67780 7255 67846 7262
rect 67780 7221 67796 7255
rect 67830 7221 67846 7255
rect 67780 7210 67846 7221
rect 67618 7209 67846 7210
rect 67146 7180 67846 7209
rect 67146 7179 67728 7180
rect 66872 7147 66948 7152
rect 66869 7091 66879 7147
rect 66932 7146 66948 7147
rect 66932 7091 67198 7146
rect 66872 7086 67198 7091
rect 66993 7044 67084 7049
rect 66993 6955 67003 7044
rect 67076 6955 67084 7044
rect 66993 6943 67084 6955
rect 67030 6549 67084 6943
rect 67144 6634 67198 7086
rect 67266 7066 67300 7179
rect 67662 7138 67728 7179
rect 67662 7104 67678 7138
rect 67712 7104 67728 7138
rect 67662 7097 67728 7104
rect 68090 7070 68125 7303
rect 67736 7066 68125 7070
rect 67260 7054 67306 7066
rect 67260 6678 67266 7054
rect 67300 6678 67306 7054
rect 67260 6666 67306 6678
rect 67378 7054 67424 7066
rect 67378 6678 67384 7054
rect 67418 6678 67424 7054
rect 67378 6666 67424 6678
rect 67496 7054 67542 7066
rect 67496 6678 67502 7054
rect 67536 6705 67542 7054
rect 67613 7054 67659 7066
rect 67613 6878 67619 7054
rect 67653 6878 67659 7054
rect 67613 6871 67659 6878
rect 67731 7054 68125 7066
rect 67731 6878 67737 7054
rect 67771 7044 68125 7054
rect 67771 7041 67984 7044
rect 67771 6878 67777 7041
rect 67950 6973 67984 7041
rect 68111 6973 68125 7044
rect 68413 7002 68495 12503
rect 67950 6952 68125 6973
rect 67613 6866 67662 6871
rect 67731 6866 67777 6878
rect 67619 6705 67662 6866
rect 67536 6678 67662 6705
rect 67496 6666 67662 6678
rect 67502 6662 67662 6666
rect 67144 6628 67375 6634
rect 67144 6594 67325 6628
rect 67359 6594 67375 6628
rect 67144 6578 67375 6594
rect 67427 6628 67493 6634
rect 67427 6594 67443 6628
rect 67477 6594 67493 6628
rect 67427 6549 67493 6594
rect 67030 6541 67493 6549
rect 67030 6509 67494 6541
rect 67586 6525 67662 6662
rect 67582 6465 67592 6525
rect 67654 6465 67664 6525
rect 66504 6453 66811 6454
rect 65361 6448 65677 6453
rect 66391 6448 66811 6453
rect 65361 6437 65744 6448
rect 65361 6410 65693 6437
rect 65361 6281 65395 6410
rect 65677 6403 65693 6410
rect 65727 6403 65744 6437
rect 65677 6397 65744 6403
rect 66324 6437 66811 6448
rect 67590 6439 67660 6465
rect 66324 6403 66341 6437
rect 66375 6410 66811 6437
rect 66375 6403 66391 6410
rect 66504 6409 66811 6410
rect 66324 6397 66391 6403
rect 65502 6370 65558 6382
rect 65502 6336 65508 6370
rect 65542 6369 65558 6370
rect 66615 6369 66671 6381
rect 65542 6353 66009 6369
rect 65542 6336 65959 6353
rect 65502 6320 65959 6336
rect 65943 6319 65959 6320
rect 65993 6319 66009 6353
rect 65943 6312 66009 6319
rect 66061 6354 66631 6369
rect 66061 6320 66077 6354
rect 66111 6335 66631 6354
rect 66665 6335 66671 6369
rect 66111 6320 66671 6335
rect 66061 6310 66128 6320
rect 66615 6319 66671 6320
rect 66777 6281 66811 6409
rect 65355 6269 65401 6281
rect 65355 6093 65361 6269
rect 65395 6093 65401 6269
rect 65355 6081 65401 6093
rect 65473 6269 65519 6281
rect 65473 6093 65479 6269
rect 65513 6093 65519 6269
rect 65473 6081 65519 6093
rect 65775 6269 65821 6281
rect 65478 5787 65512 6081
rect 65775 5893 65781 6269
rect 65815 5893 65821 6269
rect 65775 5881 65821 5893
rect 65893 6269 65939 6281
rect 65893 5893 65899 6269
rect 65933 5893 65939 6269
rect 65893 5881 65939 5893
rect 66011 6269 66057 6281
rect 66011 5893 66017 6269
rect 66051 5893 66057 6269
rect 66011 5881 66057 5893
rect 66129 6269 66175 6281
rect 66129 5893 66135 6269
rect 66169 5893 66175 6269
rect 66129 5881 66175 5893
rect 66247 6269 66293 6281
rect 66247 5893 66253 6269
rect 66287 5893 66293 6269
rect 66653 6269 66699 6281
rect 66653 6093 66659 6269
rect 66693 6093 66699 6269
rect 66653 6081 66699 6093
rect 66771 6269 66817 6281
rect 66771 6093 66777 6269
rect 66811 6093 66817 6269
rect 66771 6081 66817 6093
rect 66247 5881 66293 5893
rect 66135 5787 66169 5881
rect 66659 5787 66692 6081
rect 65478 5755 66692 5787
rect 65844 5731 66250 5755
rect 65844 5608 65956 5731
rect 66130 5608 66250 5731
rect 65844 5564 66250 5608
rect 65858 4737 66303 4743
rect 65858 4537 65870 4737
rect 66291 4537 66303 4737
rect 65858 4531 66026 4537
rect 66016 4463 66026 4531
rect 66158 4531 66303 4537
rect 66158 4463 66168 4531
rect 66026 4423 66158 4463
rect 66025 4357 66158 4423
rect 64199 4041 64876 4044
rect 61785 3878 61831 3890
rect 63723 4029 63769 4041
rect 61083 3836 61117 3878
rect 61319 3836 61353 3878
rect 61083 3808 61353 3836
rect 61437 3837 61471 3878
rect 61673 3837 61707 3878
rect 61437 3808 61707 3837
rect 61083 3760 61117 3808
rect 61083 3730 61146 3760
rect 61111 3638 61146 3730
rect 61618 3700 61718 3721
rect 61618 3646 61632 3700
rect 61697 3646 61718 3700
rect 61618 3641 61718 3646
rect 61791 3695 61825 3878
rect 61791 3641 61900 3695
rect 61111 3602 61338 3638
rect 61111 3495 61146 3602
rect 61272 3568 61338 3602
rect 61272 3534 61288 3568
rect 61322 3534 61338 3568
rect 61619 3626 61716 3641
rect 61619 3559 61676 3626
rect 61272 3528 61338 3534
rect 61513 3523 61782 3559
rect 61513 3495 61546 3523
rect 61749 3495 61782 3523
rect 61866 3495 61900 3641
rect 63558 3692 63662 3700
rect 63558 3591 63568 3692
rect 63654 3609 63664 3692
rect 63723 3653 63729 4029
rect 63763 3653 63769 4029
rect 63723 3641 63769 3653
rect 63841 4029 63887 4041
rect 63841 3653 63847 4029
rect 63881 3653 63887 4029
rect 63841 3641 63887 3653
rect 63959 4029 64005 4041
rect 63959 3653 63965 4029
rect 63999 3680 64005 4029
rect 64076 4029 64122 4041
rect 64076 3853 64082 4029
rect 64116 3853 64122 4029
rect 64076 3846 64122 3853
rect 64194 4029 64876 4041
rect 64194 3853 64200 4029
rect 64234 4016 64876 4029
rect 64234 3853 64240 4016
rect 64484 3936 64876 4016
rect 65354 4314 66827 4357
rect 65354 4011 65388 4314
rect 65720 4211 65754 4314
rect 65956 4211 65990 4314
rect 66192 4211 66226 4314
rect 66428 4211 66462 4314
rect 65714 4199 65760 4211
rect 65230 3999 65276 4011
rect 64076 3841 64125 3846
rect 64194 3841 64240 3853
rect 64082 3680 64125 3841
rect 65230 3823 65236 3999
rect 65270 3823 65276 3999
rect 65230 3811 65276 3823
rect 65348 3999 65394 4011
rect 65348 3823 65354 3999
rect 65388 3823 65394 3999
rect 65348 3811 65394 3823
rect 65466 3999 65512 4011
rect 65466 3823 65472 3999
rect 65506 3823 65512 3999
rect 65466 3811 65512 3823
rect 65584 3999 65630 4011
rect 65714 3999 65720 4199
rect 65584 3823 65590 3999
rect 65624 3823 65720 3999
rect 65754 3823 65760 4199
rect 65584 3811 65630 3823
rect 65714 3811 65760 3823
rect 65832 4199 65878 4211
rect 65832 3823 65838 4199
rect 65872 3823 65878 4199
rect 65832 3811 65878 3823
rect 65950 4199 65996 4211
rect 65950 3823 65956 4199
rect 65990 3823 65996 4199
rect 65950 3811 65996 3823
rect 66068 4199 66114 4211
rect 66068 3823 66074 4199
rect 66108 3823 66114 4199
rect 66068 3811 66114 3823
rect 66186 4199 66232 4211
rect 66186 3823 66192 4199
rect 66226 3823 66232 4199
rect 66186 3811 66232 3823
rect 66304 4199 66350 4211
rect 66304 3823 66310 4199
rect 66344 3823 66350 4199
rect 66304 3811 66350 3823
rect 66422 4199 66468 4211
rect 66422 3823 66428 4199
rect 66462 3999 66468 4199
rect 66793 4011 66827 4314
rect 67334 4234 67470 4254
rect 67334 4172 67370 4234
rect 67430 4172 67470 4234
rect 67334 4144 67470 4172
rect 67030 4114 68007 4144
rect 66551 3999 66597 4011
rect 66462 3823 66557 3999
rect 66591 3823 66597 3999
rect 66422 3811 66468 3823
rect 66551 3811 66597 3823
rect 66669 3999 66715 4011
rect 66669 3823 66675 3999
rect 66709 3823 66715 3999
rect 66669 3811 66715 3823
rect 66787 3999 66833 4011
rect 66787 3823 66793 3999
rect 66827 3823 66833 3999
rect 66787 3811 66833 3823
rect 66905 3999 66951 4011
rect 67030 4008 67062 4114
rect 67266 4008 67298 4114
rect 67502 4008 67534 4114
rect 67738 4008 67770 4114
rect 67973 4008 68007 4114
rect 66905 3823 66911 3999
rect 66945 3823 66951 3999
rect 66905 3811 66951 3823
rect 67023 3996 67069 4008
rect 67023 3820 67029 3996
rect 67063 3820 67069 3996
rect 65236 3777 65270 3811
rect 65838 3777 65872 3811
rect 66074 3777 66108 3811
rect 65236 3742 65395 3777
rect 65838 3742 66108 3777
rect 66675 3777 66709 3811
rect 66911 3777 66945 3811
rect 67023 3808 67069 3820
rect 67141 3996 67187 4008
rect 67141 3820 67147 3996
rect 67181 3820 67187 3996
rect 67141 3808 67187 3820
rect 67259 3996 67305 4008
rect 67259 3820 67265 3996
rect 67299 3820 67305 3996
rect 67259 3808 67305 3820
rect 67377 3996 67423 4008
rect 67377 3820 67383 3996
rect 67417 3820 67423 3996
rect 67377 3808 67423 3820
rect 67495 3996 67541 4008
rect 67495 3820 67501 3996
rect 67535 3820 67541 3996
rect 67495 3808 67541 3820
rect 67613 3996 67659 4008
rect 67613 3820 67619 3996
rect 67653 3820 67659 3996
rect 67613 3808 67659 3820
rect 67731 3996 67777 4008
rect 67731 3820 67737 3996
rect 67771 3820 67777 3996
rect 67731 3808 67777 3820
rect 67849 3996 67895 4008
rect 67849 3820 67855 3996
rect 67889 3820 67895 3996
rect 67849 3808 67895 3820
rect 67967 3996 68013 4008
rect 67967 3820 67973 3996
rect 68007 3820 68013 3996
rect 67967 3808 68013 3820
rect 68085 3996 68131 4008
rect 68085 3820 68091 3996
rect 68125 3820 68131 3996
rect 68085 3808 68131 3820
rect 66675 3742 66945 3777
rect 63999 3653 64125 3680
rect 63959 3641 64125 3653
rect 63965 3637 64125 3641
rect 63654 3603 63838 3609
rect 63654 3591 63788 3603
rect 63558 3569 63788 3591
rect 63822 3569 63838 3603
rect 63558 3553 63838 3569
rect 63890 3603 63956 3609
rect 63890 3569 63906 3603
rect 63940 3569 63956 3603
rect 63890 3524 63956 3569
rect 63335 3518 63956 3524
rect 60987 3483 61033 3495
rect 60987 3307 60993 3483
rect 61027 3307 61033 3483
rect 60987 3295 61033 3307
rect 61105 3483 61151 3495
rect 61105 3307 61111 3483
rect 61145 3307 61151 3483
rect 61105 3295 61151 3307
rect 61223 3483 61269 3495
rect 61223 3307 61229 3483
rect 61263 3307 61269 3483
rect 61223 3295 61269 3307
rect 61341 3483 61387 3495
rect 61341 3307 61347 3483
rect 61381 3428 61387 3483
rect 61506 3483 61552 3495
rect 61506 3428 61512 3483
rect 61381 3340 61512 3428
rect 61381 3307 61387 3340
rect 61341 3295 61387 3307
rect 61506 3307 61512 3340
rect 61546 3307 61552 3483
rect 61506 3295 61552 3307
rect 61624 3483 61670 3495
rect 61624 3307 61630 3483
rect 61664 3307 61670 3483
rect 61624 3295 61670 3307
rect 61742 3483 61788 3495
rect 61742 3307 61748 3483
rect 61782 3307 61788 3483
rect 61742 3295 61788 3307
rect 61860 3483 61906 3495
rect 61860 3307 61866 3483
rect 61900 3307 61906 3483
rect 63330 3458 63340 3518
rect 63425 3516 63956 3518
rect 63425 3484 63957 3516
rect 64049 3500 64125 3637
rect 63425 3458 63435 3484
rect 63335 3451 63430 3458
rect 64045 3440 64055 3500
rect 64117 3440 64127 3500
rect 64782 3468 65223 3531
rect 65290 3468 65300 3531
rect 61860 3295 61906 3307
rect 60993 3256 61027 3295
rect 61229 3256 61263 3295
rect 60993 3220 61263 3256
rect 61630 3257 61663 3295
rect 61866 3257 61899 3295
rect 61630 3221 61899 3257
rect 60993 3219 61159 3220
rect 61027 3140 61159 3219
rect 61017 3032 61027 3140
rect 61159 3032 61169 3140
rect 61048 2895 61054 3032
rect 61121 2895 61127 3032
rect 61048 2883 61127 2895
rect 57631 2658 58608 2688
rect 60825 2686 60888 2703
rect 60750 2682 60888 2686
rect 57631 2552 57663 2658
rect 57867 2552 57899 2658
rect 58103 2552 58135 2658
rect 58339 2552 58371 2658
rect 58574 2552 58608 2658
rect 58918 2648 60888 2682
rect 58916 2619 60888 2648
rect 58916 2603 58962 2619
rect 60750 2617 60888 2619
rect 57624 2540 57670 2552
rect 57624 2364 57630 2540
rect 57664 2364 57670 2540
rect 57624 2352 57670 2364
rect 57742 2540 57788 2552
rect 57742 2364 57748 2540
rect 57782 2364 57788 2540
rect 57742 2352 57788 2364
rect 57860 2540 57906 2552
rect 57860 2364 57866 2540
rect 57900 2364 57906 2540
rect 57860 2352 57906 2364
rect 57978 2540 58024 2552
rect 57978 2364 57984 2540
rect 58018 2364 58024 2540
rect 57978 2352 58024 2364
rect 58096 2540 58142 2552
rect 58096 2364 58102 2540
rect 58136 2364 58142 2540
rect 58096 2352 58142 2364
rect 58214 2540 58260 2552
rect 58214 2364 58220 2540
rect 58254 2364 58260 2540
rect 58214 2352 58260 2364
rect 58332 2540 58378 2552
rect 58332 2364 58338 2540
rect 58372 2364 58378 2540
rect 58332 2352 58378 2364
rect 58450 2540 58496 2552
rect 58450 2364 58456 2540
rect 58490 2364 58496 2540
rect 58450 2352 58496 2364
rect 58568 2540 58614 2552
rect 58568 2364 58574 2540
rect 58608 2364 58614 2540
rect 58568 2352 58614 2364
rect 58686 2540 58732 2552
rect 58686 2364 58692 2540
rect 58726 2364 58732 2540
rect 58686 2352 58732 2364
rect 57747 2258 57783 2352
rect 57983 2258 58019 2352
rect 58219 2259 58255 2352
rect 58381 2304 58447 2311
rect 58381 2270 58397 2304
rect 58431 2270 58447 2304
rect 58381 2259 58447 2270
rect 58219 2258 58447 2259
rect 57747 2229 58447 2258
rect 57747 2228 58329 2229
rect 57867 2115 57901 2228
rect 58263 2187 58329 2228
rect 58263 2153 58279 2187
rect 58313 2153 58329 2187
rect 58263 2146 58329 2153
rect 58691 2134 58726 2352
rect 58915 2151 58962 2603
rect 61811 2610 61890 2622
rect 61811 2495 61817 2610
rect 61884 2495 61890 2610
rect 59874 2387 59884 2495
rect 60016 2387 60026 2495
rect 61772 2387 61782 2495
rect 61914 2387 61924 2495
rect 59884 2347 60016 2387
rect 61782 2347 61914 2387
rect 59883 2281 60016 2347
rect 61781 2281 61914 2347
rect 59212 2238 60685 2281
rect 58915 2135 58961 2151
rect 58880 2134 58961 2135
rect 58691 2119 58961 2134
rect 58337 2115 58961 2119
rect 57861 2103 57907 2115
rect 57596 1625 57606 1743
rect 57724 1711 57734 1743
rect 57861 1727 57867 2103
rect 57901 1727 57907 2103
rect 57861 1715 57907 1727
rect 57979 2103 58025 2115
rect 57979 1727 57985 2103
rect 58019 1727 58025 2103
rect 57979 1715 58025 1727
rect 58097 2103 58143 2115
rect 58097 1727 58103 2103
rect 58137 1751 58143 2103
rect 58214 2103 58260 2115
rect 58214 1927 58220 2103
rect 58254 1927 58260 2103
rect 58214 1915 58260 1927
rect 58332 2103 58961 2115
rect 58332 1927 58338 2103
rect 58372 2091 58961 2103
rect 58372 2090 58614 2091
rect 58372 1927 58378 2090
rect 58880 2089 58961 2091
rect 59212 1935 59246 2238
rect 59578 2135 59612 2238
rect 59814 2135 59848 2238
rect 60050 2135 60084 2238
rect 60286 2135 60320 2238
rect 59572 2123 59618 2135
rect 58332 1915 58378 1927
rect 59088 1923 59134 1935
rect 58220 1799 58255 1915
rect 58351 1799 58459 1809
rect 58220 1751 58351 1799
rect 58459 1768 58608 1774
rect 58137 1727 58351 1751
rect 58097 1715 58351 1727
rect 58103 1711 58351 1715
rect 57724 1683 57739 1711
rect 57724 1677 57976 1683
rect 57724 1643 57926 1677
rect 57960 1643 57976 1677
rect 57724 1627 57976 1643
rect 58028 1677 58094 1683
rect 58028 1643 58044 1677
rect 58078 1643 58094 1677
rect 58277 1667 58351 1711
rect 58596 1701 58608 1768
rect 59088 1747 59094 1923
rect 59128 1747 59134 1923
rect 59088 1735 59134 1747
rect 59206 1923 59252 1935
rect 59206 1747 59212 1923
rect 59246 1747 59252 1923
rect 59206 1735 59252 1747
rect 59324 1923 59370 1935
rect 59324 1747 59330 1923
rect 59364 1747 59370 1923
rect 59324 1735 59370 1747
rect 59442 1923 59488 1935
rect 59572 1923 59578 2123
rect 59442 1747 59448 1923
rect 59482 1747 59578 1923
rect 59612 1747 59618 2123
rect 59442 1735 59488 1747
rect 59572 1735 59618 1747
rect 59690 2123 59736 2135
rect 59690 1747 59696 2123
rect 59730 1747 59736 2123
rect 59690 1735 59736 1747
rect 59808 2123 59854 2135
rect 59808 1747 59814 2123
rect 59848 1747 59854 2123
rect 59808 1735 59854 1747
rect 59926 2123 59972 2135
rect 59926 1747 59932 2123
rect 59966 1747 59972 2123
rect 59926 1735 59972 1747
rect 60044 2123 60090 2135
rect 60044 1747 60050 2123
rect 60084 1747 60090 2123
rect 60044 1735 60090 1747
rect 60162 2123 60208 2135
rect 60162 1747 60168 2123
rect 60202 1747 60208 2123
rect 60162 1735 60208 1747
rect 60280 2123 60326 2135
rect 60280 1747 60286 2123
rect 60320 1923 60326 2123
rect 60651 1935 60685 2238
rect 61110 2238 62583 2281
rect 61110 1935 61144 2238
rect 61476 2135 61510 2238
rect 61712 2135 61746 2238
rect 61948 2135 61982 2238
rect 62184 2135 62218 2238
rect 61470 2123 61516 2135
rect 60409 1923 60455 1935
rect 60320 1747 60415 1923
rect 60449 1747 60455 1923
rect 60280 1735 60326 1747
rect 60409 1735 60455 1747
rect 60527 1923 60573 1935
rect 60527 1747 60533 1923
rect 60567 1747 60573 1923
rect 60527 1735 60573 1747
rect 60645 1923 60691 1935
rect 60645 1747 60651 1923
rect 60685 1747 60691 1923
rect 60645 1735 60691 1747
rect 60763 1923 60809 1935
rect 60763 1747 60769 1923
rect 60803 1747 60809 1923
rect 60763 1735 60809 1747
rect 60986 1923 61032 1935
rect 60986 1747 60992 1923
rect 61026 1747 61032 1923
rect 60986 1735 61032 1747
rect 61104 1923 61150 1935
rect 61104 1747 61110 1923
rect 61144 1747 61150 1923
rect 61104 1735 61150 1747
rect 61222 1923 61268 1935
rect 61222 1747 61228 1923
rect 61262 1747 61268 1923
rect 61222 1735 61268 1747
rect 61340 1923 61386 1935
rect 61470 1923 61476 2123
rect 61340 1747 61346 1923
rect 61380 1747 61476 1923
rect 61510 1747 61516 2123
rect 61340 1735 61386 1747
rect 61470 1735 61516 1747
rect 61588 2123 61634 2135
rect 61588 1747 61594 2123
rect 61628 1747 61634 2123
rect 61588 1735 61634 1747
rect 61706 2123 61752 2135
rect 61706 1747 61712 2123
rect 61746 1747 61752 2123
rect 61706 1735 61752 1747
rect 61824 2123 61870 2135
rect 61824 1747 61830 2123
rect 61864 1747 61870 2123
rect 61824 1735 61870 1747
rect 61942 2123 61988 2135
rect 61942 1747 61948 2123
rect 61982 1747 61988 2123
rect 61942 1735 61988 1747
rect 62060 2123 62106 2135
rect 62060 1747 62066 2123
rect 62100 1747 62106 2123
rect 62060 1735 62106 1747
rect 62178 2123 62224 2135
rect 62178 1747 62184 2123
rect 62218 1923 62224 2123
rect 62549 1935 62583 2238
rect 62307 1923 62353 1935
rect 62218 1747 62313 1923
rect 62347 1747 62353 1923
rect 62178 1735 62224 1747
rect 62307 1735 62353 1747
rect 62425 1923 62471 1935
rect 62425 1747 62431 1923
rect 62465 1747 62471 1923
rect 62425 1735 62471 1747
rect 62543 1923 62589 1935
rect 62543 1747 62549 1923
rect 62583 1747 62589 1923
rect 62543 1735 62589 1747
rect 62661 1923 62707 1935
rect 62661 1747 62667 1923
rect 62701 1747 62707 1923
rect 62661 1735 62707 1747
rect 58459 1695 58608 1701
rect 59094 1701 59128 1735
rect 59696 1701 59730 1735
rect 59932 1701 59966 1735
rect 58351 1657 58459 1667
rect 59094 1666 59253 1701
rect 59696 1666 59966 1701
rect 60533 1701 60567 1735
rect 60769 1701 60803 1735
rect 60533 1666 60803 1701
rect 60992 1701 61026 1735
rect 61594 1701 61628 1735
rect 61830 1701 61864 1735
rect 60992 1666 61151 1701
rect 61594 1666 61864 1701
rect 62431 1701 62465 1735
rect 62667 1701 62701 1735
rect 62431 1666 62701 1701
rect 57724 1625 57739 1627
rect 57639 1611 57739 1625
rect 57639 1568 57739 1569
rect 57260 1547 57739 1568
rect 58028 1547 58094 1643
rect 57260 1499 58094 1547
rect 57260 1470 57739 1499
rect 57260 1468 57365 1470
rect 57639 1469 57739 1470
rect 57093 1283 57103 1362
rect 57196 1283 57206 1362
rect 58095 1346 58174 1358
rect 57104 109 57197 1283
rect 58095 1254 58101 1346
rect 58022 1234 58101 1254
rect 58168 1254 58174 1346
rect 58168 1234 58242 1254
rect 58022 1126 58066 1234
rect 58198 1126 58242 1234
rect 58022 1084 58242 1126
rect 57626 1054 58603 1084
rect 57626 948 57658 1054
rect 57862 948 57894 1054
rect 58098 948 58130 1054
rect 58334 948 58366 1054
rect 58569 948 58603 1054
rect 57619 936 57665 948
rect 57619 760 57625 936
rect 57659 760 57665 936
rect 57619 748 57665 760
rect 57737 936 57783 948
rect 57737 760 57743 936
rect 57777 760 57783 936
rect 57737 748 57783 760
rect 57855 936 57901 948
rect 57855 760 57861 936
rect 57895 760 57901 936
rect 57855 748 57901 760
rect 57973 936 58019 948
rect 57973 760 57979 936
rect 58013 760 58019 936
rect 57973 748 58019 760
rect 58091 936 58137 948
rect 58091 760 58097 936
rect 58131 760 58137 936
rect 58091 748 58137 760
rect 58209 936 58255 948
rect 58209 760 58215 936
rect 58249 760 58255 936
rect 58209 748 58255 760
rect 58327 936 58373 948
rect 58327 760 58333 936
rect 58367 760 58373 936
rect 58327 748 58373 760
rect 58445 936 58491 948
rect 58445 760 58451 936
rect 58485 760 58491 936
rect 58445 748 58491 760
rect 58563 936 58609 948
rect 58563 760 58569 936
rect 58603 760 58609 936
rect 58563 748 58609 760
rect 58681 936 58727 948
rect 58681 760 58687 936
rect 58721 760 58727 936
rect 58681 748 58727 760
rect 59219 882 59253 1666
rect 59932 1604 59966 1666
rect 59521 1566 60263 1604
rect 59521 1442 59555 1566
rect 59757 1442 59791 1566
rect 59993 1442 60027 1566
rect 60229 1442 60263 1566
rect 60519 1459 60529 1525
rect 60592 1459 60602 1525
rect 59515 1430 59561 1442
rect 59515 1054 59521 1430
rect 59555 1054 59561 1430
rect 59515 1042 59561 1054
rect 59633 1430 59679 1442
rect 59633 1054 59639 1430
rect 59673 1054 59679 1430
rect 59633 1042 59679 1054
rect 59751 1430 59797 1442
rect 59751 1054 59757 1430
rect 59791 1054 59797 1430
rect 59751 1042 59797 1054
rect 59869 1430 59915 1442
rect 59869 1054 59875 1430
rect 59909 1054 59915 1430
rect 59869 1042 59915 1054
rect 59987 1430 60033 1442
rect 59987 1054 59993 1430
rect 60027 1054 60033 1430
rect 59987 1042 60033 1054
rect 60105 1430 60151 1442
rect 60105 1054 60111 1430
rect 60145 1054 60151 1430
rect 60105 1042 60151 1054
rect 60223 1430 60269 1442
rect 60223 1054 60229 1430
rect 60263 1054 60269 1430
rect 60223 1042 60269 1054
rect 60635 883 60669 1666
rect 60362 882 60669 883
rect 59219 877 59535 882
rect 60249 877 60669 882
rect 59219 866 59602 877
rect 59219 839 59551 866
rect 57742 654 57778 748
rect 57978 654 58014 748
rect 58214 655 58250 748
rect 58376 700 58442 707
rect 58376 666 58392 700
rect 58426 666 58442 700
rect 58376 655 58442 666
rect 58214 654 58442 655
rect 57742 625 58442 654
rect 57742 624 58324 625
rect 57862 511 57896 624
rect 58258 583 58324 624
rect 58258 549 58274 583
rect 58308 549 58324 583
rect 58258 542 58324 549
rect 58686 515 58721 748
rect 59219 710 59253 839
rect 59535 832 59551 839
rect 59585 832 59602 866
rect 59535 826 59602 832
rect 60182 866 60669 877
rect 60182 832 60199 866
rect 60233 839 60669 866
rect 60233 832 60249 839
rect 60362 838 60669 839
rect 60182 826 60249 832
rect 59360 799 59416 811
rect 59360 765 59366 799
rect 59400 798 59416 799
rect 60473 798 60529 810
rect 59400 782 59867 798
rect 59400 765 59817 782
rect 59360 749 59817 765
rect 59801 748 59817 749
rect 59851 748 59867 782
rect 59801 741 59867 748
rect 59919 783 60489 798
rect 59919 749 59935 783
rect 59969 764 60489 783
rect 60523 764 60529 798
rect 59969 749 60529 764
rect 59919 739 59986 749
rect 60473 748 60529 749
rect 60635 710 60669 838
rect 61117 882 61151 1666
rect 61830 1604 61864 1666
rect 61419 1566 62161 1604
rect 61419 1442 61453 1566
rect 61655 1442 61689 1566
rect 61891 1442 61925 1566
rect 62127 1442 62161 1566
rect 61413 1430 61459 1442
rect 61413 1054 61419 1430
rect 61453 1054 61459 1430
rect 61413 1042 61459 1054
rect 61531 1430 61577 1442
rect 61531 1054 61537 1430
rect 61571 1054 61577 1430
rect 61531 1042 61577 1054
rect 61649 1430 61695 1442
rect 61649 1054 61655 1430
rect 61689 1054 61695 1430
rect 61649 1042 61695 1054
rect 61767 1430 61813 1442
rect 61767 1054 61773 1430
rect 61807 1054 61813 1430
rect 61767 1042 61813 1054
rect 61885 1430 61931 1442
rect 61885 1054 61891 1430
rect 61925 1054 61931 1430
rect 61885 1042 61931 1054
rect 62003 1430 62049 1442
rect 62003 1054 62009 1430
rect 62043 1054 62049 1430
rect 62003 1042 62049 1054
rect 62121 1430 62167 1442
rect 62121 1054 62127 1430
rect 62161 1054 62167 1430
rect 62121 1042 62167 1054
rect 62533 883 62567 1666
rect 63794 1634 63930 1654
rect 63794 1572 63830 1634
rect 63890 1572 63930 1634
rect 63794 1544 63930 1572
rect 63490 1514 64467 1544
rect 62145 882 62214 883
rect 62260 882 62567 883
rect 61117 877 61433 882
rect 62145 878 62567 882
rect 61117 866 61500 877
rect 61117 839 61449 866
rect 61117 710 61151 839
rect 61433 832 61449 839
rect 61483 832 61500 866
rect 61433 826 61500 832
rect 62078 867 62567 878
rect 62078 833 62095 867
rect 62129 839 62567 867
rect 62129 833 62145 839
rect 62260 838 62567 839
rect 62078 827 62145 833
rect 61258 799 61314 811
rect 61258 765 61264 799
rect 61298 798 61314 799
rect 62371 798 62427 810
rect 61298 782 61765 798
rect 61298 765 61715 782
rect 61258 749 61715 765
rect 61699 748 61715 749
rect 61749 748 61765 782
rect 61699 741 61765 748
rect 61817 783 62387 798
rect 61817 749 61833 783
rect 61867 764 62387 783
rect 62421 764 62427 798
rect 61867 749 62427 764
rect 61817 739 61884 749
rect 62371 748 62427 749
rect 62533 710 62567 838
rect 62648 1488 62715 1512
rect 62648 1454 62665 1488
rect 62699 1454 62715 1488
rect 58332 511 58721 515
rect 57856 499 57902 511
rect 57856 123 57862 499
rect 57896 123 57902 499
rect 57856 111 57902 123
rect 57974 499 58020 511
rect 57974 123 57980 499
rect 58014 123 58020 499
rect 57974 111 58020 123
rect 58092 499 58138 511
rect 58092 123 58098 499
rect 58132 147 58138 499
rect 58209 499 58255 511
rect 58209 323 58215 499
rect 58249 323 58255 499
rect 58209 311 58255 323
rect 58327 499 58721 511
rect 59213 698 59259 710
rect 59213 522 59219 698
rect 59253 522 59259 698
rect 59213 510 59259 522
rect 59331 698 59377 710
rect 59331 522 59337 698
rect 59371 522 59377 698
rect 59331 510 59377 522
rect 59633 698 59679 710
rect 58327 323 58333 499
rect 58367 486 58721 499
rect 58367 323 58373 486
rect 58643 483 58721 486
rect 58643 431 58653 483
rect 58716 431 58726 483
rect 58648 425 58721 431
rect 58327 311 58373 323
rect 58215 195 58250 311
rect 59336 216 59370 510
rect 59633 322 59639 698
rect 59673 322 59679 698
rect 59633 310 59679 322
rect 59751 698 59797 710
rect 59751 322 59757 698
rect 59791 322 59797 698
rect 59751 310 59797 322
rect 59869 698 59915 710
rect 59869 322 59875 698
rect 59909 322 59915 698
rect 59869 310 59915 322
rect 59987 698 60033 710
rect 59987 322 59993 698
rect 60027 322 60033 698
rect 59987 310 60033 322
rect 60105 698 60151 710
rect 60105 322 60111 698
rect 60145 322 60151 698
rect 60511 698 60557 710
rect 60511 522 60517 698
rect 60551 522 60557 698
rect 60511 510 60557 522
rect 60629 698 60675 710
rect 60629 522 60635 698
rect 60669 522 60675 698
rect 60629 510 60675 522
rect 61111 698 61157 710
rect 61111 522 61117 698
rect 61151 522 61157 698
rect 61111 510 61157 522
rect 61229 698 61275 710
rect 61229 522 61235 698
rect 61269 522 61275 698
rect 61229 510 61275 522
rect 61531 698 61577 710
rect 60105 310 60151 322
rect 59993 216 60027 310
rect 60517 216 60550 510
rect 58346 195 58454 205
rect 58215 147 58346 195
rect 59336 184 60550 216
rect 61234 216 61268 510
rect 61531 322 61537 698
rect 61571 322 61577 698
rect 61531 310 61577 322
rect 61649 698 61695 710
rect 61649 322 61655 698
rect 61689 322 61695 698
rect 61649 310 61695 322
rect 61767 698 61813 710
rect 61767 322 61773 698
rect 61807 322 61813 698
rect 61767 310 61813 322
rect 61885 698 61931 710
rect 61885 322 61891 698
rect 61925 322 61931 698
rect 61885 310 61931 322
rect 62003 698 62049 710
rect 62003 322 62009 698
rect 62043 322 62049 698
rect 62409 698 62455 710
rect 62409 522 62415 698
rect 62449 522 62455 698
rect 62409 510 62455 522
rect 62527 698 62573 710
rect 62527 522 62533 698
rect 62567 522 62573 698
rect 62527 510 62573 522
rect 62003 310 62049 322
rect 61891 216 61925 310
rect 62415 216 62448 510
rect 61234 184 62448 216
rect 58454 151 58599 157
rect 58132 123 58346 147
rect 58092 111 58346 123
rect 57104 107 57689 109
rect 58098 107 58346 111
rect 57104 79 57734 107
rect 57104 73 57971 79
rect 57104 39 57921 73
rect 57955 39 57971 73
rect 57104 23 57971 39
rect 58023 73 58089 79
rect 58023 39 58039 73
rect 58073 39 58089 73
rect 58272 63 58346 107
rect 58587 84 58599 151
rect 59829 99 59961 184
rect 61727 99 61859 184
rect 58454 78 58599 84
rect 58346 53 58454 63
rect 57104 7 57734 23
rect 57104 3 57689 7
rect 57104 2 57205 3
rect 57634 -46 57734 -35
rect 57598 -152 57608 -46
rect 57720 -57 57734 -46
rect 58023 -57 58089 39
rect 59819 -9 59829 99
rect 59961 -9 59971 99
rect 61717 -9 61727 99
rect 61859 -9 61869 99
rect 62648 71 62715 1454
rect 63490 1408 63522 1514
rect 63726 1408 63758 1514
rect 63962 1408 63994 1514
rect 64198 1408 64230 1514
rect 64433 1408 64467 1514
rect 63483 1396 63529 1408
rect 63483 1220 63489 1396
rect 63523 1220 63529 1396
rect 63483 1208 63529 1220
rect 63601 1396 63647 1408
rect 63601 1220 63607 1396
rect 63641 1220 63647 1396
rect 63601 1208 63647 1220
rect 63719 1396 63765 1408
rect 63719 1220 63725 1396
rect 63759 1220 63765 1396
rect 63719 1208 63765 1220
rect 63837 1396 63883 1408
rect 63837 1220 63843 1396
rect 63877 1220 63883 1396
rect 63837 1208 63883 1220
rect 63955 1396 64001 1408
rect 63955 1220 63961 1396
rect 63995 1220 64001 1396
rect 63955 1208 64001 1220
rect 64073 1396 64119 1408
rect 64073 1220 64079 1396
rect 64113 1220 64119 1396
rect 64073 1208 64119 1220
rect 64191 1396 64237 1408
rect 64191 1220 64197 1396
rect 64231 1220 64237 1396
rect 64191 1208 64237 1220
rect 64309 1396 64355 1408
rect 64309 1220 64315 1396
rect 64349 1220 64355 1396
rect 64309 1208 64355 1220
rect 64427 1396 64473 1408
rect 64427 1220 64433 1396
rect 64467 1220 64473 1396
rect 64427 1208 64473 1220
rect 64545 1396 64591 1408
rect 64545 1220 64551 1396
rect 64585 1220 64591 1396
rect 64545 1208 64591 1220
rect 63606 1114 63642 1208
rect 63842 1114 63878 1208
rect 64078 1115 64114 1208
rect 64240 1160 64306 1167
rect 64240 1126 64256 1160
rect 64290 1126 64306 1160
rect 64240 1115 64306 1126
rect 64078 1114 64306 1115
rect 63606 1085 64306 1114
rect 63606 1084 64188 1085
rect 62776 1025 62932 1031
rect 62776 927 62788 1025
rect 62920 927 62932 1025
rect 63726 971 63760 1084
rect 64122 1043 64188 1084
rect 64122 1009 64138 1043
rect 64172 1009 64188 1043
rect 64122 1002 64188 1009
rect 64550 975 64585 1208
rect 64196 974 64731 975
rect 64782 974 64877 3468
rect 65361 2958 65395 3742
rect 66074 3680 66108 3742
rect 65663 3642 66405 3680
rect 65473 3471 65483 3539
rect 65538 3471 65548 3539
rect 65663 3518 65697 3642
rect 65899 3518 65933 3642
rect 66135 3518 66169 3642
rect 66371 3518 66405 3642
rect 65657 3506 65703 3518
rect 65657 3130 65663 3506
rect 65697 3130 65703 3506
rect 65657 3118 65703 3130
rect 65775 3506 65821 3518
rect 65775 3130 65781 3506
rect 65815 3130 65821 3506
rect 65775 3118 65821 3130
rect 65893 3506 65939 3518
rect 65893 3130 65899 3506
rect 65933 3130 65939 3506
rect 65893 3118 65939 3130
rect 66011 3506 66057 3518
rect 66011 3130 66017 3506
rect 66051 3130 66057 3506
rect 66011 3118 66057 3130
rect 66129 3506 66175 3518
rect 66129 3130 66135 3506
rect 66169 3130 66175 3506
rect 66129 3118 66175 3130
rect 66247 3506 66293 3518
rect 66247 3130 66253 3506
rect 66287 3130 66293 3506
rect 66247 3118 66293 3130
rect 66365 3506 66411 3518
rect 66365 3130 66371 3506
rect 66405 3130 66411 3506
rect 66531 3301 66605 3313
rect 66527 3210 66537 3301
rect 66599 3210 66609 3301
rect 66531 3198 66605 3210
rect 66365 3118 66411 3130
rect 66777 2959 66811 3742
rect 67146 3714 67182 3808
rect 67382 3714 67418 3808
rect 67618 3715 67654 3808
rect 67780 3760 67846 3767
rect 67780 3726 67796 3760
rect 67830 3726 67846 3760
rect 67780 3715 67846 3726
rect 67618 3714 67846 3715
rect 67146 3685 67846 3714
rect 67146 3684 67728 3685
rect 66872 3652 66948 3657
rect 66869 3596 66879 3652
rect 66932 3651 66948 3652
rect 66932 3596 67198 3651
rect 66872 3591 67198 3596
rect 66993 3549 67084 3554
rect 66993 3460 67003 3549
rect 67076 3460 67084 3549
rect 66993 3448 67084 3460
rect 67030 3054 67084 3448
rect 67144 3139 67198 3591
rect 67266 3571 67300 3684
rect 67662 3643 67728 3684
rect 67662 3609 67678 3643
rect 67712 3609 67728 3643
rect 67662 3602 67728 3609
rect 68090 3575 68125 3808
rect 67736 3571 68125 3575
rect 67260 3559 67306 3571
rect 67260 3183 67266 3559
rect 67300 3183 67306 3559
rect 67260 3171 67306 3183
rect 67378 3559 67424 3571
rect 67378 3183 67384 3559
rect 67418 3183 67424 3559
rect 67378 3171 67424 3183
rect 67496 3559 67542 3571
rect 67496 3183 67502 3559
rect 67536 3210 67542 3559
rect 67613 3559 67659 3571
rect 67613 3383 67619 3559
rect 67653 3383 67659 3559
rect 67613 3376 67659 3383
rect 67731 3559 68125 3571
rect 67731 3383 67737 3559
rect 67771 3546 68125 3559
rect 67771 3383 67777 3546
rect 67950 3457 68125 3546
rect 67994 3456 68125 3457
rect 67613 3371 67662 3376
rect 67731 3371 67777 3383
rect 67619 3210 67662 3371
rect 67536 3183 67662 3210
rect 67496 3171 67662 3183
rect 67502 3167 67662 3171
rect 67144 3133 67375 3139
rect 67144 3099 67325 3133
rect 67359 3099 67375 3133
rect 67144 3083 67375 3099
rect 67427 3133 67493 3139
rect 67427 3099 67443 3133
rect 67477 3099 67493 3133
rect 67427 3054 67493 3099
rect 67030 3046 67493 3054
rect 67030 3014 67494 3046
rect 67586 3030 67662 3167
rect 67582 2970 67592 3030
rect 67654 2970 67664 3030
rect 66504 2958 66811 2959
rect 65361 2953 65677 2958
rect 66391 2953 66811 2958
rect 65361 2942 65744 2953
rect 65361 2915 65693 2942
rect 65361 2786 65395 2915
rect 65677 2908 65693 2915
rect 65727 2908 65744 2942
rect 65677 2902 65744 2908
rect 66324 2942 66811 2953
rect 67590 2944 67660 2970
rect 66324 2908 66341 2942
rect 66375 2915 66811 2942
rect 66375 2908 66391 2915
rect 66504 2914 66811 2915
rect 66324 2902 66391 2908
rect 65502 2875 65558 2887
rect 65502 2841 65508 2875
rect 65542 2874 65558 2875
rect 66615 2874 66671 2886
rect 65542 2858 66009 2874
rect 65542 2841 65959 2858
rect 65502 2825 65959 2841
rect 65943 2824 65959 2825
rect 65993 2824 66009 2858
rect 65943 2817 66009 2824
rect 66061 2859 66631 2874
rect 66061 2825 66077 2859
rect 66111 2840 66631 2859
rect 66665 2840 66671 2874
rect 66111 2825 66671 2840
rect 66061 2815 66128 2825
rect 66615 2824 66671 2825
rect 66777 2786 66811 2914
rect 65355 2774 65401 2786
rect 65355 2598 65361 2774
rect 65395 2598 65401 2774
rect 65355 2586 65401 2598
rect 65473 2774 65519 2786
rect 65473 2598 65479 2774
rect 65513 2598 65519 2774
rect 65473 2586 65519 2598
rect 65775 2774 65821 2786
rect 65478 2292 65512 2586
rect 65775 2398 65781 2774
rect 65815 2398 65821 2774
rect 65775 2386 65821 2398
rect 65893 2774 65939 2786
rect 65893 2398 65899 2774
rect 65933 2398 65939 2774
rect 65893 2386 65939 2398
rect 66011 2774 66057 2786
rect 66011 2398 66017 2774
rect 66051 2398 66057 2774
rect 66011 2386 66057 2398
rect 66129 2774 66175 2786
rect 66129 2398 66135 2774
rect 66169 2398 66175 2774
rect 66129 2386 66175 2398
rect 66247 2774 66293 2786
rect 66247 2398 66253 2774
rect 66287 2398 66293 2774
rect 66653 2774 66699 2786
rect 66653 2598 66659 2774
rect 66693 2598 66699 2774
rect 66653 2586 66699 2598
rect 66771 2774 66817 2786
rect 66771 2598 66777 2774
rect 66811 2598 66817 2774
rect 66771 2586 66817 2598
rect 66247 2386 66293 2398
rect 66135 2292 66169 2386
rect 66659 2292 66692 2586
rect 65478 2260 66692 2292
rect 65844 2236 66250 2260
rect 65844 2113 65956 2236
rect 66130 2113 66250 2236
rect 65844 2069 66250 2113
rect 64196 971 64877 974
rect 62776 921 62932 927
rect 63720 959 63766 971
rect 63168 704 63278 705
rect 63166 703 63544 704
rect 63166 698 63545 703
rect 63160 608 63170 698
rect 63254 608 63545 698
rect 63166 604 63545 608
rect 63168 603 63278 604
rect 63468 603 63545 604
rect 63490 454 63544 603
rect 63720 583 63726 959
rect 63760 583 63766 959
rect 63720 571 63766 583
rect 63838 959 63884 971
rect 63838 583 63844 959
rect 63878 583 63884 959
rect 63838 571 63884 583
rect 63956 959 64002 971
rect 63956 583 63962 959
rect 63996 610 64002 959
rect 64073 959 64119 971
rect 64073 783 64079 959
rect 64113 783 64119 959
rect 64073 776 64119 783
rect 64191 959 64877 971
rect 64191 783 64197 959
rect 64231 946 64877 959
rect 64231 783 64237 946
rect 64481 866 64877 946
rect 64073 771 64122 776
rect 64191 771 64237 783
rect 64079 610 64122 771
rect 68012 748 68125 3456
rect 68410 3423 68498 7002
rect 68536 6959 68654 12588
rect 68536 6932 68656 6959
rect 68409 3399 68499 3423
rect 68409 3331 68420 3399
rect 68486 3331 68499 3399
rect 68409 3319 68499 3331
rect 68171 3300 68316 3313
rect 68171 3209 68186 3300
rect 68296 3209 68316 3300
rect 68171 3200 68316 3209
rect 64449 744 68125 748
rect 63996 583 64122 610
rect 63956 571 64122 583
rect 63962 567 64122 571
rect 63600 551 63673 556
rect 63594 487 63604 551
rect 63670 539 63680 551
rect 63670 533 63835 539
rect 63670 499 63785 533
rect 63819 499 63835 533
rect 63670 487 63835 499
rect 63600 483 63835 487
rect 63887 533 63953 539
rect 63887 499 63903 533
rect 63937 499 63953 533
rect 63887 454 63953 499
rect 63490 446 63953 454
rect 63490 414 63954 446
rect 64046 430 64122 567
rect 64446 630 68125 744
rect 64042 370 64052 430
rect 64114 370 64124 430
rect 57720 -105 58089 -57
rect 57720 -135 57734 -105
rect 57720 -152 57730 -135
rect 58022 -208 58088 -105
rect 59851 -144 59857 -9
rect 59924 -144 59930 -9
rect 59851 -156 59930 -144
rect 62648 -208 62714 71
rect 58020 -288 62714 -208
rect 64446 -723 64611 630
rect 65858 389 66303 395
rect 65858 189 65870 389
rect 66291 189 66303 389
rect 65858 183 66026 189
rect 66016 115 66026 183
rect 66158 183 66303 189
rect 68537 260 68656 6932
rect 68537 254 68660 260
rect 68537 188 68555 254
rect 68648 188 68660 254
rect 66158 115 66168 183
rect 68537 182 68660 188
rect 68537 180 68656 182
rect 68714 172 68804 13507
rect 68851 3318 68934 13682
rect 68976 6452 69056 13783
rect 69100 9594 69192 13901
rect 69513 12797 69655 15421
rect 70709 15431 70909 15437
rect 70709 15397 70721 15431
rect 70897 15397 70909 15431
rect 70709 15350 70909 15397
rect 70509 15344 70909 15350
rect 70365 15310 70521 15344
rect 70897 15310 70909 15344
rect 70365 14547 70422 15310
rect 70509 15304 70909 15310
rect 70509 15226 70909 15232
rect 70509 15192 70521 15226
rect 70897 15192 70909 15226
rect 70509 15186 70909 15192
rect 70509 15108 70909 15114
rect 70509 15074 70521 15108
rect 70897 15074 70909 15108
rect 70509 15068 70909 15074
rect 70509 14990 70909 14996
rect 70509 14956 70521 14990
rect 70897 14956 70909 14990
rect 70509 14950 70909 14956
rect 70509 14877 70909 14883
rect 70509 14843 70521 14877
rect 70897 14843 71035 14877
rect 70509 14837 70909 14843
rect 70509 14759 70909 14765
rect 70509 14725 70521 14759
rect 70897 14725 70909 14759
rect 70509 14719 70909 14725
rect 70509 14641 70909 14647
rect 70509 14607 70521 14641
rect 70897 14607 70909 14641
rect 70509 14601 70909 14607
rect 70265 14537 70422 14547
rect 70325 14457 70422 14537
rect 70509 14523 70909 14529
rect 70509 14489 70521 14523
rect 70897 14489 70909 14523
rect 70509 14483 70909 14489
rect 70265 14447 70422 14457
rect 70365 14169 70422 14447
rect 70509 14405 70909 14411
rect 70509 14371 70521 14405
rect 70897 14371 70909 14405
rect 70509 14365 70909 14371
rect 70509 14287 70909 14293
rect 70509 14253 70521 14287
rect 70897 14253 70909 14287
rect 70509 14247 70909 14253
rect 70509 14169 70909 14175
rect 70365 14135 70521 14169
rect 70897 14135 70909 14169
rect 70365 13578 70422 14135
rect 70509 14129 70909 14135
rect 70509 14050 70909 14056
rect 70509 14016 70521 14050
rect 70897 14016 70909 14050
rect 70509 14010 70909 14016
rect 70509 13932 70909 13938
rect 70509 13898 70521 13932
rect 70897 13898 70909 13932
rect 70509 13892 70909 13898
rect 70509 13814 70909 13820
rect 70509 13780 70521 13814
rect 70897 13780 70909 13814
rect 70509 13774 70909 13780
rect 70509 13696 70909 13702
rect 70993 13696 71035 14843
rect 71095 14699 71162 15751
rect 71195 15684 71280 15696
rect 71195 15613 71208 15684
rect 71271 15613 71280 15684
rect 71195 15604 71280 15613
rect 71672 14952 71719 15751
rect 71842 14952 72042 14957
rect 71672 14951 72042 14952
rect 71672 14918 71854 14951
rect 71095 14665 71112 14699
rect 71146 14665 71162 14699
rect 71095 14649 71162 14665
rect 71483 14717 71568 14729
rect 71483 14649 71491 14717
rect 71556 14649 71568 14717
rect 71483 14637 71568 14649
rect 71198 14599 71283 14611
rect 71198 14529 71208 14599
rect 71270 14529 71283 14599
rect 71198 14519 71283 14529
rect 71672 14480 71719 14918
rect 71842 14917 71854 14918
rect 72030 14917 72042 14951
rect 71842 14911 72042 14917
rect 71842 14833 72042 14839
rect 71842 14799 71854 14833
rect 72030 14799 72461 14833
rect 71842 14765 72042 14799
rect 71842 14759 72242 14765
rect 71842 14725 71854 14759
rect 72230 14725 72242 14759
rect 71842 14719 72242 14725
rect 71842 14641 72242 14647
rect 71842 14607 71854 14641
rect 72230 14607 72242 14641
rect 71842 14601 72242 14607
rect 71842 14523 72242 14529
rect 72315 14523 72381 14538
rect 71842 14489 71854 14523
rect 72230 14522 72381 14523
rect 72230 14489 72331 14522
rect 71842 14483 72242 14489
rect 72315 14488 72331 14489
rect 72365 14488 72381 14522
rect 71672 14464 71782 14480
rect 72315 14472 72381 14488
rect 72409 14535 72461 14799
rect 72409 14523 72539 14535
rect 71672 14430 71732 14464
rect 71766 14430 71782 14464
rect 71672 14414 71782 14430
rect 72409 14457 72483 14523
rect 72535 14457 72539 14523
rect 72409 14443 72539 14457
rect 71842 14405 72242 14411
rect 71842 14371 71854 14405
rect 72230 14371 72242 14405
rect 71842 14365 72242 14371
rect 71322 14358 71394 14364
rect 71322 14299 71328 14358
rect 71388 14299 71394 14358
rect 71325 14295 71392 14299
rect 71328 14289 71388 14295
rect 71842 14287 72242 14293
rect 71842 14253 71854 14287
rect 72230 14253 72242 14287
rect 71842 14247 72242 14253
rect 71842 14209 72042 14247
rect 72409 14209 72461 14443
rect 71842 14175 71854 14209
rect 72030 14175 72461 14209
rect 71842 14169 72042 14175
rect 71671 14091 71718 14092
rect 71842 14091 72042 14097
rect 71671 14057 71854 14091
rect 72030 14057 72042 14091
rect 70509 13662 70521 13696
rect 70897 13662 71121 13696
rect 70509 13656 70909 13662
rect 70709 13578 70909 13583
rect 70365 13577 70909 13578
rect 70365 13543 70721 13577
rect 70897 13543 70909 13577
rect 70365 13541 70909 13543
rect 70709 13537 70909 13541
rect 70709 13459 70909 13465
rect 70709 13425 70721 13459
rect 70897 13425 70909 13459
rect 70709 13419 70909 13425
rect 71055 13389 71121 13662
rect 71055 13355 71071 13389
rect 71105 13355 71121 13389
rect 70709 13341 70909 13347
rect 70709 13307 70721 13341
rect 70897 13307 70909 13341
rect 71055 13339 71121 13355
rect 70709 13301 70909 13307
rect 70709 13223 70909 13229
rect 71671 13223 71718 14057
rect 71842 14051 72042 14057
rect 70709 13189 70721 13223
rect 70897 13192 71718 13223
rect 70897 13191 71815 13192
rect 72930 13191 74426 13193
rect 70897 13189 74426 13191
rect 70709 13188 74426 13189
rect 70709 13183 70909 13188
rect 71263 13042 74426 13188
rect 71720 13041 74426 13042
rect 72930 13040 74426 13041
rect 72960 13039 73352 13040
rect 69513 12786 71399 12797
rect 69511 12784 71399 12786
rect 69511 12727 71323 12784
rect 71391 12727 71399 12784
rect 69511 12716 71399 12727
rect 70709 12642 70909 12647
rect 70709 12641 71719 12642
rect 70709 12607 70721 12641
rect 70897 12607 71719 12641
rect 70709 12601 70909 12607
rect 70709 12523 70909 12529
rect 70709 12489 70721 12523
rect 70897 12489 70909 12523
rect 70709 12483 70909 12489
rect 70709 12405 70909 12411
rect 70709 12371 70721 12405
rect 70897 12371 70909 12405
rect 70709 12365 70909 12371
rect 70709 12287 70909 12293
rect 70709 12253 70721 12287
rect 70897 12253 70909 12287
rect 70709 12206 70909 12253
rect 70509 12200 70909 12206
rect 70365 12166 70521 12200
rect 70897 12166 70909 12200
rect 70365 11403 70422 12166
rect 70509 12160 70909 12166
rect 70509 12082 70909 12088
rect 70509 12048 70521 12082
rect 70897 12048 70909 12082
rect 70509 12042 70909 12048
rect 70509 11964 70909 11970
rect 70509 11930 70521 11964
rect 70897 11930 70909 11964
rect 70509 11924 70909 11930
rect 70509 11846 70909 11852
rect 70509 11812 70521 11846
rect 70897 11812 70909 11846
rect 70509 11806 70909 11812
rect 70509 11733 70909 11739
rect 70509 11699 70521 11733
rect 70897 11699 71035 11733
rect 70509 11693 70909 11699
rect 70509 11615 70909 11621
rect 70509 11581 70521 11615
rect 70897 11581 70909 11615
rect 70509 11575 70909 11581
rect 70509 11497 70909 11503
rect 70509 11463 70521 11497
rect 70897 11463 70909 11497
rect 70509 11457 70909 11463
rect 70265 11393 70422 11403
rect 70325 11313 70422 11393
rect 70509 11379 70909 11385
rect 70509 11345 70521 11379
rect 70897 11345 70909 11379
rect 70509 11339 70909 11345
rect 70265 11303 70422 11313
rect 70365 11025 70422 11303
rect 70509 11261 70909 11267
rect 70509 11227 70521 11261
rect 70897 11227 70909 11261
rect 70509 11221 70909 11227
rect 70509 11143 70909 11149
rect 70509 11109 70521 11143
rect 70897 11109 70909 11143
rect 70509 11103 70909 11109
rect 70509 11025 70909 11031
rect 70365 10991 70521 11025
rect 70897 10991 70909 11025
rect 70365 10434 70422 10991
rect 70509 10985 70909 10991
rect 70509 10906 70909 10912
rect 70509 10872 70521 10906
rect 70897 10872 70909 10906
rect 70509 10866 70909 10872
rect 70509 10788 70909 10794
rect 70509 10754 70521 10788
rect 70897 10754 70909 10788
rect 70509 10748 70909 10754
rect 70509 10670 70909 10676
rect 70509 10636 70521 10670
rect 70897 10636 70909 10670
rect 70509 10630 70909 10636
rect 70509 10552 70909 10558
rect 70993 10552 71035 11699
rect 71095 11555 71162 12607
rect 71195 12540 71280 12552
rect 71195 12469 71208 12540
rect 71271 12469 71280 12540
rect 71195 12460 71280 12469
rect 71672 11808 71719 12607
rect 71842 11808 72042 11813
rect 71672 11807 72042 11808
rect 71672 11774 71854 11807
rect 71095 11521 71112 11555
rect 71146 11521 71162 11555
rect 71095 11505 71162 11521
rect 71483 11573 71568 11585
rect 71483 11505 71491 11573
rect 71556 11505 71568 11573
rect 71483 11493 71568 11505
rect 71198 11455 71283 11467
rect 71198 11385 71208 11455
rect 71270 11385 71283 11455
rect 71198 11375 71283 11385
rect 71672 11336 71719 11774
rect 71842 11773 71854 11774
rect 72030 11773 72042 11807
rect 71842 11767 72042 11773
rect 71842 11689 72042 11695
rect 71842 11655 71854 11689
rect 72030 11655 72461 11689
rect 71842 11621 72042 11655
rect 71842 11615 72242 11621
rect 71842 11581 71854 11615
rect 72230 11581 72242 11615
rect 71842 11575 72242 11581
rect 71842 11497 72242 11503
rect 71842 11463 71854 11497
rect 72230 11463 72242 11497
rect 71842 11457 72242 11463
rect 71842 11379 72242 11385
rect 72315 11379 72381 11394
rect 71842 11345 71854 11379
rect 72230 11378 72381 11379
rect 72230 11345 72331 11378
rect 71842 11339 72242 11345
rect 72315 11344 72331 11345
rect 72365 11344 72381 11378
rect 71672 11320 71782 11336
rect 72315 11328 72381 11344
rect 72409 11391 72461 11655
rect 72409 11379 72539 11391
rect 71672 11286 71732 11320
rect 71766 11286 71782 11320
rect 71672 11270 71782 11286
rect 72409 11313 72483 11379
rect 72535 11313 72539 11379
rect 72409 11299 72539 11313
rect 71842 11261 72242 11267
rect 71842 11227 71854 11261
rect 72230 11227 72242 11261
rect 71842 11221 72242 11227
rect 71322 11214 71394 11220
rect 71322 11155 71328 11214
rect 71388 11155 71394 11214
rect 71325 11151 71392 11155
rect 71328 11145 71388 11151
rect 71842 11143 72242 11149
rect 71842 11109 71854 11143
rect 72230 11109 72242 11143
rect 71842 11103 72242 11109
rect 71842 11065 72042 11103
rect 72409 11065 72461 11299
rect 71842 11031 71854 11065
rect 72030 11031 72461 11065
rect 71842 11025 72042 11031
rect 71671 10947 71718 10948
rect 71842 10947 72042 10953
rect 71671 10913 71854 10947
rect 72030 10913 72042 10947
rect 70509 10518 70521 10552
rect 70897 10518 71121 10552
rect 70509 10512 70909 10518
rect 70709 10434 70909 10439
rect 70365 10433 70909 10434
rect 70365 10399 70721 10433
rect 70897 10399 70909 10433
rect 70365 10397 70909 10399
rect 70709 10393 70909 10397
rect 70709 10315 70909 10321
rect 70709 10281 70721 10315
rect 70897 10281 70909 10315
rect 70709 10275 70909 10281
rect 71055 10245 71121 10518
rect 71055 10211 71071 10245
rect 71105 10211 71121 10245
rect 70709 10197 70909 10203
rect 70709 10163 70721 10197
rect 70897 10163 70909 10197
rect 71055 10195 71121 10211
rect 70709 10157 70909 10163
rect 70709 10079 70909 10085
rect 71671 10079 71718 10913
rect 71842 10907 72042 10913
rect 70709 10045 70721 10079
rect 70897 10047 71718 10079
rect 70897 10045 72874 10047
rect 73034 10045 74207 10047
rect 70709 10044 74207 10045
rect 70709 10039 70909 10044
rect 71263 9898 74207 10044
rect 71399 9897 74207 9898
rect 72959 9895 74207 9897
rect 69100 9582 71404 9594
rect 69100 9525 71327 9582
rect 71395 9525 71404 9582
rect 69100 9513 71404 9525
rect 71487 9582 71571 9597
rect 71487 9525 71495 9582
rect 71563 9525 71571 9582
rect 71487 9523 71571 9525
rect 71495 9515 71563 9523
rect 70713 9440 70913 9445
rect 70713 9439 71723 9440
rect 70713 9405 70725 9439
rect 70901 9405 71723 9439
rect 70713 9399 70913 9405
rect 70713 9321 70913 9327
rect 70713 9287 70725 9321
rect 70901 9287 70913 9321
rect 70713 9281 70913 9287
rect 70713 9203 70913 9209
rect 70713 9169 70725 9203
rect 70901 9169 70913 9203
rect 70713 9163 70913 9169
rect 70713 9085 70913 9091
rect 70713 9051 70725 9085
rect 70901 9051 70913 9085
rect 70713 9004 70913 9051
rect 70513 8998 70913 9004
rect 70369 8964 70525 8998
rect 70901 8964 70913 8998
rect 70369 8201 70426 8964
rect 70513 8958 70913 8964
rect 70513 8880 70913 8886
rect 70513 8846 70525 8880
rect 70901 8846 70913 8880
rect 70513 8840 70913 8846
rect 70513 8762 70913 8768
rect 70513 8728 70525 8762
rect 70901 8728 70913 8762
rect 70513 8722 70913 8728
rect 70513 8644 70913 8650
rect 70513 8610 70525 8644
rect 70901 8610 70913 8644
rect 70513 8604 70913 8610
rect 70513 8531 70913 8537
rect 70513 8497 70525 8531
rect 70901 8497 71039 8531
rect 70513 8491 70913 8497
rect 70513 8413 70913 8419
rect 70513 8379 70525 8413
rect 70901 8379 70913 8413
rect 70513 8373 70913 8379
rect 70513 8295 70913 8301
rect 70513 8261 70525 8295
rect 70901 8261 70913 8295
rect 70513 8255 70913 8261
rect 70269 8191 70426 8201
rect 70329 8111 70426 8191
rect 70513 8177 70913 8183
rect 70513 8143 70525 8177
rect 70901 8143 70913 8177
rect 70513 8137 70913 8143
rect 70269 8101 70426 8111
rect 70369 7823 70426 8101
rect 70513 8059 70913 8065
rect 70513 8025 70525 8059
rect 70901 8025 70913 8059
rect 70513 8019 70913 8025
rect 70513 7941 70913 7947
rect 70513 7907 70525 7941
rect 70901 7907 70913 7941
rect 70513 7901 70913 7907
rect 70513 7823 70913 7829
rect 70369 7789 70525 7823
rect 70901 7789 70913 7823
rect 70369 7232 70426 7789
rect 70513 7783 70913 7789
rect 70513 7704 70913 7710
rect 70513 7670 70525 7704
rect 70901 7670 70913 7704
rect 70513 7664 70913 7670
rect 70513 7586 70913 7592
rect 70513 7552 70525 7586
rect 70901 7552 70913 7586
rect 70513 7546 70913 7552
rect 70513 7468 70913 7474
rect 70513 7434 70525 7468
rect 70901 7434 70913 7468
rect 70513 7428 70913 7434
rect 70513 7350 70913 7356
rect 70997 7350 71039 8497
rect 71099 8353 71166 9405
rect 71199 9338 71284 9350
rect 71199 9267 71212 9338
rect 71275 9267 71284 9338
rect 71199 9258 71284 9267
rect 71676 8606 71723 9405
rect 71846 8606 72046 8611
rect 71676 8605 72046 8606
rect 71676 8572 71858 8605
rect 71099 8319 71116 8353
rect 71150 8319 71166 8353
rect 71099 8303 71166 8319
rect 71487 8371 71572 8383
rect 71487 8303 71495 8371
rect 71560 8303 71572 8371
rect 71487 8291 71572 8303
rect 71202 8253 71287 8265
rect 71202 8183 71212 8253
rect 71274 8183 71287 8253
rect 71202 8173 71287 8183
rect 71676 8134 71723 8572
rect 71846 8571 71858 8572
rect 72034 8571 72046 8605
rect 71846 8565 72046 8571
rect 71846 8487 72046 8493
rect 71846 8453 71858 8487
rect 72034 8453 72465 8487
rect 71846 8419 72046 8453
rect 71846 8413 72246 8419
rect 71846 8379 71858 8413
rect 72234 8379 72246 8413
rect 71846 8373 72246 8379
rect 71846 8295 72246 8301
rect 71846 8261 71858 8295
rect 72234 8261 72246 8295
rect 71846 8255 72246 8261
rect 71846 8177 72246 8183
rect 72319 8177 72385 8192
rect 71846 8143 71858 8177
rect 72234 8176 72385 8177
rect 72234 8143 72335 8176
rect 71846 8137 72246 8143
rect 72319 8142 72335 8143
rect 72369 8142 72385 8176
rect 71676 8118 71786 8134
rect 72319 8126 72385 8142
rect 72413 8189 72465 8453
rect 72413 8177 72543 8189
rect 71676 8084 71736 8118
rect 71770 8084 71786 8118
rect 71676 8068 71786 8084
rect 72413 8111 72487 8177
rect 72539 8111 72543 8177
rect 72413 8097 72543 8111
rect 71846 8059 72246 8065
rect 71846 8025 71858 8059
rect 72234 8025 72246 8059
rect 71846 8019 72246 8025
rect 71326 8012 71398 8018
rect 71326 7953 71332 8012
rect 71392 7953 71398 8012
rect 71329 7949 71396 7953
rect 71332 7943 71392 7949
rect 71846 7941 72246 7947
rect 71846 7907 71858 7941
rect 72234 7907 72246 7941
rect 71846 7901 72246 7907
rect 71846 7863 72046 7901
rect 72413 7863 72465 8097
rect 71846 7829 71858 7863
rect 72034 7829 72465 7863
rect 71846 7823 72046 7829
rect 71675 7745 71722 7746
rect 71846 7745 72046 7751
rect 71675 7711 71858 7745
rect 72034 7711 72046 7745
rect 70513 7316 70525 7350
rect 70901 7316 71125 7350
rect 70513 7310 70913 7316
rect 70713 7232 70913 7237
rect 70369 7231 70913 7232
rect 70369 7197 70725 7231
rect 70901 7197 70913 7231
rect 70369 7195 70913 7197
rect 70713 7191 70913 7195
rect 70713 7113 70913 7119
rect 70713 7079 70725 7113
rect 70901 7079 70913 7113
rect 70713 7073 70913 7079
rect 71059 7043 71125 7316
rect 71059 7009 71075 7043
rect 71109 7009 71125 7043
rect 70713 6995 70913 7001
rect 70713 6961 70725 6995
rect 70901 6961 70913 6995
rect 71059 6993 71125 7009
rect 70713 6955 70913 6961
rect 70713 6877 70913 6883
rect 71675 6877 71722 7711
rect 71846 7705 72046 7711
rect 70713 6843 70725 6877
rect 70901 6847 71722 6877
rect 70901 6846 71791 6847
rect 72962 6846 73911 6849
rect 70901 6843 73911 6846
rect 70713 6842 73911 6843
rect 70713 6837 70913 6842
rect 71267 6697 73911 6842
rect 71267 6696 71413 6697
rect 71722 6696 73911 6697
rect 72962 6695 73911 6696
rect 73016 6693 73911 6695
rect 68976 6451 71359 6452
rect 68976 6438 71403 6451
rect 68976 6381 71327 6438
rect 71395 6381 71403 6438
rect 68976 6379 71403 6381
rect 68976 6371 71395 6379
rect 70713 6296 70913 6301
rect 70713 6295 71723 6296
rect 70713 6261 70725 6295
rect 70901 6261 71723 6295
rect 70713 6255 70913 6261
rect 70713 6177 70913 6183
rect 70713 6143 70725 6177
rect 70901 6143 70913 6177
rect 70713 6137 70913 6143
rect 70713 6059 70913 6065
rect 70713 6025 70725 6059
rect 70901 6025 70913 6059
rect 70713 6019 70913 6025
rect 70713 5941 70913 5947
rect 70713 5907 70725 5941
rect 70901 5907 70913 5941
rect 70713 5860 70913 5907
rect 70513 5854 70913 5860
rect 70369 5820 70525 5854
rect 70901 5820 70913 5854
rect 70369 5057 70426 5820
rect 70513 5814 70913 5820
rect 70513 5736 70913 5742
rect 70513 5702 70525 5736
rect 70901 5702 70913 5736
rect 70513 5696 70913 5702
rect 70513 5618 70913 5624
rect 70513 5584 70525 5618
rect 70901 5584 70913 5618
rect 70513 5578 70913 5584
rect 70513 5500 70913 5506
rect 70513 5466 70525 5500
rect 70901 5466 70913 5500
rect 70513 5460 70913 5466
rect 70513 5387 70913 5393
rect 70513 5353 70525 5387
rect 70901 5353 71039 5387
rect 70513 5347 70913 5353
rect 70513 5269 70913 5275
rect 70513 5235 70525 5269
rect 70901 5235 70913 5269
rect 70513 5229 70913 5235
rect 70513 5151 70913 5157
rect 70513 5117 70525 5151
rect 70901 5117 70913 5151
rect 70513 5111 70913 5117
rect 70269 5047 70426 5057
rect 70329 4967 70426 5047
rect 70513 5033 70913 5039
rect 70513 4999 70525 5033
rect 70901 4999 70913 5033
rect 70513 4993 70913 4999
rect 70269 4957 70426 4967
rect 70369 4679 70426 4957
rect 70513 4915 70913 4921
rect 70513 4881 70525 4915
rect 70901 4881 70913 4915
rect 70513 4875 70913 4881
rect 70513 4797 70913 4803
rect 70513 4763 70525 4797
rect 70901 4763 70913 4797
rect 70513 4757 70913 4763
rect 70513 4679 70913 4685
rect 70369 4645 70525 4679
rect 70901 4645 70913 4679
rect 70369 4088 70426 4645
rect 70513 4639 70913 4645
rect 70513 4560 70913 4566
rect 70513 4526 70525 4560
rect 70901 4526 70913 4560
rect 70513 4520 70913 4526
rect 70513 4442 70913 4448
rect 70513 4408 70525 4442
rect 70901 4408 70913 4442
rect 70513 4402 70913 4408
rect 70513 4324 70913 4330
rect 70513 4290 70525 4324
rect 70901 4290 70913 4324
rect 70513 4284 70913 4290
rect 70513 4206 70913 4212
rect 70997 4206 71039 5353
rect 71099 5209 71166 6261
rect 71199 6194 71284 6206
rect 71199 6123 71212 6194
rect 71275 6123 71284 6194
rect 71199 6114 71284 6123
rect 71676 5462 71723 6261
rect 71846 5462 72046 5467
rect 71676 5461 72046 5462
rect 71676 5428 71858 5461
rect 71099 5175 71116 5209
rect 71150 5175 71166 5209
rect 71099 5159 71166 5175
rect 71487 5227 71572 5239
rect 71487 5159 71495 5227
rect 71560 5159 71572 5227
rect 71487 5147 71572 5159
rect 71202 5109 71287 5121
rect 71202 5039 71212 5109
rect 71274 5039 71287 5109
rect 71202 5029 71287 5039
rect 71676 4990 71723 5428
rect 71846 5427 71858 5428
rect 72034 5427 72046 5461
rect 71846 5421 72046 5427
rect 71846 5343 72046 5349
rect 71846 5309 71858 5343
rect 72034 5309 72465 5343
rect 71846 5275 72046 5309
rect 71846 5269 72246 5275
rect 71846 5235 71858 5269
rect 72234 5235 72246 5269
rect 71846 5229 72246 5235
rect 71846 5151 72246 5157
rect 71846 5117 71858 5151
rect 72234 5117 72246 5151
rect 71846 5111 72246 5117
rect 71846 5033 72246 5039
rect 72319 5033 72385 5048
rect 71846 4999 71858 5033
rect 72234 5032 72385 5033
rect 72234 4999 72335 5032
rect 71846 4993 72246 4999
rect 72319 4998 72335 4999
rect 72369 4998 72385 5032
rect 71676 4974 71786 4990
rect 72319 4982 72385 4998
rect 72413 5045 72465 5309
rect 72413 5033 72543 5045
rect 71676 4940 71736 4974
rect 71770 4940 71786 4974
rect 71676 4924 71786 4940
rect 72413 4967 72487 5033
rect 72539 4967 72543 5033
rect 72413 4953 72543 4967
rect 71846 4915 72246 4921
rect 71846 4881 71858 4915
rect 72234 4881 72246 4915
rect 71846 4875 72246 4881
rect 71326 4868 71398 4874
rect 71326 4809 71332 4868
rect 71392 4809 71398 4868
rect 71329 4805 71396 4809
rect 71332 4799 71392 4805
rect 71846 4797 72246 4803
rect 71846 4763 71858 4797
rect 72234 4763 72246 4797
rect 71846 4757 72246 4763
rect 71846 4719 72046 4757
rect 72413 4719 72465 4953
rect 71846 4685 71858 4719
rect 72034 4685 72465 4719
rect 71846 4679 72046 4685
rect 71675 4601 71722 4602
rect 71846 4601 72046 4607
rect 71675 4567 71858 4601
rect 72034 4567 72046 4601
rect 70513 4172 70525 4206
rect 70901 4172 71125 4206
rect 70513 4166 70913 4172
rect 70713 4088 70913 4093
rect 70369 4087 70913 4088
rect 70369 4053 70725 4087
rect 70901 4053 70913 4087
rect 70369 4051 70913 4053
rect 70713 4047 70913 4051
rect 70713 3969 70913 3975
rect 70713 3935 70725 3969
rect 70901 3935 70913 3969
rect 70713 3929 70913 3935
rect 71059 3899 71125 4172
rect 71059 3865 71075 3899
rect 71109 3865 71125 3899
rect 70713 3851 70913 3857
rect 70713 3817 70725 3851
rect 70901 3817 70913 3851
rect 71059 3849 71125 3865
rect 70713 3811 70913 3817
rect 70713 3733 70913 3739
rect 71675 3733 71722 4567
rect 71846 4561 72046 4567
rect 70713 3699 70725 3733
rect 70901 3702 71722 3733
rect 70901 3701 71815 3702
rect 72962 3701 73354 3702
rect 70901 3699 73651 3701
rect 70713 3698 73651 3699
rect 70713 3693 70913 3698
rect 71267 3552 73651 3698
rect 71722 3551 73651 3552
rect 73323 3549 73651 3551
rect 71315 3318 71399 3319
rect 68851 3306 71401 3318
rect 68851 3249 71323 3306
rect 71391 3249 71401 3306
rect 68851 3239 71401 3249
rect 71483 3306 71567 3321
rect 71483 3249 71491 3306
rect 71559 3249 71567 3306
rect 71483 3247 71567 3249
rect 71491 3239 71559 3247
rect 70709 3164 70909 3169
rect 70709 3163 71719 3164
rect 70709 3129 70721 3163
rect 70897 3129 71719 3163
rect 70709 3123 70909 3129
rect 70709 3045 70909 3051
rect 70709 3011 70721 3045
rect 70897 3011 70909 3045
rect 70709 3005 70909 3011
rect 70709 2927 70909 2933
rect 70709 2893 70721 2927
rect 70897 2893 70909 2927
rect 70709 2887 70909 2893
rect 70709 2809 70909 2815
rect 70709 2775 70721 2809
rect 70897 2775 70909 2809
rect 70709 2728 70909 2775
rect 70509 2722 70909 2728
rect 70365 2688 70521 2722
rect 70897 2688 70909 2722
rect 70365 1925 70422 2688
rect 70509 2682 70909 2688
rect 70509 2604 70909 2610
rect 70509 2570 70521 2604
rect 70897 2570 70909 2604
rect 70509 2564 70909 2570
rect 70509 2486 70909 2492
rect 70509 2452 70521 2486
rect 70897 2452 70909 2486
rect 70509 2446 70909 2452
rect 70509 2368 70909 2374
rect 70509 2334 70521 2368
rect 70897 2334 70909 2368
rect 70509 2328 70909 2334
rect 70509 2255 70909 2261
rect 70509 2221 70521 2255
rect 70897 2221 71035 2255
rect 70509 2215 70909 2221
rect 70509 2137 70909 2143
rect 70509 2103 70521 2137
rect 70897 2103 70909 2137
rect 70509 2097 70909 2103
rect 70509 2019 70909 2025
rect 70509 1985 70521 2019
rect 70897 1985 70909 2019
rect 70509 1979 70909 1985
rect 70265 1915 70422 1925
rect 70325 1835 70422 1915
rect 70509 1901 70909 1907
rect 70509 1867 70521 1901
rect 70897 1867 70909 1901
rect 70509 1861 70909 1867
rect 70265 1825 70422 1835
rect 70365 1547 70422 1825
rect 70509 1783 70909 1789
rect 70509 1749 70521 1783
rect 70897 1749 70909 1783
rect 70509 1743 70909 1749
rect 70509 1665 70909 1671
rect 70509 1631 70521 1665
rect 70897 1631 70909 1665
rect 70509 1625 70909 1631
rect 70509 1547 70909 1553
rect 70365 1513 70521 1547
rect 70897 1513 70909 1547
rect 70365 956 70422 1513
rect 70509 1507 70909 1513
rect 70509 1428 70909 1434
rect 70509 1394 70521 1428
rect 70897 1394 70909 1428
rect 70509 1388 70909 1394
rect 70509 1310 70909 1316
rect 70509 1276 70521 1310
rect 70897 1276 70909 1310
rect 70509 1270 70909 1276
rect 70509 1192 70909 1198
rect 70509 1158 70521 1192
rect 70897 1158 70909 1192
rect 70509 1152 70909 1158
rect 70509 1074 70909 1080
rect 70993 1074 71035 2221
rect 71095 2077 71162 3129
rect 71195 3062 71280 3074
rect 71195 2991 71208 3062
rect 71271 2991 71280 3062
rect 71195 2982 71280 2991
rect 71672 2330 71719 3129
rect 71842 2330 72042 2335
rect 71672 2329 72042 2330
rect 71672 2296 71854 2329
rect 71095 2043 71112 2077
rect 71146 2043 71162 2077
rect 71095 2027 71162 2043
rect 71483 2095 71568 2107
rect 71483 2027 71491 2095
rect 71556 2027 71568 2095
rect 71483 2015 71568 2027
rect 71198 1977 71283 1989
rect 71198 1907 71208 1977
rect 71270 1907 71283 1977
rect 71198 1897 71283 1907
rect 71672 1858 71719 2296
rect 71842 2295 71854 2296
rect 72030 2295 72042 2329
rect 71842 2289 72042 2295
rect 71842 2211 72042 2217
rect 71842 2177 71854 2211
rect 72030 2177 72461 2211
rect 71842 2143 72042 2177
rect 71842 2137 72242 2143
rect 71842 2103 71854 2137
rect 72230 2103 72242 2137
rect 71842 2097 72242 2103
rect 71842 2019 72242 2025
rect 71842 1985 71854 2019
rect 72230 1985 72242 2019
rect 71842 1979 72242 1985
rect 71842 1901 72242 1907
rect 72315 1901 72381 1916
rect 71842 1867 71854 1901
rect 72230 1900 72381 1901
rect 72230 1867 72331 1900
rect 71842 1861 72242 1867
rect 72315 1866 72331 1867
rect 72365 1866 72381 1900
rect 71672 1842 71782 1858
rect 72315 1850 72381 1866
rect 72409 1913 72461 2177
rect 72409 1901 72539 1913
rect 71672 1808 71732 1842
rect 71766 1808 71782 1842
rect 71672 1792 71782 1808
rect 72409 1835 72483 1901
rect 72535 1835 72539 1901
rect 72409 1821 72539 1835
rect 71842 1783 72242 1789
rect 71842 1749 71854 1783
rect 72230 1749 72242 1783
rect 71842 1743 72242 1749
rect 71322 1736 71394 1742
rect 71322 1677 71328 1736
rect 71388 1677 71394 1736
rect 71325 1673 71392 1677
rect 71328 1667 71388 1673
rect 71842 1665 72242 1671
rect 71842 1631 71854 1665
rect 72230 1631 72242 1665
rect 71842 1625 72242 1631
rect 71842 1587 72042 1625
rect 72409 1587 72461 1821
rect 71842 1553 71854 1587
rect 72030 1553 72461 1587
rect 71842 1547 72042 1553
rect 71671 1469 71718 1470
rect 71842 1469 72042 1475
rect 71671 1435 71854 1469
rect 72030 1435 72042 1469
rect 70509 1040 70521 1074
rect 70897 1040 71121 1074
rect 70509 1034 70909 1040
rect 70709 956 70909 961
rect 70365 955 70909 956
rect 70365 921 70721 955
rect 70897 921 70909 955
rect 70365 919 70909 921
rect 70709 915 70909 919
rect 70709 837 70909 843
rect 70709 803 70721 837
rect 70897 803 70909 837
rect 70709 797 70909 803
rect 71055 767 71121 1040
rect 71055 733 71071 767
rect 71105 733 71121 767
rect 70709 719 70909 725
rect 70709 685 70721 719
rect 70897 685 70909 719
rect 71055 717 71121 733
rect 70709 679 70909 685
rect 70709 601 70909 607
rect 71671 601 71718 1435
rect 71842 1429 72042 1435
rect 70709 567 70721 601
rect 70897 571 71718 601
rect 72958 571 73391 572
rect 70897 567 73391 571
rect 70709 566 73391 567
rect 70709 561 70909 566
rect 71263 421 73391 566
rect 72958 420 73391 421
rect 73206 418 73391 420
rect 71315 172 71399 175
rect 68714 162 71401 172
rect 66026 75 66158 115
rect 68714 105 71323 162
rect 71391 105 71401 162
rect 68714 95 71401 105
rect 71483 162 71567 172
rect 71483 105 71491 162
rect 71559 105 71567 162
rect 71483 103 71567 105
rect 71491 95 71559 103
rect 68714 94 68804 95
rect 66025 9 66158 75
rect 70709 20 70909 25
rect 70709 19 71719 20
rect 65354 -34 66827 9
rect 70709 -15 70721 19
rect 70897 -15 71719 19
rect 70709 -21 70909 -15
rect 65354 -337 65388 -34
rect 65720 -137 65754 -34
rect 65956 -137 65990 -34
rect 66192 -137 66226 -34
rect 66428 -137 66462 -34
rect 65714 -149 65760 -137
rect 65230 -349 65276 -337
rect 65230 -525 65236 -349
rect 65270 -525 65276 -349
rect 65230 -537 65276 -525
rect 65348 -349 65394 -337
rect 65348 -525 65354 -349
rect 65388 -525 65394 -349
rect 65348 -537 65394 -525
rect 65466 -349 65512 -337
rect 65466 -525 65472 -349
rect 65506 -525 65512 -349
rect 65466 -537 65512 -525
rect 65584 -349 65630 -337
rect 65714 -349 65720 -149
rect 65584 -525 65590 -349
rect 65624 -525 65720 -349
rect 65754 -525 65760 -149
rect 65584 -537 65630 -525
rect 65714 -537 65760 -525
rect 65832 -149 65878 -137
rect 65832 -525 65838 -149
rect 65872 -525 65878 -149
rect 65832 -537 65878 -525
rect 65950 -149 65996 -137
rect 65950 -525 65956 -149
rect 65990 -525 65996 -149
rect 65950 -537 65996 -525
rect 66068 -149 66114 -137
rect 66068 -525 66074 -149
rect 66108 -525 66114 -149
rect 66068 -537 66114 -525
rect 66186 -149 66232 -137
rect 66186 -525 66192 -149
rect 66226 -525 66232 -149
rect 66186 -537 66232 -525
rect 66304 -149 66350 -137
rect 66304 -525 66310 -149
rect 66344 -525 66350 -149
rect 66304 -537 66350 -525
rect 66422 -149 66468 -137
rect 66422 -525 66428 -149
rect 66462 -349 66468 -149
rect 66793 -337 66827 -34
rect 67334 -114 67470 -94
rect 67334 -176 67370 -114
rect 67430 -176 67470 -114
rect 70709 -99 70909 -93
rect 70709 -133 70721 -99
rect 70897 -133 70909 -99
rect 70709 -139 70909 -133
rect 67334 -204 67470 -176
rect 67030 -234 68007 -204
rect 66551 -349 66597 -337
rect 66462 -525 66557 -349
rect 66591 -525 66597 -349
rect 66422 -537 66468 -525
rect 66551 -537 66597 -525
rect 66669 -349 66715 -337
rect 66669 -525 66675 -349
rect 66709 -525 66715 -349
rect 66669 -537 66715 -525
rect 66787 -349 66833 -337
rect 66787 -525 66793 -349
rect 66827 -525 66833 -349
rect 66787 -537 66833 -525
rect 66905 -349 66951 -337
rect 67030 -340 67062 -234
rect 67266 -340 67298 -234
rect 67502 -340 67534 -234
rect 67738 -340 67770 -234
rect 67973 -340 68007 -234
rect 70709 -217 70909 -211
rect 70709 -251 70721 -217
rect 70897 -251 70909 -217
rect 70709 -257 70909 -251
rect 70709 -335 70909 -329
rect 66905 -525 66911 -349
rect 66945 -525 66951 -349
rect 66905 -537 66951 -525
rect 67023 -352 67069 -340
rect 67023 -528 67029 -352
rect 67063 -528 67069 -352
rect 65236 -571 65270 -537
rect 65838 -571 65872 -537
rect 66074 -571 66108 -537
rect 65236 -606 65395 -571
rect 65838 -606 66108 -571
rect 66675 -571 66709 -537
rect 66911 -571 66945 -537
rect 67023 -540 67069 -528
rect 67141 -352 67187 -340
rect 67141 -528 67147 -352
rect 67181 -528 67187 -352
rect 67141 -540 67187 -528
rect 67259 -352 67305 -340
rect 67259 -528 67265 -352
rect 67299 -528 67305 -352
rect 67259 -540 67305 -528
rect 67377 -352 67423 -340
rect 67377 -528 67383 -352
rect 67417 -528 67423 -352
rect 67377 -540 67423 -528
rect 67495 -352 67541 -340
rect 67495 -528 67501 -352
rect 67535 -528 67541 -352
rect 67495 -540 67541 -528
rect 67613 -352 67659 -340
rect 67613 -528 67619 -352
rect 67653 -528 67659 -352
rect 67613 -540 67659 -528
rect 67731 -352 67777 -340
rect 67731 -528 67737 -352
rect 67771 -528 67777 -352
rect 67731 -540 67777 -528
rect 67849 -352 67895 -340
rect 67849 -528 67855 -352
rect 67889 -528 67895 -352
rect 67849 -540 67895 -528
rect 67967 -352 68013 -340
rect 67967 -528 67973 -352
rect 68007 -528 68013 -352
rect 67967 -540 68013 -528
rect 68085 -352 68131 -340
rect 68085 -528 68091 -352
rect 68125 -528 68131 -352
rect 70709 -369 70721 -335
rect 70897 -369 70909 -335
rect 70709 -416 70909 -369
rect 70509 -422 70909 -416
rect 68085 -540 68131 -528
rect 70365 -456 70521 -422
rect 70897 -456 70909 -422
rect 66675 -606 66945 -571
rect 56696 -874 64611 -723
rect 65204 -687 65301 -681
rect 65204 -758 65216 -687
rect 65289 -691 65301 -687
rect 65290 -754 65301 -691
rect 65289 -758 65301 -754
rect 65204 -764 65301 -758
rect 56775 -876 64611 -874
rect 64782 -817 65246 -816
rect 64782 -880 65223 -817
rect 65290 -880 65300 -817
rect 64782 -883 65246 -880
rect 62268 -952 63556 -951
rect 55800 -1300 56593 -1220
rect 55550 -1313 56593 -1300
rect 55510 -1325 56593 -1313
rect 55045 -1438 55079 -1325
rect 55515 -1329 56593 -1325
rect 59194 -953 63680 -952
rect 59194 -962 63681 -953
rect 59194 -1052 63584 -962
rect 63668 -1052 63681 -962
rect 59194 -1058 63681 -1052
rect 59194 -1059 63680 -1058
rect 55441 -1363 55507 -1356
rect 55441 -1397 55457 -1363
rect 55491 -1397 55507 -1363
rect 55441 -1438 55507 -1397
rect 54925 -1439 55507 -1438
rect 54925 -1468 55625 -1439
rect 54925 -1562 54961 -1468
rect 55161 -1562 55197 -1468
rect 55397 -1469 55625 -1468
rect 55397 -1562 55433 -1469
rect 55559 -1480 55625 -1469
rect 55559 -1514 55575 -1480
rect 55609 -1514 55625 -1480
rect 55559 -1521 55625 -1514
rect 55869 -1562 55904 -1329
rect 54802 -1574 54848 -1562
rect 54802 -1750 54808 -1574
rect 54842 -1750 54848 -1574
rect 54802 -1762 54848 -1750
rect 54920 -1574 54966 -1562
rect 54920 -1750 54926 -1574
rect 54960 -1750 54966 -1574
rect 54920 -1762 54966 -1750
rect 55038 -1574 55084 -1562
rect 55038 -1750 55044 -1574
rect 55078 -1750 55084 -1574
rect 55038 -1762 55084 -1750
rect 55156 -1574 55202 -1562
rect 55156 -1750 55162 -1574
rect 55196 -1750 55202 -1574
rect 55156 -1762 55202 -1750
rect 55274 -1574 55320 -1562
rect 55274 -1750 55280 -1574
rect 55314 -1750 55320 -1574
rect 55274 -1762 55320 -1750
rect 55392 -1574 55438 -1562
rect 55392 -1750 55398 -1574
rect 55432 -1750 55438 -1574
rect 55392 -1762 55438 -1750
rect 55510 -1574 55556 -1562
rect 55510 -1750 55516 -1574
rect 55550 -1750 55556 -1574
rect 55510 -1762 55556 -1750
rect 55628 -1574 55674 -1562
rect 55628 -1750 55634 -1574
rect 55668 -1750 55674 -1574
rect 55628 -1762 55674 -1750
rect 55746 -1574 55792 -1562
rect 55746 -1750 55752 -1574
rect 55786 -1750 55792 -1574
rect 55746 -1762 55792 -1750
rect 55864 -1574 55910 -1562
rect 55864 -1750 55870 -1574
rect 55904 -1750 55910 -1574
rect 55864 -1762 55910 -1750
rect 54809 -1868 54841 -1762
rect 55045 -1868 55077 -1762
rect 55281 -1868 55313 -1762
rect 55517 -1868 55549 -1762
rect 55752 -1868 55786 -1762
rect 54809 -1898 55786 -1868
rect 55113 -1926 55249 -1898
rect 55113 -1988 55149 -1926
rect 55209 -1988 55249 -1926
rect 55113 -2008 55249 -1988
rect 33761 -2190 35303 -2189
rect 47682 -2190 48106 -2189
rect 33761 -2266 33773 -2190
rect 33867 -2195 48106 -2190
rect 33867 -2199 41414 -2195
rect 33867 -2266 36374 -2199
rect 33761 -2268 36374 -2266
rect 36470 -2268 41414 -2199
rect 33761 -2269 41414 -2268
rect 41514 -2269 48106 -2195
rect 33761 -2272 48106 -2269
rect 33763 -2274 48106 -2272
rect 48620 -2161 54584 -2086
rect 34629 -2275 47728 -2274
rect 34249 -2305 47795 -2303
rect 48620 -2305 48701 -2161
rect 59194 -2200 59350 -1059
rect 63801 -1211 63937 -1191
rect 63801 -1273 63837 -1211
rect 63897 -1273 63937 -1211
rect 63801 -1301 63937 -1273
rect 63497 -1331 64474 -1301
rect 63497 -1437 63529 -1331
rect 63733 -1437 63765 -1331
rect 63969 -1437 64001 -1331
rect 64205 -1437 64237 -1331
rect 64440 -1437 64474 -1331
rect 63490 -1449 63536 -1437
rect 63490 -1625 63496 -1449
rect 63530 -1625 63536 -1449
rect 63490 -1637 63536 -1625
rect 63608 -1449 63654 -1437
rect 63608 -1625 63614 -1449
rect 63648 -1625 63654 -1449
rect 63608 -1637 63654 -1625
rect 63726 -1449 63772 -1437
rect 63726 -1625 63732 -1449
rect 63766 -1625 63772 -1449
rect 63726 -1637 63772 -1625
rect 63844 -1449 63890 -1437
rect 63844 -1625 63850 -1449
rect 63884 -1625 63890 -1449
rect 63844 -1637 63890 -1625
rect 63962 -1449 64008 -1437
rect 63962 -1625 63968 -1449
rect 64002 -1625 64008 -1449
rect 63962 -1637 64008 -1625
rect 64080 -1449 64126 -1437
rect 64080 -1625 64086 -1449
rect 64120 -1625 64126 -1449
rect 64080 -1637 64126 -1625
rect 64198 -1449 64244 -1437
rect 64198 -1625 64204 -1449
rect 64238 -1625 64244 -1449
rect 64198 -1637 64244 -1625
rect 64316 -1449 64362 -1437
rect 64316 -1625 64322 -1449
rect 64356 -1625 64362 -1449
rect 64316 -1637 64362 -1625
rect 64434 -1449 64480 -1437
rect 64434 -1625 64440 -1449
rect 64474 -1625 64480 -1449
rect 64434 -1637 64480 -1625
rect 64552 -1449 64598 -1437
rect 64552 -1625 64558 -1449
rect 64592 -1625 64598 -1449
rect 64552 -1637 64598 -1625
rect 62511 -1696 63095 -1695
rect 34249 -2311 48701 -2305
rect 34249 -2397 34260 -2311
rect 34359 -2397 48701 -2311
rect 34249 -2405 48701 -2397
rect 34629 -2406 48701 -2405
rect 48729 -2281 59350 -2200
rect 59388 -1705 63096 -1696
rect 59388 -1795 62999 -1705
rect 63083 -1795 63096 -1705
rect 63613 -1731 63649 -1637
rect 63849 -1731 63885 -1637
rect 64085 -1730 64121 -1637
rect 64247 -1685 64313 -1678
rect 64247 -1719 64263 -1685
rect 64297 -1719 64313 -1685
rect 64247 -1730 64313 -1719
rect 64085 -1731 64313 -1730
rect 63613 -1760 64313 -1731
rect 63613 -1761 64195 -1760
rect 59388 -1801 63096 -1795
rect 59388 -1802 63095 -1801
rect 59388 -1803 61573 -1802
rect 48729 -2282 54419 -2281
rect 34352 -2445 35303 -2444
rect 34352 -2446 47744 -2445
rect 48729 -2446 48813 -2282
rect 59388 -2323 59544 -1803
rect 63733 -1874 63767 -1761
rect 64129 -1802 64195 -1761
rect 64129 -1836 64145 -1802
rect 64179 -1836 64195 -1802
rect 64129 -1843 64195 -1836
rect 64557 -1870 64592 -1637
rect 64782 -1870 64877 -883
rect 65361 -1390 65395 -606
rect 66074 -668 66108 -606
rect 65663 -706 66405 -668
rect 65473 -877 65483 -809
rect 65538 -877 65548 -809
rect 65663 -830 65697 -706
rect 65899 -830 65933 -706
rect 66135 -830 66169 -706
rect 66371 -830 66405 -706
rect 65657 -842 65703 -830
rect 65657 -1218 65663 -842
rect 65697 -1218 65703 -842
rect 65657 -1230 65703 -1218
rect 65775 -842 65821 -830
rect 65775 -1218 65781 -842
rect 65815 -1218 65821 -842
rect 65775 -1230 65821 -1218
rect 65893 -842 65939 -830
rect 65893 -1218 65899 -842
rect 65933 -1218 65939 -842
rect 65893 -1230 65939 -1218
rect 66011 -842 66057 -830
rect 66011 -1218 66017 -842
rect 66051 -1218 66057 -842
rect 66011 -1230 66057 -1218
rect 66129 -842 66175 -830
rect 66129 -1218 66135 -842
rect 66169 -1218 66175 -842
rect 66129 -1230 66175 -1218
rect 66247 -842 66293 -830
rect 66247 -1218 66253 -842
rect 66287 -1218 66293 -842
rect 66247 -1230 66293 -1218
rect 66365 -842 66411 -830
rect 66365 -1218 66371 -842
rect 66405 -1218 66411 -842
rect 66531 -1047 66605 -1035
rect 66527 -1138 66537 -1047
rect 66599 -1138 66609 -1047
rect 66531 -1150 66605 -1138
rect 66365 -1230 66411 -1218
rect 66777 -1389 66811 -606
rect 67146 -634 67182 -540
rect 67382 -634 67418 -540
rect 67618 -633 67654 -540
rect 67780 -588 67846 -581
rect 67780 -622 67796 -588
rect 67830 -622 67846 -588
rect 67780 -633 67846 -622
rect 67618 -634 67846 -633
rect 67146 -663 67846 -634
rect 67146 -664 67728 -663
rect 66872 -696 66948 -691
rect 66869 -752 66879 -696
rect 66932 -697 66948 -696
rect 66932 -752 67198 -697
rect 66872 -757 67198 -752
rect 66993 -799 67084 -794
rect 66993 -888 67003 -799
rect 67076 -888 67084 -799
rect 66993 -900 67084 -888
rect 67030 -1294 67084 -900
rect 67144 -1209 67198 -757
rect 67266 -777 67300 -664
rect 67662 -705 67728 -664
rect 67662 -739 67678 -705
rect 67712 -739 67728 -705
rect 67662 -746 67728 -739
rect 68090 -773 68125 -540
rect 67736 -777 68125 -773
rect 67260 -789 67306 -777
rect 67260 -1165 67266 -789
rect 67300 -1165 67306 -789
rect 67260 -1177 67306 -1165
rect 67378 -789 67424 -777
rect 67378 -1165 67384 -789
rect 67418 -1165 67424 -789
rect 67378 -1177 67424 -1165
rect 67496 -789 67542 -777
rect 67496 -1165 67502 -789
rect 67536 -1138 67542 -789
rect 67613 -789 67659 -777
rect 67613 -965 67619 -789
rect 67653 -965 67659 -789
rect 67613 -972 67659 -965
rect 67731 -788 68125 -777
rect 67731 -789 67968 -788
rect 67731 -965 67737 -789
rect 67771 -802 67968 -789
rect 67771 -965 67777 -802
rect 67950 -876 67968 -802
rect 68110 -876 68125 -788
rect 67950 -891 68125 -876
rect 67613 -977 67662 -972
rect 67731 -977 67777 -965
rect 67619 -1138 67662 -977
rect 67536 -1165 67662 -1138
rect 67496 -1177 67662 -1165
rect 67502 -1181 67662 -1177
rect 67144 -1215 67375 -1209
rect 67144 -1249 67325 -1215
rect 67359 -1249 67375 -1215
rect 67144 -1265 67375 -1249
rect 67427 -1215 67493 -1209
rect 67427 -1249 67443 -1215
rect 67477 -1249 67493 -1215
rect 67427 -1294 67493 -1249
rect 67030 -1302 67493 -1294
rect 67030 -1334 67494 -1302
rect 67586 -1318 67662 -1181
rect 70365 -1219 70422 -456
rect 70509 -462 70909 -456
rect 70509 -540 70909 -534
rect 70509 -574 70521 -540
rect 70897 -574 70909 -540
rect 70509 -580 70909 -574
rect 70509 -658 70909 -652
rect 70509 -692 70521 -658
rect 70897 -692 70909 -658
rect 70509 -698 70909 -692
rect 70509 -776 70909 -770
rect 70509 -810 70521 -776
rect 70897 -810 70909 -776
rect 70509 -816 70909 -810
rect 70509 -889 70909 -883
rect 70509 -923 70521 -889
rect 70897 -923 71035 -889
rect 70509 -929 70909 -923
rect 70509 -1007 70909 -1001
rect 70509 -1041 70521 -1007
rect 70897 -1041 70909 -1007
rect 70509 -1047 70909 -1041
rect 70509 -1125 70909 -1119
rect 70509 -1159 70521 -1125
rect 70897 -1159 70909 -1125
rect 70509 -1165 70909 -1159
rect 70265 -1229 70422 -1219
rect 70325 -1309 70422 -1229
rect 70509 -1243 70909 -1237
rect 70509 -1277 70521 -1243
rect 70897 -1277 70909 -1243
rect 70509 -1283 70909 -1277
rect 67582 -1378 67592 -1318
rect 67654 -1378 67664 -1318
rect 70265 -1319 70422 -1309
rect 66504 -1390 66811 -1389
rect 65361 -1395 65677 -1390
rect 66391 -1395 66811 -1390
rect 65361 -1406 65744 -1395
rect 65361 -1433 65693 -1406
rect 65361 -1562 65395 -1433
rect 65677 -1440 65693 -1433
rect 65727 -1440 65744 -1406
rect 65677 -1446 65744 -1440
rect 66324 -1406 66811 -1395
rect 67590 -1404 67660 -1378
rect 66324 -1440 66341 -1406
rect 66375 -1433 66811 -1406
rect 66375 -1440 66391 -1433
rect 66504 -1434 66811 -1433
rect 66324 -1446 66391 -1440
rect 65502 -1473 65558 -1461
rect 65502 -1507 65508 -1473
rect 65542 -1474 65558 -1473
rect 66615 -1474 66671 -1462
rect 65542 -1490 66009 -1474
rect 65542 -1507 65959 -1490
rect 65502 -1523 65959 -1507
rect 65943 -1524 65959 -1523
rect 65993 -1524 66009 -1490
rect 65943 -1531 66009 -1524
rect 66061 -1489 66631 -1474
rect 66061 -1523 66077 -1489
rect 66111 -1508 66631 -1489
rect 66665 -1508 66671 -1474
rect 66111 -1523 66671 -1508
rect 66061 -1533 66128 -1523
rect 66615 -1524 66671 -1523
rect 66777 -1562 66811 -1434
rect 65355 -1574 65401 -1562
rect 65355 -1750 65361 -1574
rect 65395 -1750 65401 -1574
rect 65355 -1762 65401 -1750
rect 65473 -1574 65519 -1562
rect 65473 -1750 65479 -1574
rect 65513 -1750 65519 -1574
rect 65473 -1762 65519 -1750
rect 65775 -1574 65821 -1562
rect 64203 -1874 64877 -1870
rect 63727 -1886 63773 -1874
rect 34352 -2448 48813 -2446
rect 34352 -2454 41222 -2448
rect 34352 -2520 34377 -2454
rect 34521 -2520 41222 -2454
rect 41314 -2520 48813 -2448
rect 34352 -2529 48813 -2520
rect 34629 -2530 48813 -2529
rect 47721 -2531 48813 -2530
rect 48841 -2405 59544 -2323
rect 33949 -2579 35303 -2578
rect 48841 -2579 48919 -2405
rect 59388 -2406 59544 -2405
rect 59593 -2012 59998 -2010
rect 59593 -2014 63291 -2012
rect 59593 -2021 63665 -2014
rect 59593 -2111 63168 -2021
rect 63252 -2111 63665 -2021
rect 59593 -2116 63665 -2111
rect 59593 -2117 63291 -2116
rect 59593 -2118 59998 -2117
rect 59593 -2446 59749 -2118
rect 63611 -2306 63665 -2116
rect 63727 -2262 63733 -1886
rect 63767 -2262 63773 -1886
rect 63727 -2274 63773 -2262
rect 63845 -1886 63891 -1874
rect 63845 -2262 63851 -1886
rect 63885 -2262 63891 -1886
rect 63845 -2274 63891 -2262
rect 63963 -1886 64009 -1874
rect 63963 -2262 63969 -1886
rect 64003 -2235 64009 -1886
rect 64080 -1886 64126 -1874
rect 64080 -2062 64086 -1886
rect 64120 -2062 64126 -1886
rect 64080 -2069 64126 -2062
rect 64198 -1886 64877 -1874
rect 64198 -2062 64204 -1886
rect 64238 -1899 64877 -1886
rect 64238 -2062 64244 -1899
rect 64488 -1979 64877 -1899
rect 64080 -2074 64129 -2069
rect 64198 -2074 64244 -2062
rect 65478 -2056 65512 -1762
rect 65775 -1950 65781 -1574
rect 65815 -1950 65821 -1574
rect 65775 -1962 65821 -1950
rect 65893 -1574 65939 -1562
rect 65893 -1950 65899 -1574
rect 65933 -1950 65939 -1574
rect 65893 -1962 65939 -1950
rect 66011 -1574 66057 -1562
rect 66011 -1950 66017 -1574
rect 66051 -1950 66057 -1574
rect 66011 -1962 66057 -1950
rect 66129 -1574 66175 -1562
rect 66129 -1950 66135 -1574
rect 66169 -1950 66175 -1574
rect 66129 -1962 66175 -1950
rect 66247 -1574 66293 -1562
rect 66247 -1950 66253 -1574
rect 66287 -1950 66293 -1574
rect 66653 -1574 66699 -1562
rect 66653 -1750 66659 -1574
rect 66693 -1750 66699 -1574
rect 66653 -1762 66699 -1750
rect 66771 -1574 66817 -1562
rect 66771 -1750 66777 -1574
rect 66811 -1750 66817 -1574
rect 66771 -1762 66817 -1750
rect 70365 -1597 70422 -1319
rect 70509 -1361 70909 -1355
rect 70509 -1395 70521 -1361
rect 70897 -1395 70909 -1361
rect 70509 -1401 70909 -1395
rect 70509 -1479 70909 -1473
rect 70509 -1513 70521 -1479
rect 70897 -1513 70909 -1479
rect 70509 -1519 70909 -1513
rect 70509 -1597 70909 -1591
rect 70365 -1631 70521 -1597
rect 70897 -1631 70909 -1597
rect 66247 -1962 66293 -1950
rect 66135 -2056 66169 -1962
rect 66659 -2056 66692 -1762
rect 64086 -2235 64129 -2074
rect 65478 -2088 66692 -2056
rect 64003 -2262 64129 -2235
rect 63963 -2274 64129 -2262
rect 63969 -2278 64129 -2274
rect 63611 -2312 63842 -2306
rect 63611 -2346 63792 -2312
rect 63826 -2346 63842 -2312
rect 63611 -2362 63842 -2346
rect 63894 -2312 63960 -2306
rect 63894 -2346 63910 -2312
rect 63944 -2346 63960 -2312
rect 33949 -2594 48919 -2579
rect 33949 -2665 33962 -2594
rect 34076 -2665 48919 -2594
rect 33949 -2680 48919 -2665
rect 48947 -2455 59749 -2446
rect 48947 -2523 54654 -2455
rect 54723 -2523 59749 -2455
rect 48947 -2530 59749 -2523
rect 59796 -2367 59952 -2365
rect 63480 -2367 63543 -2366
rect 59796 -2370 63555 -2367
rect 59796 -2445 63481 -2370
rect 63542 -2391 63555 -2370
rect 63894 -2391 63960 -2346
rect 63542 -2399 63960 -2391
rect 63542 -2431 63961 -2399
rect 64053 -2415 64129 -2278
rect 65844 -2112 66250 -2088
rect 65844 -2235 65956 -2112
rect 66130 -2235 66250 -2112
rect 70365 -2188 70422 -1631
rect 70509 -1637 70909 -1631
rect 70509 -1716 70909 -1710
rect 70509 -1750 70521 -1716
rect 70897 -1750 70909 -1716
rect 70509 -1756 70909 -1750
rect 70509 -1834 70909 -1828
rect 70509 -1868 70521 -1834
rect 70897 -1868 70909 -1834
rect 70509 -1874 70909 -1868
rect 70509 -1952 70909 -1946
rect 70509 -1986 70521 -1952
rect 70897 -1986 70909 -1952
rect 70509 -1992 70909 -1986
rect 70509 -2070 70909 -2064
rect 70993 -2070 71035 -923
rect 71095 -1067 71162 -15
rect 71195 -82 71280 -70
rect 71195 -153 71208 -82
rect 71271 -153 71280 -82
rect 71195 -162 71280 -153
rect 71672 -814 71719 -15
rect 71842 -814 72042 -809
rect 71672 -815 72042 -814
rect 71672 -848 71854 -815
rect 71095 -1101 71112 -1067
rect 71146 -1101 71162 -1067
rect 71095 -1117 71162 -1101
rect 71483 -1049 71568 -1037
rect 71483 -1117 71491 -1049
rect 71556 -1117 71568 -1049
rect 71483 -1129 71568 -1117
rect 71198 -1167 71283 -1155
rect 71198 -1237 71208 -1167
rect 71270 -1237 71283 -1167
rect 71198 -1247 71283 -1237
rect 71672 -1286 71719 -848
rect 71842 -849 71854 -848
rect 72030 -849 72042 -815
rect 71842 -855 72042 -849
rect 71842 -933 72042 -927
rect 71842 -967 71854 -933
rect 72030 -967 72461 -933
rect 71842 -1001 72042 -967
rect 71842 -1007 72242 -1001
rect 71842 -1041 71854 -1007
rect 72230 -1041 72242 -1007
rect 71842 -1047 72242 -1041
rect 71842 -1125 72242 -1119
rect 71842 -1159 71854 -1125
rect 72230 -1159 72242 -1125
rect 71842 -1165 72242 -1159
rect 71842 -1243 72242 -1237
rect 72315 -1243 72381 -1228
rect 71842 -1277 71854 -1243
rect 72230 -1244 72381 -1243
rect 72230 -1277 72331 -1244
rect 71842 -1283 72242 -1277
rect 72315 -1278 72331 -1277
rect 72365 -1278 72381 -1244
rect 71672 -1302 71782 -1286
rect 72315 -1294 72381 -1278
rect 72409 -1231 72461 -967
rect 72409 -1243 72539 -1231
rect 71672 -1336 71732 -1302
rect 71766 -1336 71782 -1302
rect 71672 -1352 71782 -1336
rect 72409 -1309 72483 -1243
rect 72535 -1309 72539 -1243
rect 72409 -1323 72539 -1309
rect 71842 -1361 72242 -1355
rect 71842 -1395 71854 -1361
rect 72230 -1395 72242 -1361
rect 71842 -1401 72242 -1395
rect 71322 -1408 71394 -1402
rect 71322 -1467 71328 -1408
rect 71388 -1467 71394 -1408
rect 71325 -1471 71392 -1467
rect 71328 -1477 71388 -1471
rect 71842 -1479 72242 -1473
rect 71842 -1513 71854 -1479
rect 72230 -1513 72242 -1479
rect 71842 -1519 72242 -1513
rect 71842 -1557 72042 -1519
rect 72409 -1557 72461 -1323
rect 71842 -1591 71854 -1557
rect 72030 -1591 72461 -1557
rect 71842 -1597 72042 -1591
rect 71671 -1675 71718 -1674
rect 71842 -1675 72042 -1669
rect 71671 -1709 71854 -1675
rect 72030 -1709 72042 -1675
rect 70509 -2104 70521 -2070
rect 70897 -2104 71121 -2070
rect 70509 -2110 70909 -2104
rect 70709 -2188 70909 -2183
rect 70365 -2189 70909 -2188
rect 70365 -2223 70721 -2189
rect 70897 -2223 70909 -2189
rect 70365 -2225 70909 -2223
rect 70709 -2229 70909 -2225
rect 65844 -2279 66250 -2235
rect 70709 -2307 70909 -2301
rect 70709 -2341 70721 -2307
rect 70897 -2341 70909 -2307
rect 70709 -2347 70909 -2341
rect 71055 -2377 71121 -2104
rect 71055 -2411 71071 -2377
rect 71105 -2411 71121 -2377
rect 63542 -2445 63555 -2431
rect 59796 -2455 63555 -2445
rect 33949 -2681 47803 -2680
rect 34629 -2682 47803 -2681
rect 33764 -2717 33904 -2716
rect 33764 -2718 35303 -2717
rect 36475 -2718 36681 -2716
rect 48947 -2718 49042 -2530
rect 33764 -2720 49042 -2718
rect 31375 -2768 31387 -2734
rect 31563 -2767 31901 -2734
rect 33761 -2726 49042 -2720
rect 31563 -2768 31575 -2767
rect 31375 -2774 31575 -2768
rect 33761 -2809 33773 -2726
rect 33880 -2732 49042 -2726
rect 33880 -2798 36506 -2732
rect 36650 -2798 49042 -2732
rect 33880 -2809 49042 -2798
rect 33761 -2815 49042 -2809
rect 33764 -2819 49042 -2815
rect 49070 -2580 53926 -2579
rect 59796 -2580 59952 -2455
rect 64049 -2475 64059 -2415
rect 64121 -2475 64131 -2415
rect 70709 -2425 70909 -2419
rect 70709 -2459 70721 -2425
rect 70897 -2459 70909 -2425
rect 71055 -2427 71121 -2411
rect 70709 -2465 70909 -2459
rect 49070 -2680 59952 -2580
rect 70709 -2543 70909 -2537
rect 71671 -2543 71718 -1709
rect 71842 -1715 72042 -1709
rect 70709 -2577 70721 -2543
rect 70897 -2577 71718 -2543
rect 70709 -2578 72913 -2577
rect 70709 -2583 70909 -2578
rect 71263 -2579 72913 -2578
rect 33764 -2820 33904 -2819
rect 34629 -2820 47572 -2819
rect 31375 -2852 31575 -2846
rect 30150 -2868 30350 -2862
rect 29804 -2902 30162 -2868
rect 30338 -2902 30350 -2868
rect 30150 -2908 30350 -2902
rect 30384 -2886 31387 -2852
rect 31563 -2886 31575 -2852
rect 49070 -2857 49160 -2680
rect 71263 -2697 73103 -2579
rect 72955 -2818 73103 -2697
rect 30150 -2986 30350 -2980
rect 30384 -2986 30419 -2886
rect 31375 -2892 31575 -2886
rect 36212 -2877 49160 -2857
rect 36212 -2931 36220 -2877
rect 36315 -2931 49160 -2877
rect 36212 -2938 49160 -2931
rect 72956 -2851 73103 -2818
rect 30150 -3020 30162 -2986
rect 30338 -3020 30419 -2986
rect 31053 -2950 31167 -2938
rect 30150 -3026 30350 -3020
rect 31053 -3052 31059 -2950
rect 31161 -3052 31167 -2950
rect 31053 -3064 31167 -3052
rect 72956 -3178 73105 -2851
rect 29541 -3179 73105 -3178
rect 29309 -3277 73105 -3179
rect 29309 -3282 29815 -3277
rect 29373 -3283 29815 -3282
rect 73208 -3341 73391 418
rect 29541 -3344 73391 -3341
rect 29148 -3428 73391 -3344
rect 29148 -3432 29829 -3428
rect 29218 -3434 29829 -3432
rect 28987 -3489 29807 -3485
rect 73479 -3489 73651 3549
rect 28987 -3587 73652 -3489
rect 28987 -3588 29807 -3587
rect 29038 -3592 29807 -3588
rect 28826 -3648 29602 -3647
rect 73729 -3648 73911 6693
rect 28826 -3745 73911 -3648
rect 28826 -3749 29602 -3745
rect 28833 -3754 29602 -3749
rect 28648 -3806 29664 -3804
rect 74004 -3806 74207 9895
rect 28648 -3896 74210 -3806
rect 28648 -3898 29664 -3896
rect 74281 -3957 74426 13040
rect 29541 -3959 74427 -3957
rect 28465 -4050 74427 -3959
rect 28465 -4052 29710 -4050
rect 28465 -4054 28581 -4052
rect 28309 -4111 29656 -4110
rect 74502 -4111 74653 16173
rect 28309 -4201 74653 -4111
rect 28309 -4203 29656 -4201
rect 28137 -4247 29692 -4243
rect 74716 -4247 74819 19315
rect 28137 -4337 74819 -4247
rect 28137 -4340 29692 -4337
rect 28137 -4341 28253 -4340
<< via1 >>
rect 38149 25093 38280 25215
rect 40041 24711 40173 24819
rect 42523 24765 42655 24873
rect 42924 24775 42980 24789
rect 42924 24741 42940 24775
rect 42940 24741 42974 24775
rect 42974 24741 42980 24775
rect 42924 24723 42980 24741
rect 43670 24765 43802 24873
rect 41794 24651 41860 24667
rect 41794 24617 41810 24651
rect 41810 24617 41844 24651
rect 41844 24617 41860 24651
rect 41794 24601 41860 24617
rect 46554 24708 46686 24816
rect 49036 24762 49168 24870
rect 4280 22234 4360 22240
rect 4280 22180 4284 22234
rect 4284 22180 4356 22234
rect 4356 22180 4360 22234
rect 7424 22234 7504 22240
rect 7424 22180 7428 22234
rect 7428 22180 7500 22234
rect 7500 22180 7504 22234
rect 10556 22230 10636 22236
rect 10556 22176 10560 22230
rect 10560 22176 10632 22230
rect 10632 22176 10636 22230
rect 13700 22230 13780 22236
rect 13700 22176 13704 22230
rect 13704 22176 13776 22230
rect 13776 22176 13780 22230
rect 16902 22234 16982 22240
rect 16902 22180 16906 22234
rect 16906 22180 16978 22234
rect 16978 22180 16982 22234
rect 20046 22234 20126 22240
rect 20046 22180 20050 22234
rect 20050 22180 20122 22234
rect 20122 22180 20126 22234
rect 23178 22230 23258 22236
rect 23178 22176 23182 22230
rect 23182 22176 23254 22230
rect 23254 22176 23258 22230
rect 2748 21167 2827 21234
rect 4352 21294 4422 21297
rect 4352 21239 4358 21294
rect 4358 21239 4418 21294
rect 4418 21239 4422 21294
rect 4352 21235 4422 21239
rect 5436 21293 5507 21297
rect 5436 21238 5443 21293
rect 5443 21238 5503 21293
rect 5503 21238 5507 21293
rect 5436 21234 5507 21238
rect 4122 21163 4181 21177
rect 4122 21129 4134 21163
rect 4134 21129 4168 21163
rect 4168 21129 4181 21163
rect 4122 21117 4181 21129
rect 4472 21009 4540 21014
rect 4472 20954 4476 21009
rect 4476 20954 4536 21009
rect 4536 20954 4540 21009
rect 4472 20949 4540 20954
rect 26322 22230 26402 22236
rect 26322 22176 26326 22230
rect 26326 22176 26398 22230
rect 26398 22176 26402 22230
rect 5694 21178 5751 21182
rect 5694 21118 5698 21178
rect 5698 21118 5747 21178
rect 5747 21118 5751 21178
rect 5694 21114 5751 21118
rect 7496 21294 7566 21297
rect 7496 21239 7502 21294
rect 7502 21239 7562 21294
rect 7562 21239 7566 21294
rect 7496 21235 7566 21239
rect 8580 21293 8651 21297
rect 8580 21238 8587 21293
rect 8587 21238 8647 21293
rect 8647 21238 8651 21293
rect 8580 21234 8651 21238
rect 7266 21163 7325 21177
rect 7266 21129 7278 21163
rect 7278 21129 7312 21163
rect 7312 21129 7325 21163
rect 7266 21117 7325 21129
rect 6012 20801 6065 20858
rect 7616 21009 7684 21014
rect 7616 20954 7620 21009
rect 7620 20954 7680 21009
rect 7680 20954 7684 21009
rect 7616 20949 7684 20954
rect 8838 21178 8895 21182
rect 8838 21118 8842 21178
rect 8842 21118 8891 21178
rect 8891 21118 8895 21178
rect 8838 21114 8895 21118
rect 10628 21290 10698 21293
rect 10628 21235 10634 21290
rect 10634 21235 10694 21290
rect 10694 21235 10698 21290
rect 10628 21231 10698 21235
rect 11712 21289 11783 21293
rect 11712 21234 11719 21289
rect 11719 21234 11779 21289
rect 11779 21234 11783 21289
rect 11712 21230 11783 21234
rect 10398 21159 10457 21173
rect 10398 21125 10410 21159
rect 10410 21125 10444 21159
rect 10444 21125 10457 21159
rect 10398 21113 10457 21125
rect 8838 21010 8895 21014
rect 8838 20950 8842 21010
rect 8842 20950 8891 21010
rect 8891 20950 8895 21010
rect 8838 20946 8895 20950
rect 4280 19976 4284 20022
rect 4284 19976 4342 20022
rect 4342 19976 4346 20022
rect 4280 19970 4346 19976
rect 7424 19976 7428 20022
rect 7428 19976 7486 20022
rect 7486 19976 7490 20022
rect 7424 19970 7490 19976
rect 10748 21005 10816 21010
rect 10748 20950 10752 21005
rect 10752 20950 10812 21005
rect 10812 20950 10816 21005
rect 10748 20945 10816 20950
rect 11970 21174 12027 21178
rect 11970 21114 11974 21174
rect 11974 21114 12023 21174
rect 12023 21114 12027 21174
rect 11970 21110 12027 21114
rect 13772 21290 13842 21293
rect 13772 21235 13778 21290
rect 13778 21235 13838 21290
rect 13838 21235 13842 21290
rect 13772 21231 13842 21235
rect 14856 21289 14927 21293
rect 14856 21234 14863 21289
rect 14863 21234 14923 21289
rect 14923 21234 14927 21289
rect 14856 21230 14927 21234
rect 13542 21159 13601 21173
rect 13542 21125 13554 21159
rect 13554 21125 13588 21159
rect 13588 21125 13601 21159
rect 13542 21113 13601 21125
rect 11970 21006 12027 21010
rect 11970 20946 11974 21006
rect 11974 20946 12023 21006
rect 12023 20946 12027 21006
rect 11970 20942 12027 20946
rect 9146 20672 9210 20731
rect 13892 21005 13960 21010
rect 13892 20950 13896 21005
rect 13896 20950 13956 21005
rect 13956 20950 13960 21005
rect 13892 20945 13960 20950
rect 16974 21294 17044 21297
rect 16974 21239 16980 21294
rect 16980 21239 17040 21294
rect 17040 21239 17044 21294
rect 16974 21235 17044 21239
rect 18058 21293 18129 21297
rect 18058 21238 18065 21293
rect 18065 21238 18125 21293
rect 18125 21238 18129 21293
rect 18058 21234 18129 21238
rect 16744 21163 16803 21177
rect 16744 21129 16756 21163
rect 16756 21129 16790 21163
rect 16790 21129 16803 21163
rect 16744 21117 16803 21129
rect 15114 21006 15171 21010
rect 15114 20946 15118 21006
rect 15118 20946 15167 21006
rect 15167 20946 15171 21006
rect 15114 20942 15171 20946
rect 12290 20509 12346 20578
rect 12084 20100 12141 20167
rect 17094 21009 17162 21014
rect 17094 20954 17098 21009
rect 17098 20954 17158 21009
rect 17158 20954 17162 21009
rect 17094 20949 17162 20954
rect 18316 21178 18373 21182
rect 18316 21118 18320 21178
rect 18320 21118 18369 21178
rect 18369 21118 18373 21178
rect 18316 21114 18373 21118
rect 20118 21294 20188 21297
rect 20118 21239 20124 21294
rect 20124 21239 20184 21294
rect 20184 21239 20188 21294
rect 20118 21235 20188 21239
rect 21202 21293 21273 21297
rect 21202 21238 21209 21293
rect 21209 21238 21269 21293
rect 21269 21238 21273 21293
rect 21202 21234 21273 21238
rect 19888 21163 19947 21177
rect 19888 21129 19900 21163
rect 19900 21129 19934 21163
rect 19934 21129 19947 21163
rect 19888 21117 19947 21129
rect 18316 21010 18373 21014
rect 18316 20950 18320 21010
rect 18320 20950 18369 21010
rect 18369 20950 18373 21010
rect 18316 20946 18373 20950
rect 15509 20359 15571 20427
rect 15223 20241 15292 20302
rect 18408 20468 18462 20526
rect 20238 21009 20306 21014
rect 20238 20954 20242 21009
rect 20242 20954 20302 21009
rect 20302 20954 20306 21009
rect 20238 20949 20306 20954
rect 24704 21343 24764 21396
rect 23250 21290 23320 21293
rect 23250 21235 23256 21290
rect 23256 21235 23316 21290
rect 23316 21235 23320 21290
rect 23250 21231 23320 21235
rect 24334 21289 24405 21293
rect 24334 21234 24341 21289
rect 24341 21234 24401 21289
rect 24401 21234 24405 21289
rect 24334 21230 24405 21234
rect 23020 21159 23079 21173
rect 23020 21125 23032 21159
rect 23032 21125 23066 21159
rect 23066 21125 23079 21159
rect 23020 21113 23079 21125
rect 21460 21010 21517 21014
rect 21460 20950 21464 21010
rect 21464 20950 21513 21010
rect 21513 20950 21517 21010
rect 21460 20946 21517 20950
rect 18687 20222 18746 20279
rect 21540 20574 21604 20631
rect 23370 21005 23438 21010
rect 23370 20950 23374 21005
rect 23374 20950 23434 21005
rect 23434 20950 23438 21005
rect 23370 20945 23438 20950
rect 27738 21381 27792 21443
rect 27952 21436 28039 21443
rect 27952 21392 28039 21436
rect 27952 21386 28039 21392
rect 24592 21174 24649 21178
rect 24592 21114 24596 21174
rect 24596 21114 24645 21174
rect 24645 21114 24649 21174
rect 24592 21110 24649 21114
rect 26394 21290 26464 21293
rect 26394 21235 26400 21290
rect 26400 21235 26460 21290
rect 26460 21235 26464 21290
rect 26394 21231 26464 21235
rect 27478 21289 27549 21293
rect 27478 21234 27485 21289
rect 27485 21234 27545 21289
rect 27545 21234 27549 21289
rect 27478 21230 27549 21234
rect 26164 21159 26223 21173
rect 26164 21125 26176 21159
rect 26176 21125 26210 21159
rect 26210 21125 26223 21159
rect 26164 21113 26223 21125
rect 24592 21006 24649 21010
rect 24592 20946 24596 21006
rect 24596 20946 24645 21006
rect 24645 20946 24649 21006
rect 24592 20942 24649 20946
rect 24684 20712 24754 20772
rect 21813 20096 21872 20162
rect 10556 19972 10560 20018
rect 10560 19972 10618 20018
rect 10618 19972 10622 20018
rect 10556 19966 10622 19972
rect 13700 19972 13704 20018
rect 13704 19972 13762 20018
rect 13762 19972 13766 20018
rect 13700 19966 13766 19972
rect 16902 19976 16906 20022
rect 16906 19976 16964 20022
rect 16964 19976 16968 20022
rect 16902 19970 16968 19976
rect 20046 19976 20050 20022
rect 20050 19976 20108 20022
rect 20108 19976 20112 20022
rect 20046 19970 20112 19976
rect 23178 19972 23182 20018
rect 23182 19972 23240 20018
rect 23240 19972 23244 20018
rect 23178 19966 23244 19972
rect 8942 19875 9012 19951
rect 26514 21005 26582 21010
rect 26514 20950 26518 21005
rect 26518 20950 26578 21005
rect 26578 20950 26582 21005
rect 26514 20945 26582 20950
rect 27736 21290 27793 21294
rect 27736 21230 27740 21290
rect 27740 21230 27789 21290
rect 27789 21230 27793 21290
rect 27736 21226 27793 21230
rect 27736 21006 27793 21010
rect 27736 20946 27740 21006
rect 27740 20946 27789 21006
rect 27789 20946 27793 21006
rect 27957 20998 28037 21009
rect 27957 20954 28037 20998
rect 27957 20947 28037 20954
rect 27736 20942 27793 20946
rect 27739 20706 27793 20768
rect 27739 20571 27793 20633
rect 27956 20622 28038 20663
rect 27956 20611 28038 20622
rect 27737 20459 27791 20521
rect 27949 20512 28039 20521
rect 27949 20468 27950 20512
rect 27950 20468 28039 20512
rect 27949 20464 28039 20468
rect 27737 20334 27791 20396
rect 27945 20385 28046 20392
rect 27945 20341 27949 20385
rect 27949 20341 28042 20385
rect 28042 20341 28046 20385
rect 27945 20339 28046 20341
rect 42460 23954 42559 24051
rect 40321 23648 40429 23780
rect 28535 20861 28595 20865
rect 28535 20820 28541 20861
rect 28541 20820 28591 20861
rect 28591 20820 28595 20861
rect 28535 20813 28595 20820
rect 28883 20572 28958 20640
rect 27732 20093 27786 20155
rect 29020 20154 29090 20222
rect 32926 20169 33084 20306
rect 27945 20147 28045 20150
rect 27945 20103 27949 20147
rect 27949 20103 28042 20147
rect 28042 20103 28045 20147
rect 27945 20098 28045 20103
rect 26322 19972 26326 20018
rect 26326 19972 26384 20018
rect 26384 19972 26388 20018
rect 26322 19966 26388 19972
rect 24932 19801 25005 19882
rect 27735 19871 27789 19933
rect 27945 19923 28043 19929
rect 27945 19879 27948 19923
rect 27948 19879 28041 19923
rect 28041 19879 28043 19923
rect 27945 19875 28043 19879
rect 28779 19724 28832 19793
rect -1493 19498 -1401 19562
rect -1493 19383 -1401 19447
rect -1493 19262 -1401 19326
rect -1493 19143 -1401 19207
rect -1493 19029 -1401 19093
rect -1493 18915 -1401 18979
rect -1492 18800 -1400 18864
rect -1492 18686 -1400 18750
rect 15050 18561 15104 18615
rect 27826 18577 27886 18636
rect 28671 19300 28724 19365
rect 4638 16975 4690 17027
rect 14956 18468 15010 18522
rect 16588 18376 16642 18430
rect 5806 16975 5858 17027
rect 16413 18281 16467 18335
rect 18049 18191 18103 18245
rect 6974 16975 7026 17027
rect 17911 18097 17965 18151
rect 19551 18003 19605 18057
rect 19372 17909 19426 17963
rect 8142 16975 8194 17027
rect 21007 17819 21061 17873
rect 20879 17724 20933 17778
rect 9316 16973 9368 17025
rect 22460 17633 22514 17687
rect 22329 17538 22383 17592
rect 10484 16973 10536 17025
rect 23905 17447 23959 17501
rect 23795 17354 23849 17408
rect 11652 16973 11704 17025
rect 12820 16973 12872 17025
rect 14498 16777 14558 16839
rect 15946 16777 16006 16839
rect 17444 16775 17504 16837
rect 18892 16775 18952 16837
rect 20412 16777 20472 16839
rect 21860 16777 21920 16839
rect 23358 16775 23418 16837
rect 24806 16775 24866 16837
rect 5109 15651 5161 15703
rect 6277 15651 6329 15703
rect 7445 15651 7497 15703
rect 8613 15651 8665 15703
rect 9787 15649 9839 15701
rect 10955 15649 11007 15701
rect 12123 15649 12175 15701
rect 13291 15649 13343 15701
rect 14716 15942 14802 16030
rect 14830 15813 14916 15901
rect 14274 15627 14336 15635
rect 14274 15581 14278 15627
rect 14278 15581 14330 15627
rect 14330 15581 14336 15627
rect 14274 15575 14336 15581
rect 16180 15960 16234 16014
rect 16292 15830 16346 15884
rect 15722 15627 15784 15635
rect 15722 15581 15726 15627
rect 15726 15581 15778 15627
rect 15778 15581 15784 15627
rect 15722 15575 15784 15581
rect 17677 15962 17731 16016
rect 17789 15824 17843 15878
rect 17220 15625 17282 15633
rect 17220 15579 17224 15625
rect 17224 15579 17276 15625
rect 17276 15579 17282 15625
rect 17220 15573 17282 15579
rect 19125 15955 19179 16009
rect 19241 15830 19295 15884
rect 18668 15625 18730 15633
rect 18668 15579 18672 15625
rect 18672 15579 18724 15625
rect 18724 15579 18730 15625
rect 18668 15573 18730 15579
rect 20644 15960 20698 16014
rect 20757 15830 20811 15884
rect 20188 15627 20250 15635
rect 20188 15581 20192 15627
rect 20192 15581 20244 15627
rect 20244 15581 20250 15627
rect 20188 15575 20250 15581
rect 1778 15096 1858 15102
rect 1778 15042 1782 15096
rect 1782 15042 1854 15096
rect 1854 15042 1858 15096
rect 1850 14156 1920 14159
rect 1850 14101 1856 14156
rect 1856 14101 1916 14156
rect 1916 14101 1920 14156
rect 1850 14097 1920 14101
rect 2934 14155 3005 14159
rect 2934 14100 2941 14155
rect 2941 14100 3001 14155
rect 3001 14100 3005 14155
rect 2934 14096 3005 14100
rect 1620 14025 1679 14039
rect 1620 13991 1632 14025
rect 1632 13991 1666 14025
rect 1666 13991 1679 14025
rect 1620 13979 1679 13991
rect 1970 13871 2038 13876
rect 1970 13816 1974 13871
rect 1974 13816 2034 13871
rect 2034 13816 2038 13871
rect 1970 13811 2038 13816
rect 4922 15096 5002 15102
rect 4922 15042 4926 15096
rect 4926 15042 4998 15096
rect 4998 15042 5002 15096
rect 3192 14040 3249 14044
rect 3192 13980 3196 14040
rect 3196 13980 3245 14040
rect 3245 13980 3249 14040
rect 3192 13976 3249 13980
rect 4994 14156 5064 14159
rect 4994 14101 5000 14156
rect 5000 14101 5060 14156
rect 5060 14101 5064 14156
rect 4994 14097 5064 14101
rect 6078 14155 6149 14159
rect 6078 14100 6085 14155
rect 6085 14100 6145 14155
rect 6145 14100 6149 14155
rect 6078 14096 6149 14100
rect 4764 14025 4823 14039
rect 4764 13991 4776 14025
rect 4776 13991 4810 14025
rect 4810 13991 4823 14025
rect 4764 13979 4823 13991
rect 3192 13872 3249 13876
rect 3192 13812 3196 13872
rect 3196 13812 3245 13872
rect 3245 13812 3249 13872
rect 3192 13808 3249 13812
rect 1778 12838 1782 12884
rect 1782 12838 1840 12884
rect 1840 12838 1844 12884
rect 1778 12832 1844 12838
rect 1778 12362 1858 12368
rect 1778 12308 1782 12362
rect 1782 12308 1854 12362
rect 1854 12308 1858 12362
rect 80 11232 191 11361
rect 1850 11422 1920 11425
rect 1850 11367 1856 11422
rect 1856 11367 1916 11422
rect 1916 11367 1920 11422
rect 1850 11363 1920 11367
rect 2934 11421 3005 11425
rect 2934 11366 2941 11421
rect 2941 11366 3001 11421
rect 3001 11366 3005 11421
rect 2934 11362 3005 11366
rect 1620 11291 1679 11305
rect 1620 11257 1632 11291
rect 1632 11257 1666 11291
rect 1666 11257 1679 11291
rect 1620 11245 1679 11257
rect 1970 11137 2038 11142
rect 1970 11082 1974 11137
rect 1974 11082 2034 11137
rect 2034 11082 2038 11137
rect 1970 11077 2038 11082
rect -547 10879 -425 10936
rect 142 10867 201 10937
rect 5114 13871 5182 13876
rect 5114 13816 5118 13871
rect 5118 13816 5178 13871
rect 5178 13816 5182 13871
rect 5114 13811 5182 13816
rect 22094 15957 22148 16011
rect 22205 15825 22259 15879
rect 21636 15627 21698 15635
rect 21636 15581 21640 15627
rect 21640 15581 21692 15627
rect 21692 15581 21698 15627
rect 21636 15575 21698 15581
rect 23588 15958 23642 16012
rect 23703 15826 23757 15881
rect 23134 15625 23196 15633
rect 23134 15579 23138 15625
rect 23138 15579 23190 15625
rect 23190 15579 23196 15625
rect 23134 15573 23196 15579
rect 25630 16122 25701 16181
rect 25346 16021 25415 16085
rect 24582 15625 24644 15633
rect 24582 15579 24586 15625
rect 24586 15579 24638 15625
rect 24638 15579 24644 15625
rect 24582 15573 24644 15579
rect 8054 15092 8134 15098
rect 8054 15038 8058 15092
rect 8058 15038 8130 15092
rect 8130 15038 8134 15092
rect 6336 14040 6393 14044
rect 6336 13980 6340 14040
rect 6340 13980 6389 14040
rect 6389 13980 6393 14040
rect 6336 13976 6393 13980
rect 8126 14152 8196 14155
rect 8126 14097 8132 14152
rect 8132 14097 8192 14152
rect 8192 14097 8196 14152
rect 8126 14093 8196 14097
rect 9210 14151 9281 14155
rect 9210 14096 9217 14151
rect 9217 14096 9277 14151
rect 9277 14096 9281 14151
rect 9210 14092 9281 14096
rect 7896 14021 7955 14035
rect 7896 13987 7908 14021
rect 7908 13987 7942 14021
rect 7942 13987 7955 14021
rect 7896 13975 7955 13987
rect 6336 13872 6393 13876
rect 6336 13812 6340 13872
rect 6340 13812 6389 13872
rect 6389 13812 6393 13872
rect 6336 13808 6393 13812
rect 4922 12838 4926 12884
rect 4926 12838 4984 12884
rect 4984 12838 4988 12884
rect 4922 12832 4988 12838
rect 8246 13867 8314 13872
rect 8246 13812 8250 13867
rect 8250 13812 8310 13867
rect 8310 13812 8314 13867
rect 8246 13807 8314 13812
rect 11198 15092 11278 15098
rect 11198 15038 11202 15092
rect 11202 15038 11274 15092
rect 11274 15038 11278 15092
rect 9468 14036 9525 14040
rect 9468 13976 9472 14036
rect 9472 13976 9521 14036
rect 9521 13976 9525 14036
rect 9468 13972 9525 13976
rect 11270 14152 11340 14155
rect 11270 14097 11276 14152
rect 11276 14097 11336 14152
rect 11336 14097 11340 14152
rect 11270 14093 11340 14097
rect 12354 14151 12425 14155
rect 12354 14096 12361 14151
rect 12361 14096 12421 14151
rect 12421 14096 12425 14151
rect 12354 14092 12425 14096
rect 11040 14021 11099 14035
rect 11040 13987 11052 14021
rect 11052 13987 11086 14021
rect 11086 13987 11099 14021
rect 11040 13975 11099 13987
rect 9468 13868 9525 13872
rect 9468 13808 9472 13868
rect 9472 13808 9521 13868
rect 9521 13808 9525 13868
rect 9468 13804 9525 13808
rect 8054 12834 8058 12880
rect 8058 12834 8116 12880
rect 8116 12834 8120 12880
rect 8054 12828 8120 12834
rect 14400 15096 14480 15102
rect 14400 15042 14404 15096
rect 14404 15042 14476 15096
rect 14476 15042 14480 15096
rect 12612 14036 12669 14040
rect 12612 13976 12616 14036
rect 12616 13976 12665 14036
rect 12665 13976 12669 14036
rect 12612 13972 12669 13976
rect 14472 14156 14542 14159
rect 14472 14101 14478 14156
rect 14478 14101 14538 14156
rect 14538 14101 14542 14156
rect 14472 14097 14542 14101
rect 15556 14155 15627 14159
rect 15556 14100 15563 14155
rect 15563 14100 15623 14155
rect 15623 14100 15627 14155
rect 15556 14096 15627 14100
rect 14242 14025 14301 14039
rect 14242 13991 14254 14025
rect 14254 13991 14288 14025
rect 14288 13991 14301 14025
rect 14242 13979 14301 13991
rect 11198 12834 11202 12880
rect 11202 12834 11260 12880
rect 11260 12834 11264 12880
rect 11198 12828 11264 12834
rect 17544 15096 17624 15102
rect 17544 15042 17548 15096
rect 17548 15042 17620 15096
rect 17620 15042 17624 15096
rect 15814 14040 15871 14044
rect 15814 13980 15818 14040
rect 15818 13980 15867 14040
rect 15867 13980 15871 14040
rect 15814 13976 15871 13980
rect 17616 14156 17686 14159
rect 17616 14101 17622 14156
rect 17622 14101 17682 14156
rect 17682 14101 17686 14156
rect 17616 14097 17686 14101
rect 18700 14155 18771 14159
rect 18700 14100 18707 14155
rect 18707 14100 18767 14155
rect 18767 14100 18771 14155
rect 18700 14096 18771 14100
rect 17386 14025 17445 14039
rect 17386 13991 17398 14025
rect 17398 13991 17432 14025
rect 17432 13991 17445 14025
rect 17386 13979 17445 13991
rect 14400 12838 14404 12884
rect 14404 12838 14462 12884
rect 14462 12838 14466 12884
rect 14400 12832 14466 12838
rect 17736 13871 17804 13876
rect 17736 13816 17740 13871
rect 17740 13816 17800 13871
rect 17800 13816 17804 13871
rect 17736 13811 17804 13816
rect 20676 15092 20756 15098
rect 20676 15038 20680 15092
rect 20680 15038 20752 15092
rect 20752 15038 20756 15092
rect 18958 14040 19015 14044
rect 18958 13980 18962 14040
rect 18962 13980 19011 14040
rect 19011 13980 19015 14040
rect 18958 13976 19015 13980
rect 20748 14152 20818 14155
rect 20748 14097 20754 14152
rect 20754 14097 20814 14152
rect 20814 14097 20818 14152
rect 20748 14093 20818 14097
rect 21832 14151 21903 14155
rect 21832 14096 21839 14151
rect 21839 14096 21899 14151
rect 21899 14096 21903 14151
rect 21832 14092 21903 14096
rect 20518 14021 20577 14035
rect 20518 13987 20530 14021
rect 20530 13987 20564 14021
rect 20564 13987 20577 14021
rect 20518 13975 20577 13987
rect 18958 13872 19015 13876
rect 18958 13812 18962 13872
rect 18962 13812 19011 13872
rect 19011 13812 19015 13872
rect 18958 13808 19015 13812
rect 17544 12838 17548 12884
rect 17548 12838 17606 12884
rect 17606 12838 17610 12884
rect 17544 12832 17610 12838
rect 20868 13867 20936 13872
rect 20868 13812 20872 13867
rect 20872 13812 20932 13867
rect 20932 13812 20936 13867
rect 20868 13807 20936 13812
rect 23820 15092 23900 15098
rect 23820 15038 23824 15092
rect 23824 15038 23896 15092
rect 23896 15038 23900 15092
rect 22090 14036 22147 14040
rect 22090 13976 22094 14036
rect 22094 13976 22143 14036
rect 22143 13976 22147 14036
rect 22090 13972 22147 13976
rect 23892 14152 23962 14155
rect 23892 14097 23898 14152
rect 23898 14097 23958 14152
rect 23958 14097 23962 14152
rect 23892 14093 23962 14097
rect 24976 14151 25047 14155
rect 24976 14096 24983 14151
rect 24983 14096 25043 14151
rect 25043 14096 25047 14151
rect 24976 14092 25047 14096
rect 23662 14021 23721 14035
rect 23662 13987 23674 14021
rect 23674 13987 23708 14021
rect 23708 13987 23721 14021
rect 23662 13975 23721 13987
rect 22090 13868 22147 13872
rect 22090 13808 22094 13868
rect 22094 13808 22143 13868
rect 22143 13808 22147 13868
rect 22090 13804 22147 13808
rect 20676 12834 20680 12880
rect 20680 12834 20738 12880
rect 20738 12834 20742 12880
rect 20676 12828 20742 12834
rect 24012 13867 24080 13872
rect 24012 13812 24016 13867
rect 24016 13812 24076 13867
rect 24076 13812 24080 13867
rect 24012 13807 24080 13812
rect 25234 14036 25291 14040
rect 25234 13976 25238 14036
rect 25238 13976 25287 14036
rect 25287 13976 25291 14036
rect 25234 13972 25291 13976
rect 25828 14070 25911 14158
rect 25234 13868 25291 13872
rect 25234 13808 25238 13868
rect 25238 13808 25287 13868
rect 25287 13808 25291 13868
rect 25234 13804 25291 13808
rect 23820 12834 23824 12880
rect 23824 12834 23882 12880
rect 23882 12834 23886 12880
rect 23820 12828 23886 12834
rect 4922 12362 5002 12368
rect 4922 12308 4926 12362
rect 4926 12308 4998 12362
rect 4998 12308 5002 12362
rect 3192 11306 3249 11310
rect 3192 11246 3196 11306
rect 3196 11246 3245 11306
rect 3245 11246 3249 11306
rect 3192 11242 3249 11246
rect 4994 11422 5064 11425
rect 4994 11367 5000 11422
rect 5000 11367 5060 11422
rect 5060 11367 5064 11422
rect 4994 11363 5064 11367
rect 6078 11421 6149 11425
rect 6078 11366 6085 11421
rect 6085 11366 6145 11421
rect 6145 11366 6149 11421
rect 6078 11362 6149 11366
rect 4764 11291 4823 11305
rect 4764 11257 4776 11291
rect 4776 11257 4810 11291
rect 4810 11257 4823 11291
rect 4764 11245 4823 11257
rect 3192 11138 3249 11142
rect 3192 11078 3196 11138
rect 3196 11078 3245 11138
rect 3245 11078 3249 11138
rect 3192 11074 3249 11078
rect -783 10687 -661 10744
rect 141 10682 202 10745
rect -1048 10459 -926 10516
rect 141 10459 203 10525
rect -1255 10274 -1133 10331
rect 140 10271 203 10329
rect 1778 10104 1782 10150
rect 1782 10104 1840 10150
rect 1840 10104 1844 10150
rect 1778 10098 1844 10104
rect -1515 9927 -1393 9984
rect 140 9925 204 9986
rect 3520 10859 3591 10930
rect 5114 11137 5182 11142
rect 5114 11082 5118 11137
rect 5118 11082 5178 11137
rect 5178 11082 5182 11137
rect 5114 11077 5182 11082
rect 8054 12358 8134 12364
rect 8054 12304 8058 12358
rect 8058 12304 8130 12358
rect 8130 12304 8134 12358
rect 6336 11306 6393 11310
rect 6336 11246 6340 11306
rect 6340 11246 6389 11306
rect 6389 11246 6393 11306
rect 6336 11242 6393 11246
rect 8126 11418 8196 11421
rect 8126 11363 8132 11418
rect 8132 11363 8192 11418
rect 8192 11363 8196 11418
rect 8126 11359 8196 11363
rect 9210 11417 9281 11421
rect 9210 11362 9217 11417
rect 9217 11362 9277 11417
rect 9277 11362 9281 11417
rect 9210 11358 9281 11362
rect 7896 11287 7955 11301
rect 7896 11253 7908 11287
rect 7908 11253 7942 11287
rect 7942 11253 7955 11287
rect 7896 11241 7955 11253
rect 6336 11138 6393 11142
rect 6336 11078 6340 11138
rect 6340 11078 6389 11138
rect 6389 11078 6393 11138
rect 6336 11074 6393 11078
rect 4922 10104 4926 10150
rect 4926 10104 4984 10150
rect 4984 10104 4988 10150
rect 4922 10098 4988 10104
rect 8246 11133 8314 11138
rect 8246 11078 8250 11133
rect 8250 11078 8310 11133
rect 8310 11078 8314 11133
rect 8246 11073 8314 11078
rect 9468 11418 9525 11422
rect 9468 11358 9472 11418
rect 9472 11358 9521 11418
rect 9521 11358 9525 11418
rect 9468 11354 9525 11358
rect 11198 12358 11278 12364
rect 11198 12304 11202 12358
rect 11202 12304 11274 12358
rect 11274 12304 11278 12358
rect 9468 11302 9525 11306
rect 9468 11242 9472 11302
rect 9472 11242 9521 11302
rect 9521 11242 9525 11302
rect 9468 11238 9525 11242
rect 11270 11418 11340 11421
rect 11270 11363 11276 11418
rect 11276 11363 11336 11418
rect 11336 11363 11340 11418
rect 11270 11359 11340 11363
rect 12354 11417 12425 11421
rect 12354 11362 12361 11417
rect 12361 11362 12421 11417
rect 12421 11362 12425 11417
rect 12354 11358 12425 11362
rect 11040 11287 11099 11301
rect 11040 11253 11052 11287
rect 11052 11253 11086 11287
rect 11086 11253 11099 11287
rect 11040 11241 11099 11253
rect 9468 11134 9525 11138
rect 9468 11074 9472 11134
rect 9472 11074 9521 11134
rect 9521 11074 9525 11134
rect 9468 11070 9525 11074
rect 6650 10678 6720 10771
rect 8054 10100 8058 10146
rect 8058 10100 8116 10146
rect 8116 10100 8120 10146
rect 8054 10094 8120 10100
rect 11390 11133 11458 11138
rect 11390 11078 11394 11133
rect 11394 11078 11454 11133
rect 11454 11078 11458 11133
rect 11390 11073 11458 11078
rect 14400 12362 14480 12368
rect 14400 12308 14404 12362
rect 14404 12308 14476 12362
rect 14476 12308 14480 12362
rect 12612 11302 12669 11306
rect 12612 11242 12616 11302
rect 12616 11242 12665 11302
rect 12665 11242 12669 11302
rect 12612 11238 12669 11242
rect 14472 11422 14542 11425
rect 14472 11367 14478 11422
rect 14478 11367 14538 11422
rect 14538 11367 14542 11422
rect 14472 11363 14542 11367
rect 15556 11421 15627 11425
rect 15556 11366 15563 11421
rect 15563 11366 15623 11421
rect 15623 11366 15627 11421
rect 15556 11362 15627 11366
rect 14242 11291 14301 11305
rect 14242 11257 14254 11291
rect 14254 11257 14288 11291
rect 14288 11257 14301 11291
rect 14242 11245 14301 11257
rect 12612 11134 12669 11138
rect 12612 11074 12616 11134
rect 12616 11074 12665 11134
rect 12665 11074 12669 11134
rect 12612 11070 12669 11074
rect 9783 10445 9879 10540
rect 11198 10100 11202 10146
rect 11202 10100 11260 10146
rect 11260 10100 11264 10146
rect 11198 10094 11264 10100
rect 14592 11137 14660 11142
rect 14592 11082 14596 11137
rect 14596 11082 14656 11137
rect 14656 11082 14660 11137
rect 14592 11077 14660 11082
rect 17544 12362 17624 12368
rect 17544 12308 17548 12362
rect 17548 12308 17620 12362
rect 17620 12308 17624 12362
rect 15814 11306 15871 11310
rect 15814 11246 15818 11306
rect 15818 11246 15867 11306
rect 15867 11246 15871 11306
rect 15814 11242 15871 11246
rect 17616 11422 17686 11425
rect 17616 11367 17622 11422
rect 17622 11367 17682 11422
rect 17682 11367 17686 11422
rect 17616 11363 17686 11367
rect 18700 11421 18771 11425
rect 18700 11366 18707 11421
rect 18707 11366 18767 11421
rect 18767 11366 18771 11421
rect 18700 11362 18771 11366
rect 17386 11291 17445 11305
rect 17386 11257 17398 11291
rect 17398 11257 17432 11291
rect 17432 11257 17445 11291
rect 17386 11245 17445 11257
rect 15814 11138 15871 11142
rect 15814 11078 15818 11138
rect 15818 11078 15867 11138
rect 15867 11078 15871 11138
rect 15814 11074 15871 11078
rect 13001 10267 13079 10336
rect 14400 10104 14404 10150
rect 14404 10104 14462 10150
rect 14462 10104 14466 10150
rect 14400 10098 14466 10104
rect -1730 9758 -1608 9815
rect 138 9754 202 9814
rect 17736 11137 17804 11142
rect 17736 11082 17740 11137
rect 17740 11082 17800 11137
rect 17800 11082 17804 11137
rect 17736 11077 17804 11082
rect 20676 12358 20756 12364
rect 20676 12304 20680 12358
rect 20680 12304 20752 12358
rect 20752 12304 20756 12358
rect 18958 11306 19015 11310
rect 18958 11246 18962 11306
rect 18962 11246 19011 11306
rect 19011 11246 19015 11306
rect 18958 11242 19015 11246
rect 20748 11418 20818 11421
rect 20748 11363 20754 11418
rect 20754 11363 20814 11418
rect 20814 11363 20818 11418
rect 20748 11359 20818 11363
rect 21832 11417 21903 11421
rect 21832 11362 21839 11417
rect 21839 11362 21899 11417
rect 21899 11362 21903 11417
rect 21832 11358 21903 11362
rect 20518 11287 20577 11301
rect 20518 11253 20530 11287
rect 20530 11253 20564 11287
rect 20564 11253 20577 11287
rect 20518 11241 20577 11253
rect 18958 11138 19015 11142
rect 18958 11078 18962 11138
rect 18962 11078 19011 11138
rect 19011 11078 19015 11138
rect 18958 11074 19015 11078
rect 17544 10104 17548 10150
rect 17548 10104 17606 10150
rect 17606 10104 17610 10150
rect 17544 10098 17610 10104
rect 16159 9924 16226 9992
rect 20868 11133 20936 11138
rect 20868 11078 20872 11133
rect 20872 11078 20932 11133
rect 20932 11078 20936 11133
rect 20868 11073 20936 11078
rect 23820 12358 23900 12364
rect 23820 12304 23824 12358
rect 23824 12304 23896 12358
rect 23896 12304 23900 12358
rect 22090 11302 22147 11306
rect 22090 11242 22094 11302
rect 22094 11242 22143 11302
rect 22143 11242 22147 11302
rect 22090 11238 22147 11242
rect 23892 11418 23962 11421
rect 23892 11363 23898 11418
rect 23898 11363 23958 11418
rect 23958 11363 23962 11418
rect 23892 11359 23962 11363
rect 24976 11417 25047 11421
rect 24976 11362 24983 11417
rect 24983 11362 25043 11417
rect 25043 11362 25047 11417
rect 24976 11358 25047 11362
rect 23662 11287 23721 11301
rect 23662 11253 23674 11287
rect 23674 11253 23708 11287
rect 23708 11253 23721 11287
rect 23662 11241 23721 11253
rect 22090 11134 22147 11138
rect 22090 11074 22094 11134
rect 22094 11074 22143 11134
rect 22143 11074 22147 11134
rect 22090 11070 22147 11074
rect 19294 10046 19362 10118
rect 20676 10100 20680 10146
rect 20680 10100 20738 10146
rect 20738 10100 20742 10146
rect 20676 10094 20742 10100
rect 24012 11133 24080 11138
rect 24012 11078 24016 11133
rect 24016 11078 24076 11133
rect 24076 11078 24080 11133
rect 24012 11073 24080 11078
rect 25234 11302 25291 11306
rect 25234 11242 25238 11302
rect 25238 11242 25287 11302
rect 25287 11242 25291 11302
rect 25234 11238 25291 11242
rect 25234 11134 25291 11138
rect 25234 11074 25238 11134
rect 25238 11074 25287 11134
rect 25287 11074 25291 11134
rect 25234 11070 25291 11074
rect 22408 10100 22472 10177
rect 23820 10100 23824 10146
rect 23824 10100 23882 10146
rect 23882 10100 23886 10146
rect 23820 10094 23886 10100
rect -1991 9398 -1869 9455
rect 136 9399 203 9460
rect 1788 9630 1868 9636
rect 1788 9576 1792 9630
rect 1792 9576 1864 9630
rect 1864 9576 1868 9630
rect 1860 8690 1930 8693
rect 1860 8635 1866 8690
rect 1866 8635 1926 8690
rect 1926 8635 1930 8690
rect 1860 8631 1930 8635
rect 2944 8689 3015 8693
rect 2944 8634 2951 8689
rect 2951 8634 3011 8689
rect 3011 8634 3015 8689
rect 2944 8630 3015 8634
rect 1630 8559 1689 8573
rect 1630 8525 1642 8559
rect 1642 8525 1676 8559
rect 1676 8525 1689 8559
rect 1630 8513 1689 8525
rect 1980 8405 2048 8410
rect 1980 8350 1984 8405
rect 1984 8350 2044 8405
rect 2044 8350 2048 8405
rect 1980 8345 2048 8350
rect 3202 8690 3259 8694
rect 3202 8630 3206 8690
rect 3206 8630 3255 8690
rect 3255 8630 3259 8690
rect 3202 8626 3259 8630
rect 4932 9630 5012 9636
rect 4932 9576 4936 9630
rect 4936 9576 5008 9630
rect 5008 9576 5012 9630
rect 3202 8574 3259 8578
rect 3202 8514 3206 8574
rect 3206 8514 3255 8574
rect 3255 8514 3259 8574
rect 3202 8510 3259 8514
rect 5004 8690 5074 8693
rect 5004 8635 5010 8690
rect 5010 8635 5070 8690
rect 5070 8635 5074 8690
rect 5004 8631 5074 8635
rect 6088 8689 6159 8693
rect 6088 8634 6095 8689
rect 6095 8634 6155 8689
rect 6155 8634 6159 8689
rect 6088 8630 6159 8634
rect 4774 8559 4833 8573
rect 4774 8525 4786 8559
rect 4786 8525 4820 8559
rect 4820 8525 4833 8559
rect 4774 8513 4833 8525
rect 3202 8406 3259 8410
rect 3202 8346 3206 8406
rect 3206 8346 3255 8406
rect 3255 8346 3259 8406
rect 3202 8342 3259 8346
rect 1788 7372 1792 7418
rect 1792 7372 1850 7418
rect 1850 7372 1854 7418
rect 1788 7366 1854 7372
rect 5124 8405 5192 8410
rect 5124 8350 5128 8405
rect 5128 8350 5188 8405
rect 5188 8350 5192 8405
rect 5124 8345 5192 8350
rect 6346 8690 6403 8694
rect 6346 8630 6350 8690
rect 6350 8630 6399 8690
rect 6399 8630 6403 8690
rect 6346 8626 6403 8630
rect 8064 9626 8144 9632
rect 8064 9572 8068 9626
rect 8068 9572 8140 9626
rect 8140 9572 8144 9626
rect 11208 9626 11288 9632
rect 11208 9572 11212 9626
rect 11212 9572 11284 9626
rect 11284 9572 11288 9626
rect 6346 8574 6403 8578
rect 6346 8514 6350 8574
rect 6350 8514 6399 8574
rect 6399 8514 6403 8574
rect 6346 8510 6403 8514
rect 8136 8686 8206 8689
rect 8136 8631 8142 8686
rect 8142 8631 8202 8686
rect 8202 8631 8206 8686
rect 8136 8627 8206 8631
rect 9220 8685 9291 8689
rect 9220 8630 9227 8685
rect 9227 8630 9287 8685
rect 9287 8630 9291 8685
rect 9220 8626 9291 8630
rect 7906 8555 7965 8569
rect 7906 8521 7918 8555
rect 7918 8521 7952 8555
rect 7952 8521 7965 8555
rect 7906 8509 7965 8521
rect 6346 8406 6403 8410
rect 6346 8346 6350 8406
rect 6350 8346 6399 8406
rect 6399 8346 6403 8406
rect 6346 8342 6403 8346
rect 4932 7372 4936 7418
rect 4936 7372 4994 7418
rect 4994 7372 4998 7418
rect 4932 7366 4998 7372
rect 8256 8401 8324 8406
rect 8256 8346 8260 8401
rect 8260 8346 8320 8401
rect 8320 8346 8324 8401
rect 8256 8341 8324 8346
rect 9478 8686 9535 8690
rect 9478 8626 9482 8686
rect 9482 8626 9531 8686
rect 9531 8626 9535 8686
rect 9478 8622 9535 8626
rect 9478 8570 9535 8574
rect 9478 8510 9482 8570
rect 9482 8510 9531 8570
rect 9531 8510 9535 8570
rect 9478 8506 9535 8510
rect 9478 8402 9535 8406
rect 9478 8342 9482 8402
rect 9482 8342 9531 8402
rect 9531 8342 9535 8402
rect 9478 8338 9535 8342
rect 8064 7368 8068 7414
rect 8068 7368 8126 7414
rect 8126 7368 8130 7414
rect 8064 7362 8130 7368
rect 11280 8686 11350 8689
rect 11280 8631 11286 8686
rect 11286 8631 11346 8686
rect 11346 8631 11350 8686
rect 11280 8627 11350 8631
rect 12364 8685 12435 8689
rect 12364 8630 12371 8685
rect 12371 8630 12431 8685
rect 12431 8630 12435 8685
rect 12364 8626 12435 8630
rect 11050 8555 11109 8569
rect 11050 8521 11062 8555
rect 11062 8521 11096 8555
rect 11096 8521 11109 8555
rect 11050 8509 11109 8521
rect 11400 8401 11468 8406
rect 11400 8346 11404 8401
rect 11404 8346 11464 8401
rect 11464 8346 11468 8401
rect 11400 8341 11468 8346
rect 12622 8686 12679 8690
rect 12622 8626 12626 8686
rect 12626 8626 12675 8686
rect 12675 8626 12679 8686
rect 12622 8622 12679 8626
rect 14410 9630 14490 9636
rect 14410 9576 14414 9630
rect 14414 9576 14486 9630
rect 14486 9576 14490 9630
rect 12622 8570 12679 8574
rect 12622 8510 12626 8570
rect 12626 8510 12675 8570
rect 12675 8510 12679 8570
rect 12622 8506 12679 8510
rect 14482 8690 14552 8693
rect 14482 8635 14488 8690
rect 14488 8635 14548 8690
rect 14548 8635 14552 8690
rect 14482 8631 14552 8635
rect 15566 8689 15637 8693
rect 15566 8634 15573 8689
rect 15573 8634 15633 8689
rect 15633 8634 15637 8689
rect 15566 8630 15637 8634
rect 14252 8559 14311 8573
rect 14252 8525 14264 8559
rect 14264 8525 14298 8559
rect 14298 8525 14311 8559
rect 14252 8513 14311 8525
rect 12622 8402 12679 8406
rect 12622 8342 12626 8402
rect 12626 8342 12675 8402
rect 12675 8342 12679 8402
rect 12622 8338 12679 8342
rect 11208 7368 11212 7414
rect 11212 7368 11270 7414
rect 11270 7368 11274 7414
rect 11208 7362 11274 7368
rect 14602 8405 14670 8410
rect 14602 8350 14606 8405
rect 14606 8350 14666 8405
rect 14666 8350 14670 8405
rect 14602 8345 14670 8350
rect 15824 8690 15881 8694
rect 15824 8630 15828 8690
rect 15828 8630 15877 8690
rect 15877 8630 15881 8690
rect 15824 8626 15881 8630
rect 25837 11029 25904 11099
rect 17554 9630 17634 9636
rect 17554 9576 17558 9630
rect 17558 9576 17630 9630
rect 17630 9576 17634 9630
rect 15824 8574 15881 8578
rect 15824 8514 15828 8574
rect 15828 8514 15877 8574
rect 15877 8514 15881 8574
rect 15824 8510 15881 8514
rect 17626 8690 17696 8693
rect 17626 8635 17632 8690
rect 17632 8635 17692 8690
rect 17692 8635 17696 8690
rect 17626 8631 17696 8635
rect 18710 8689 18781 8693
rect 18710 8634 18717 8689
rect 18717 8634 18777 8689
rect 18777 8634 18781 8689
rect 18710 8630 18781 8634
rect 17396 8559 17455 8573
rect 17396 8525 17408 8559
rect 17408 8525 17442 8559
rect 17442 8525 17455 8559
rect 17396 8513 17455 8525
rect 15824 8406 15881 8410
rect 15824 8346 15828 8406
rect 15828 8346 15877 8406
rect 15877 8346 15881 8406
rect 15824 8342 15881 8346
rect 14410 7372 14414 7418
rect 14414 7372 14472 7418
rect 14472 7372 14476 7418
rect 14410 7366 14476 7372
rect 3283 6731 3359 6751
rect 3283 6695 3359 6731
rect 3283 6677 3359 6695
rect 17746 8405 17814 8410
rect 17746 8350 17750 8405
rect 17750 8350 17810 8405
rect 17810 8350 17814 8405
rect 17746 8345 17814 8350
rect 18968 8690 19025 8694
rect 18968 8630 18972 8690
rect 18972 8630 19021 8690
rect 19021 8630 19025 8690
rect 18968 8626 19025 8630
rect 20686 9626 20766 9632
rect 20686 9572 20690 9626
rect 20690 9572 20762 9626
rect 20762 9572 20766 9626
rect 18968 8574 19025 8578
rect 18968 8514 18972 8574
rect 18972 8514 19021 8574
rect 19021 8514 19025 8574
rect 18968 8510 19025 8514
rect 20758 8686 20828 8689
rect 20758 8631 20764 8686
rect 20764 8631 20824 8686
rect 20824 8631 20828 8686
rect 20758 8627 20828 8631
rect 21842 8685 21913 8689
rect 21842 8630 21849 8685
rect 21849 8630 21909 8685
rect 21909 8630 21913 8685
rect 21842 8626 21913 8630
rect 20528 8555 20587 8569
rect 20528 8521 20540 8555
rect 20540 8521 20574 8555
rect 20574 8521 20587 8555
rect 20528 8509 20587 8521
rect 18968 8406 19025 8410
rect 18968 8346 18972 8406
rect 18972 8346 19021 8406
rect 19021 8346 19025 8406
rect 18968 8342 19025 8346
rect 17554 7372 17558 7418
rect 17558 7372 17616 7418
rect 17616 7372 17620 7418
rect 17554 7366 17620 7372
rect 4021 6731 4097 6751
rect 4021 6695 4097 6731
rect 4021 6677 4097 6695
rect 20878 8401 20946 8406
rect 20878 8346 20882 8401
rect 20882 8346 20942 8401
rect 20942 8346 20946 8401
rect 20878 8341 20946 8346
rect 22100 8686 22157 8690
rect 22100 8626 22104 8686
rect 22104 8626 22153 8686
rect 22153 8626 22157 8686
rect 22100 8622 22157 8626
rect 23830 9626 23910 9632
rect 23830 9572 23834 9626
rect 23834 9572 23906 9626
rect 23906 9572 23910 9626
rect 22100 8570 22157 8574
rect 22100 8510 22104 8570
rect 22104 8510 22153 8570
rect 22153 8510 22157 8570
rect 22100 8506 22157 8510
rect 23902 8686 23972 8689
rect 23902 8631 23908 8686
rect 23908 8631 23968 8686
rect 23968 8631 23972 8686
rect 23902 8627 23972 8631
rect 24986 8685 25057 8689
rect 24986 8630 24993 8685
rect 24993 8630 25053 8685
rect 25053 8630 25057 8685
rect 24986 8626 25057 8630
rect 23672 8555 23731 8569
rect 23672 8521 23684 8555
rect 23684 8521 23718 8555
rect 23718 8521 23731 8555
rect 23672 8509 23731 8521
rect 22100 8402 22157 8406
rect 22100 8342 22104 8402
rect 22104 8342 22153 8402
rect 22153 8342 22157 8402
rect 22100 8338 22157 8342
rect 20686 7368 20690 7414
rect 20690 7368 20748 7414
rect 20748 7368 20752 7414
rect 20686 7362 20752 7368
rect 4759 6731 4835 6751
rect 4759 6695 4835 6731
rect 4759 6677 4835 6695
rect 5497 6731 5573 6751
rect 5497 6695 5573 6731
rect 5497 6677 5573 6695
rect 24022 8401 24090 8406
rect 24022 8346 24026 8401
rect 24026 8346 24086 8401
rect 24086 8346 24090 8401
rect 24022 8341 24090 8346
rect 25244 8686 25301 8690
rect 25244 8626 25248 8686
rect 25248 8626 25297 8686
rect 25297 8626 25301 8686
rect 25244 8622 25301 8626
rect 25244 8570 25301 8574
rect 25244 8510 25248 8570
rect 25248 8510 25297 8570
rect 25297 8510 25301 8570
rect 25244 8506 25301 8510
rect 25244 8402 25301 8406
rect 25244 8342 25248 8402
rect 25248 8342 25297 8402
rect 25297 8342 25301 8402
rect 25244 8338 25301 8342
rect 23830 7368 23834 7414
rect 23834 7368 23892 7414
rect 23892 7368 23896 7414
rect 23830 7362 23896 7368
rect 6237 6731 6313 6751
rect 6237 6695 6313 6731
rect 6237 6677 6313 6695
rect 6979 6731 7055 6751
rect 6979 6695 7055 6731
rect 6979 6677 7055 6695
rect 7717 6731 7793 6751
rect 7717 6695 7793 6731
rect 7717 6677 7793 6695
rect 8455 6733 8531 6753
rect 8455 6697 8531 6733
rect 8455 6679 8531 6697
rect 10061 6690 10115 6698
rect 10061 6652 10067 6690
rect 10067 6652 10105 6690
rect 10105 6652 10115 6690
rect 10061 6644 10115 6652
rect 12129 6688 12183 6696
rect 12129 6650 12135 6688
rect 12135 6650 12173 6688
rect 12173 6650 12183 6688
rect 14198 6690 14252 6698
rect 12129 6642 12183 6650
rect 14198 6652 14204 6690
rect 14204 6652 14242 6690
rect 14242 6652 14252 6690
rect 14198 6644 14252 6652
rect 16266 6688 16320 6696
rect 16266 6650 16272 6688
rect 16272 6650 16310 6688
rect 16310 6650 16320 6688
rect 18335 6688 18389 6696
rect 16266 6642 16320 6650
rect 18335 6650 18341 6688
rect 18341 6650 18379 6688
rect 18379 6650 18389 6688
rect 18335 6642 18389 6650
rect 20403 6686 20457 6694
rect 20403 6648 20409 6686
rect 20409 6648 20447 6686
rect 20447 6648 20457 6686
rect 22472 6688 22526 6696
rect 20403 6640 20457 6648
rect 3333 5863 3435 5869
rect 3333 5809 3345 5863
rect 3345 5809 3423 5863
rect 3423 5809 3435 5863
rect 3333 5803 3435 5809
rect 4071 5863 4173 5869
rect 4071 5809 4083 5863
rect 4083 5809 4161 5863
rect 4161 5809 4173 5863
rect 4071 5803 4173 5809
rect 4809 5863 4911 5869
rect 4809 5809 4821 5863
rect 4821 5809 4899 5863
rect 4899 5809 4911 5863
rect 4809 5803 4911 5809
rect 5547 5863 5649 5869
rect 5547 5809 5559 5863
rect 5559 5809 5637 5863
rect 5637 5809 5649 5863
rect 5547 5803 5649 5809
rect 6287 5863 6389 5869
rect 6287 5809 6299 5863
rect 6299 5809 6377 5863
rect 6377 5809 6389 5863
rect 6287 5803 6389 5809
rect 7029 5863 7131 5869
rect 7029 5809 7041 5863
rect 7041 5809 7119 5863
rect 7119 5809 7131 5863
rect 7029 5803 7131 5809
rect 7767 5863 7869 5869
rect 7767 5809 7779 5863
rect 7779 5809 7857 5863
rect 7857 5809 7869 5863
rect 7767 5803 7869 5809
rect 8505 5865 8607 5871
rect 8505 5811 8517 5865
rect 8517 5811 8595 5865
rect 8595 5811 8607 5865
rect 8505 5805 8607 5811
rect 9481 5836 9535 5890
rect 22472 6650 22478 6688
rect 22478 6650 22516 6688
rect 22516 6650 22526 6688
rect 22472 6642 22526 6650
rect 24540 6686 24594 6694
rect 24540 6648 24546 6686
rect 24546 6648 24584 6686
rect 24584 6648 24594 6686
rect 24540 6640 24594 6648
rect 10857 5830 10923 5896
rect 483 4566 563 4635
rect 257 4405 352 4483
rect 3 4213 84 4287
rect -1993 3398 -1872 3408
rect -1993 3361 -1976 3398
rect -1976 3361 -1883 3398
rect -1883 3361 -1872 3398
rect -1993 3349 -1872 3361
rect -1520 3158 -1404 3173
rect -1520 3122 -1506 3158
rect -1506 3122 -1414 3158
rect -1414 3122 -1404 3158
rect -1520 3110 -1404 3122
rect -1258 3044 -1137 3060
rect -1258 3001 -1246 3044
rect -1246 3001 -1166 3044
rect -1166 3001 -1137 3044
rect -1258 2993 -1137 3001
rect -1049 2933 -925 2945
rect -1049 2876 -1030 2933
rect -1030 2876 -952 2933
rect -952 2876 -925 2933
rect -1049 2863 -925 2876
rect 10111 4468 10173 4474
rect 10111 4426 10117 4468
rect 10117 4426 10167 4468
rect 10167 4426 10173 4468
rect 10111 4416 10173 4426
rect -550 -479 -446 -317
rect 11549 5834 11603 5888
rect 12925 5828 12991 5894
rect 12179 4466 12241 4472
rect 12179 4424 12185 4466
rect 12185 4424 12235 4466
rect 12235 4424 12241 4466
rect 12179 4414 12241 4424
rect 13618 5836 13672 5890
rect 14994 5830 15060 5896
rect 14248 4468 14310 4474
rect 14248 4426 14254 4468
rect 14254 4426 14304 4468
rect 14304 4426 14310 4468
rect 14248 4416 14310 4426
rect 15686 5834 15740 5888
rect 17062 5828 17128 5894
rect 16316 4466 16378 4472
rect 16316 4424 16322 4466
rect 16322 4424 16372 4466
rect 16372 4424 16378 4466
rect 16316 4414 16378 4424
rect 17755 5834 17809 5888
rect 19131 5828 19197 5894
rect 18385 4466 18447 4472
rect 18385 4424 18391 4466
rect 18391 4424 18441 4466
rect 18441 4424 18447 4466
rect 18385 4414 18447 4424
rect 19823 5832 19877 5886
rect 21199 5826 21265 5892
rect 20453 4464 20515 4470
rect 20453 4422 20459 4464
rect 20459 4422 20509 4464
rect 20509 4422 20515 4464
rect 20453 4412 20515 4422
rect 21892 5834 21946 5888
rect 23268 5828 23334 5894
rect 22522 4466 22584 4472
rect 22522 4424 22528 4466
rect 22528 4424 22578 4466
rect 22578 4424 22584 4466
rect 22522 4414 22584 4424
rect 23960 5832 24014 5886
rect 27829 18374 27889 18436
rect 27836 18184 27896 18246
rect 28564 18177 28616 18252
rect 27836 17995 27896 18064
rect 28461 17987 28515 18064
rect 27848 17814 27909 17877
rect 28360 17806 28414 17876
rect 27851 17614 27922 17686
rect 28258 17600 28311 17675
rect 27851 17154 27905 17209
rect 28157 17152 28211 17216
rect 27801 16747 27857 16801
rect 28052 16731 28118 16807
rect 30505 13083 30571 13149
rect 30701 13097 30761 13161
rect 30761 13097 30762 13161
rect 29703 12331 29757 12341
rect 29703 12293 29711 12331
rect 29711 12293 29749 12331
rect 29749 12293 29757 12331
rect 29703 12287 29757 12293
rect 31927 12393 31985 12399
rect 31927 12343 31933 12393
rect 31933 12343 31975 12393
rect 31975 12343 31985 12393
rect 31927 12337 31985 12343
rect 30511 11707 30565 11761
rect 31074 11441 31153 11518
rect 30503 11015 30569 11081
rect 30699 11028 30759 11090
rect 29701 10263 29755 10273
rect 29701 10225 29709 10263
rect 29709 10225 29747 10263
rect 29747 10225 29755 10263
rect 29701 10219 29755 10225
rect 31925 10325 31983 10331
rect 31925 10275 31931 10325
rect 31931 10275 31973 10325
rect 31973 10275 31983 10325
rect 31925 10269 31983 10275
rect 30509 9639 30563 9693
rect 31077 9375 31148 9449
rect 30505 8946 30571 9012
rect 30702 8961 30761 9021
rect 30761 8961 30762 9021
rect 29703 8194 29757 8204
rect 29703 8156 29711 8194
rect 29711 8156 29749 8194
rect 29749 8156 29757 8194
rect 29703 8150 29757 8156
rect 31927 8256 31985 8262
rect 31927 8206 31933 8256
rect 31933 8206 31975 8256
rect 31975 8206 31985 8256
rect 31927 8200 31985 8206
rect 30511 7570 30565 7624
rect 31084 7307 31147 7372
rect 32549 9228 32615 9302
rect 27321 7099 27389 7157
rect 32416 7143 32478 7207
rect 27074 6806 27130 6863
rect 26851 6502 26912 6555
rect 26667 6340 26737 6398
rect 26467 6190 26535 6248
rect 26281 6031 26339 6085
rect 25336 5826 25402 5892
rect 25628 5832 25688 5885
rect 26047 5841 26111 5901
rect 25346 5696 25417 5704
rect 25346 5636 25348 5696
rect 25348 5636 25414 5696
rect 25414 5636 25417 5696
rect 25346 5627 25417 5636
rect 25636 5635 25688 5693
rect 24590 4464 24652 4470
rect 24590 4422 24596 4464
rect 24596 4422 24646 4464
rect 24646 4422 24652 4464
rect 24590 4412 24652 4422
rect 142 3398 221 3411
rect 142 3354 151 3398
rect 151 3354 205 3398
rect 205 3354 221 3398
rect 142 3348 221 3354
rect 30503 6878 30569 6944
rect 30701 6892 30756 6953
rect 29701 6126 29755 6136
rect 29701 6088 29709 6126
rect 29709 6088 29747 6126
rect 29747 6088 29755 6126
rect 29701 6082 29755 6088
rect 31925 6188 31983 6194
rect 31925 6138 31931 6188
rect 31931 6138 31973 6188
rect 31973 6138 31983 6188
rect 31925 6132 31983 6138
rect 30509 5502 30563 5556
rect 31076 5240 31149 5304
rect 30503 4809 30569 4875
rect 30700 4823 30756 4884
rect 29701 4057 29755 4067
rect 29701 4019 29709 4057
rect 29709 4019 29747 4057
rect 29747 4019 29755 4057
rect 29701 4013 29755 4019
rect 31925 4119 31983 4125
rect 31925 4069 31931 4119
rect 31931 4069 31973 4119
rect 31973 4069 31983 4119
rect 31925 4063 31983 4069
rect 30509 3433 30563 3487
rect 138 3150 217 3161
rect 138 3106 150 3150
rect 150 3106 204 3150
rect 204 3106 217 3150
rect 138 3098 217 3106
rect 136 3034 215 3048
rect 136 2990 149 3034
rect 149 2990 203 3034
rect 203 2990 215 3034
rect 136 2985 215 2990
rect 134 2910 211 2921
rect 134 2866 149 2910
rect 149 2866 203 2910
rect 203 2866 211 2910
rect 134 2860 211 2866
rect 1508 2378 1588 2384
rect 1508 2324 1512 2378
rect 1512 2324 1584 2378
rect 1584 2324 1588 2378
rect 117 1438 174 1442
rect 117 1378 121 1438
rect 121 1378 170 1438
rect 170 1378 174 1438
rect 117 1374 174 1378
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 121 1262 170 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 361 1437 432 1441
rect 361 1382 365 1437
rect 365 1382 425 1437
rect 425 1382 432 1437
rect 361 1378 432 1382
rect 1446 1438 1516 1441
rect 1446 1383 1450 1438
rect 1450 1383 1510 1438
rect 1510 1383 1516 1438
rect 1446 1379 1516 1383
rect 1687 1307 1746 1321
rect 1687 1273 1700 1307
rect 1700 1273 1734 1307
rect 1734 1273 1746 1307
rect 1687 1261 1746 1273
rect 1328 1153 1396 1158
rect 1328 1098 1332 1153
rect 1332 1098 1392 1153
rect 1392 1098 1396 1153
rect 1328 1093 1396 1098
rect 4652 2378 4732 2384
rect 4652 2324 4656 2378
rect 4656 2324 4728 2378
rect 4728 2324 4732 2378
rect 3261 1438 3318 1442
rect 3261 1378 3265 1438
rect 3265 1378 3314 1438
rect 3314 1378 3318 1438
rect 3261 1374 3318 1378
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3265 1262 3314 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 1522 120 1526 166
rect 1526 120 1584 166
rect 1584 120 1588 166
rect 1522 114 1588 120
rect -285 -317 -181 -155
rect -792 -766 -688 -604
rect 3505 1437 3576 1441
rect 3505 1382 3509 1437
rect 3509 1382 3569 1437
rect 3569 1382 3576 1437
rect 3505 1378 3576 1382
rect 4590 1438 4660 1441
rect 4590 1383 4594 1438
rect 4594 1383 4654 1438
rect 4654 1383 4660 1438
rect 4590 1379 4660 1383
rect 4831 1307 4890 1321
rect 4831 1273 4844 1307
rect 4844 1273 4878 1307
rect 4878 1273 4890 1307
rect 4831 1261 4890 1273
rect 4472 1153 4540 1158
rect 4472 1098 4476 1153
rect 4476 1098 4536 1153
rect 4536 1098 4540 1153
rect 4472 1093 4540 1098
rect 7784 2382 7864 2388
rect 7784 2328 7788 2382
rect 7788 2328 7860 2382
rect 7860 2328 7864 2382
rect 6393 1442 6450 1446
rect 6393 1382 6397 1442
rect 6397 1382 6446 1442
rect 6446 1382 6450 1442
rect 6393 1378 6450 1382
rect 6393 1326 6450 1330
rect 6393 1266 6397 1326
rect 6397 1266 6446 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 6637 1441 6708 1445
rect 6637 1386 6641 1441
rect 6641 1386 6701 1441
rect 6701 1386 6708 1441
rect 6637 1382 6708 1386
rect 7722 1442 7792 1445
rect 7722 1387 7726 1442
rect 7726 1387 7786 1442
rect 7786 1387 7792 1442
rect 7722 1383 7792 1387
rect 7963 1311 8022 1325
rect 7963 1277 7976 1311
rect 7976 1277 8010 1311
rect 8010 1277 8022 1311
rect 7963 1265 8022 1277
rect 7604 1157 7672 1162
rect 7604 1102 7608 1157
rect 7608 1102 7668 1157
rect 7668 1102 7672 1157
rect 7604 1097 7672 1102
rect 10928 2382 11008 2388
rect 10928 2328 10932 2382
rect 10932 2328 11004 2382
rect 11004 2328 11008 2382
rect 9537 1442 9594 1446
rect 9537 1382 9541 1442
rect 9541 1382 9590 1442
rect 9590 1382 9594 1442
rect 9537 1378 9594 1382
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9541 1266 9590 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 4666 120 4670 166
rect 4670 120 4728 166
rect 4728 120 4732 166
rect 4666 114 4732 120
rect 7798 124 7802 170
rect 7802 124 7860 170
rect 7860 124 7864 170
rect 7798 118 7864 124
rect 9781 1441 9852 1445
rect 9781 1386 9785 1441
rect 9785 1386 9845 1441
rect 9845 1386 9852 1441
rect 9781 1382 9852 1386
rect 10866 1442 10936 1445
rect 10866 1387 10870 1442
rect 10870 1387 10930 1442
rect 10930 1387 10936 1442
rect 10866 1383 10936 1387
rect 11107 1311 11166 1325
rect 11107 1277 11120 1311
rect 11120 1277 11154 1311
rect 11154 1277 11166 1311
rect 11107 1265 11166 1277
rect 10748 1157 10816 1162
rect 10748 1102 10752 1157
rect 10752 1102 10812 1157
rect 10812 1102 10816 1157
rect 10748 1097 10816 1102
rect 14130 2378 14210 2384
rect 14130 2324 14134 2378
rect 14134 2324 14206 2378
rect 14206 2324 14210 2378
rect 12739 1438 12796 1442
rect 12739 1378 12743 1438
rect 12743 1378 12792 1438
rect 12792 1378 12796 1438
rect 12739 1374 12796 1378
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12743 1262 12792 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 10942 124 10946 170
rect 10946 124 11004 170
rect 11004 124 11008 170
rect 10942 118 11008 124
rect 12983 1437 13054 1441
rect 12983 1382 12987 1437
rect 12987 1382 13047 1437
rect 13047 1382 13054 1437
rect 12983 1378 13054 1382
rect 14068 1438 14138 1441
rect 14068 1383 14072 1438
rect 14072 1383 14132 1438
rect 14132 1383 14138 1438
rect 14068 1379 14138 1383
rect 14309 1307 14368 1321
rect 14309 1273 14322 1307
rect 14322 1273 14356 1307
rect 14356 1273 14368 1307
rect 14309 1261 14368 1273
rect 17274 2378 17354 2384
rect 17274 2324 17278 2378
rect 17278 2324 17350 2378
rect 17350 2324 17354 2378
rect 15883 1438 15940 1442
rect 15883 1378 15887 1438
rect 15887 1378 15936 1438
rect 15936 1378 15940 1438
rect 15883 1374 15940 1378
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15887 1262 15936 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 13950 1153 14018 1158
rect 13950 1098 13954 1153
rect 13954 1098 14014 1153
rect 14014 1098 14018 1153
rect 13950 1093 14018 1098
rect 14144 120 14148 166
rect 14148 120 14206 166
rect 14206 120 14210 166
rect 14144 114 14210 120
rect 1540 -1514 1620 -1508
rect 1540 -1568 1544 -1514
rect 1544 -1568 1616 -1514
rect 1616 -1568 1620 -1514
rect 149 -2454 206 -2450
rect 149 -2514 153 -2454
rect 153 -2514 202 -2454
rect 202 -2514 206 -2454
rect 149 -2518 206 -2514
rect 149 -2634 206 -2566
rect 393 -2455 464 -2451
rect 393 -2510 397 -2455
rect 397 -2510 457 -2455
rect 457 -2510 464 -2455
rect 393 -2514 464 -2510
rect 1478 -2454 1548 -2451
rect 1478 -2509 1482 -2454
rect 1482 -2509 1542 -2454
rect 1542 -2509 1548 -2454
rect 1478 -2513 1548 -2509
rect 1719 -2585 1778 -2571
rect 1719 -2619 1732 -2585
rect 1732 -2619 1766 -2585
rect 1766 -2619 1778 -2585
rect 1719 -2631 1778 -2619
rect 1360 -2739 1428 -2734
rect 1360 -2794 1364 -2739
rect 1364 -2794 1424 -2739
rect 1424 -2794 1428 -2739
rect 1360 -2799 1428 -2794
rect 4684 -1514 4764 -1508
rect 4684 -1568 4688 -1514
rect 4688 -1568 4760 -1514
rect 4760 -1568 4764 -1514
rect 3293 -2454 3350 -2450
rect 3293 -2514 3297 -2454
rect 3297 -2514 3346 -2454
rect 3346 -2514 3350 -2454
rect 3293 -2518 3350 -2514
rect 3293 -2634 3350 -2566
rect 1554 -3772 1558 -3726
rect 1558 -3772 1616 -3726
rect 1616 -3772 1620 -3726
rect 1554 -3778 1620 -3772
rect 3537 -2455 3608 -2451
rect 3537 -2510 3541 -2455
rect 3541 -2510 3601 -2455
rect 3601 -2510 3608 -2455
rect 3537 -2514 3608 -2510
rect 4622 -2454 4692 -2451
rect 4622 -2509 4626 -2454
rect 4626 -2509 4686 -2454
rect 4686 -2509 4692 -2454
rect 4622 -2513 4692 -2509
rect 4863 -2585 4922 -2571
rect 4863 -2619 4876 -2585
rect 4876 -2619 4910 -2585
rect 4910 -2619 4922 -2585
rect 4863 -2631 4922 -2619
rect 7816 -1510 7896 -1504
rect 7816 -1564 7820 -1510
rect 7820 -1564 7892 -1510
rect 7892 -1564 7896 -1510
rect 6425 -2450 6482 -2446
rect 6425 -2510 6429 -2450
rect 6429 -2510 6478 -2450
rect 6478 -2510 6482 -2450
rect 6425 -2514 6482 -2510
rect 4504 -2739 4572 -2734
rect 4504 -2794 4508 -2739
rect 4508 -2794 4568 -2739
rect 4568 -2794 4572 -2739
rect 4504 -2799 4572 -2794
rect 6425 -2630 6482 -2562
rect 6669 -2451 6740 -2447
rect 6669 -2506 6673 -2451
rect 6673 -2506 6733 -2451
rect 6733 -2506 6740 -2451
rect 6669 -2510 6740 -2506
rect 7754 -2450 7824 -2447
rect 7754 -2505 7758 -2450
rect 7758 -2505 7818 -2450
rect 7818 -2505 7824 -2450
rect 7754 -2509 7824 -2505
rect 7995 -2581 8054 -2567
rect 7995 -2615 8008 -2581
rect 8008 -2615 8042 -2581
rect 8042 -2615 8054 -2581
rect 7995 -2627 8054 -2615
rect 16127 1437 16198 1441
rect 16127 1382 16131 1437
rect 16131 1382 16191 1437
rect 16191 1382 16198 1437
rect 16127 1378 16198 1382
rect 17212 1438 17282 1441
rect 17212 1383 17216 1438
rect 17216 1383 17276 1438
rect 17276 1383 17282 1438
rect 17212 1379 17282 1383
rect 17453 1307 17512 1321
rect 17453 1273 17466 1307
rect 17466 1273 17500 1307
rect 17500 1273 17512 1307
rect 17453 1261 17512 1273
rect 17094 1153 17162 1158
rect 17094 1098 17098 1153
rect 17098 1098 17158 1153
rect 17158 1098 17162 1153
rect 17094 1093 17162 1098
rect 20406 2382 20486 2388
rect 20406 2328 20410 2382
rect 20410 2328 20482 2382
rect 20482 2328 20486 2382
rect 19015 1442 19072 1446
rect 19015 1382 19019 1442
rect 19019 1382 19068 1442
rect 19068 1382 19072 1442
rect 19015 1378 19072 1382
rect 19015 1326 19072 1330
rect 19015 1266 19019 1326
rect 19019 1266 19068 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 19259 1441 19330 1445
rect 19259 1386 19263 1441
rect 19263 1386 19323 1441
rect 19323 1386 19330 1441
rect 19259 1382 19330 1386
rect 20344 1442 20414 1445
rect 20344 1387 20348 1442
rect 20348 1387 20408 1442
rect 20408 1387 20414 1442
rect 20344 1383 20414 1387
rect 20585 1311 20644 1325
rect 20585 1277 20598 1311
rect 20598 1277 20632 1311
rect 20632 1277 20644 1311
rect 20585 1265 20644 1277
rect 20226 1157 20294 1162
rect 20226 1102 20230 1157
rect 20230 1102 20290 1157
rect 20290 1102 20294 1157
rect 20226 1097 20294 1102
rect 23550 2382 23630 2388
rect 23550 2328 23554 2382
rect 23554 2328 23626 2382
rect 23626 2328 23630 2382
rect 22159 1442 22216 1446
rect 22159 1382 22163 1442
rect 22163 1382 22212 1442
rect 22212 1382 22216 1442
rect 22159 1378 22216 1382
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22163 1266 22212 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 17288 120 17292 166
rect 17292 120 17350 166
rect 17350 120 17354 166
rect 17288 114 17354 120
rect 10960 -1510 11040 -1504
rect 10960 -1564 10964 -1510
rect 10964 -1564 11036 -1510
rect 11036 -1564 11040 -1510
rect 9569 -2450 9626 -2446
rect 9569 -2510 9573 -2450
rect 9573 -2510 9622 -2450
rect 9622 -2510 9626 -2450
rect 9569 -2514 9626 -2510
rect 7636 -2735 7704 -2730
rect 7636 -2790 7640 -2735
rect 7640 -2790 7700 -2735
rect 7700 -2790 7704 -2735
rect 7636 -2795 7704 -2790
rect 9569 -2630 9626 -2562
rect 4698 -3772 4702 -3726
rect 4702 -3772 4760 -3726
rect 4760 -3772 4764 -3726
rect 4698 -3778 4764 -3772
rect 9813 -2451 9884 -2447
rect 9813 -2506 9817 -2451
rect 9817 -2506 9877 -2451
rect 9877 -2506 9884 -2451
rect 9813 -2510 9884 -2506
rect 10898 -2450 10968 -2447
rect 10898 -2505 10902 -2450
rect 10902 -2505 10962 -2450
rect 10962 -2505 10968 -2450
rect 10898 -2509 10968 -2505
rect 11139 -2581 11198 -2567
rect 11139 -2615 11152 -2581
rect 11152 -2615 11186 -2581
rect 11186 -2615 11198 -2581
rect 11139 -2627 11198 -2615
rect 22403 1441 22474 1445
rect 22403 1386 22407 1441
rect 22407 1386 22467 1441
rect 22467 1386 22474 1441
rect 22403 1382 22474 1386
rect 23488 1442 23558 1445
rect 23488 1387 23492 1442
rect 23492 1387 23552 1442
rect 23552 1387 23558 1442
rect 23488 1383 23558 1387
rect 23729 1311 23788 1325
rect 23729 1277 23742 1311
rect 23742 1277 23776 1311
rect 23776 1277 23788 1311
rect 23729 1265 23788 1277
rect 23370 1157 23438 1162
rect 23370 1102 23374 1157
rect 23374 1102 23434 1157
rect 23434 1102 23438 1157
rect 23370 1097 23438 1102
rect 20420 124 20424 170
rect 20424 124 20482 170
rect 20482 124 20486 170
rect 20420 118 20486 124
rect 23564 124 23568 170
rect 23568 124 23626 170
rect 23626 124 23630 170
rect 23564 118 23630 124
rect 14162 -1514 14242 -1508
rect 14162 -1568 14166 -1514
rect 14166 -1568 14238 -1514
rect 14238 -1568 14242 -1514
rect 12771 -2454 12828 -2450
rect 12771 -2514 12775 -2454
rect 12775 -2514 12824 -2454
rect 12824 -2514 12828 -2454
rect 12771 -2518 12828 -2514
rect 10780 -2735 10848 -2730
rect 10780 -2790 10784 -2735
rect 10784 -2790 10844 -2735
rect 10844 -2790 10848 -2735
rect 10780 -2795 10848 -2790
rect 12771 -2634 12828 -2566
rect 7830 -3768 7834 -3722
rect 7834 -3768 7892 -3722
rect 7892 -3768 7896 -3722
rect 7830 -3774 7896 -3768
rect 10974 -3768 10978 -3722
rect 10978 -3768 11036 -3722
rect 11036 -3768 11040 -3722
rect 10974 -3774 11040 -3768
rect 13015 -2455 13086 -2451
rect 13015 -2510 13019 -2455
rect 13019 -2510 13079 -2455
rect 13079 -2510 13086 -2455
rect 13015 -2514 13086 -2510
rect 14100 -2454 14170 -2451
rect 14100 -2509 14104 -2454
rect 14104 -2509 14164 -2454
rect 14164 -2509 14170 -2454
rect 14100 -2513 14170 -2509
rect 14341 -2585 14400 -2571
rect 14341 -2619 14354 -2585
rect 14354 -2619 14388 -2585
rect 14388 -2619 14400 -2585
rect 14341 -2631 14400 -2619
rect 17306 -1514 17386 -1508
rect 17306 -1568 17310 -1514
rect 17310 -1568 17382 -1514
rect 17382 -1568 17386 -1514
rect 15915 -2454 15972 -2450
rect 15915 -2514 15919 -2454
rect 15919 -2514 15968 -2454
rect 15968 -2514 15972 -2454
rect 15915 -2518 15972 -2514
rect 13982 -2739 14050 -2734
rect 13982 -2794 13986 -2739
rect 13986 -2794 14046 -2739
rect 14046 -2794 14050 -2739
rect 13982 -2799 14050 -2794
rect 15915 -2634 15972 -2566
rect 14176 -3772 14180 -3726
rect 14180 -3772 14238 -3726
rect 14238 -3772 14242 -3726
rect 14176 -3778 14242 -3772
rect 16159 -2455 16230 -2451
rect 16159 -2510 16163 -2455
rect 16163 -2510 16223 -2455
rect 16223 -2510 16230 -2455
rect 16159 -2514 16230 -2510
rect 17244 -2454 17314 -2451
rect 17244 -2509 17248 -2454
rect 17248 -2509 17308 -2454
rect 17308 -2509 17314 -2454
rect 17244 -2513 17314 -2509
rect 17485 -2585 17544 -2571
rect 17485 -2619 17498 -2585
rect 17498 -2619 17532 -2585
rect 17532 -2619 17544 -2585
rect 17485 -2631 17544 -2619
rect 17126 -2739 17194 -2734
rect 17126 -2794 17130 -2739
rect 17130 -2794 17190 -2739
rect 17190 -2794 17194 -2739
rect 17126 -2799 17194 -2794
rect 20438 -1510 20518 -1504
rect 20438 -1564 20442 -1510
rect 20442 -1564 20514 -1510
rect 20514 -1564 20518 -1510
rect 19047 -2450 19104 -2446
rect 19047 -2510 19051 -2450
rect 19051 -2510 19100 -2450
rect 19100 -2510 19104 -2450
rect 19047 -2514 19104 -2510
rect 19047 -2630 19104 -2562
rect 19291 -2451 19362 -2447
rect 19291 -2506 19295 -2451
rect 19295 -2506 19355 -2451
rect 19355 -2506 19362 -2451
rect 19291 -2510 19362 -2506
rect 20376 -2450 20446 -2447
rect 20376 -2505 20380 -2450
rect 20380 -2505 20440 -2450
rect 20440 -2505 20446 -2450
rect 20376 -2509 20446 -2505
rect 20617 -2581 20676 -2567
rect 20617 -2615 20630 -2581
rect 20630 -2615 20664 -2581
rect 20664 -2615 20676 -2581
rect 20617 -2627 20676 -2615
rect 23582 -1510 23662 -1504
rect 23582 -1564 23586 -1510
rect 23586 -1564 23658 -1510
rect 23658 -1564 23662 -1510
rect 22191 -2450 22248 -2446
rect 22191 -2510 22195 -2450
rect 22195 -2510 22244 -2450
rect 22244 -2510 22248 -2450
rect 22191 -2514 22248 -2510
rect 22191 -2630 22248 -2562
rect 20258 -2735 20326 -2730
rect 20258 -2790 20262 -2735
rect 20262 -2790 20322 -2735
rect 20322 -2790 20326 -2735
rect 20258 -2795 20326 -2790
rect 17320 -3772 17324 -3726
rect 17324 -3772 17382 -3726
rect 17382 -3772 17386 -3726
rect 17320 -3778 17386 -3772
rect 20452 -3768 20456 -3722
rect 20456 -3768 20514 -3722
rect 20514 -3768 20518 -3722
rect 20452 -3774 20518 -3768
rect 22435 -2451 22506 -2447
rect 22435 -2506 22439 -2451
rect 22439 -2506 22499 -2451
rect 22499 -2506 22506 -2451
rect 22435 -2510 22506 -2506
rect 23520 -2450 23590 -2447
rect 23520 -2505 23524 -2450
rect 23524 -2505 23584 -2450
rect 23584 -2505 23590 -2450
rect 23520 -2509 23590 -2505
rect 23761 -2581 23820 -2567
rect 23761 -2615 23774 -2581
rect 23774 -2615 23808 -2581
rect 23808 -2615 23820 -2581
rect 23761 -2627 23820 -2615
rect 23402 -2735 23470 -2730
rect 23402 -2790 23406 -2735
rect 23406 -2790 23466 -2735
rect 23466 -2790 23470 -2735
rect 23402 -2795 23470 -2790
rect 23596 -3768 23600 -3722
rect 23600 -3768 23658 -3722
rect 23658 -3768 23662 -3722
rect 23596 -3774 23662 -3768
rect 31079 3172 31144 3238
rect 30501 2741 30567 2807
rect 30699 2755 30755 2817
rect 29699 1989 29753 1999
rect 29699 1951 29707 1989
rect 29707 1951 29745 1989
rect 29745 1951 29753 1989
rect 29699 1945 29753 1951
rect 31923 2051 31981 2057
rect 31923 2001 31929 2051
rect 31929 2001 31971 2051
rect 31971 2001 31981 2051
rect 31923 1995 31981 2001
rect 30507 1365 30561 1419
rect 31079 1101 31144 1171
rect 30503 672 30569 738
rect 30703 687 30755 747
rect 29701 -80 29755 -70
rect 29701 -118 29709 -80
rect 29709 -118 29747 -80
rect 29747 -118 29755 -80
rect 29701 -124 29755 -118
rect 31925 -18 31983 -12
rect 31925 -68 31931 -18
rect 31931 -68 31973 -18
rect 31973 -68 31983 -18
rect 31925 -74 31983 -68
rect 30509 -704 30563 -650
rect 31076 -968 31149 -898
rect 33107 13195 33168 13247
rect 41869 23365 42001 23473
rect 39307 23087 39419 23193
rect 40055 23061 40187 23169
rect 43616 23977 43681 24031
rect 49437 24772 49493 24786
rect 49437 24738 49453 24772
rect 49453 24738 49487 24772
rect 49487 24738 49493 24772
rect 49437 24720 49493 24738
rect 50183 24762 50315 24870
rect 48307 24648 48373 24664
rect 48307 24614 48323 24648
rect 48323 24614 48357 24648
rect 48357 24614 48373 24648
rect 48307 24598 48373 24614
rect 53088 24703 53220 24811
rect 55570 24757 55702 24865
rect 44711 23965 44779 24040
rect 43011 23363 43143 23471
rect 41868 22718 42000 22826
rect 43766 22718 43898 22826
rect 39590 21956 39708 22074
rect 40335 21998 40443 22130
rect 45190 23607 45426 23751
rect 48973 23951 49072 24048
rect 46834 23645 46942 23777
rect 39087 21614 39180 21693
rect 40050 21457 40182 21565
rect 42513 21840 42576 21856
rect 42513 21806 42542 21840
rect 42542 21806 42576 21840
rect 42513 21790 42576 21806
rect 45325 22059 45437 22061
rect 45325 21955 45443 22059
rect 45331 21953 45443 21955
rect 40637 20762 40700 20814
rect 40330 20394 40438 20526
rect 39592 20179 39704 20285
rect 41813 20322 41945 20430
rect 43711 20322 43843 20430
rect 48382 23362 48514 23470
rect 45820 23084 45932 23190
rect 46568 23058 46700 23166
rect 50129 23974 50194 24028
rect 55971 24767 56027 24781
rect 55971 24733 55987 24767
rect 55987 24733 56021 24767
rect 56021 24733 56027 24767
rect 55971 24715 56027 24733
rect 56717 24757 56849 24865
rect 54841 24643 54907 24659
rect 54841 24609 54857 24643
rect 54857 24609 54891 24643
rect 54891 24609 54907 24643
rect 54841 24593 54907 24609
rect 59646 24707 59778 24815
rect 62128 24761 62260 24869
rect 51224 23962 51292 24037
rect 49524 23360 49656 23468
rect 48381 22715 48513 22823
rect 50279 22715 50411 22823
rect 46103 21953 46221 22071
rect 46848 21995 46956 22127
rect 51727 23601 51960 23758
rect 55507 23946 55606 24043
rect 53368 23640 53476 23772
rect 45600 21611 45693 21690
rect 46563 21454 46695 21562
rect 49026 21837 49089 21853
rect 49026 21803 49055 21837
rect 49055 21803 49089 21837
rect 49026 21787 49089 21803
rect 51859 22054 51971 22056
rect 51859 21950 51977 22054
rect 51865 21948 51977 21950
rect 47150 20759 47213 20811
rect 46843 20391 46951 20523
rect 46105 20176 46217 20282
rect 48326 20319 48458 20427
rect 50224 20319 50356 20427
rect 54916 23357 55048 23465
rect 52354 23079 52466 23185
rect 53102 23053 53234 23161
rect 56663 23969 56728 24023
rect 62529 24771 62585 24785
rect 62529 24737 62545 24771
rect 62545 24737 62579 24771
rect 62579 24737 62585 24771
rect 62529 24719 62585 24737
rect 63275 24761 63407 24869
rect 61399 24647 61465 24663
rect 61399 24613 61415 24647
rect 61415 24613 61449 24647
rect 61449 24613 61465 24647
rect 61399 24597 61465 24613
rect 57758 23957 57826 24032
rect 56058 23355 56190 23463
rect 54915 22710 55047 22818
rect 56813 22710 56945 22818
rect 52637 21948 52755 22066
rect 53382 21990 53490 22122
rect 58287 23596 58534 23759
rect 62065 23950 62164 24047
rect 59926 23644 60034 23776
rect 52134 21606 52227 21685
rect 53097 21449 53229 21557
rect 55560 21832 55623 21848
rect 55560 21798 55589 21832
rect 55589 21798 55623 21832
rect 55560 21782 55623 21798
rect 58417 22058 58529 22060
rect 58417 21954 58535 22058
rect 58423 21952 58535 21954
rect 53684 20754 53747 20806
rect 53377 20386 53485 20518
rect 52639 20171 52751 20277
rect 54860 20314 54992 20422
rect 56758 20314 56890 20422
rect 61474 23361 61606 23469
rect 58912 23083 59024 23189
rect 59660 23057 59792 23165
rect 63221 23973 63286 24027
rect 64316 23961 64384 24036
rect 62616 23359 62748 23467
rect 61473 22714 61605 22822
rect 63371 22714 63503 22822
rect 59195 21952 59313 22070
rect 59940 21994 60048 22126
rect 58692 21610 58785 21689
rect 59655 21453 59787 21561
rect 62118 21836 62181 21852
rect 62118 21802 62147 21836
rect 62147 21802 62181 21836
rect 62118 21786 62181 21802
rect 60242 20758 60305 20810
rect 59935 20390 60043 20522
rect 59197 20175 59309 20281
rect 61418 20318 61550 20426
rect 63316 20318 63448 20426
rect 45026 19907 45154 19985
rect 51539 19723 51650 19834
rect 58127 19533 58261 19651
rect 39618 19157 39750 19265
rect 40440 19167 40496 19181
rect 40440 19133 40446 19167
rect 40446 19133 40480 19167
rect 40480 19133 40496 19167
rect 40440 19115 40496 19133
rect 40765 19157 40897 19265
rect 39739 18369 39804 18423
rect 40277 17755 40409 17863
rect 41560 19043 41626 19059
rect 41560 19009 41576 19043
rect 41576 19009 41610 19043
rect 41610 19009 41626 19043
rect 41560 18993 41626 19009
rect 43247 19103 43379 19211
rect 46176 19153 46308 19261
rect 46998 19163 47054 19177
rect 46998 19129 47004 19163
rect 47004 19129 47038 19163
rect 47038 19129 47054 19163
rect 46998 19111 47054 19129
rect 47323 19153 47455 19261
rect 40861 18346 40960 18443
rect 42991 18040 43099 18172
rect 45199 18353 45267 18428
rect 46297 18365 46362 18419
rect 44513 17996 44737 18132
rect 41419 17757 41551 17865
rect 43233 17453 43365 17561
rect 44001 17479 44113 17585
rect 39522 17110 39654 17218
rect 41420 17110 41552 17218
rect 42977 16390 43085 16522
rect 40844 16232 40907 16248
rect 40844 16198 40878 16232
rect 40878 16198 40907 16232
rect 40844 16182 40907 16198
rect 43712 16348 43830 16466
rect 44495 17462 44496 17568
rect 44496 17462 44607 17568
rect 46835 17751 46967 17859
rect 48118 19039 48184 19055
rect 48118 19005 48134 19039
rect 48134 19005 48168 19039
rect 48168 19005 48184 19039
rect 48118 18989 48184 19005
rect 49805 19099 49937 19207
rect 52710 19158 52842 19266
rect 53532 19168 53588 19182
rect 53532 19134 53538 19168
rect 53538 19134 53572 19168
rect 53572 19134 53588 19168
rect 53532 19116 53588 19134
rect 53857 19158 53989 19266
rect 47419 18342 47518 18439
rect 49549 18036 49657 18168
rect 51733 18358 51801 18433
rect 52831 18370 52896 18424
rect 51056 17990 51306 18146
rect 47977 17753 48109 17861
rect 49791 17449 49923 17557
rect 50559 17475 50671 17581
rect 46080 17106 46212 17214
rect 47978 17106 48110 17214
rect 44496 16454 44608 16456
rect 44490 16350 44608 16454
rect 49535 16386 49643 16518
rect 44490 16348 44602 16350
rect 44240 16006 44333 16085
rect 43238 15849 43370 15957
rect 42720 15154 42783 15206
rect 39577 14714 39709 14822
rect 41475 14714 41607 14822
rect 42982 14786 43090 14918
rect 43716 14571 43828 14677
rect 47402 16228 47465 16244
rect 47402 16194 47436 16228
rect 47436 16194 47465 16228
rect 47402 16178 47465 16194
rect 50270 16344 50388 16462
rect 51053 17559 51165 17564
rect 51053 17462 51059 17559
rect 51059 17462 51162 17559
rect 51162 17462 51165 17559
rect 51053 17458 51165 17462
rect 53369 17756 53501 17864
rect 54652 19044 54718 19060
rect 54652 19010 54668 19044
rect 54668 19010 54702 19044
rect 54702 19010 54718 19044
rect 54652 18994 54718 19010
rect 56339 19104 56471 19212
rect 59223 19161 59355 19269
rect 60045 19171 60101 19185
rect 60045 19137 60051 19171
rect 60051 19137 60085 19171
rect 60085 19137 60101 19171
rect 60045 19119 60101 19137
rect 60370 19161 60502 19269
rect 53953 18347 54052 18444
rect 56083 18041 56191 18173
rect 58246 18361 58314 18436
rect 59344 18373 59409 18427
rect 57605 17998 57833 18135
rect 54511 17758 54643 17866
rect 56325 17454 56457 17562
rect 57093 17480 57205 17586
rect 52614 17111 52746 17219
rect 54512 17111 54644 17219
rect 51054 16450 51166 16452
rect 51048 16346 51166 16450
rect 56069 16391 56177 16523
rect 51048 16344 51160 16346
rect 50798 16002 50891 16081
rect 49796 15845 49928 15953
rect 49278 15150 49341 15202
rect 46135 14710 46267 14818
rect 48033 14710 48165 14818
rect 49540 14782 49648 14914
rect 50274 14567 50386 14673
rect 53936 16233 53999 16249
rect 53936 16199 53970 16233
rect 53970 16199 53999 16233
rect 53936 16183 53999 16199
rect 56804 16349 56922 16467
rect 57587 17563 57699 17569
rect 57587 17471 57595 17563
rect 57595 17471 57693 17563
rect 57693 17471 57699 17563
rect 57587 17463 57699 17471
rect 59882 17759 60014 17867
rect 61165 19047 61231 19063
rect 61165 19013 61181 19047
rect 61181 19013 61215 19047
rect 61215 19013 61231 19047
rect 61165 18997 61231 19013
rect 62852 19107 62984 19215
rect 60466 18350 60565 18447
rect 62596 18044 62704 18176
rect 64118 17998 64350 18129
rect 61024 17761 61156 17869
rect 62838 17457 62970 17565
rect 63606 17483 63718 17589
rect 59127 17114 59259 17222
rect 61025 17114 61157 17222
rect 57588 16455 57700 16457
rect 57582 16351 57700 16455
rect 62582 16394 62690 16526
rect 57582 16349 57694 16351
rect 57332 16007 57425 16086
rect 56330 15850 56462 15958
rect 55812 15155 55875 15207
rect 52669 14715 52801 14823
rect 54567 14715 54699 14823
rect 56074 14787 56182 14919
rect 56808 14572 56920 14678
rect 60449 16236 60512 16252
rect 60449 16202 60483 16236
rect 60483 16202 60512 16236
rect 60449 16186 60512 16202
rect 63317 16352 63435 16470
rect 71327 22147 71395 22204
rect 71495 22200 71563 22204
rect 71495 22151 71499 22200
rect 71499 22151 71559 22200
rect 71559 22151 71563 22200
rect 71495 22147 71563 22151
rect 64101 16458 64213 16460
rect 64095 16354 64213 16458
rect 64095 16352 64207 16354
rect 63845 16010 63938 16089
rect 62843 15853 62975 15961
rect 62325 15158 62388 15210
rect 59182 14718 59314 14826
rect 61080 14718 61212 14826
rect 62587 14790 62695 14922
rect 70269 20809 70329 20813
rect 70269 20737 70275 20809
rect 70275 20737 70329 20809
rect 70269 20733 70329 20737
rect 71212 21956 71275 21960
rect 71212 21896 71216 21956
rect 71216 21896 71271 21956
rect 71271 21896 71275 21956
rect 71212 21889 71275 21896
rect 71495 20989 71560 20993
rect 71495 20929 71500 20989
rect 71500 20929 71555 20989
rect 71555 20929 71560 20989
rect 71495 20925 71560 20929
rect 71212 20871 71274 20875
rect 71212 20811 71215 20871
rect 71215 20811 71270 20871
rect 71270 20811 71274 20871
rect 71212 20805 71274 20811
rect 72487 20795 72539 20799
rect 72487 20737 72533 20795
rect 72533 20737 72539 20795
rect 72487 20733 72539 20737
rect 71332 20621 71392 20634
rect 71332 20587 71346 20621
rect 71346 20587 71380 20621
rect 71380 20587 71392 20621
rect 71332 20575 71392 20587
rect 68248 19149 68316 19159
rect 68248 19086 68260 19149
rect 68260 19086 68309 19149
rect 68309 19086 68316 19149
rect 68248 19076 68316 19086
rect 71327 19003 71395 19060
rect 71495 19056 71563 19060
rect 71495 19007 71499 19056
rect 71499 19007 71559 19056
rect 71559 19007 71563 19056
rect 71495 19003 71563 19007
rect 70269 17665 70329 17669
rect 70269 17593 70275 17665
rect 70275 17593 70329 17665
rect 70269 17589 70329 17593
rect 71212 18812 71275 18816
rect 71212 18752 71216 18812
rect 71216 18752 71271 18812
rect 71271 18752 71275 18812
rect 71212 18745 71275 18752
rect 71495 17845 71560 17849
rect 71495 17785 71500 17845
rect 71500 17785 71555 17845
rect 71555 17785 71560 17845
rect 71495 17781 71560 17785
rect 71212 17727 71274 17731
rect 71212 17667 71215 17727
rect 71215 17667 71270 17727
rect 71270 17667 71274 17727
rect 71212 17661 71274 17667
rect 72487 17651 72539 17655
rect 72487 17593 72533 17651
rect 72533 17593 72539 17651
rect 72487 17589 72539 17593
rect 71332 17477 71392 17490
rect 71332 17443 71346 17477
rect 71346 17443 71380 17477
rect 71380 17443 71392 17477
rect 71332 17431 71392 17443
rect 71323 15871 71391 15928
rect 71491 15924 71559 15928
rect 71491 15875 71495 15924
rect 71495 15875 71555 15924
rect 71555 15875 71559 15924
rect 71491 15871 71559 15875
rect 63321 14575 63433 14681
rect 64375 13504 64526 13505
rect 64365 13415 64526 13504
rect 64375 13414 64526 13415
rect 57855 13258 58004 13346
rect 51328 13111 51484 13199
rect 57731 13155 57817 13164
rect 57731 13097 57742 13155
rect 57742 13097 57810 13155
rect 57810 13097 57817 13155
rect 57731 13089 57817 13097
rect 44758 12942 44887 13039
rect 51208 13036 51295 13043
rect 51208 12980 51217 13036
rect 51217 12980 51288 13036
rect 51288 12980 51295 13036
rect 51208 12973 51295 12980
rect 68502 12784 68646 12865
rect 44633 12703 44726 12710
rect 44633 12658 44641 12703
rect 44641 12658 44720 12703
rect 44720 12658 44726 12703
rect 44633 12649 44726 12658
rect 41911 12313 41971 12375
rect 48460 12312 48520 12374
rect 55114 12333 55174 12395
rect 33107 11105 33164 11159
rect 42133 11163 42195 11171
rect 42133 11117 42139 11163
rect 42139 11117 42191 11163
rect 42191 11117 42195 11163
rect 42133 11111 42195 11117
rect 33893 10779 33977 10837
rect 34131 10449 34199 10452
rect 34131 10404 34138 10449
rect 34138 10404 34195 10449
rect 34195 10404 34199 10449
rect 34131 10400 34199 10404
rect 35247 10413 35307 10475
rect 38237 10236 38271 10268
rect 38271 10236 38338 10268
rect 38338 10236 38369 10268
rect 38237 10160 38369 10236
rect 40719 10286 40753 10322
rect 40753 10286 40820 10322
rect 40820 10286 40851 10322
rect 40719 10214 40851 10286
rect 33775 9226 33865 9318
rect 35469 9263 35531 9271
rect 35469 9217 35475 9263
rect 35475 9217 35527 9263
rect 35527 9217 35531 9263
rect 35469 9211 35531 9217
rect 41120 10224 41176 10238
rect 41120 10190 41136 10224
rect 41136 10190 41170 10224
rect 41170 10190 41176 10224
rect 41120 10172 41176 10190
rect 41866 10288 41895 10322
rect 41895 10288 41962 10322
rect 41962 10288 41998 10322
rect 41866 10214 41998 10288
rect 39990 10100 40056 10116
rect 39990 10066 40006 10100
rect 40006 10066 40040 10100
rect 40040 10066 40056 10100
rect 39990 10050 40056 10066
rect 40656 9403 40755 9500
rect 38517 9196 38625 9229
rect 33103 9042 33166 9103
rect 38517 9129 38612 9196
rect 38612 9129 38625 9196
rect 38517 9097 38625 9129
rect 37009 8519 37121 8625
rect 35239 7828 35299 7890
rect 37008 7511 37120 7513
rect 37008 7407 37126 7511
rect 37014 7405 37126 7407
rect 33103 6978 33166 7039
rect 40065 8825 40197 8922
rect 40065 8814 40098 8825
rect 40098 8814 40165 8825
rect 40165 8814 40197 8825
rect 37503 8536 37615 8642
rect 38251 8585 38283 8618
rect 38283 8585 38350 8618
rect 38350 8585 38383 8618
rect 38251 8510 38383 8585
rect 41812 9426 41877 9480
rect 48682 11162 48744 11170
rect 48682 11116 48688 11162
rect 48688 11116 48740 11162
rect 48740 11116 48744 11162
rect 48682 11110 48744 11116
rect 48116 10681 48173 10735
rect 55336 11183 55398 11191
rect 55336 11137 55342 11183
rect 55342 11137 55394 11183
rect 55394 11137 55398 11183
rect 55336 11131 55398 11137
rect 44786 10324 44820 10356
rect 44820 10324 44887 10356
rect 44887 10324 44918 10356
rect 44786 10248 44918 10324
rect 47268 10375 47303 10410
rect 47303 10375 47370 10410
rect 47370 10375 47400 10410
rect 47268 10302 47400 10375
rect 47669 10312 47725 10326
rect 47669 10278 47685 10312
rect 47685 10278 47719 10312
rect 47719 10278 47725 10312
rect 47669 10260 47725 10278
rect 48415 10377 48447 10410
rect 48447 10377 48514 10410
rect 48514 10377 48547 10410
rect 48415 10302 48547 10377
rect 46539 10188 46605 10204
rect 46539 10154 46555 10188
rect 46555 10154 46589 10188
rect 46589 10154 46605 10188
rect 46539 10138 46605 10154
rect 47205 9491 47304 9588
rect 45066 9278 45174 9317
rect 45066 9211 45158 9278
rect 45158 9211 45174 9278
rect 45066 9185 45174 9211
rect 41207 8827 41339 8920
rect 41207 8812 41236 8827
rect 41236 8812 41303 8827
rect 41303 8812 41339 8827
rect 43558 8607 43670 8713
rect 40064 8167 40196 8275
rect 41962 8243 41995 8275
rect 41995 8243 42062 8275
rect 42062 8243 42094 8275
rect 41962 8167 42094 8243
rect 37786 7405 37904 7523
rect 38531 7546 38639 7579
rect 38531 7479 38627 7546
rect 38627 7479 38639 7546
rect 38531 7447 38639 7479
rect 37283 7063 37376 7142
rect 33932 6597 34019 6701
rect 33102 4907 33169 4974
rect 33108 2846 33164 2900
rect 34729 6600 34806 6696
rect 35461 6678 35523 6686
rect 35461 6632 35467 6678
rect 35467 6632 35519 6678
rect 35519 6632 35523 6678
rect 35461 6626 35523 6632
rect 38246 6979 38281 7014
rect 38281 6979 38348 7014
rect 38348 6979 38378 7014
rect 38246 6906 38378 6979
rect 40709 7289 40772 7305
rect 40709 7255 40738 7289
rect 40738 7255 40772 7289
rect 40709 7239 40772 7255
rect 38833 6211 38896 6263
rect 38526 5938 38634 5975
rect 38526 5871 38625 5938
rect 38625 5871 38634 5938
rect 38526 5843 38634 5871
rect 37788 5628 37900 5734
rect 40009 5785 40141 5879
rect 40009 5771 40038 5785
rect 40038 5771 40105 5785
rect 40105 5771 40141 5785
rect 41907 5771 42039 5879
rect 35220 4550 35280 4612
rect 38229 4456 38259 4488
rect 38259 4456 38326 4488
rect 38326 4456 38361 4488
rect 38229 4380 38361 4456
rect 40711 4511 40739 4542
rect 40739 4511 40806 4542
rect 40806 4511 40843 4542
rect 40711 4434 40843 4511
rect 41112 4444 41168 4458
rect 41112 4410 41128 4444
rect 41128 4410 41162 4444
rect 41162 4410 41168 4444
rect 41112 4392 41168 4410
rect 41858 4508 41895 4542
rect 41895 4508 41962 4542
rect 41962 4508 41990 4542
rect 41858 4434 41990 4508
rect 39982 4320 40048 4336
rect 39982 4286 39998 4320
rect 39998 4286 40032 4320
rect 40032 4286 40048 4320
rect 39982 4270 40048 4286
rect 35442 3400 35504 3408
rect 35442 3354 35448 3400
rect 35448 3354 35500 3400
rect 35500 3354 35504 3400
rect 35442 3348 35504 3354
rect 40648 3623 40747 3720
rect 38509 3409 38617 3449
rect 38509 3342 38602 3409
rect 38602 3342 38617 3409
rect 38509 3317 38617 3342
rect 37001 2739 37113 2845
rect 35236 1790 35296 1852
rect 40057 3048 40189 3142
rect 40057 3034 40079 3048
rect 40079 3034 40146 3048
rect 40146 3034 40189 3048
rect 37495 2756 37607 2862
rect 38243 2803 38280 2838
rect 38280 2803 38347 2838
rect 38347 2803 38375 2838
rect 38243 2730 38375 2803
rect 41804 3646 41869 3700
rect 46614 8921 46746 9010
rect 46614 8902 46643 8921
rect 46643 8902 46710 8921
rect 46710 8902 46746 8921
rect 44052 8624 44164 8730
rect 44800 8672 44834 8706
rect 44834 8672 44901 8706
rect 44901 8672 44932 8706
rect 44800 8598 44932 8672
rect 48361 9514 48426 9568
rect 49456 9502 49524 9577
rect 47756 8913 47888 9008
rect 47756 8900 47782 8913
rect 47782 8900 47849 8913
rect 47849 8900 47888 8913
rect 46613 8255 46745 8363
rect 48511 8330 48549 8363
rect 48549 8330 48616 8363
rect 48616 8330 48643 8363
rect 48511 8255 48643 8330
rect 44335 7493 44453 7611
rect 45080 7628 45188 7667
rect 45080 7561 45176 7628
rect 45176 7561 45188 7628
rect 45080 7535 45188 7561
rect 43832 7151 43925 7230
rect 44795 7072 44826 7102
rect 44826 7072 44893 7102
rect 44893 7072 44927 7102
rect 44795 6994 44927 7072
rect 47258 7377 47321 7393
rect 47258 7343 47287 7377
rect 47287 7343 47321 7377
rect 47258 7327 47321 7343
rect 45382 6299 45445 6351
rect 45075 6027 45183 6063
rect 45075 5960 45173 6027
rect 45173 5960 45183 6027
rect 45075 5931 45183 5960
rect 44337 5716 44449 5822
rect 46558 5870 46690 5967
rect 46558 5859 46587 5870
rect 46587 5859 46654 5870
rect 46654 5859 46690 5870
rect 48456 5859 48588 5967
rect 49525 6801 49645 6890
rect 44780 4454 44814 4486
rect 44814 4454 44881 4486
rect 44881 4454 44912 4486
rect 44780 4378 44912 4454
rect 47262 4507 47295 4540
rect 47295 4507 47362 4540
rect 47362 4507 47394 4540
rect 47262 4432 47394 4507
rect 47663 4442 47719 4456
rect 47663 4408 47679 4442
rect 47679 4408 47713 4442
rect 47713 4408 47719 4442
rect 47663 4390 47719 4408
rect 48409 4507 48443 4540
rect 48443 4507 48510 4540
rect 48510 4507 48541 4540
rect 48409 4432 48541 4507
rect 46533 4318 46599 4334
rect 46533 4284 46549 4318
rect 46549 4284 46583 4318
rect 46583 4284 46599 4318
rect 46533 4268 46599 4284
rect 42899 3634 42967 3709
rect 47199 3621 47298 3718
rect 45060 3403 45168 3447
rect 45060 3336 45152 3403
rect 45152 3336 45168 3403
rect 45060 3315 45168 3336
rect 41199 3043 41331 3140
rect 41199 3032 41232 3043
rect 41232 3032 41299 3043
rect 41299 3032 41331 3043
rect 40056 2387 40188 2495
rect 41954 2462 41986 2495
rect 41986 2462 42053 2495
rect 42053 2462 42086 2495
rect 41954 2387 42086 2462
rect 37778 1625 37896 1743
rect 38523 1759 38631 1799
rect 38523 1692 38610 1759
rect 38610 1692 38631 1759
rect 38523 1667 38631 1692
rect 37275 1283 37368 1362
rect 33774 957 33861 1038
rect 34127 969 34208 1032
rect 33108 778 33164 832
rect 33108 -1284 33164 -1230
rect 30501 -1396 30567 -1330
rect 30698 -1383 30757 -1318
rect 29699 -2148 29753 -2138
rect 29699 -2186 29707 -2148
rect 29707 -2186 29745 -2148
rect 29745 -2186 29753 -2148
rect 29699 -2192 29753 -2186
rect 31923 -2086 31981 -2080
rect 31923 -2136 31929 -2086
rect 31929 -2136 31971 -2086
rect 31971 -2136 31981 -2086
rect 31923 -2142 31981 -2136
rect 35458 640 35520 648
rect 35458 594 35464 640
rect 35464 594 35516 640
rect 35516 594 35520 640
rect 35458 588 35520 594
rect 38238 1204 38269 1234
rect 38269 1204 38336 1234
rect 38336 1204 38370 1234
rect 38238 1126 38370 1204
rect 40701 1509 40764 1525
rect 40701 1475 40730 1509
rect 40730 1475 40764 1509
rect 40701 1459 40764 1475
rect 38825 431 38888 483
rect 38518 167 38626 195
rect 38518 100 38610 167
rect 38610 100 38626 167
rect 38518 63 38626 100
rect 37780 -152 37892 -46
rect 40001 -1 40133 99
rect 40001 -9 40031 -1
rect 40031 -9 40098 -1
rect 40098 -9 40133 -1
rect 41899 -9 42031 99
rect 43552 2737 43664 2843
rect 42168 -723 42230 -717
rect 42168 -769 42174 -723
rect 42174 -769 42226 -723
rect 42226 -769 42230 -723
rect 42168 -777 42230 -769
rect 41229 -1042 41305 -956
rect 41460 -1174 41589 -1083
rect 46608 3045 46740 3140
rect 46608 3032 46637 3045
rect 46637 3032 46704 3045
rect 46704 3032 46740 3045
rect 44046 2754 44158 2860
rect 44794 2810 44825 2836
rect 44825 2810 44892 2836
rect 44892 2810 44926 2836
rect 44794 2728 44926 2810
rect 48355 3644 48420 3698
rect 51440 10254 51473 10288
rect 51473 10254 51540 10288
rect 51540 10254 51572 10288
rect 51440 10180 51572 10254
rect 53922 10310 53954 10342
rect 53954 10310 54021 10342
rect 54021 10310 54054 10342
rect 53922 10234 54054 10310
rect 54323 10244 54379 10258
rect 54323 10210 54339 10244
rect 54339 10210 54373 10244
rect 54373 10210 54379 10244
rect 54323 10192 54379 10210
rect 55069 10309 55101 10342
rect 55101 10309 55168 10342
rect 55168 10309 55201 10342
rect 55069 10234 55201 10309
rect 53193 10120 53259 10136
rect 53193 10086 53209 10120
rect 53209 10086 53243 10120
rect 53243 10086 53259 10120
rect 53193 10070 53259 10086
rect 53859 9423 53958 9520
rect 51720 9212 51828 9249
rect 51720 9145 51808 9212
rect 51808 9145 51828 9212
rect 51720 9117 51828 9145
rect 50211 7531 50323 7533
rect 50211 7427 50329 7531
rect 50217 7426 50329 7427
rect 50217 7425 50329 7426
rect 53268 8849 53400 8942
rect 53268 8834 53296 8849
rect 53296 8834 53363 8849
rect 53363 8834 53400 8849
rect 50706 8556 50818 8662
rect 51454 8606 51488 8638
rect 51488 8606 51555 8638
rect 51555 8606 51586 8638
rect 51454 8530 51586 8606
rect 55015 9446 55080 9500
rect 58065 10323 58093 10356
rect 58093 10323 58160 10356
rect 58160 10323 58197 10356
rect 58065 10248 58197 10323
rect 60547 10375 60577 10410
rect 60577 10375 60644 10410
rect 60644 10375 60679 10410
rect 60547 10302 60679 10375
rect 60948 10312 61004 10326
rect 60948 10278 60964 10312
rect 60964 10278 60998 10312
rect 60998 10278 61004 10312
rect 60948 10260 61004 10278
rect 61694 10381 61726 10410
rect 61726 10381 61793 10410
rect 61793 10381 61826 10410
rect 61694 10302 61826 10381
rect 59818 10188 59884 10204
rect 59818 10154 59834 10188
rect 59834 10154 59868 10188
rect 59868 10154 59884 10188
rect 59818 10138 59884 10154
rect 60484 9491 60583 9588
rect 58345 9288 58453 9317
rect 58345 9221 58440 9288
rect 58440 9221 58453 9288
rect 58345 9185 58453 9221
rect 54410 8852 54542 8940
rect 54410 8832 54442 8852
rect 54442 8832 54509 8852
rect 54509 8832 54542 8852
rect 56837 8607 56949 8713
rect 53267 8187 53399 8295
rect 55165 8258 55195 8295
rect 55195 8258 55262 8295
rect 55262 8258 55297 8295
rect 55165 8187 55297 8258
rect 50989 7425 51107 7543
rect 51734 7561 51842 7599
rect 51734 7494 51825 7561
rect 51825 7494 51842 7561
rect 51734 7467 51842 7494
rect 50486 7083 50579 7162
rect 51449 7003 51483 7034
rect 51483 7003 51550 7034
rect 51550 7003 51581 7034
rect 51449 6926 51581 7003
rect 53912 7309 53975 7325
rect 53912 7275 53941 7309
rect 53941 7275 53975 7309
rect 53912 7259 53975 7275
rect 52036 6231 52099 6283
rect 51729 5956 51837 5995
rect 51729 5889 51827 5956
rect 51827 5889 51837 5956
rect 51729 5863 51837 5889
rect 50991 5648 51103 5754
rect 53212 5804 53344 5899
rect 53212 5791 53236 5804
rect 53236 5791 53303 5804
rect 53303 5791 53344 5804
rect 55110 5791 55242 5899
rect 56163 5503 56286 5512
rect 56163 5404 56172 5503
rect 56172 5404 56278 5503
rect 56278 5404 56286 5503
rect 56163 5398 56286 5404
rect 51435 4451 51465 4487
rect 51465 4451 51532 4487
rect 51532 4451 51567 4487
rect 51435 4379 51567 4451
rect 53917 4511 53950 4541
rect 53950 4511 54017 4541
rect 54017 4511 54049 4541
rect 53917 4433 54049 4511
rect 54318 4443 54374 4457
rect 54318 4409 54334 4443
rect 54334 4409 54368 4443
rect 54368 4409 54374 4443
rect 54318 4391 54374 4409
rect 55064 4508 55099 4541
rect 55099 4508 55166 4541
rect 55166 4508 55196 4541
rect 55064 4433 55196 4508
rect 53188 4319 53254 4335
rect 53188 4285 53204 4319
rect 53204 4285 53238 4319
rect 53238 4285 53254 4319
rect 53188 4269 53254 4285
rect 53854 3622 53953 3719
rect 51715 3412 51823 3448
rect 51715 3345 51813 3412
rect 51813 3345 51823 3412
rect 51715 3316 51823 3345
rect 47750 3034 47882 3138
rect 47750 3030 47778 3034
rect 47778 3030 47845 3034
rect 47845 3030 47882 3034
rect 50140 2736 50344 2849
rect 50292 2735 50344 2736
rect 46607 2385 46739 2493
rect 48505 2461 48542 2493
rect 48542 2461 48609 2493
rect 48609 2461 48637 2493
rect 48505 2385 48637 2461
rect 44329 1623 44447 1741
rect 45074 1758 45182 1797
rect 45074 1691 45168 1758
rect 45168 1691 45182 1758
rect 45074 1665 45182 1691
rect 43826 1281 43919 1360
rect 44789 1199 44825 1232
rect 44825 1199 44892 1232
rect 44892 1199 44921 1232
rect 44789 1124 44921 1199
rect 47252 1507 47315 1523
rect 47252 1473 47281 1507
rect 47281 1473 47315 1507
rect 47252 1457 47315 1473
rect 45376 429 45439 481
rect 45069 158 45177 193
rect 45069 91 45157 158
rect 45157 91 45177 158
rect 45069 61 45177 91
rect 44331 -154 44443 -48
rect 46552 -2 46684 97
rect 46552 -11 46579 -2
rect 46579 -11 46646 -2
rect 46646 -11 46684 -2
rect 48450 -11 48582 97
rect 48722 -718 48784 -712
rect 48722 -764 48728 -718
rect 48728 -764 48780 -718
rect 48780 -764 48784 -718
rect 48722 -772 48784 -764
rect 41946 -1981 42006 -1919
rect 30507 -2772 30561 -2718
rect 53263 3049 53395 3141
rect 53263 3033 53289 3049
rect 53289 3033 53356 3049
rect 53356 3033 53395 3049
rect 50701 2755 50813 2861
rect 51449 2805 51485 2837
rect 51485 2805 51552 2837
rect 51552 2805 51581 2837
rect 51449 2729 51581 2805
rect 55010 3645 55075 3699
rect 59893 8908 60025 9010
rect 59893 8902 59917 8908
rect 59917 8902 59984 8908
rect 59984 8902 60025 8908
rect 57331 8624 57443 8730
rect 58079 8672 58116 8706
rect 58116 8672 58183 8706
rect 58183 8672 58211 8706
rect 58079 8598 58211 8672
rect 61640 9514 61705 9568
rect 62618 9502 62686 9577
rect 61035 8910 61167 9008
rect 61035 8900 61060 8910
rect 61060 8900 61127 8910
rect 61127 8900 61167 8910
rect 59892 8255 60024 8363
rect 61790 8327 61823 8363
rect 61823 8327 61890 8363
rect 61890 8327 61922 8363
rect 61790 8255 61922 8327
rect 57614 7493 57732 7611
rect 58359 7627 58467 7667
rect 58359 7560 58445 7627
rect 58445 7560 58467 7627
rect 58359 7535 58467 7560
rect 57111 7151 57204 7230
rect 56632 6724 56728 6824
rect 58074 7064 58108 7102
rect 58108 7064 58175 7102
rect 58175 7064 58206 7102
rect 58074 6994 58206 7064
rect 60537 7377 60600 7393
rect 60537 7343 60566 7377
rect 60566 7343 60600 7377
rect 60537 7327 60600 7343
rect 58661 6299 58724 6351
rect 58354 6022 58462 6063
rect 58354 5955 58451 6022
rect 58451 5955 58462 6022
rect 58354 5931 58462 5955
rect 57616 5716 57728 5822
rect 59837 5870 59969 5967
rect 59837 5859 59867 5870
rect 59867 5859 59934 5870
rect 59934 5859 59969 5870
rect 61735 5859 61867 5967
rect 63767 12166 63827 12228
rect 66024 12123 66156 12157
rect 66024 12049 66156 12123
rect 67368 11758 67428 11820
rect 63112 11081 63191 11155
rect 63264 10945 63345 11041
rect 65221 11180 65288 11243
rect 63989 11016 64051 11024
rect 63989 10970 63995 11016
rect 63995 10970 64047 11016
rect 64047 10970 64051 11016
rect 63989 10964 64051 10970
rect 65221 11054 65288 11117
rect 63762 9595 63822 9657
rect 65481 11108 65536 11125
rect 65481 11074 65486 11108
rect 65486 11074 65520 11108
rect 65520 11074 65536 11108
rect 65481 11057 65536 11074
rect 66535 10796 66597 10887
rect 66877 11227 66930 11238
rect 66877 11193 66886 11227
rect 66886 11193 66920 11227
rect 66920 11193 66930 11227
rect 66877 11182 66930 11193
rect 67001 11046 67074 11135
rect 67990 11072 68102 11130
rect 67774 10801 67882 10882
rect 67590 10608 67652 10616
rect 67590 10562 67596 10608
rect 67596 10562 67648 10608
rect 67648 10562 67652 10608
rect 67590 10556 67652 10562
rect 65954 9813 66128 9822
rect 65954 9711 65973 9813
rect 65973 9711 66108 9813
rect 66108 9711 66128 9813
rect 65954 9699 66128 9711
rect 63411 8633 63493 8714
rect 63984 8445 64046 8453
rect 63984 8399 63990 8445
rect 63990 8399 64042 8445
rect 64042 8399 64046 8445
rect 63984 8393 64046 8399
rect 66026 8032 66158 8066
rect 66026 7958 66158 8032
rect 67370 7667 67430 7729
rect 65223 7089 65290 7152
rect 63762 6562 63822 6624
rect 63516 5726 63605 5813
rect 57272 5503 57395 5512
rect 57272 5404 57281 5503
rect 57281 5404 57387 5503
rect 57387 5404 57395 5503
rect 57272 5398 57395 5404
rect 65223 6963 65290 7026
rect 63984 5412 64046 5420
rect 63984 5366 63990 5412
rect 63990 5366 64042 5412
rect 64042 5366 64046 5412
rect 63984 5360 64046 5366
rect 63833 4642 63893 4704
rect 58057 4456 58089 4488
rect 58089 4456 58156 4488
rect 58156 4456 58189 4488
rect 58057 4380 58189 4456
rect 60539 4504 60568 4542
rect 60568 4504 60635 4542
rect 60635 4504 60671 4542
rect 60539 4434 60671 4504
rect 60940 4444 60996 4458
rect 60940 4410 60956 4444
rect 60956 4410 60990 4444
rect 60990 4410 60996 4444
rect 60940 4392 60996 4410
rect 61686 4510 61716 4542
rect 61716 4510 61783 4542
rect 61783 4510 61818 4542
rect 61686 4434 61818 4510
rect 59810 4320 59876 4336
rect 59810 4286 59826 4320
rect 59826 4286 59860 4320
rect 59860 4286 59876 4320
rect 59810 4270 59876 4286
rect 56105 3633 56173 3708
rect 60476 3623 60575 3720
rect 58337 3417 58445 3449
rect 58337 3350 58429 3417
rect 58429 3350 58445 3417
rect 58337 3317 58445 3350
rect 54405 3052 54537 3139
rect 54405 3031 54435 3052
rect 54435 3031 54502 3052
rect 54502 3031 54537 3052
rect 53262 2386 53394 2494
rect 55160 2463 55196 2494
rect 55196 2463 55263 2494
rect 55263 2463 55292 2494
rect 55160 2386 55292 2463
rect 50984 1624 51102 1742
rect 51729 1761 51837 1798
rect 51729 1694 51824 1761
rect 51824 1694 51837 1761
rect 51729 1666 51837 1694
rect 50481 1282 50574 1361
rect 51444 1197 51480 1233
rect 51480 1197 51547 1233
rect 51547 1197 51576 1233
rect 51444 1125 51576 1197
rect 53907 1508 53970 1524
rect 53907 1474 53936 1508
rect 53936 1474 53970 1508
rect 53907 1458 53970 1474
rect 52031 430 52094 482
rect 51724 152 51832 194
rect 51724 85 51827 152
rect 51827 85 51832 152
rect 51724 62 51832 85
rect 50169 -97 50271 -85
rect 50169 -165 50188 -97
rect 50188 -165 50258 -97
rect 50258 -165 50271 -97
rect 50169 -172 50271 -165
rect 50986 -153 51098 -47
rect 53207 -1 53339 98
rect 53207 -10 53229 -1
rect 53229 -10 53296 -1
rect 53296 -10 53339 -1
rect 55105 -10 55237 98
rect 56829 2739 56941 2845
rect 55371 -730 55433 -724
rect 55371 -776 55377 -730
rect 55377 -776 55429 -730
rect 55429 -776 55433 -730
rect 55371 -784 55433 -776
rect 48500 -1976 48560 -1914
rect 54657 -1181 54726 -1092
rect 56828 1731 56940 1733
rect 56828 1627 56946 1731
rect 56834 1625 56946 1627
rect 59885 3053 60017 3142
rect 59885 3034 59920 3053
rect 59920 3034 59987 3053
rect 59987 3034 60017 3053
rect 57323 2756 57435 2862
rect 58071 2806 58104 2838
rect 58104 2806 58171 2838
rect 58171 2806 58203 2838
rect 58071 2730 58203 2806
rect 65483 7017 65538 7034
rect 65483 6983 65488 7017
rect 65488 6983 65522 7017
rect 65522 6983 65538 7017
rect 65483 6966 65538 6983
rect 66537 6705 66599 6796
rect 66879 7136 66932 7147
rect 66879 7102 66888 7136
rect 66888 7102 66922 7136
rect 66922 7102 66932 7136
rect 66879 7091 66932 7102
rect 67003 6955 67076 7044
rect 67592 6517 67654 6525
rect 67592 6471 67598 6517
rect 67598 6471 67650 6517
rect 67650 6471 67654 6517
rect 67592 6465 67654 6471
rect 65956 5722 66130 5731
rect 65956 5620 65975 5722
rect 65975 5620 66110 5722
rect 66110 5620 66130 5722
rect 65956 5608 66130 5620
rect 66026 4537 66158 4571
rect 66026 4463 66158 4537
rect 61632 3646 61697 3700
rect 63568 3591 63654 3692
rect 67370 4172 67430 4234
rect 63340 3458 63425 3518
rect 64055 3492 64117 3500
rect 64055 3446 64061 3492
rect 64061 3446 64113 3492
rect 64113 3446 64117 3492
rect 64055 3440 64117 3446
rect 65223 3468 65290 3531
rect 61027 3044 61159 3140
rect 61027 3032 61054 3044
rect 61054 3032 61121 3044
rect 61121 3032 61159 3044
rect 59884 2387 60016 2495
rect 61782 2461 61817 2495
rect 61817 2461 61884 2495
rect 61884 2461 61914 2495
rect 61782 2387 61914 2461
rect 57606 1625 57724 1743
rect 58351 1768 58459 1799
rect 58351 1701 58447 1768
rect 58447 1701 58459 1768
rect 58351 1667 58459 1701
rect 57103 1283 57196 1362
rect 58066 1197 58101 1234
rect 58101 1197 58168 1234
rect 58168 1197 58198 1234
rect 58066 1126 58198 1197
rect 60529 1509 60592 1525
rect 60529 1475 60558 1509
rect 60558 1475 60592 1509
rect 60529 1459 60592 1475
rect 63830 1572 63890 1634
rect 58653 431 58716 483
rect 58346 151 58454 195
rect 58346 84 58438 151
rect 58438 84 58454 151
rect 58346 63 58454 84
rect 57608 -152 57720 -46
rect 59829 5 59961 99
rect 59829 -9 59857 5
rect 59857 -9 59924 5
rect 59924 -9 59961 5
rect 61727 -9 61859 99
rect 62795 936 62912 1017
rect 65483 3522 65538 3539
rect 65483 3488 65488 3522
rect 65488 3488 65522 3522
rect 65522 3488 65538 3522
rect 65483 3471 65538 3488
rect 66537 3210 66599 3301
rect 66879 3641 66932 3652
rect 66879 3607 66888 3641
rect 66888 3607 66922 3641
rect 66922 3607 66932 3641
rect 66879 3596 66932 3607
rect 67003 3460 67076 3549
rect 67592 3022 67654 3030
rect 67592 2976 67598 3022
rect 67598 2976 67650 3022
rect 67650 2976 67654 3022
rect 67592 2970 67654 2976
rect 65956 2227 66130 2236
rect 65956 2125 65975 2227
rect 65975 2125 66110 2227
rect 66110 2125 66130 2227
rect 65956 2113 66130 2125
rect 63170 608 63254 698
rect 68186 3288 68296 3300
rect 68186 3216 68192 3288
rect 68192 3216 68287 3288
rect 68287 3216 68296 3288
rect 68186 3209 68296 3216
rect 63604 487 63670 551
rect 64052 422 64114 430
rect 64052 376 64058 422
rect 64058 376 64110 422
rect 64110 376 64114 422
rect 64052 370 64114 376
rect 66026 189 66158 223
rect 66026 115 66158 189
rect 70265 14533 70325 14537
rect 70265 14461 70271 14533
rect 70271 14461 70325 14533
rect 70265 14457 70325 14461
rect 71208 15680 71271 15684
rect 71208 15620 71212 15680
rect 71212 15620 71267 15680
rect 71267 15620 71271 15680
rect 71208 15613 71271 15620
rect 71491 14713 71556 14717
rect 71491 14653 71496 14713
rect 71496 14653 71551 14713
rect 71551 14653 71556 14713
rect 71491 14649 71556 14653
rect 71208 14595 71270 14599
rect 71208 14535 71211 14595
rect 71211 14535 71266 14595
rect 71266 14535 71270 14595
rect 71208 14529 71270 14535
rect 72483 14519 72535 14523
rect 72483 14461 72529 14519
rect 72529 14461 72535 14519
rect 72483 14457 72535 14461
rect 71328 14345 71388 14358
rect 71328 14311 71342 14345
rect 71342 14311 71376 14345
rect 71376 14311 71388 14345
rect 71328 14299 71388 14311
rect 71323 12727 71391 12784
rect 70265 11389 70325 11393
rect 70265 11317 70271 11389
rect 70271 11317 70325 11389
rect 70265 11313 70325 11317
rect 71208 12536 71271 12540
rect 71208 12476 71212 12536
rect 71212 12476 71267 12536
rect 71267 12476 71271 12536
rect 71208 12469 71271 12476
rect 71491 11569 71556 11573
rect 71491 11509 71496 11569
rect 71496 11509 71551 11569
rect 71551 11509 71556 11569
rect 71491 11505 71556 11509
rect 71208 11451 71270 11455
rect 71208 11391 71211 11451
rect 71211 11391 71266 11451
rect 71266 11391 71270 11451
rect 71208 11385 71270 11391
rect 72483 11375 72535 11379
rect 72483 11317 72529 11375
rect 72529 11317 72535 11375
rect 72483 11313 72535 11317
rect 71328 11201 71388 11214
rect 71328 11167 71342 11201
rect 71342 11167 71376 11201
rect 71376 11167 71388 11201
rect 71328 11155 71388 11167
rect 71327 9525 71395 9582
rect 71495 9578 71563 9582
rect 71495 9529 71499 9578
rect 71499 9529 71559 9578
rect 71559 9529 71563 9578
rect 71495 9525 71563 9529
rect 70269 8187 70329 8191
rect 70269 8115 70275 8187
rect 70275 8115 70329 8187
rect 70269 8111 70329 8115
rect 71212 9334 71275 9338
rect 71212 9274 71216 9334
rect 71216 9274 71271 9334
rect 71271 9274 71275 9334
rect 71212 9267 71275 9274
rect 71495 8367 71560 8371
rect 71495 8307 71500 8367
rect 71500 8307 71555 8367
rect 71555 8307 71560 8367
rect 71495 8303 71560 8307
rect 71212 8249 71274 8253
rect 71212 8189 71215 8249
rect 71215 8189 71270 8249
rect 71270 8189 71274 8249
rect 71212 8183 71274 8189
rect 72487 8173 72539 8177
rect 72487 8115 72533 8173
rect 72533 8115 72539 8173
rect 72487 8111 72539 8115
rect 71332 7999 71392 8012
rect 71332 7965 71346 7999
rect 71346 7965 71380 7999
rect 71380 7965 71392 7999
rect 71332 7953 71392 7965
rect 71327 6381 71395 6438
rect 70269 5043 70329 5047
rect 70269 4971 70275 5043
rect 70275 4971 70329 5043
rect 70269 4967 70329 4971
rect 71212 6190 71275 6194
rect 71212 6130 71216 6190
rect 71216 6130 71271 6190
rect 71271 6130 71275 6190
rect 71212 6123 71275 6130
rect 71495 5223 71560 5227
rect 71495 5163 71500 5223
rect 71500 5163 71555 5223
rect 71555 5163 71560 5223
rect 71495 5159 71560 5163
rect 71212 5105 71274 5109
rect 71212 5045 71215 5105
rect 71215 5045 71270 5105
rect 71270 5045 71274 5105
rect 71212 5039 71274 5045
rect 72487 5029 72539 5033
rect 72487 4971 72533 5029
rect 72533 4971 72539 5029
rect 72487 4967 72539 4971
rect 71332 4855 71392 4868
rect 71332 4821 71346 4855
rect 71346 4821 71380 4855
rect 71380 4821 71392 4855
rect 71332 4809 71392 4821
rect 71323 3249 71391 3306
rect 71491 3302 71559 3306
rect 71491 3253 71495 3302
rect 71495 3253 71555 3302
rect 71555 3253 71559 3302
rect 71491 3249 71559 3253
rect 70265 1911 70325 1915
rect 70265 1839 70271 1911
rect 70271 1839 70325 1911
rect 70265 1835 70325 1839
rect 71208 3058 71271 3062
rect 71208 2998 71212 3058
rect 71212 2998 71267 3058
rect 71267 2998 71271 3058
rect 71208 2991 71271 2998
rect 71491 2091 71556 2095
rect 71491 2031 71496 2091
rect 71496 2031 71551 2091
rect 71551 2031 71556 2091
rect 71491 2027 71556 2031
rect 71208 1973 71270 1977
rect 71208 1913 71211 1973
rect 71211 1913 71266 1973
rect 71266 1913 71270 1973
rect 71208 1907 71270 1913
rect 72483 1897 72535 1901
rect 72483 1839 72529 1897
rect 72529 1839 72535 1897
rect 72483 1835 72535 1839
rect 71328 1723 71388 1736
rect 71328 1689 71342 1723
rect 71342 1689 71376 1723
rect 71376 1689 71388 1723
rect 71328 1677 71388 1689
rect 71323 105 71391 162
rect 71491 158 71559 162
rect 71491 109 71495 158
rect 71495 109 71555 158
rect 71555 109 71559 158
rect 71491 105 71559 109
rect 67370 -176 67430 -114
rect 65223 -754 65289 -691
rect 65289 -754 65290 -691
rect 65223 -880 65290 -817
rect 63584 -1052 63668 -962
rect 55149 -1988 55209 -1926
rect 36374 -2268 36470 -2199
rect 41414 -2269 41514 -2195
rect 63837 -1273 63897 -1211
rect 34260 -2397 34359 -2311
rect 62999 -1795 63083 -1705
rect 65483 -826 65538 -809
rect 65483 -860 65488 -826
rect 65488 -860 65522 -826
rect 65522 -860 65538 -826
rect 65483 -877 65538 -860
rect 66537 -1138 66599 -1047
rect 66879 -707 66932 -696
rect 66879 -741 66888 -707
rect 66888 -741 66922 -707
rect 66922 -741 66932 -707
rect 66879 -752 66932 -741
rect 67003 -888 67076 -799
rect 67968 -876 68110 -788
rect 70265 -1233 70325 -1229
rect 70265 -1305 70271 -1233
rect 70271 -1305 70325 -1233
rect 70265 -1309 70325 -1305
rect 67592 -1326 67654 -1318
rect 67592 -1372 67598 -1326
rect 67598 -1372 67650 -1326
rect 67650 -1372 67654 -1326
rect 67592 -1378 67654 -1372
rect 41222 -2520 41314 -2448
rect 63168 -2111 63252 -2021
rect 54654 -2523 54723 -2455
rect 63481 -2445 63542 -2370
rect 65956 -2121 66130 -2112
rect 65956 -2223 65975 -2121
rect 65975 -2223 66110 -2121
rect 66110 -2223 66130 -2121
rect 65956 -2235 66130 -2223
rect 71208 -86 71271 -82
rect 71208 -146 71212 -86
rect 71212 -146 71267 -86
rect 71267 -146 71271 -86
rect 71208 -153 71271 -146
rect 71491 -1053 71556 -1049
rect 71491 -1113 71496 -1053
rect 71496 -1113 71551 -1053
rect 71551 -1113 71556 -1053
rect 71491 -1117 71556 -1113
rect 71208 -1171 71270 -1167
rect 71208 -1231 71211 -1171
rect 71211 -1231 71266 -1171
rect 71266 -1231 71270 -1171
rect 71208 -1237 71270 -1231
rect 72483 -1247 72535 -1243
rect 72483 -1305 72529 -1247
rect 72529 -1305 72535 -1247
rect 72483 -1309 72535 -1305
rect 71328 -1421 71388 -1408
rect 71328 -1455 71342 -1421
rect 71342 -1455 71376 -1421
rect 71376 -1455 71388 -1421
rect 71328 -1467 71388 -1455
rect 64059 -2423 64121 -2415
rect 64059 -2469 64065 -2423
rect 64065 -2469 64117 -2423
rect 64117 -2469 64121 -2423
rect 64059 -2475 64121 -2469
rect 36220 -2931 36315 -2877
rect 31078 -3033 31142 -2968
<< metal2 >>
rect 38134 25215 38293 25235
rect 38134 25093 38149 25215
rect 38280 25093 38293 25215
rect 4272 22268 4372 22278
rect 4272 22166 4372 22176
rect 7416 22268 7516 22278
rect 7416 22166 7516 22176
rect 10548 22264 10648 22274
rect 10548 22162 10648 22172
rect 13692 22264 13792 22274
rect 13692 22162 13792 22172
rect 16894 22268 16994 22278
rect 16894 22166 16994 22176
rect 20038 22268 20138 22278
rect 20038 22166 20138 22176
rect 23170 22264 23270 22274
rect 23170 22162 23270 22172
rect 26314 22264 26414 22274
rect 26314 22162 26414 22172
rect 27738 21445 27792 21453
rect 24704 21443 27803 21445
rect 24704 21396 27738 21443
rect 24764 21381 27738 21396
rect 27792 21381 27803 21443
rect 27724 21380 27803 21381
rect 27948 21444 28042 21454
rect 27738 21371 27792 21380
rect 27948 21371 28042 21381
rect 24704 21333 24764 21343
rect 5425 21307 5518 21309
rect 8569 21307 8662 21309
rect 18047 21307 18140 21309
rect 21191 21307 21284 21309
rect 4343 21303 10710 21307
rect 11701 21303 11794 21305
rect 14845 21303 14938 21305
rect 16965 21303 23373 21307
rect 24323 21303 24416 21305
rect 27467 21303 27560 21305
rect 27736 21303 27793 21304
rect 4343 21302 24590 21303
rect 26385 21302 27801 21303
rect 4343 21297 27804 21302
rect 2735 21242 2840 21252
rect 4343 21235 4352 21297
rect 4422 21235 5436 21297
rect 4343 21234 5436 21235
rect 5507 21235 7496 21297
rect 7566 21235 8580 21297
rect 5507 21234 8580 21235
rect 8651 21293 16974 21297
rect 8651 21234 10628 21293
rect 4343 21231 10628 21234
rect 10698 21231 11712 21293
rect 4343 21230 11712 21231
rect 11783 21231 13772 21293
rect 13842 21231 14856 21293
rect 11783 21230 14856 21231
rect 14927 21235 16974 21293
rect 17044 21235 18058 21297
rect 14927 21234 18058 21235
rect 18129 21235 20118 21297
rect 20188 21235 21202 21297
rect 18129 21234 21202 21235
rect 21273 21294 27804 21297
rect 21273 21293 27736 21294
rect 21273 21234 23250 21293
rect 14927 21231 23250 21234
rect 23320 21231 24334 21293
rect 14927 21230 24334 21231
rect 24405 21231 26394 21293
rect 26464 21231 27478 21293
rect 24405 21230 27478 21231
rect 27549 21230 27736 21293
rect 4343 21226 27736 21230
rect 27793 21226 27804 21294
rect 4343 21223 27804 21226
rect 8831 21219 15182 21223
rect 21450 21222 27804 21223
rect 21560 21219 27804 21222
rect 11960 21218 13854 21219
rect 24582 21218 26428 21219
rect 27726 21218 27804 21219
rect 27736 21216 27793 21218
rect 18316 21190 18373 21192
rect 18288 21187 18384 21190
rect 2735 21142 2840 21152
rect 4122 21182 5762 21187
rect 4122 21177 5694 21182
rect 4181 21117 5694 21177
rect 4122 21114 5694 21117
rect 5751 21114 5762 21182
rect 4122 21108 5762 21114
rect 7266 21182 9128 21187
rect 7266 21177 8838 21182
rect 7325 21117 8838 21177
rect 7266 21114 8838 21117
rect 8895 21114 9128 21182
rect 7266 21108 9128 21114
rect 4122 21107 4181 21108
rect 7266 21107 7325 21108
rect 5683 21024 5762 21034
rect 5666 21022 5683 21023
rect 4461 21014 5683 21022
rect 4461 20949 4472 21014
rect 4540 20949 5683 21014
rect 4461 20938 5683 20949
rect 8838 21023 8895 21024
rect 8810 21022 8906 21023
rect 7605 21014 8906 21022
rect 7605 20949 7616 21014
rect 7684 20949 8838 21014
rect 7605 20946 8838 20949
rect 8895 20946 8906 21014
rect 7605 20938 8906 20946
rect 8838 20936 8895 20938
rect 5683 20925 5762 20935
rect 2744 20890 2837 20900
rect 2734 20814 2744 20877
rect 9047 20877 9128 21108
rect 10398 21178 12038 21183
rect 10398 21173 11970 21178
rect 10457 21113 11970 21173
rect 10398 21110 11970 21113
rect 12027 21110 12038 21178
rect 10398 21104 12038 21110
rect 13542 21173 15449 21183
rect 13601 21113 15449 21173
rect 13542 21104 15449 21113
rect 16744 21182 18384 21187
rect 16744 21177 18316 21182
rect 16803 21117 18316 21177
rect 16744 21114 18316 21117
rect 18373 21114 18384 21182
rect 16744 21108 18384 21114
rect 16744 21107 16803 21108
rect 18288 21105 18384 21108
rect 19888 21177 21706 21187
rect 24592 21186 24649 21188
rect 24564 21183 24660 21186
rect 19947 21117 21706 21177
rect 19888 21108 21706 21117
rect 19888 21107 19947 21108
rect 18316 21104 18373 21105
rect 10398 21103 10457 21104
rect 13542 21103 13601 21104
rect 11970 21019 12027 21020
rect 15114 21019 15171 21020
rect 11942 21018 12038 21019
rect 15086 21018 15182 21019
rect 10737 21010 12038 21018
rect 10737 20945 10748 21010
rect 10816 20945 11970 21010
rect 10737 20942 11970 20945
rect 12027 20942 12038 21010
rect 10737 20934 12038 20942
rect 13880 21010 15182 21018
rect 13880 20945 13892 21010
rect 13960 20945 15114 21010
rect 13880 20942 15114 20945
rect 15171 20942 15182 21010
rect 13880 20934 15182 20942
rect 11970 20932 12027 20934
rect 13880 20877 13961 20934
rect 15114 20932 15171 20934
rect 2837 20858 6065 20877
rect 2837 20814 6012 20858
rect 2734 20801 6012 20814
rect 2734 20787 6065 20801
rect 9047 20798 13961 20877
rect 15359 20855 15449 21104
rect 21649 21064 21706 21108
rect 23020 21178 24660 21183
rect 23020 21173 24592 21178
rect 23079 21113 24592 21173
rect 23020 21110 24592 21113
rect 24649 21110 24660 21178
rect 23020 21104 24660 21110
rect 23020 21103 23079 21104
rect 24564 21101 24660 21104
rect 26164 21173 27804 21183
rect 26223 21169 27804 21173
rect 26223 21113 27738 21169
rect 27794 21113 27804 21169
rect 26164 21104 27804 21113
rect 26164 21103 26223 21104
rect 27738 21103 27794 21104
rect 24592 21100 24649 21101
rect 18316 21023 18373 21024
rect 21460 21023 21517 21024
rect 18288 21022 18384 21023
rect 21432 21022 21528 21023
rect 17083 21014 18384 21022
rect 17083 20949 17094 21014
rect 17162 20949 18316 21014
rect 17083 20946 18316 20949
rect 18373 20946 18384 21014
rect 17083 20938 18384 20946
rect 18750 21014 21528 21022
rect 21649 21019 21864 21064
rect 24592 21019 24649 21020
rect 27736 21019 27793 21020
rect 18750 20949 20238 21014
rect 20306 20949 21460 21014
rect 18750 20946 21460 20949
rect 21517 20946 21528 21014
rect 18750 20938 21528 20946
rect 18316 20936 18373 20938
rect 18750 20855 18829 20938
rect 21460 20936 21517 20938
rect 15359 20787 18829 20855
rect 21792 20893 21864 21019
rect 24564 21018 24660 21019
rect 27708 21018 27804 21019
rect 23359 21010 24660 21018
rect 23359 20945 23370 21010
rect 23438 20945 24592 21010
rect 23359 20942 24592 20945
rect 24649 20942 24660 21010
rect 23359 20934 24660 20942
rect 24971 21010 27804 21018
rect 24971 20945 26514 21010
rect 26582 20945 27736 21010
rect 24971 20942 27736 20945
rect 27793 20942 27804 21010
rect 24971 20934 27804 20942
rect 27948 21013 28044 21023
rect 24592 20932 24649 20934
rect 24971 20893 25046 20934
rect 27736 20932 27793 20934
rect 27948 20929 28044 20939
rect 21792 20828 25046 20893
rect 28530 20867 28598 20877
rect 28530 20801 28598 20811
rect 24684 20772 24754 20782
rect 9146 20731 9210 20741
rect 24677 20712 24684 20769
rect 27739 20769 27793 20778
rect 24754 20768 27804 20769
rect 24754 20712 27739 20768
rect 24677 20706 27739 20712
rect 27793 20706 27804 20768
rect 24677 20705 27804 20706
rect 24684 20702 24754 20705
rect 27739 20696 27793 20705
rect 9146 20662 9210 20672
rect 27951 20667 28043 20677
rect 21540 20634 21604 20641
rect 27739 20634 27793 20643
rect 21540 20633 27804 20634
rect 21540 20631 27739 20633
rect 12290 20578 12346 20588
rect 21604 20574 27739 20631
rect 21540 20571 27739 20574
rect 27793 20571 27804 20633
rect 27951 20600 28043 20610
rect 28877 20640 28966 20650
rect 21540 20570 27804 20571
rect 28877 20572 28883 20640
rect 28958 20572 28966 20640
rect 21540 20564 21604 20570
rect 27739 20561 27793 20570
rect 12290 20499 12346 20509
rect 18408 20526 18462 20536
rect 27737 20522 27791 20531
rect 27946 20522 28046 20532
rect 18462 20521 27802 20522
rect 18462 20468 27737 20521
rect 18408 20459 27737 20468
rect 27791 20459 27802 20521
rect 18408 20458 27802 20459
rect 27946 20464 27949 20466
rect 28039 20464 28046 20466
rect 27737 20449 27791 20458
rect 27946 20456 28046 20464
rect 27949 20454 28039 20456
rect 15509 20427 15571 20437
rect 27737 20397 27791 20406
rect 27575 20396 27802 20397
rect 15509 20349 15571 20359
rect 15695 20334 27737 20396
rect 27791 20334 27802 20396
rect 15695 20333 27802 20334
rect 27941 20395 28050 20405
rect 15223 20302 15292 20312
rect 15695 20298 15763 20333
rect 27737 20324 27791 20333
rect 27941 20326 28050 20336
rect 15292 20241 15763 20298
rect 15223 20234 15763 20241
rect 18687 20279 18746 20289
rect 15223 20231 15292 20234
rect 18687 20212 18746 20222
rect 21651 20203 22098 20267
rect 12084 20167 12141 20177
rect 21651 20162 21715 20203
rect 12141 20100 21715 20162
rect 12084 20098 21715 20100
rect 21813 20162 21872 20172
rect 12084 20090 12141 20098
rect 22034 20163 22098 20203
rect 27732 20163 27786 20165
rect 22034 20155 27803 20163
rect 22034 20098 27732 20155
rect 21813 20086 21872 20096
rect 27721 20093 27732 20098
rect 27786 20098 27803 20155
rect 27940 20154 28050 20164
rect 27786 20093 27797 20098
rect 27721 20092 27797 20093
rect 27732 20083 27786 20092
rect 27940 20084 28050 20094
rect 4276 20024 4352 20034
rect 4276 19956 4352 19966
rect 7420 20024 7496 20034
rect 7420 19956 7496 19966
rect 10552 20020 10628 20030
rect 8942 19951 9012 19961
rect 10552 19952 10628 19962
rect 13696 20020 13772 20030
rect 13696 19952 13772 19962
rect 16898 20024 16974 20034
rect 16898 19956 16974 19966
rect 20042 20024 20118 20034
rect 20042 19956 20118 19966
rect 23174 20020 23250 20030
rect 23174 19952 23250 19962
rect 26318 20020 26394 20030
rect 26318 19952 26394 19962
rect 27735 19934 27789 19941
rect 27682 19933 27800 19934
rect 9012 19875 24873 19924
rect 27682 19923 27735 19933
rect 8942 19870 24873 19875
rect 8942 19865 9012 19870
rect 24810 19865 24873 19870
rect 24932 19882 25005 19892
rect 24810 19762 24874 19865
rect 24932 19791 25005 19801
rect 25144 19871 27735 19923
rect 27789 19871 27800 19933
rect 25144 19870 27800 19871
rect 27943 19933 28047 19943
rect 25144 19762 25208 19870
rect 27735 19861 27789 19870
rect 27943 19862 28047 19872
rect 28779 19801 28832 19803
rect 24810 19734 25208 19762
rect 28769 19793 28839 19801
rect 28769 19724 28779 19793
rect 28832 19724 28839 19793
rect 306 19573 546 19574
rect 28769 19573 28839 19724
rect -397 19572 546 19573
rect 843 19572 2347 19573
rect 28105 19572 28839 19573
rect -397 19571 28839 19572
rect -1506 19562 28839 19571
rect -1506 19498 -1493 19562
rect -1401 19498 28839 19562
rect -1506 19492 28839 19498
rect -1506 19491 5791 19492
rect -1506 19489 -384 19491
rect 140 19490 1173 19491
rect 28051 19490 28839 19492
rect -1493 19488 -1401 19489
rect 306 19458 546 19459
rect -397 19457 546 19458
rect 843 19457 2347 19458
rect -397 19456 28732 19457
rect -1506 19447 28732 19456
rect -1506 19383 -1493 19447
rect -1401 19383 28732 19447
rect -1506 19377 28732 19383
rect -1506 19376 5791 19377
rect -1506 19374 -384 19376
rect 140 19375 1173 19376
rect 28051 19375 28732 19377
rect -1493 19373 -1401 19374
rect 28662 19365 28732 19375
rect 306 19337 546 19338
rect -397 19336 546 19337
rect 843 19336 2347 19337
rect -397 19335 28625 19336
rect -1506 19326 28625 19335
rect -1506 19262 -1493 19326
rect -1401 19262 28625 19326
rect 28662 19300 28671 19365
rect 28724 19300 28732 19365
rect 28662 19291 28732 19300
rect 28671 19290 28724 19291
rect -1506 19256 28625 19262
rect -1506 19255 5791 19256
rect -1506 19253 -384 19255
rect 140 19254 1173 19255
rect 28051 19254 28625 19256
rect 28092 19253 28625 19254
rect -1493 19252 -1401 19253
rect 306 19218 546 19219
rect -397 19217 546 19218
rect 843 19217 2347 19218
rect -397 19216 28523 19217
rect -1506 19207 28523 19216
rect -1506 19143 -1493 19207
rect -1401 19143 28523 19207
rect -1506 19137 28523 19143
rect -1506 19136 5791 19137
rect -1506 19134 -384 19136
rect 140 19135 1173 19136
rect 28051 19135 28523 19137
rect -1493 19133 -1401 19134
rect 306 19104 546 19105
rect -397 19103 546 19104
rect 843 19103 2347 19104
rect -397 19102 28421 19103
rect -1506 19093 28421 19102
rect -1506 19029 -1493 19093
rect -1401 19029 28421 19093
rect -1506 19023 28421 19029
rect -1506 19022 5791 19023
rect -1506 19020 -384 19022
rect 140 19021 1173 19022
rect 28051 19021 28421 19023
rect -1493 19019 -1401 19020
rect 306 18990 546 18991
rect -397 18989 546 18990
rect 843 18989 2347 18990
rect 28082 18989 28319 18990
rect -397 18988 28319 18989
rect -1506 18979 28319 18988
rect -1506 18915 -1493 18979
rect -1401 18915 28319 18979
rect -1506 18909 28319 18915
rect -1506 18908 5791 18909
rect -1506 18906 -384 18908
rect 140 18907 1173 18908
rect 28051 18907 28319 18909
rect -1493 18905 -1401 18906
rect 306 18875 546 18876
rect -397 18874 546 18875
rect 843 18874 2348 18875
rect -397 18873 28216 18874
rect -1505 18864 28216 18873
rect -1505 18800 -1492 18864
rect -1400 18800 28216 18864
rect -1505 18794 28216 18800
rect -1505 18793 5792 18794
rect -1505 18791 -384 18793
rect 140 18792 1173 18793
rect -1492 18790 -1400 18791
rect 306 18761 546 18762
rect -397 18760 546 18761
rect 843 18760 2348 18761
rect -1492 18759 -1400 18760
rect -397 18759 28118 18760
rect -1505 18750 28118 18759
rect -1505 18686 -1492 18750
rect -1400 18686 28118 18750
rect -1505 18680 28118 18686
rect -1505 18679 5792 18680
rect -1505 18677 -384 18679
rect 140 18678 1173 18679
rect -1492 18676 -1400 18677
rect 27826 18636 27886 18646
rect 15050 18615 27826 18625
rect 15104 18577 27826 18615
rect 27826 18567 27886 18577
rect 15050 18551 15104 18561
rect 14956 18522 15010 18532
rect 14956 18458 15010 18468
rect 4622 17048 4712 17058
rect 4622 16947 4712 16957
rect 5790 17048 5880 17058
rect 5790 16947 5880 16957
rect 6958 17048 7048 17058
rect 6958 16947 7048 16957
rect 8126 17048 8216 17058
rect 8126 16947 8216 16957
rect 9300 17046 9390 17056
rect 9300 16945 9390 16955
rect 10468 17046 10558 17056
rect 10468 16945 10558 16955
rect 11636 17046 11726 17056
rect 11636 16945 11726 16955
rect 12804 17046 12894 17056
rect 12804 16945 12894 16955
rect 14498 16839 14558 16849
rect 14498 16767 14558 16777
rect 14958 16121 15008 18458
rect 14730 16071 15008 16121
rect 14731 16040 14781 16071
rect 14716 16030 14802 16040
rect 14716 15932 14802 15942
rect 14830 15911 14915 15912
rect 14830 15902 14916 15911
rect 14915 15901 14916 15902
rect 15051 15901 15101 18551
rect 16588 18439 16642 18440
rect 27829 18439 27889 18446
rect 16585 18436 27889 18439
rect 16585 18430 27829 18436
rect 16585 18376 16588 18430
rect 16642 18376 27829 18430
rect 16585 18374 27829 18376
rect 16413 18335 16467 18345
rect 15946 16839 16006 16849
rect 15946 16767 16006 16777
rect 16413 16104 16467 18281
rect 16180 16050 16467 16104
rect 16180 16014 16234 16050
rect 16180 15950 16234 15960
rect 14916 15813 15101 15901
rect 16288 15897 16349 15907
rect 16588 15884 16642 18374
rect 27829 18364 27889 18374
rect 18049 18250 18103 18255
rect 27836 18250 27896 18256
rect 18048 18246 27896 18250
rect 18048 18245 27836 18246
rect 18048 18191 18049 18245
rect 18103 18191 27836 18245
rect 18048 18184 27836 18191
rect 17911 18151 17965 18161
rect 17444 16837 17504 16847
rect 17444 16765 17504 16775
rect 17677 16017 17731 16026
rect 17911 16017 17965 18097
rect 17677 16016 17965 16017
rect 17731 15962 17965 16016
rect 17677 15952 17731 15962
rect 16349 15830 16642 15884
rect 17788 15888 17848 15898
rect 18049 15878 18103 18184
rect 27836 18174 27896 18184
rect 19551 18064 19605 18067
rect 27836 18064 27896 18074
rect 19551 18057 27836 18064
rect 19605 18003 27836 18057
rect 19551 17995 27836 18003
rect 19551 17993 19606 17995
rect 19372 17963 19426 17973
rect 18892 16837 18952 16847
rect 18892 16765 18952 16775
rect 19125 16009 19179 16019
rect 19372 16009 19426 17909
rect 19179 15955 19426 16009
rect 19125 15945 19179 15955
rect 14915 15812 14916 15813
rect 14830 15803 14916 15812
rect 16288 15808 16349 15818
rect 17848 15824 18103 15878
rect 19238 15895 19298 15905
rect 19552 15884 19606 17993
rect 27836 17985 27896 17995
rect 21007 17877 21061 17883
rect 27848 17877 27909 17887
rect 21007 17873 27848 17877
rect 21061 17819 27848 17873
rect 21007 17814 27848 17819
rect 20879 17778 20933 17788
rect 20412 16839 20472 16849
rect 20412 16767 20472 16777
rect 20644 16014 20722 16024
rect 20879 16014 20933 17724
rect 20698 15960 20933 16014
rect 20644 15959 20933 15960
rect 20644 15950 20722 15959
rect 19298 15830 19606 15884
rect 20750 15897 20817 15907
rect 21007 15884 21061 17814
rect 27848 17804 27909 17814
rect 22460 17687 22514 17697
rect 27851 17686 27922 17696
rect 22514 17633 27851 17686
rect 22460 17614 27851 17633
rect 22329 17592 22383 17602
rect 21860 16839 21920 16849
rect 21860 16767 21920 16777
rect 22094 16011 22148 16021
rect 22329 16011 22383 17538
rect 22148 15957 22383 16011
rect 22094 15947 22148 15957
rect 20817 15830 21061 15884
rect 22202 15891 22266 15901
rect 22460 15879 22514 17614
rect 27851 17604 27922 17614
rect 23905 17501 23959 17511
rect 23795 17416 23849 17418
rect 23795 17408 23850 17416
rect 23849 17354 23850 17408
rect 23358 16837 23418 16847
rect 23358 16765 23418 16775
rect 23588 16012 23642 16022
rect 23795 16012 23850 17354
rect 23642 15958 23850 16012
rect 23588 15948 23642 15958
rect 17788 15810 17848 15820
rect 19238 15810 19298 15820
rect 20750 15809 20817 15819
rect 22266 15825 22514 15879
rect 23692 15899 23768 15909
rect 23905 15882 23959 17447
rect 27316 17210 27430 17211
rect 27316 17209 27647 17210
rect 27851 17209 27905 17219
rect 27316 17154 27851 17209
rect 24806 16837 24866 16847
rect 24806 16765 24866 16775
rect 25630 16181 25701 16191
rect 25630 16112 25701 16122
rect 25346 16085 25415 16095
rect 25346 16011 25415 16021
rect 27316 15882 27395 17154
rect 27851 17144 27905 17154
rect 27800 16802 27858 16812
rect 27800 16736 27858 16746
rect 28052 16807 28118 18680
rect 28149 17216 28216 18794
rect 28249 17675 28319 18907
rect 28351 17876 28421 19021
rect 28453 18064 28523 19135
rect 28555 18252 28625 19253
rect 28555 18177 28564 18252
rect 28616 18177 28625 18252
rect 28555 18170 28625 18177
rect 28564 18167 28616 18170
rect 28453 17987 28461 18064
rect 28515 17987 28523 18064
rect 28453 17980 28523 17987
rect 28461 17977 28515 17980
rect 28351 17806 28360 17876
rect 28414 17806 28421 17876
rect 28351 17798 28421 17806
rect 28360 17796 28414 17798
rect 28249 17600 28258 17675
rect 28311 17600 28319 17675
rect 28249 17573 28319 17600
rect 28149 17152 28157 17216
rect 28211 17152 28216 17216
rect 28149 17144 28216 17152
rect 28157 17142 28211 17144
rect 28052 16721 28118 16731
rect 23898 15881 27395 15882
rect 23768 15826 27395 15881
rect 22202 15807 22266 15817
rect 23898 15825 27395 15826
rect 14830 15802 14915 15803
rect 23692 15802 23768 15812
rect 5087 15721 5177 15731
rect 5087 15620 5177 15630
rect 6255 15721 6345 15731
rect 6255 15620 6345 15630
rect 7423 15721 7513 15731
rect 7423 15620 7513 15630
rect 8591 15721 8681 15731
rect 8591 15620 8681 15630
rect 9765 15719 9855 15729
rect 9765 15618 9855 15628
rect 10933 15719 11023 15729
rect 10933 15618 11023 15628
rect 12101 15719 12191 15729
rect 12101 15618 12191 15628
rect 13269 15719 13359 15729
rect 14274 15643 14336 15645
rect 15722 15643 15784 15645
rect 20188 15643 20250 15645
rect 21636 15643 21698 15645
rect 13269 15618 13359 15628
rect 14272 15635 14336 15643
rect 14272 15633 14274 15635
rect 14272 15561 14336 15571
rect 15720 15635 15784 15643
rect 17220 15641 17282 15643
rect 18668 15641 18730 15643
rect 15720 15633 15722 15635
rect 15720 15561 15784 15571
rect 17218 15633 17282 15641
rect 17218 15631 17220 15633
rect 17218 15559 17282 15569
rect 18666 15633 18730 15641
rect 18666 15631 18668 15633
rect 18666 15559 18730 15569
rect 20186 15635 20250 15643
rect 20186 15633 20188 15635
rect 20186 15561 20250 15571
rect 21634 15635 21698 15643
rect 23134 15641 23196 15643
rect 24582 15641 24644 15643
rect 21634 15633 21636 15635
rect 21634 15561 21698 15571
rect 23132 15633 23196 15641
rect 23132 15631 23134 15633
rect 23132 15559 23196 15569
rect 24580 15633 24644 15641
rect 24580 15631 24582 15633
rect 24580 15559 24644 15569
rect 1770 15130 1870 15140
rect 1770 15028 1870 15038
rect 4914 15130 5014 15140
rect 4914 15028 5014 15038
rect 8046 15126 8146 15136
rect 8046 15024 8146 15034
rect 11190 15126 11290 15136
rect 11190 15024 11290 15034
rect 14392 15130 14492 15140
rect 14392 15028 14492 15038
rect 17536 15130 17636 15140
rect 17536 15028 17636 15038
rect 20668 15126 20768 15136
rect 20668 15024 20768 15034
rect 23812 15126 23912 15136
rect 23812 15024 23912 15034
rect 2923 14169 3016 14171
rect 6067 14169 6160 14171
rect 15545 14169 15638 14171
rect 18689 14169 18782 14171
rect 1841 14165 3260 14169
rect 4985 14165 6404 14169
rect 9199 14165 9292 14167
rect 12343 14165 12436 14167
rect 14463 14165 15882 14169
rect 17607 14165 19026 14169
rect 21821 14165 21914 14167
rect 24965 14165 25058 14167
rect 1841 14159 25927 14165
rect 1841 14097 1850 14159
rect 1920 14097 2934 14159
rect 1841 14096 2934 14097
rect 3005 14097 4994 14159
rect 5064 14097 6078 14159
rect 3005 14096 6078 14097
rect 6149 14155 14472 14159
rect 6149 14096 8126 14155
rect 1841 14093 8126 14096
rect 8196 14093 9210 14155
rect 1841 14092 9210 14093
rect 9281 14093 11270 14155
rect 11340 14093 12354 14155
rect 9281 14092 12354 14093
rect 12425 14097 14472 14155
rect 14542 14097 15556 14159
rect 12425 14096 15556 14097
rect 15627 14097 17616 14159
rect 17686 14097 18700 14159
rect 15627 14096 18700 14097
rect 18771 14158 25927 14159
rect 18771 14155 25828 14158
rect 18771 14096 20748 14155
rect 12425 14093 20748 14096
rect 20818 14093 21832 14155
rect 12425 14092 21832 14093
rect 21903 14093 23892 14155
rect 23962 14093 24976 14155
rect 21903 14092 24976 14093
rect 25047 14092 25828 14155
rect 1841 14081 25828 14092
rect 25911 14081 25927 14158
rect 25828 14060 25911 14070
rect 1620 14044 3260 14049
rect 1620 14039 3192 14044
rect 1679 13979 3192 14039
rect 1620 13976 3192 13979
rect 3249 13976 3260 14044
rect 1620 13970 3260 13976
rect 1620 13969 1679 13970
rect 3164 13967 3260 13970
rect 4764 14044 6404 14049
rect 9440 14045 9536 14048
rect 12584 14045 12680 14048
rect 4764 14039 6336 14044
rect 4823 13979 6336 14039
rect 4764 13976 6336 13979
rect 6393 13976 6404 14044
rect 4764 13970 6404 13976
rect 4764 13969 4823 13970
rect 6308 13967 6404 13970
rect 7896 14040 9536 14045
rect 7896 14035 9468 14040
rect 7955 13975 9468 14035
rect 7896 13972 9468 13975
rect 9525 13972 9536 14040
rect 3192 13966 3249 13967
rect 6336 13966 6393 13967
rect 7896 13966 9536 13972
rect 7896 13965 7955 13966
rect 9440 13963 9536 13966
rect 11040 14040 12680 14045
rect 11040 14035 12612 14040
rect 11099 13975 12612 14035
rect 11040 13972 12612 13975
rect 12669 13972 12680 14040
rect 11040 13966 12680 13972
rect 14242 14044 15882 14049
rect 14242 14039 15814 14044
rect 14301 13979 15814 14039
rect 14242 13976 15814 13979
rect 15871 13976 15882 14044
rect 14242 13970 15882 13976
rect 14242 13969 14301 13970
rect 15786 13967 15882 13970
rect 17386 14044 19026 14049
rect 22090 14048 22147 14050
rect 22062 14045 22158 14048
rect 25206 14045 25302 14048
rect 17386 14039 18958 14044
rect 17445 13979 18958 14039
rect 17386 13976 18958 13979
rect 19015 13976 19026 14044
rect 17386 13970 19026 13976
rect 20518 14040 22158 14045
rect 20518 14035 22090 14040
rect 20577 13975 22090 14035
rect 20518 13972 22090 13975
rect 22147 13972 22158 14040
rect 17386 13969 17445 13970
rect 15814 13966 15871 13967
rect 20518 13966 22158 13972
rect 11040 13965 11099 13966
rect 12584 13963 12680 13966
rect 20518 13965 20577 13966
rect 22062 13963 22158 13966
rect 23662 14040 25302 14045
rect 23662 14035 25234 14040
rect 23721 13975 25234 14035
rect 23662 13972 25234 13975
rect 25291 13972 25302 14040
rect 23662 13966 25302 13972
rect 23662 13965 23721 13966
rect 25206 13963 25302 13966
rect 9468 13962 9525 13963
rect 12612 13962 12669 13963
rect 22090 13962 22147 13963
rect 25234 13962 25291 13963
rect 3192 13885 3249 13886
rect 6336 13885 6393 13886
rect 18958 13885 19015 13886
rect 3164 13884 3260 13885
rect 6308 13884 6404 13885
rect 18930 13884 19026 13885
rect 1959 13876 3260 13884
rect 1959 13811 1970 13876
rect 2038 13811 3192 13876
rect 1959 13808 3192 13811
rect 3249 13808 3260 13876
rect 1959 13800 3260 13808
rect 5103 13876 6404 13884
rect 9468 13881 9525 13882
rect 9440 13880 9536 13881
rect 5103 13811 5114 13876
rect 5182 13811 6336 13876
rect 5103 13808 6336 13811
rect 6393 13808 6404 13876
rect 5103 13800 6404 13808
rect 8235 13872 9536 13880
rect 8235 13807 8246 13872
rect 8314 13807 9468 13872
rect 8235 13804 9468 13807
rect 9525 13804 9536 13872
rect 3192 13798 3249 13800
rect 6336 13798 6393 13800
rect 8235 13796 9536 13804
rect 17725 13876 19026 13884
rect 22090 13881 22147 13882
rect 25234 13881 25291 13882
rect 22062 13880 22158 13881
rect 25206 13880 25302 13881
rect 17725 13811 17736 13876
rect 17804 13811 18958 13876
rect 17725 13808 18958 13811
rect 19015 13808 19026 13876
rect 17725 13800 19026 13808
rect 20857 13872 22158 13880
rect 20857 13807 20868 13872
rect 20936 13807 22090 13872
rect 20857 13804 22090 13807
rect 22147 13804 22158 13872
rect 18958 13798 19015 13800
rect 20857 13796 22158 13804
rect 24001 13872 25302 13880
rect 24001 13807 24012 13872
rect 24080 13807 25234 13872
rect 24001 13804 25234 13807
rect 25291 13804 25302 13872
rect 24001 13796 25302 13804
rect 9468 13794 9525 13796
rect 22090 13794 22147 13796
rect 25234 13794 25291 13796
rect 1774 12886 1850 12896
rect 1774 12818 1850 12828
rect 4918 12886 4994 12896
rect 4918 12818 4994 12828
rect 8050 12882 8126 12892
rect 8050 12814 8126 12824
rect 11194 12882 11270 12892
rect 11194 12814 11270 12824
rect 14396 12886 14472 12896
rect 14396 12818 14472 12828
rect 17540 12886 17616 12896
rect 17540 12818 17616 12828
rect 20672 12882 20748 12892
rect 20672 12814 20748 12824
rect 23816 12882 23892 12892
rect 23816 12814 23892 12824
rect 1770 12396 1870 12406
rect 1770 12294 1870 12304
rect 4914 12396 5014 12406
rect 4914 12294 5014 12304
rect 8046 12392 8146 12402
rect 8046 12290 8146 12300
rect 11190 12392 11290 12402
rect 11190 12290 11290 12300
rect 14392 12396 14492 12406
rect 14392 12294 14492 12304
rect 17536 12396 17636 12406
rect 17536 12294 17636 12304
rect 20668 12392 20768 12402
rect 20668 12290 20768 12300
rect 23812 12392 23912 12402
rect 23812 12290 23912 12300
rect 2923 11435 3016 11437
rect 6067 11435 6160 11437
rect 15545 11435 15638 11437
rect 1841 11434 3257 11435
rect 4985 11434 6401 11435
rect 14463 11434 19023 11435
rect 1841 11431 8179 11434
rect 9199 11431 9292 11433
rect 12343 11431 12436 11433
rect 14463 11431 19026 11434
rect 21821 11431 21914 11433
rect 24965 11431 25058 11433
rect 28877 11432 28966 20572
rect 32913 20318 33097 20328
rect 27778 11431 28966 11432
rect 1841 11430 9533 11431
rect 11261 11430 12677 11431
rect 14463 11430 28966 11431
rect 1841 11429 9536 11430
rect 11261 11429 28966 11430
rect 1841 11425 28966 11429
rect -307 11361 241 11377
rect -307 11337 80 11361
rect -310 11232 80 11337
rect 191 11232 241 11361
rect 1841 11363 1850 11425
rect 1920 11363 2934 11425
rect 1841 11362 2934 11363
rect 3005 11363 4994 11425
rect 5064 11363 6078 11425
rect 3005 11362 6078 11363
rect 6149 11422 14472 11425
rect 6149 11421 9468 11422
rect 6149 11362 8126 11421
rect 1841 11359 8126 11362
rect 8196 11359 9210 11421
rect 1841 11358 9210 11359
rect 9281 11358 9468 11421
rect 1841 11354 9468 11358
rect 9525 11421 14472 11422
rect 9525 11359 11270 11421
rect 11340 11359 12354 11421
rect 9525 11358 12354 11359
rect 12425 11363 14472 11421
rect 14542 11363 15556 11425
rect 12425 11362 15556 11363
rect 15627 11363 17616 11425
rect 17686 11363 18700 11425
rect 15627 11362 18700 11363
rect 18771 11421 28966 11425
rect 18771 11362 20748 11421
rect 12425 11359 20748 11362
rect 20818 11359 21832 11421
rect 12425 11358 21832 11359
rect 21903 11359 23892 11421
rect 23962 11359 24976 11421
rect 21903 11358 24976 11359
rect 25047 11358 28966 11421
rect 9525 11354 28966 11358
rect 1841 11351 28966 11354
rect 6372 11347 12680 11351
rect 18948 11350 28966 11351
rect 18958 11348 28966 11350
rect 18995 11347 28966 11348
rect 25392 11346 28966 11347
rect 27778 11345 28966 11346
rect 28877 11344 28966 11345
rect 29011 20222 29100 20239
rect 29011 20154 29020 20222
rect 29090 20154 29100 20222
rect 3192 11318 3249 11320
rect 15814 11318 15871 11320
rect 3164 11315 3260 11318
rect 1620 11310 3260 11315
rect 1620 11305 3192 11310
rect 1679 11245 3192 11305
rect 1620 11242 3192 11245
rect 3249 11242 3260 11310
rect 1620 11236 3260 11242
rect 1620 11235 1679 11236
rect 3164 11233 3260 11236
rect 4764 11310 6404 11315
rect 9468 11314 9525 11316
rect 15786 11315 15882 11318
rect 9440 11311 9536 11314
rect 12584 11311 12680 11314
rect 4764 11305 6336 11310
rect 4823 11245 6336 11305
rect 4764 11242 6336 11245
rect 6393 11242 6404 11310
rect 4764 11236 6404 11242
rect 4764 11235 4823 11236
rect 6308 11233 6404 11236
rect 7896 11306 9536 11311
rect 7896 11301 9468 11306
rect 7955 11241 9468 11301
rect 7896 11238 9468 11241
rect 9525 11238 9536 11306
rect 3192 11232 3249 11233
rect 6336 11232 6393 11233
rect 7896 11232 9536 11238
rect -310 11220 241 11232
rect 7896 11231 7955 11232
rect 9440 11229 9536 11232
rect 11040 11306 12680 11311
rect 11040 11301 12612 11306
rect 11099 11241 12612 11301
rect 11040 11238 12612 11241
rect 12669 11238 12680 11306
rect 11040 11232 12680 11238
rect 14242 11310 15882 11315
rect 14242 11305 15814 11310
rect 14301 11245 15814 11305
rect 14242 11242 15814 11245
rect 15871 11242 15882 11310
rect 14242 11236 15882 11242
rect 14242 11235 14301 11236
rect 15786 11233 15882 11236
rect 17386 11310 19026 11315
rect 22090 11314 22147 11316
rect 25234 11314 25291 11316
rect 22062 11311 22158 11314
rect 25206 11311 25302 11314
rect 17386 11305 18958 11310
rect 17445 11245 18958 11305
rect 17386 11242 18958 11245
rect 19015 11242 19026 11310
rect 17386 11236 19026 11242
rect 17386 11235 17445 11236
rect 18930 11233 19026 11236
rect 20518 11306 22158 11311
rect 20518 11301 22090 11306
rect 20577 11241 22090 11301
rect 20518 11238 22090 11241
rect 22147 11238 22158 11306
rect 15814 11232 15871 11233
rect 18958 11232 19015 11233
rect 20518 11232 22158 11238
rect 11040 11231 11099 11232
rect 12584 11229 12680 11232
rect 20518 11231 20577 11232
rect 22062 11229 22158 11232
rect 23662 11306 25302 11311
rect 23662 11301 25234 11306
rect 23721 11241 25234 11301
rect 23662 11238 25234 11241
rect 25291 11238 25302 11306
rect 23662 11232 25302 11238
rect 23662 11231 23721 11232
rect 25206 11229 25302 11232
rect 9468 11228 9525 11229
rect 12612 11228 12669 11229
rect 22090 11228 22147 11229
rect 25234 11228 25291 11229
rect -570 10936 -404 10951
rect -570 10879 -547 10936
rect -425 10879 -404 10936
rect -570 10806 -404 10879
rect -783 10753 -661 10754
rect -806 10744 -640 10753
rect -806 10687 -783 10744
rect -661 10687 -640 10744
rect -1068 10516 -900 10540
rect -1068 10459 -1048 10516
rect -926 10459 -900 10516
rect -1278 10331 -1112 10348
rect -1278 10274 -1255 10331
rect -1133 10274 -1112 10331
rect -1540 9984 -1372 10006
rect -1540 9927 -1515 9984
rect -1393 9927 -1372 9984
rect -1749 9815 -1583 9834
rect -1749 9758 -1730 9815
rect -1608 9758 -1583 9815
rect -2011 9455 -1843 9481
rect -2011 9398 -1991 9455
rect -1869 9398 -1843 9455
rect -2011 3408 -1843 9398
rect -2011 3349 -1993 3408
rect -1872 3349 -1843 3408
rect -2011 3336 -1843 3349
rect -1749 3282 -1583 9758
rect -1749 3217 -1727 3282
rect -1616 3217 -1583 3282
rect -1749 3204 -1583 3217
rect -1540 3173 -1372 9927
rect -1540 3110 -1520 3173
rect -1404 3110 -1372 3173
rect -1540 3087 -1372 3110
rect -1278 3060 -1112 10274
rect -1278 2993 -1258 3060
rect -1137 2993 -1112 3060
rect -1278 2974 -1112 2993
rect -1068 2945 -900 10459
rect -1068 2863 -1049 2945
rect -925 2863 -900 2945
rect -1068 2846 -900 2863
rect -806 2840 -640 10687
rect -806 2757 -791 2840
rect -659 2757 -640 2840
rect -806 2736 -640 2757
rect -572 2722 -404 10806
rect -572 2637 -545 2722
rect -428 2637 -404 2722
rect -572 2615 -404 2637
rect -310 1165 -144 11220
rect 3192 11151 3249 11152
rect 6336 11151 6393 11152
rect 15814 11151 15871 11152
rect 18958 11151 19015 11152
rect 3164 11150 3260 11151
rect 6308 11150 6404 11151
rect 15786 11150 15882 11151
rect 18930 11150 19026 11151
rect 1959 11142 3260 11150
rect 1959 11077 1970 11142
rect 2038 11077 3192 11142
rect 1959 11074 3192 11077
rect 3249 11074 3260 11142
rect 1959 11066 3260 11074
rect 5103 11142 6404 11150
rect 9468 11147 9525 11148
rect 12612 11147 12669 11148
rect 9440 11146 9536 11147
rect 12584 11146 12680 11147
rect 5103 11077 5114 11142
rect 5182 11077 6336 11142
rect 5103 11074 6336 11077
rect 6393 11074 6404 11142
rect 5103 11066 6404 11074
rect 8235 11138 9536 11146
rect 8235 11073 8246 11138
rect 8314 11073 9468 11138
rect 8235 11070 9468 11073
rect 9525 11070 9536 11138
rect 3192 11064 3249 11066
rect 6336 11064 6393 11066
rect 8235 11062 9536 11070
rect 11379 11138 12680 11146
rect 11379 11073 11390 11138
rect 11458 11073 12612 11138
rect 11379 11070 12612 11073
rect 12669 11070 12680 11138
rect 11379 11062 12680 11070
rect 14581 11142 15882 11150
rect 14581 11077 14592 11142
rect 14660 11077 15814 11142
rect 14581 11074 15814 11077
rect 15871 11074 15882 11142
rect 14581 11066 15882 11074
rect 17725 11142 19026 11150
rect 22090 11147 22147 11148
rect 25234 11147 25291 11148
rect 22062 11146 22158 11147
rect 25206 11146 25302 11147
rect 17725 11077 17736 11142
rect 17804 11077 18958 11142
rect 17725 11074 18958 11077
rect 19015 11074 19026 11142
rect 17725 11066 19026 11074
rect 20857 11138 22158 11146
rect 20857 11073 20868 11138
rect 20936 11073 22090 11138
rect 20857 11070 22090 11073
rect 22147 11070 22158 11138
rect 15814 11064 15871 11066
rect 18958 11064 19015 11066
rect 20857 11062 22158 11070
rect 24001 11138 25302 11146
rect 24001 11073 24012 11138
rect 24080 11073 25234 11138
rect 24001 11070 25234 11073
rect 25291 11070 25302 11138
rect 25837 11106 25904 11109
rect 29011 11107 29100 20154
rect 32913 20147 33097 20157
rect 38134 18434 38293 25093
rect 42512 24884 42665 24894
rect 40030 24830 40183 24840
rect 43659 24884 43812 24894
rect 42924 24789 42980 24799
rect 42512 24745 42665 24755
rect 40030 24691 40183 24701
rect 42799 24723 42924 24785
rect 42980 24723 42981 24785
rect 49025 24881 49178 24891
rect 43659 24745 43812 24755
rect 46543 24827 46696 24837
rect 41794 24674 41860 24677
rect 40868 24667 41860 24674
rect 40868 24601 41794 24667
rect 40301 23638 40311 23791
rect 40440 23638 40450 23791
rect 38827 23203 39040 23204
rect 39308 23203 39424 23204
rect 38827 23193 39424 23203
rect 38827 23181 39307 23193
rect 38827 23078 38849 23181
rect 38991 23087 39307 23181
rect 39419 23087 39424 23193
rect 38991 23078 39424 23087
rect 38827 23061 39424 23078
rect 40044 23180 40197 23190
rect 38827 23060 39040 23061
rect 40044 23041 40197 23051
rect 38809 22082 38947 22086
rect 38803 22081 39052 22082
rect 39590 22081 39708 22084
rect 38803 22076 39708 22081
rect 38803 21950 38809 22076
rect 38947 22074 39708 22076
rect 38947 21956 39590 22074
rect 40315 21988 40325 22141
rect 40454 21988 40464 22141
rect 38947 21950 39708 21956
rect 38803 21946 39708 21950
rect 38809 21940 38947 21946
rect 39077 21702 39192 21712
rect 39077 21595 39192 21605
rect 39587 20295 39703 21946
rect 40039 21576 40192 21586
rect 40039 21437 40192 21447
rect 40637 20818 40700 20824
rect 40868 20818 40936 24601
rect 41794 24591 41860 24601
rect 42799 24062 42859 24723
rect 42924 24713 42980 24723
rect 50172 24881 50325 24891
rect 49437 24786 49493 24796
rect 49025 24742 49178 24752
rect 46543 24688 46696 24698
rect 49312 24720 49437 24782
rect 49493 24720 49494 24782
rect 55559 24876 55712 24886
rect 50172 24742 50325 24752
rect 53077 24822 53230 24832
rect 48307 24671 48373 24674
rect 42721 24061 42859 24062
rect 42459 24051 42859 24061
rect 42459 23954 42460 24051
rect 42559 23954 42859 24051
rect 47381 24664 48373 24671
rect 47381 24598 48307 24664
rect 43616 24040 43681 24041
rect 44711 24040 44779 24050
rect 43615 24031 44711 24040
rect 43615 23977 43616 24031
rect 43681 23977 44711 24031
rect 43615 23966 44711 23977
rect 44711 23955 44779 23965
rect 42459 23946 42859 23954
rect 42459 23942 42768 23946
rect 45007 23777 45140 23778
rect 45007 23751 45450 23777
rect 45007 23607 45190 23751
rect 45426 23607 45450 23751
rect 46814 23635 46824 23788
rect 46953 23635 46963 23788
rect 45007 23583 45450 23607
rect 41859 23483 42012 23493
rect 41859 23344 42012 23354
rect 43001 23481 43154 23491
rect 43001 23342 43154 23352
rect 41857 22837 42010 22847
rect 41857 22698 42010 22708
rect 43755 22837 43908 22847
rect 43755 22698 43908 22708
rect 42498 21866 42576 21876
rect 42498 21770 42576 21780
rect 40632 20814 40936 20818
rect 40632 20762 40637 20814
rect 40700 20762 40936 20814
rect 40632 20756 40936 20762
rect 40637 20752 40700 20756
rect 40310 20384 40320 20537
rect 40449 20384 40459 20537
rect 41803 20440 41956 20450
rect 41803 20301 41956 20311
rect 43701 20440 43854 20450
rect 43701 20301 43854 20311
rect 39587 20285 39704 20295
rect 39587 20179 39592 20285
rect 39587 20169 39704 20179
rect 39587 20168 39703 20169
rect 45007 19985 45171 23583
rect 45253 23207 45533 23230
rect 45253 23083 45281 23207
rect 45510 23200 45533 23207
rect 45821 23200 45937 23201
rect 45510 23190 45937 23200
rect 45510 23084 45820 23190
rect 45932 23084 45937 23190
rect 45510 23083 45937 23084
rect 45253 23058 45937 23083
rect 46557 23177 46710 23187
rect 45253 23057 45533 23058
rect 46557 23038 46710 23048
rect 45313 22079 45478 22089
rect 45313 22078 45481 22079
rect 46103 22078 46221 22081
rect 45313 22071 46221 22078
rect 45313 22061 46103 22071
rect 45313 21955 45325 22061
rect 45437 22059 46103 22061
rect 45313 21953 45331 21955
rect 45443 21953 46103 22059
rect 46828 21985 46838 22138
rect 46967 21985 46977 22138
rect 45313 21946 46221 21953
rect 45319 21944 46221 21946
rect 45356 21943 46221 21944
rect 45590 21699 45705 21709
rect 45590 21592 45705 21602
rect 46100 20292 46216 21943
rect 46552 21573 46705 21583
rect 46552 21434 46705 21444
rect 47150 20815 47213 20821
rect 47381 20815 47449 24598
rect 48307 24588 48373 24598
rect 49312 24059 49372 24720
rect 49437 24710 49493 24720
rect 56706 24876 56859 24886
rect 55971 24781 56027 24791
rect 55559 24737 55712 24747
rect 53077 24683 53230 24693
rect 55846 24715 55971 24777
rect 56027 24715 56028 24777
rect 62117 24880 62270 24890
rect 56706 24737 56859 24747
rect 59635 24826 59788 24836
rect 54841 24666 54907 24669
rect 49234 24058 49372 24059
rect 48972 24048 49372 24058
rect 48972 23951 48973 24048
rect 49072 23951 49372 24048
rect 53915 24659 54907 24666
rect 53915 24593 54841 24659
rect 50129 24037 50194 24038
rect 51224 24037 51292 24047
rect 50128 24028 51224 24037
rect 50128 23974 50129 24028
rect 50194 23974 51224 24028
rect 50128 23963 51224 23974
rect 51224 23952 51292 23962
rect 48972 23943 49372 23951
rect 48972 23939 49281 23943
rect 51524 23758 51979 23777
rect 51524 23601 51727 23758
rect 51960 23601 51979 23758
rect 53348 23630 53358 23783
rect 53487 23630 53497 23783
rect 51524 23578 51979 23601
rect 48372 23480 48525 23490
rect 48372 23341 48525 23351
rect 49514 23478 49667 23488
rect 49514 23339 49667 23349
rect 48370 22834 48523 22844
rect 48370 22695 48523 22705
rect 50268 22834 50421 22844
rect 50268 22695 50421 22705
rect 49011 21863 49089 21873
rect 49011 21767 49089 21777
rect 47145 20811 47449 20815
rect 47145 20759 47150 20811
rect 47213 20759 47449 20811
rect 47145 20753 47449 20759
rect 47150 20749 47213 20753
rect 46823 20381 46833 20534
rect 46962 20381 46972 20534
rect 48316 20437 48469 20447
rect 48316 20298 48469 20308
rect 50214 20437 50367 20447
rect 50214 20298 50367 20308
rect 46100 20282 46217 20292
rect 46100 20176 46105 20282
rect 46100 20166 46217 20176
rect 46100 20165 46216 20166
rect 45007 19907 45026 19985
rect 45154 19907 45171 19985
rect 45007 19895 45171 19907
rect 51524 19834 51671 23578
rect 51907 23577 51979 23578
rect 51863 23230 52089 23231
rect 51814 23213 52089 23230
rect 51814 23073 51840 23213
rect 52058 23195 52089 23213
rect 52355 23195 52471 23196
rect 52058 23185 52471 23195
rect 52058 23079 52354 23185
rect 52466 23079 52471 23185
rect 52058 23073 52471 23079
rect 51814 23053 52471 23073
rect 53091 23172 53244 23182
rect 51814 23052 52073 23053
rect 53091 23033 53244 23043
rect 51847 22074 52012 22084
rect 51847 22073 52015 22074
rect 52637 22073 52755 22076
rect 51847 22066 52755 22073
rect 51847 22056 52637 22066
rect 51847 21950 51859 22056
rect 51971 22054 52637 22056
rect 51847 21948 51865 21950
rect 51977 21948 52637 22054
rect 53362 21980 53372 22133
rect 53501 21980 53511 22133
rect 51847 21941 52755 21948
rect 51853 21939 52755 21941
rect 51890 21938 52755 21939
rect 52124 21694 52239 21704
rect 52124 21587 52239 21597
rect 52634 20287 52750 21938
rect 53086 21568 53239 21578
rect 53086 21429 53239 21439
rect 53684 20810 53747 20816
rect 53915 20810 53983 24593
rect 54841 24583 54907 24593
rect 55846 24054 55906 24715
rect 55971 24705 56027 24715
rect 63264 24880 63417 24890
rect 62529 24785 62585 24795
rect 62117 24741 62270 24751
rect 59635 24687 59788 24697
rect 62404 24719 62529 24781
rect 62585 24719 62586 24781
rect 63264 24741 63417 24751
rect 61399 24670 61465 24673
rect 55768 24053 55906 24054
rect 55506 24043 55906 24053
rect 55506 23946 55507 24043
rect 55606 23946 55906 24043
rect 60473 24663 61465 24670
rect 60473 24597 61399 24663
rect 56663 24032 56728 24033
rect 57758 24032 57826 24042
rect 56662 24023 57758 24032
rect 56662 23969 56663 24023
rect 56728 23969 57758 24023
rect 56662 23958 57758 23969
rect 57758 23947 57826 23957
rect 55506 23938 55906 23946
rect 55506 23934 55815 23938
rect 58450 23778 58544 23779
rect 58112 23759 58544 23778
rect 58112 23596 58287 23759
rect 58534 23596 58544 23759
rect 59906 23634 59916 23787
rect 60045 23634 60055 23787
rect 58112 23582 58544 23596
rect 58112 23581 58526 23582
rect 54906 23475 55059 23485
rect 54906 23336 55059 23346
rect 56048 23473 56201 23483
rect 56048 23334 56201 23344
rect 54904 22829 55057 22839
rect 54904 22690 55057 22700
rect 56802 22829 56955 22839
rect 56802 22690 56955 22700
rect 55545 21858 55623 21868
rect 55545 21762 55623 21772
rect 53679 20806 53983 20810
rect 53679 20754 53684 20806
rect 53747 20754 53983 20806
rect 53679 20748 53983 20754
rect 53684 20744 53747 20748
rect 53357 20376 53367 20529
rect 53496 20376 53506 20529
rect 54850 20432 55003 20442
rect 54850 20293 55003 20303
rect 56748 20432 56901 20442
rect 56748 20293 56901 20303
rect 52634 20277 52751 20287
rect 52634 20171 52639 20277
rect 52634 20161 52751 20171
rect 52634 20160 52750 20161
rect 51524 19723 51539 19834
rect 51650 19723 51671 19834
rect 51524 19710 51671 19723
rect 58112 19651 58271 23581
rect 58346 23215 58642 23235
rect 58346 23070 58364 23215
rect 58616 23199 58642 23215
rect 58913 23199 59029 23200
rect 58616 23189 59029 23199
rect 58616 23083 58912 23189
rect 59024 23083 59029 23189
rect 58616 23070 59029 23083
rect 58346 23057 59029 23070
rect 59649 23176 59802 23186
rect 59649 23037 59802 23047
rect 58405 22078 58570 22088
rect 58405 22077 58573 22078
rect 59195 22077 59313 22080
rect 58405 22070 59313 22077
rect 58405 22060 59195 22070
rect 58405 21954 58417 22060
rect 58529 22058 59195 22060
rect 58405 21952 58423 21954
rect 58535 21952 59195 22058
rect 59920 21984 59930 22137
rect 60059 21984 60069 22137
rect 58405 21945 59313 21952
rect 58411 21943 59313 21945
rect 58448 21942 59313 21943
rect 58682 21698 58797 21708
rect 58682 21591 58797 21601
rect 59192 20291 59308 21942
rect 59644 21572 59797 21582
rect 59644 21433 59797 21443
rect 60242 20814 60305 20820
rect 60473 20814 60541 24597
rect 61399 24587 61465 24597
rect 62404 24058 62464 24719
rect 62529 24709 62585 24719
rect 62326 24057 62464 24058
rect 62064 24047 62464 24057
rect 62064 23950 62065 24047
rect 62164 23950 62464 24047
rect 63221 24036 63286 24037
rect 64316 24036 64384 24046
rect 63220 24027 64316 24036
rect 63220 23973 63221 24027
rect 63286 23973 64316 24027
rect 63220 23962 64316 23973
rect 64316 23951 64384 23961
rect 62064 23942 62464 23950
rect 62064 23938 62373 23942
rect 61464 23479 61617 23489
rect 61464 23340 61617 23350
rect 62606 23477 62759 23487
rect 62606 23338 62759 23348
rect 61462 22833 61615 22843
rect 61462 22694 61615 22704
rect 63360 22833 63513 22843
rect 63360 22694 63513 22704
rect 68767 22207 71240 22208
rect 68767 22120 71286 22207
rect 71319 22204 71404 22215
rect 71486 22204 71571 22215
rect 71317 22147 71327 22204
rect 71395 22147 71405 22204
rect 71485 22147 71495 22204
rect 71563 22147 71573 22204
rect 62103 21862 62181 21872
rect 62103 21766 62181 21776
rect 60237 20810 60541 20814
rect 60237 20758 60242 20810
rect 60305 20758 60541 20810
rect 60237 20752 60541 20758
rect 60242 20748 60305 20752
rect 59915 20380 59925 20533
rect 60054 20380 60064 20533
rect 61408 20436 61561 20446
rect 61408 20297 61561 20307
rect 63306 20436 63459 20446
rect 63306 20297 63459 20307
rect 59192 20281 59309 20291
rect 59192 20175 59197 20281
rect 59192 20165 59309 20175
rect 59192 20164 59308 20165
rect 58112 19533 58127 19651
rect 58261 19533 58271 19651
rect 58112 19519 58271 19533
rect 39608 19276 39761 19286
rect 40755 19276 40908 19286
rect 40440 19181 40496 19191
rect 39608 19137 39761 19147
rect 40439 19115 40440 19177
rect 40496 19115 40621 19177
rect 46166 19272 46319 19282
rect 40755 19137 40908 19147
rect 43237 19222 43390 19232
rect 40440 19105 40496 19115
rect 40561 18454 40621 19115
rect 47313 19272 47466 19282
rect 46998 19177 47054 19187
rect 46166 19133 46319 19143
rect 46997 19111 46998 19173
rect 47054 19111 47179 19173
rect 52700 19277 52853 19287
rect 47313 19133 47466 19143
rect 49795 19218 49948 19228
rect 46998 19101 47054 19111
rect 43237 19083 43390 19093
rect 41560 19066 41626 19069
rect 41560 19059 42552 19066
rect 41626 18993 42552 19059
rect 41560 18983 41626 18993
rect 40561 18453 40699 18454
rect 40561 18443 40961 18453
rect 38134 18432 38885 18434
rect 39739 18432 39804 18433
rect 38134 18423 39805 18432
rect 38134 18379 39739 18423
rect 38133 18369 39739 18379
rect 39804 18369 39805 18423
rect 38133 18358 39805 18369
rect 38133 18270 39167 18358
rect 40561 18346 40861 18443
rect 40960 18346 40961 18443
rect 40561 18338 40961 18346
rect 40652 18334 40961 18338
rect 40266 17873 40419 17883
rect 40266 17734 40419 17744
rect 41408 17875 41561 17885
rect 41408 17736 41561 17746
rect 39512 17229 39665 17239
rect 39512 17090 39665 17100
rect 41410 17229 41563 17239
rect 41410 17090 41563 17100
rect 40844 16258 40922 16268
rect 40844 16162 40922 16172
rect 42484 15210 42552 18993
rect 47119 18450 47179 19111
rect 53847 19277 54000 19287
rect 53532 19182 53588 19192
rect 52700 19138 52853 19148
rect 53531 19116 53532 19178
rect 53588 19116 53713 19178
rect 59213 19280 59366 19290
rect 53847 19138 54000 19148
rect 56329 19223 56482 19233
rect 53532 19106 53588 19116
rect 49795 19079 49948 19089
rect 48118 19062 48184 19065
rect 48118 19055 49110 19062
rect 48184 18989 49110 19055
rect 48118 18979 48184 18989
rect 47119 18449 47257 18450
rect 47119 18439 47519 18449
rect 45199 18428 45267 18438
rect 46297 18428 46362 18429
rect 45267 18419 46363 18428
rect 45267 18365 46297 18419
rect 46362 18365 46363 18419
rect 45267 18354 46363 18365
rect 45199 18343 45267 18353
rect 47119 18342 47419 18439
rect 47518 18342 47519 18439
rect 47119 18334 47519 18342
rect 47210 18330 47519 18334
rect 42970 18030 42980 18183
rect 43109 18030 43119 18183
rect 44489 18132 44900 18151
rect 44489 17996 44513 18132
rect 44737 17996 44900 18132
rect 44489 17978 44900 17996
rect 43996 17595 44112 17596
rect 44452 17595 44619 17596
rect 43996 17585 44619 17595
rect 43223 17572 43376 17582
rect 43996 17479 44001 17585
rect 44113 17568 44619 17585
rect 44113 17479 44495 17568
rect 43996 17462 44495 17479
rect 44607 17462 44619 17568
rect 43996 17453 44619 17462
rect 43223 17433 43376 17443
rect 42956 16380 42966 16533
rect 43095 16380 43105 16533
rect 43712 16473 43830 16476
rect 44455 16474 44620 16484
rect 44452 16473 44620 16474
rect 43712 16466 44620 16473
rect 43830 16456 44620 16466
rect 43830 16454 44496 16456
rect 43830 16348 44490 16454
rect 44608 16350 44620 16456
rect 44602 16348 44620 16350
rect 43712 16341 44620 16348
rect 43712 16339 44614 16341
rect 43712 16338 44577 16339
rect 43228 15968 43381 15978
rect 43228 15829 43381 15839
rect 42720 15210 42783 15216
rect 42484 15206 42788 15210
rect 42484 15154 42720 15206
rect 42783 15154 42788 15206
rect 42484 15148 42788 15154
rect 42720 15144 42783 15148
rect 39566 14832 39719 14842
rect 39566 14693 39719 14703
rect 41464 14832 41617 14842
rect 42961 14776 42971 14929
rect 43100 14776 43110 14929
rect 41464 14693 41617 14703
rect 43717 14687 43833 16338
rect 44228 16094 44343 16104
rect 44228 15987 44343 15997
rect 43716 14677 43833 14687
rect 43828 14571 43833 14677
rect 43716 14561 43833 14571
rect 43717 14560 43833 14561
rect 33107 13252 33168 13257
rect 30696 13247 33172 13252
rect 30696 13195 33107 13247
rect 33168 13195 33172 13247
rect 30696 13194 33172 13195
rect 30696 13161 30767 13194
rect 33107 13185 33168 13194
rect 30505 13149 30571 13155
rect 30696 13097 30701 13161
rect 30762 13097 30767 13161
rect 30696 13085 30767 13097
rect 44746 13099 44900 17978
rect 46824 17869 46977 17879
rect 46824 17730 46977 17740
rect 47966 17871 48119 17881
rect 47966 17732 48119 17742
rect 46070 17225 46223 17235
rect 46070 17086 46223 17096
rect 47968 17225 48121 17235
rect 47968 17086 48121 17096
rect 47402 16254 47480 16264
rect 47402 16158 47480 16168
rect 49042 15206 49110 18989
rect 53653 18455 53713 19116
rect 60360 19280 60513 19290
rect 60045 19185 60101 19195
rect 59213 19141 59366 19151
rect 60044 19119 60045 19181
rect 60101 19119 60226 19181
rect 60360 19141 60513 19151
rect 62842 19226 62995 19236
rect 60045 19109 60101 19119
rect 56329 19084 56482 19094
rect 54652 19067 54718 19070
rect 54652 19060 55644 19067
rect 54718 18994 55644 19060
rect 54652 18984 54718 18994
rect 53653 18454 53791 18455
rect 53653 18444 54053 18454
rect 51733 18433 51801 18443
rect 52831 18433 52896 18434
rect 51801 18424 52897 18433
rect 51801 18370 52831 18424
rect 52896 18370 52897 18424
rect 51801 18359 52897 18370
rect 51733 18348 51801 18358
rect 53653 18347 53953 18444
rect 54052 18347 54053 18444
rect 53653 18339 54053 18347
rect 53744 18335 54053 18339
rect 49528 18026 49538 18179
rect 49667 18026 49677 18179
rect 51041 18146 51496 18158
rect 51041 17990 51056 18146
rect 51306 17990 51496 18146
rect 51041 17973 51496 17990
rect 51311 17748 51496 17973
rect 51312 17617 51496 17748
rect 53358 17874 53511 17884
rect 53358 17735 53511 17745
rect 54500 17876 54653 17886
rect 54500 17737 54653 17747
rect 50554 17591 50670 17592
rect 51010 17591 51177 17592
rect 50554 17581 51177 17591
rect 49781 17568 49934 17578
rect 50554 17475 50559 17581
rect 50671 17564 51177 17581
rect 50671 17475 51053 17564
rect 50554 17458 51053 17475
rect 51165 17458 51177 17564
rect 50554 17449 51177 17458
rect 49781 17429 49934 17439
rect 49514 16376 49524 16529
rect 49653 16376 49663 16529
rect 50270 16469 50388 16472
rect 51013 16470 51178 16480
rect 51010 16469 51178 16470
rect 50270 16462 51178 16469
rect 50388 16452 51178 16462
rect 50388 16450 51054 16452
rect 50388 16344 51048 16450
rect 51166 16346 51178 16452
rect 51160 16344 51178 16346
rect 50270 16337 51178 16344
rect 50270 16335 51172 16337
rect 50270 16334 51135 16335
rect 49786 15964 49939 15974
rect 49786 15825 49939 15835
rect 49278 15206 49341 15212
rect 49042 15202 49346 15206
rect 49042 15150 49278 15202
rect 49341 15150 49346 15202
rect 49042 15144 49346 15150
rect 49278 15140 49341 15144
rect 46124 14828 46277 14838
rect 46124 14689 46277 14699
rect 48022 14828 48175 14838
rect 49519 14772 49529 14925
rect 49658 14772 49668 14925
rect 48022 14689 48175 14699
rect 50275 14683 50391 16334
rect 50786 16090 50901 16100
rect 50786 15983 50901 15993
rect 50274 14673 50391 14683
rect 50386 14567 50391 14673
rect 50274 14557 50391 14567
rect 50275 14556 50391 14557
rect 51311 13288 51496 17617
rect 52604 17230 52757 17240
rect 52604 17091 52757 17101
rect 54502 17230 54655 17240
rect 54502 17091 54655 17101
rect 53936 16259 54014 16269
rect 53936 16163 54014 16173
rect 55576 15211 55644 18994
rect 60166 18458 60226 19119
rect 62842 19087 62995 19097
rect 68233 19159 68333 19171
rect 68233 19076 68248 19159
rect 68316 19076 68333 19159
rect 61165 19070 61231 19073
rect 61165 19063 62157 19070
rect 61231 18997 62157 19063
rect 61165 18987 61231 18997
rect 60166 18457 60304 18458
rect 60166 18447 60566 18457
rect 58246 18436 58314 18446
rect 59344 18436 59409 18437
rect 58314 18427 59410 18436
rect 58314 18373 59344 18427
rect 59409 18373 59410 18427
rect 58314 18362 59410 18373
rect 58246 18351 58314 18361
rect 60166 18350 60466 18447
rect 60565 18350 60566 18447
rect 60166 18342 60566 18350
rect 60257 18338 60566 18342
rect 56062 18031 56072 18184
rect 56201 18031 56211 18184
rect 57584 18135 58021 18152
rect 57584 17998 57605 18135
rect 57833 17998 58021 18135
rect 57584 17978 58021 17998
rect 57088 17596 57204 17597
rect 57544 17596 57711 17597
rect 57088 17586 57711 17596
rect 56315 17573 56468 17583
rect 57088 17480 57093 17586
rect 57205 17569 57711 17586
rect 57205 17480 57587 17569
rect 57088 17463 57587 17480
rect 57699 17463 57711 17569
rect 57088 17454 57711 17463
rect 56315 17434 56468 17444
rect 56048 16381 56058 16534
rect 56187 16381 56197 16534
rect 56804 16474 56922 16477
rect 57547 16475 57712 16485
rect 57544 16474 57712 16475
rect 56804 16467 57712 16474
rect 56922 16457 57712 16467
rect 56922 16455 57588 16457
rect 56922 16349 57582 16455
rect 57700 16351 57712 16457
rect 57694 16349 57712 16351
rect 56804 16342 57712 16349
rect 56804 16340 57706 16342
rect 56804 16339 57669 16340
rect 56320 15969 56473 15979
rect 56320 15830 56473 15840
rect 55812 15211 55875 15217
rect 55576 15207 55880 15211
rect 55576 15155 55812 15207
rect 55875 15155 55880 15207
rect 55576 15149 55880 15155
rect 55812 15145 55875 15149
rect 52658 14833 52811 14843
rect 52658 14694 52811 14704
rect 54556 14833 54709 14843
rect 56053 14777 56063 14930
rect 56192 14777 56202 14930
rect 54556 14694 54709 14704
rect 56809 14688 56925 16339
rect 57320 16095 57435 16105
rect 57320 15988 57435 15998
rect 56808 14678 56925 14688
rect 56920 14572 56925 14678
rect 56808 14562 56925 14572
rect 56809 14561 56925 14562
rect 57840 13346 58019 17978
rect 59871 17877 60024 17887
rect 59871 17738 60024 17748
rect 61013 17879 61166 17889
rect 61013 17740 61166 17750
rect 59117 17233 59270 17243
rect 59117 17094 59270 17104
rect 61015 17233 61168 17243
rect 61015 17094 61168 17104
rect 60449 16262 60527 16272
rect 60449 16166 60527 16176
rect 62089 15214 62157 18997
rect 62575 18034 62585 18187
rect 62714 18034 62724 18187
rect 64465 18150 64538 18153
rect 64094 18129 64538 18150
rect 64094 17998 64118 18129
rect 64350 17998 64538 18129
rect 64094 17984 64538 17998
rect 64351 17895 64538 17984
rect 63997 17637 64259 17659
rect 63601 17599 63717 17600
rect 63997 17599 64020 17637
rect 63601 17589 64020 17599
rect 62828 17576 62981 17586
rect 63601 17483 63606 17589
rect 63718 17483 64020 17589
rect 63601 17481 64020 17483
rect 64238 17481 64259 17637
rect 63601 17457 64259 17481
rect 62828 17437 62981 17447
rect 62561 16384 62571 16537
rect 62700 16384 62710 16537
rect 63317 16477 63435 16480
rect 64060 16478 64225 16488
rect 64057 16477 64225 16478
rect 63317 16470 64225 16477
rect 63435 16460 64225 16470
rect 63435 16458 64101 16460
rect 63435 16352 64095 16458
rect 64213 16354 64225 16460
rect 64207 16352 64225 16354
rect 63317 16345 64225 16352
rect 63317 16343 64219 16345
rect 63317 16342 64182 16343
rect 62833 15972 62986 15982
rect 62833 15833 62986 15843
rect 62325 15214 62388 15220
rect 62089 15210 62393 15214
rect 62089 15158 62325 15210
rect 62388 15158 62393 15210
rect 62089 15152 62393 15158
rect 62325 15148 62388 15152
rect 59171 14836 59324 14846
rect 59171 14697 59324 14707
rect 61069 14836 61222 14846
rect 62566 14780 62576 14933
rect 62705 14780 62715 14933
rect 61069 14697 61222 14707
rect 63322 14691 63438 16342
rect 63833 16098 63948 16108
rect 63833 15991 63948 16001
rect 63321 14681 63438 14691
rect 63433 14575 63438 14681
rect 63321 14565 63438 14575
rect 63322 14564 63438 14565
rect 64352 13505 64538 17895
rect 64352 13504 64375 13505
rect 64352 13415 64365 13504
rect 64352 13414 64375 13415
rect 64526 13414 64538 13505
rect 64352 13401 64538 13414
rect 64465 13399 64538 13401
rect 51311 13199 51497 13288
rect 57840 13258 57855 13346
rect 58004 13258 58019 13346
rect 57840 13245 58019 13258
rect 51311 13111 51328 13199
rect 51484 13111 51497 13199
rect 29685 12275 29695 12353
rect 29765 12275 29775 12353
rect 30505 11761 30571 13083
rect 44746 13039 44901 13099
rect 51311 13098 51497 13111
rect 57724 13180 57823 13190
rect 57724 13068 57823 13078
rect 44746 12942 44758 13039
rect 44887 12995 44901 13039
rect 51199 13050 51299 13060
rect 44887 12942 44900 12995
rect 51199 12955 51299 12965
rect 44746 12932 44900 12942
rect 44619 12714 44737 12724
rect 44619 12636 44737 12646
rect 31915 12333 31925 12405
rect 31995 12333 32005 12405
rect 55114 12395 55174 12405
rect 41911 12375 41971 12385
rect 41911 12303 41971 12313
rect 48460 12374 48520 12384
rect 55114 12323 55174 12333
rect 48460 12302 48520 12312
rect 63767 12228 63827 12238
rect 63767 12156 63827 12166
rect 66013 12168 66166 12178
rect 66013 12029 66166 12039
rect 30505 11707 30511 11761
rect 30565 11707 30571 11761
rect 67368 11820 67428 11830
rect 67368 11748 67428 11758
rect 31064 11526 31160 11536
rect 31064 11419 31160 11429
rect 65221 11248 65288 11253
rect 65214 11243 66930 11248
rect 55336 11199 55398 11201
rect 55336 11191 55400 11199
rect 55398 11189 55400 11191
rect 42133 11179 42195 11181
rect 42133 11171 42197 11179
rect 42195 11169 42197 11171
rect 33107 11166 33164 11169
rect 27727 11106 29100 11107
rect 24001 11062 25302 11070
rect 25817 11099 29100 11106
rect 9468 11060 9525 11062
rect 12612 11060 12669 11062
rect 22090 11060 22147 11062
rect 25234 11060 25291 11062
rect 25817 11029 25837 11099
rect 25904 11029 29100 11099
rect 30690 11159 33172 11166
rect 30690 11105 33107 11159
rect 33164 11105 33172 11159
rect 30690 11095 33172 11105
rect 42133 11097 42197 11107
rect 48682 11178 48744 11180
rect 48682 11170 48746 11178
rect 48744 11168 48746 11170
rect 65214 11180 65221 11243
rect 65288 11238 66930 11243
rect 65288 11182 66877 11238
rect 65288 11180 66930 11182
rect 65214 11172 66930 11180
rect 65221 11170 65288 11172
rect 63112 11156 63191 11165
rect 55336 11117 55400 11127
rect 59163 11155 63191 11156
rect 48682 11096 48746 11106
rect 30690 11090 30766 11095
rect 25817 11020 29100 11029
rect 30503 11081 30569 11087
rect 25837 11019 25904 11020
rect 30690 11028 30699 11090
rect 30759 11028 30766 11090
rect 30690 11017 30766 11028
rect 59163 11081 63112 11155
rect 67001 11135 67074 11145
rect 65221 11126 65288 11127
rect 65481 11126 67001 11135
rect 59163 11080 63191 11081
rect 142 10937 3591 10947
rect 201 10930 3591 10937
rect 201 10867 3520 10930
rect 142 10859 3520 10867
rect 142 10857 201 10859
rect 3520 10849 3591 10859
rect 6650 10771 6720 10781
rect 140 10745 6650 10758
rect 140 10682 141 10745
rect 202 10682 6650 10745
rect 140 10678 6650 10682
rect 140 10672 6720 10678
rect 6650 10668 6720 10672
rect 9783 10542 9879 10550
rect 140 10540 9879 10542
rect 140 10525 9783 10540
rect 140 10459 141 10525
rect 203 10459 9783 10525
rect 140 10448 9783 10459
rect 9783 10435 9879 10445
rect 139 10336 13079 10346
rect 139 10329 13001 10336
rect 139 10271 140 10329
rect 203 10271 13001 10329
rect 139 10267 13001 10271
rect 139 10260 13079 10267
rect 13001 10257 13079 10260
rect 29683 10207 29693 10285
rect 29763 10207 29773 10285
rect 22408 10184 22472 10187
rect 22397 10177 22482 10184
rect 1774 10152 1850 10162
rect 1774 10084 1850 10094
rect 4918 10152 4994 10162
rect 4918 10084 4994 10094
rect 8050 10148 8126 10158
rect 8050 10080 8126 10090
rect 11194 10148 11270 10158
rect 11194 10080 11270 10090
rect 14396 10152 14472 10162
rect 14396 10084 14472 10094
rect 17540 10152 17616 10162
rect 20672 10148 20748 10158
rect 19294 10118 19362 10128
rect 17540 10084 17616 10094
rect 19284 10046 19294 10106
rect 19362 10046 19371 10106
rect 20672 10080 20748 10090
rect 22397 10100 22408 10177
rect 22472 10100 22482 10177
rect 139 10002 16224 10003
rect 139 9992 16226 10002
rect 139 9986 16159 9992
rect 139 9925 140 9986
rect 204 9925 16159 9986
rect 139 9924 16159 9925
rect 139 9914 16226 9924
rect 19284 9830 19371 10046
rect 136 9814 19371 9830
rect 136 9754 138 9814
rect 202 9754 19371 9814
rect 136 9743 19371 9754
rect 1780 9664 1880 9674
rect 1780 9562 1880 9572
rect 4924 9664 5024 9674
rect 4924 9562 5024 9572
rect 8056 9660 8156 9670
rect 8056 9558 8156 9568
rect 11200 9660 11300 9670
rect 11200 9558 11300 9568
rect 14402 9664 14502 9674
rect 14402 9562 14502 9572
rect 17546 9664 17646 9674
rect 17546 9562 17646 9572
rect 20678 9660 20778 9670
rect 20678 9558 20778 9568
rect 22397 9479 22482 10100
rect 23816 10148 23892 10158
rect 23816 10080 23892 10090
rect 30503 9693 30569 11015
rect 34107 10951 34223 10961
rect 34097 10895 34107 10941
rect 34223 10940 51000 10941
rect 59163 10940 59232 11080
rect 63112 11071 63191 11080
rect 65213 11125 67001 11126
rect 65213 11117 65481 11125
rect 65213 11054 65221 11117
rect 65288 11057 65481 11117
rect 65536 11057 67001 11125
rect 65288 11054 67001 11057
rect 63264 11041 63345 11051
rect 65213 11047 67001 11054
rect 65214 11046 65303 11047
rect 67977 11142 68115 11152
rect 67977 11050 68115 11060
rect 65221 11044 65288 11046
rect 34223 10895 59232 10940
rect 34097 10881 59232 10895
rect 59286 11033 59360 11034
rect 59286 11032 61620 11033
rect 59286 10951 63264 11032
rect 59286 10853 59360 10951
rect 61434 10950 63264 10951
rect 67001 11036 67074 11046
rect 63989 11032 64051 11034
rect 63989 11024 64053 11032
rect 64051 11022 64053 11024
rect 63989 10950 64053 10960
rect 63264 10935 63345 10945
rect 33887 10837 59360 10853
rect 33887 10779 33893 10837
rect 33977 10787 59360 10837
rect 66535 10887 67892 10897
rect 66597 10882 67892 10887
rect 66597 10801 67774 10882
rect 67882 10801 67892 10882
rect 66597 10796 67892 10801
rect 33977 10779 33988 10787
rect 33887 10768 33988 10779
rect 35247 10475 35307 10485
rect 34131 10456 34199 10462
rect 34120 10452 34211 10456
rect 34120 10400 34131 10452
rect 34199 10400 34211 10452
rect 35247 10403 35307 10413
rect 31913 10265 31923 10337
rect 31993 10265 32003 10337
rect 23822 9660 23922 9670
rect 30503 9639 30509 9693
rect 30563 9639 30569 9693
rect 23822 9558 23922 9568
rect 136 9460 22482 9479
rect 203 9399 22482 9460
rect 136 9387 22482 9399
rect 22397 9386 22482 9387
rect 31066 9456 31158 9466
rect 31066 9354 31158 9364
rect 32542 9318 33875 9330
rect 32542 9302 33775 9318
rect 32542 9228 32549 9302
rect 32615 9228 33775 9302
rect 32542 9226 33775 9228
rect 33865 9226 33875 9318
rect 32542 9218 33875 9226
rect 33775 9216 33865 9218
rect 33103 9111 33166 9113
rect 30689 9103 33174 9111
rect 30689 9042 33103 9103
rect 33166 9042 33174 9103
rect 30689 9037 33174 9042
rect 30690 9021 30767 9037
rect 33103 9032 33166 9037
rect 30505 9012 30571 9018
rect 30690 8961 30702 9021
rect 30762 8961 30767 9021
rect 30690 8949 30767 8961
rect 2933 8703 3026 8705
rect 3202 8703 3259 8704
rect 6077 8703 6170 8705
rect 6346 8703 6403 8704
rect 15555 8703 15648 8705
rect 15824 8703 15881 8704
rect 18699 8703 18792 8705
rect 18968 8703 19025 8704
rect 1851 8702 3267 8703
rect 4995 8702 6411 8703
rect 14473 8702 15889 8703
rect 17617 8702 19033 8703
rect 1851 8699 3270 8702
rect 4995 8699 6414 8702
rect 9209 8699 9302 8701
rect 9478 8699 9535 8700
rect 12353 8699 12446 8701
rect 12622 8699 12679 8700
rect 14473 8699 15892 8702
rect 17617 8699 19036 8702
rect 21831 8699 21924 8701
rect 22100 8699 22157 8700
rect 24975 8699 25068 8701
rect 25244 8699 25301 8700
rect 1851 8694 25312 8699
rect 1851 8693 3202 8694
rect 1851 8631 1860 8693
rect 1930 8631 2944 8693
rect 1851 8630 2944 8631
rect 3015 8630 3202 8693
rect 1851 8626 3202 8630
rect 3259 8693 6346 8694
rect 3259 8631 5004 8693
rect 5074 8631 6088 8693
rect 3259 8630 6088 8631
rect 6159 8630 6346 8693
rect 3259 8626 6346 8630
rect 6403 8693 15824 8694
rect 6403 8690 14482 8693
rect 6403 8689 9478 8690
rect 6403 8627 8136 8689
rect 8206 8627 9220 8689
rect 6403 8626 9220 8627
rect 9291 8626 9478 8689
rect 1851 8622 9478 8626
rect 9535 8689 12622 8690
rect 9535 8627 11280 8689
rect 11350 8627 12364 8689
rect 9535 8626 12364 8627
rect 12435 8626 12622 8689
rect 9535 8622 12622 8626
rect 12679 8631 14482 8690
rect 14552 8631 15566 8693
rect 12679 8630 15566 8631
rect 15637 8630 15824 8693
rect 12679 8626 15824 8630
rect 15881 8693 18968 8694
rect 15881 8631 17626 8693
rect 17696 8631 18710 8693
rect 15881 8630 18710 8631
rect 18781 8630 18968 8693
rect 15881 8626 18968 8630
rect 19025 8690 25312 8694
rect 19025 8689 22100 8690
rect 19025 8627 20758 8689
rect 20828 8627 21842 8689
rect 19025 8626 21842 8627
rect 21913 8626 22100 8689
rect 12679 8622 22100 8626
rect 22157 8689 25244 8690
rect 22157 8627 23902 8689
rect 23972 8627 24986 8689
rect 22157 8626 24986 8627
rect 25057 8626 25244 8689
rect 22157 8622 25244 8626
rect 25301 8622 25312 8690
rect 1851 8614 25312 8622
rect 9478 8612 9535 8614
rect 12622 8612 12679 8614
rect 22100 8612 22157 8614
rect 25244 8612 25301 8614
rect 1630 8578 3270 8583
rect 1630 8573 3202 8578
rect 1689 8513 3202 8573
rect 1630 8510 3202 8513
rect 3259 8510 3270 8578
rect 1630 8504 3270 8510
rect 1630 8503 1689 8504
rect 3174 8501 3270 8504
rect 4774 8578 6414 8583
rect 9478 8582 9535 8584
rect 12622 8582 12679 8584
rect 9450 8579 9546 8582
rect 12594 8579 12690 8582
rect 4774 8573 6346 8578
rect 4833 8513 6346 8573
rect 4774 8510 6346 8513
rect 6403 8510 6414 8578
rect 4774 8504 6414 8510
rect 4774 8503 4833 8504
rect 6318 8501 6414 8504
rect 7906 8574 9546 8579
rect 7906 8569 9478 8574
rect 7965 8509 9478 8569
rect 7906 8506 9478 8509
rect 9535 8506 9546 8574
rect 3202 8500 3259 8501
rect 6346 8500 6403 8501
rect 7906 8500 9546 8506
rect 7906 8499 7965 8500
rect 9450 8497 9546 8500
rect 11050 8574 12690 8579
rect 11050 8569 12622 8574
rect 11109 8509 12622 8569
rect 11050 8506 12622 8509
rect 12679 8506 12690 8574
rect 11050 8500 12690 8506
rect 14252 8578 15892 8583
rect 14252 8573 15824 8578
rect 14311 8513 15824 8573
rect 14252 8510 15824 8513
rect 15881 8510 15892 8578
rect 14252 8504 15892 8510
rect 14252 8503 14311 8504
rect 15796 8501 15892 8504
rect 17396 8578 19036 8583
rect 22100 8582 22157 8584
rect 25244 8582 25301 8584
rect 22072 8579 22168 8582
rect 25216 8579 25312 8582
rect 17396 8573 18968 8578
rect 17455 8513 18968 8573
rect 17396 8510 18968 8513
rect 19025 8510 19036 8578
rect 17396 8504 19036 8510
rect 17396 8503 17455 8504
rect 18940 8501 19036 8504
rect 20528 8574 22168 8579
rect 20528 8569 22100 8574
rect 20587 8509 22100 8569
rect 20528 8506 22100 8509
rect 22157 8506 22168 8574
rect 15824 8500 15881 8501
rect 18968 8500 19025 8501
rect 20528 8500 22168 8506
rect 11050 8499 11109 8500
rect 12594 8497 12690 8500
rect 20528 8499 20587 8500
rect 22072 8497 22168 8500
rect 23672 8574 25312 8579
rect 23672 8569 25244 8574
rect 23731 8509 25244 8569
rect 23672 8506 25244 8509
rect 25301 8506 25312 8574
rect 23672 8500 25312 8506
rect 23672 8499 23731 8500
rect 25216 8497 25312 8500
rect 9478 8496 9535 8497
rect 12622 8496 12679 8497
rect 22100 8496 22157 8497
rect 25244 8496 25301 8497
rect 3202 8419 3259 8420
rect 6346 8419 6403 8420
rect 15824 8419 15881 8420
rect 18968 8419 19025 8420
rect 3174 8418 3270 8419
rect 6318 8418 6414 8419
rect 15796 8418 15892 8419
rect 18940 8418 19036 8419
rect 1969 8410 3270 8418
rect 1969 8345 1980 8410
rect 2048 8345 3202 8410
rect 1969 8342 3202 8345
rect 3259 8342 3270 8410
rect 1969 8334 3270 8342
rect 5113 8410 6414 8418
rect 9478 8415 9535 8416
rect 12622 8415 12679 8416
rect 9450 8414 9546 8415
rect 12594 8414 12690 8415
rect 5113 8345 5124 8410
rect 5192 8345 6346 8410
rect 5113 8342 6346 8345
rect 6403 8342 6414 8410
rect 5113 8334 6414 8342
rect 8245 8406 9546 8414
rect 8245 8341 8256 8406
rect 8324 8341 9478 8406
rect 8245 8338 9478 8341
rect 9535 8338 9546 8406
rect 3202 8332 3259 8334
rect 6346 8332 6403 8334
rect 8245 8330 9546 8338
rect 11389 8406 12690 8414
rect 11389 8341 11400 8406
rect 11468 8341 12622 8406
rect 11389 8338 12622 8341
rect 12679 8338 12690 8406
rect 11389 8330 12690 8338
rect 14591 8410 15892 8418
rect 14591 8345 14602 8410
rect 14670 8345 15824 8410
rect 14591 8342 15824 8345
rect 15881 8342 15892 8410
rect 14591 8334 15892 8342
rect 17735 8410 19036 8418
rect 22100 8415 22157 8416
rect 25244 8415 25301 8416
rect 22072 8414 22168 8415
rect 25216 8414 25312 8415
rect 17735 8345 17746 8410
rect 17814 8345 18968 8410
rect 17735 8342 18968 8345
rect 19025 8342 19036 8410
rect 17735 8334 19036 8342
rect 20867 8406 22168 8414
rect 20867 8341 20878 8406
rect 20946 8341 22100 8406
rect 20867 8338 22100 8341
rect 22157 8338 22168 8406
rect 15824 8332 15881 8334
rect 18968 8332 19025 8334
rect 20867 8330 22168 8338
rect 24011 8406 25312 8414
rect 24011 8341 24022 8406
rect 24090 8341 25244 8406
rect 24011 8338 25244 8341
rect 25301 8338 25312 8406
rect 24011 8330 25312 8338
rect 9478 8328 9535 8330
rect 12622 8328 12679 8330
rect 22100 8328 22157 8330
rect 25244 8328 25301 8330
rect 29685 8138 29695 8216
rect 29765 8138 29775 8216
rect 30505 7624 30571 8946
rect 31915 8196 31925 8268
rect 31995 8196 32005 8268
rect 30505 7570 30511 7624
rect 30565 7570 30571 7624
rect 1784 7420 1860 7430
rect 1784 7352 1860 7362
rect 4928 7420 5004 7430
rect 4928 7352 5004 7362
rect 8060 7416 8136 7426
rect 8060 7348 8136 7358
rect 11204 7416 11280 7426
rect 11204 7348 11280 7358
rect 14406 7420 14482 7430
rect 14406 7352 14482 7362
rect 17550 7420 17626 7430
rect 17550 7352 17626 7362
rect 20682 7416 20758 7426
rect 20682 7348 20758 7358
rect 23826 7416 23902 7426
rect 23826 7348 23902 7358
rect 31072 7384 31157 7394
rect 31072 7288 31157 7298
rect 32407 7207 33286 7217
rect 27321 7158 27389 7167
rect 27506 7158 27562 7168
rect 27317 7157 27506 7158
rect 27317 7099 27321 7157
rect 27389 7099 27506 7157
rect 27317 7096 27506 7099
rect 32407 7143 32416 7207
rect 32478 7143 33286 7207
rect 32407 7131 33286 7143
rect 27321 7089 27389 7096
rect 27506 7086 27562 7096
rect 33103 7046 33166 7049
rect 30688 7039 33173 7046
rect 30688 6978 33103 7039
rect 33166 6978 33173 7039
rect 30688 6971 33173 6978
rect 30689 6953 30768 6971
rect 33103 6968 33166 6971
rect 30503 6944 30569 6950
rect 30689 6892 30701 6953
rect 30756 6892 30768 6953
rect 30689 6882 30768 6892
rect 27074 6865 27130 6873
rect 27506 6867 27562 6877
rect 27063 6863 27506 6865
rect 27063 6806 27074 6863
rect 27130 6806 27506 6863
rect 27063 6805 27506 6806
rect 27063 6804 27562 6805
rect 27074 6796 27130 6804
rect 27506 6795 27562 6804
rect 3273 6761 3367 6771
rect 3273 6667 3367 6677
rect 4011 6761 4105 6771
rect 4011 6667 4105 6677
rect 4749 6761 4843 6771
rect 4749 6667 4843 6677
rect 5487 6761 5581 6771
rect 5487 6667 5581 6677
rect 6227 6761 6321 6771
rect 6227 6667 6321 6677
rect 6969 6761 7063 6771
rect 6969 6667 7063 6677
rect 7707 6761 7801 6771
rect 7707 6667 7801 6677
rect 8445 6763 8539 6773
rect 8445 6669 8539 6679
rect 10049 6706 10127 6716
rect 10049 6626 10127 6636
rect 12117 6704 12195 6714
rect 12117 6624 12195 6634
rect 14186 6706 14264 6716
rect 14186 6626 14264 6636
rect 16254 6704 16332 6714
rect 16254 6624 16332 6634
rect 18323 6704 18401 6714
rect 18323 6624 18401 6634
rect 20391 6702 20469 6712
rect 20391 6622 20469 6632
rect 22460 6704 22538 6714
rect 22460 6624 22538 6634
rect 24528 6702 24606 6712
rect 24528 6622 24606 6632
rect 26851 6560 26912 6565
rect 27507 6561 27563 6571
rect 26849 6555 27507 6560
rect 26849 6502 26851 6555
rect 26912 6502 27507 6555
rect 26849 6499 27507 6502
rect 26851 6492 26912 6499
rect 27507 6489 27563 6499
rect 26667 6399 26737 6408
rect 27506 6400 27562 6410
rect 26662 6398 27506 6399
rect 26662 6340 26667 6398
rect 26737 6340 27506 6398
rect 26662 6338 27506 6340
rect 26667 6330 26737 6338
rect 27506 6328 27562 6338
rect 26467 6248 26535 6258
rect 27506 6249 27562 6259
rect 26464 6190 26467 6248
rect 26535 6190 27506 6248
rect 26464 6187 27506 6190
rect 26467 6180 26535 6187
rect 27506 6177 27562 6187
rect 26281 6088 26339 6095
rect 27506 6088 27562 6098
rect 26277 6085 27506 6088
rect 26277 6031 26281 6085
rect 26339 6031 27506 6085
rect 26277 6027 27506 6031
rect 26281 6021 26339 6027
rect 29683 6070 29693 6148
rect 29763 6070 29773 6148
rect 27506 6016 27562 6026
rect 10847 5905 10930 5915
rect 23264 5910 23339 5920
rect 9481 5890 10847 5896
rect 3333 5873 3435 5879
rect 4071 5873 4173 5879
rect 4809 5873 4911 5879
rect 5547 5873 5649 5879
rect 6287 5873 6389 5879
rect 7029 5873 7131 5879
rect 7767 5873 7869 5879
rect 8505 5875 8607 5881
rect 3331 5869 3435 5873
rect 3331 5803 3333 5869
rect 3331 5795 3435 5803
rect 4069 5869 4173 5873
rect 4069 5803 4071 5869
rect 4069 5795 4173 5803
rect 4807 5869 4911 5873
rect 4807 5803 4809 5869
rect 4807 5795 4911 5803
rect 5545 5869 5649 5873
rect 5545 5803 5547 5869
rect 5545 5795 5649 5803
rect 6285 5869 6389 5873
rect 6285 5803 6287 5869
rect 6285 5795 6389 5803
rect 7027 5869 7131 5873
rect 7027 5803 7029 5869
rect 7027 5795 7131 5803
rect 7765 5869 7869 5873
rect 7765 5803 7767 5869
rect 7765 5795 7869 5803
rect 8503 5871 8607 5875
rect 8503 5805 8505 5871
rect 9535 5836 10847 5890
rect 9481 5830 10847 5836
rect 12927 5894 12994 5903
rect 15000 5896 15065 5906
rect 17061 5896 17128 5906
rect 11549 5888 12925 5894
rect 12991 5893 12997 5894
rect 11603 5834 12925 5888
rect 11549 5828 12925 5834
rect 12994 5829 12997 5893
rect 13618 5890 14994 5896
rect 13672 5836 14994 5890
rect 13618 5830 14994 5836
rect 15065 5830 15066 5896
rect 19132 5894 19196 5903
rect 15686 5888 17061 5894
rect 15740 5834 17061 5888
rect 12991 5828 12997 5829
rect 15686 5828 17061 5834
rect 17128 5828 17134 5894
rect 17755 5888 19131 5894
rect 17809 5834 19131 5888
rect 17755 5828 19131 5834
rect 19197 5828 19203 5894
rect 21199 5892 21268 5902
rect 26047 5902 26111 5911
rect 27506 5902 27562 5911
rect 26046 5901 27562 5902
rect 19823 5886 21199 5892
rect 19877 5832 21199 5886
rect 10847 5815 10930 5825
rect 12927 5819 12994 5828
rect 15000 5818 15065 5828
rect 17061 5817 17128 5827
rect 19132 5818 19196 5828
rect 19823 5826 21199 5832
rect 21268 5826 21271 5892
rect 21892 5888 23264 5894
rect 21946 5834 23264 5888
rect 21892 5828 23264 5834
rect 23339 5828 23340 5894
rect 23960 5886 25336 5892
rect 24014 5832 25336 5886
rect 21199 5816 21268 5826
rect 23960 5826 25336 5832
rect 25402 5826 25408 5892
rect 25624 5886 25690 5896
rect 26046 5841 26047 5901
rect 26111 5841 27506 5901
rect 26046 5840 27506 5841
rect 26047 5831 26111 5840
rect 27506 5829 27562 5839
rect 23264 5814 23339 5824
rect 25624 5819 25690 5829
rect 8503 5797 8607 5805
rect 8505 5795 8607 5797
rect 3333 5793 3435 5795
rect 4071 5793 4173 5795
rect 4809 5793 4911 5795
rect 5547 5793 5649 5795
rect 6287 5793 6389 5795
rect 7029 5793 7131 5795
rect 7767 5793 7869 5795
rect 25346 5704 25417 5714
rect 25346 5617 25417 5627
rect 25636 5694 25688 5703
rect 27506 5697 27562 5707
rect 25636 5693 27506 5694
rect 25688 5635 27506 5693
rect 25636 5625 25688 5635
rect 27506 5625 27562 5635
rect 30503 5556 30569 6878
rect 31913 6128 31923 6200
rect 31993 6128 32003 6200
rect 30503 5502 30509 5556
rect 30563 5502 30569 5556
rect 31067 5314 31156 5324
rect 31067 5219 31156 5229
rect 33102 4978 33169 4984
rect 30690 4974 33173 4978
rect 30690 4907 33102 4974
rect 33169 4907 33173 4974
rect 30690 4903 33173 4907
rect 30690 4884 30770 4903
rect 33102 4897 33169 4903
rect 30503 4875 30569 4881
rect 30690 4823 30700 4884
rect 30756 4823 30770 4884
rect 30690 4813 30770 4823
rect 474 4640 569 4650
rect 474 4552 569 4562
rect 248 4486 358 4496
rect 248 4387 358 4397
rect 10107 4476 10179 4486
rect 10107 4396 10179 4406
rect 12175 4474 12247 4484
rect 12175 4394 12247 4404
rect 14244 4476 14316 4486
rect 14244 4396 14316 4406
rect 16312 4474 16384 4484
rect 16312 4394 16384 4404
rect 18381 4474 18453 4484
rect 18381 4394 18453 4404
rect 20449 4472 20521 4482
rect 20449 4392 20521 4402
rect 22518 4474 22590 4484
rect 22518 4394 22590 4404
rect 24586 4472 24658 4482
rect 24586 4392 24658 4402
rect -10 4290 95 4300
rect -10 4196 95 4206
rect 29683 4001 29693 4079
rect 29763 4001 29773 4079
rect 30503 3487 30569 4809
rect 31913 4059 31923 4131
rect 31993 4059 32003 4131
rect 30503 3433 30509 3487
rect 30563 3433 30569 3487
rect 22037 3423 22119 3424
rect 12384 3421 22119 3423
rect 142 3420 221 3421
rect 2821 3420 22119 3421
rect 116 3411 22119 3420
rect 116 3348 142 3411
rect 221 3348 22119 3411
rect 116 3338 22119 3348
rect 2821 3336 22119 3338
rect 6227 3288 18966 3290
rect 2926 3287 18966 3288
rect 116 3277 18966 3287
rect 116 3214 135 3277
rect 214 3214 18966 3277
rect 116 3205 18966 3214
rect 135 3204 214 3205
rect 2926 3203 18966 3205
rect 15863 3202 18966 3203
rect 6250 3173 15829 3175
rect 2926 3172 15829 3173
rect 115 3161 15829 3172
rect 115 3098 138 3161
rect 217 3098 15829 3161
rect 115 3090 15829 3098
rect 138 3088 217 3090
rect 2926 3088 15829 3090
rect 136 3057 215 3058
rect 2905 3057 12690 3060
rect 115 3048 12690 3057
rect 115 2985 136 3048
rect 215 3024 12690 3048
rect 215 2985 12697 3024
rect 115 2975 12697 2985
rect 2957 2934 6299 2935
rect 2957 2933 9488 2934
rect 115 2921 9488 2933
rect -33 2875 53 2889
rect -33 2773 -22 2875
rect 43 2818 53 2875
rect 115 2860 134 2921
rect 211 2916 9488 2921
rect 211 2860 9490 2916
rect 115 2851 9490 2860
rect 134 2850 211 2851
rect 2957 2850 9490 2851
rect 6235 2849 9490 2850
rect 43 2817 144 2818
rect 3001 2817 6343 2820
rect 43 2773 6343 2817
rect -33 2735 6343 2773
rect -33 2733 144 2735
rect 114 2684 3198 2698
rect 114 2627 130 2684
rect 214 2627 3198 2684
rect 114 2616 3198 2627
rect 1496 2412 1596 2422
rect 1496 2310 1596 2320
rect 117 1451 174 1452
rect 350 1451 443 1453
rect 109 1450 1525 1451
rect 106 1442 1525 1450
rect 106 1374 117 1442
rect 174 1441 1525 1442
rect 174 1378 361 1441
rect 432 1379 1446 1441
rect 1516 1379 1525 1441
rect 432 1378 1525 1379
rect 174 1374 1525 1378
rect 106 1367 1525 1374
rect 106 1366 184 1367
rect 117 1364 174 1366
rect 117 1334 174 1336
rect 106 1331 202 1334
rect 106 1326 1746 1331
rect 106 1258 117 1326
rect 174 1321 1746 1326
rect 174 1261 1687 1321
rect 174 1258 1746 1261
rect 106 1252 1746 1258
rect 106 1249 202 1252
rect 1687 1251 1746 1252
rect 117 1248 174 1249
rect 3116 1167 3198 2616
rect 4640 2412 4740 2422
rect 4640 2310 4740 2320
rect 3261 1451 3318 1452
rect 3494 1451 3587 1453
rect 3253 1450 4669 1451
rect 3250 1442 4669 1450
rect 3250 1374 3261 1442
rect 3318 1441 4669 1442
rect 3318 1378 3505 1441
rect 3576 1379 4590 1441
rect 4660 1379 4669 1441
rect 3576 1378 4669 1379
rect 3318 1374 4669 1378
rect 3250 1367 4669 1374
rect 3250 1366 3328 1367
rect 3261 1364 3318 1366
rect 3261 1334 3318 1336
rect 3250 1331 3346 1334
rect 3250 1326 4890 1331
rect 3250 1258 3261 1326
rect 3318 1321 4890 1326
rect 3318 1261 4831 1321
rect 3318 1258 4890 1261
rect 3250 1252 4890 1258
rect 3250 1249 3346 1252
rect 4831 1251 4890 1252
rect 3261 1248 3318 1249
rect 6266 1200 6343 2735
rect 7772 2416 7872 2426
rect 7772 2314 7872 2324
rect 6393 1455 6450 1456
rect 6626 1455 6719 1457
rect 6385 1454 7801 1455
rect 6382 1446 7801 1454
rect 6382 1378 6393 1446
rect 6450 1445 7801 1446
rect 6450 1382 6637 1445
rect 6708 1383 7722 1445
rect 7792 1383 7801 1445
rect 6708 1382 7801 1383
rect 6450 1378 7801 1382
rect 6382 1371 7801 1378
rect 6382 1370 6460 1371
rect 6393 1368 6450 1370
rect 6393 1338 6450 1340
rect 6382 1335 6478 1338
rect 6382 1330 8022 1335
rect 6382 1262 6393 1330
rect 6450 1325 8022 1330
rect 6450 1265 7963 1325
rect 6450 1262 8022 1265
rect 6382 1256 8022 1262
rect 6382 1253 6478 1256
rect 7963 1255 8022 1256
rect 6393 1252 6450 1253
rect 6265 1171 6344 1200
rect 6265 1170 6503 1171
rect 9412 1170 9490 2849
rect 10916 2416 11016 2426
rect 10916 2314 11016 2324
rect 9537 1455 9594 1456
rect 9770 1455 9863 1457
rect 9529 1454 10945 1455
rect 9526 1446 10945 1454
rect 9526 1378 9537 1446
rect 9594 1445 10945 1446
rect 9594 1382 9781 1445
rect 9852 1383 10866 1445
rect 10936 1383 10945 1445
rect 9852 1382 10945 1383
rect 9594 1378 10945 1382
rect 9526 1371 10945 1378
rect 9526 1370 9604 1371
rect 9537 1368 9594 1370
rect 9537 1338 9594 1340
rect 9526 1335 9622 1338
rect 9526 1330 11166 1335
rect 9526 1262 9537 1330
rect 9594 1325 11166 1330
rect 9594 1265 11107 1325
rect 9594 1262 11166 1265
rect 9526 1256 11166 1262
rect 9526 1253 9622 1256
rect 11107 1255 11166 1256
rect 9537 1252 9594 1253
rect 12620 1178 12697 2975
rect 14118 2412 14218 2422
rect 14118 2310 14218 2320
rect 12739 1451 12796 1452
rect 12972 1451 13065 1453
rect 12731 1450 14147 1451
rect 12728 1442 14147 1450
rect 12728 1374 12739 1442
rect 12796 1441 14147 1442
rect 12796 1378 12983 1441
rect 13054 1379 14068 1441
rect 14138 1379 14147 1441
rect 13054 1378 14147 1379
rect 12796 1374 14147 1378
rect 12728 1367 14147 1374
rect 12728 1366 12806 1367
rect 12739 1364 12796 1366
rect 12739 1334 12796 1336
rect 12728 1331 12824 1334
rect 12728 1326 14368 1331
rect 12728 1258 12739 1326
rect 12796 1321 14368 1326
rect 12796 1261 14309 1321
rect 12796 1258 14368 1261
rect 12728 1252 14368 1258
rect 12728 1249 12824 1252
rect 14309 1251 14368 1252
rect 12739 1248 12796 1249
rect 15756 1209 15829 3088
rect 17262 2412 17362 2422
rect 17262 2310 17362 2320
rect 15883 1451 15940 1452
rect 16116 1451 16209 1453
rect 15875 1450 17291 1451
rect 15872 1442 17291 1450
rect 15872 1374 15883 1442
rect 15940 1441 17291 1442
rect 15940 1378 16127 1441
rect 16198 1379 17212 1441
rect 17282 1379 17291 1441
rect 16198 1378 17291 1379
rect 15940 1374 17291 1378
rect 15872 1367 17291 1374
rect 15872 1366 15950 1367
rect 15883 1364 15940 1366
rect 15883 1334 15940 1336
rect 15872 1331 15968 1334
rect 15872 1326 17512 1331
rect 15872 1258 15883 1326
rect 15940 1321 17512 1326
rect 15940 1261 17453 1321
rect 15940 1258 17512 1261
rect 15872 1252 17512 1258
rect 15872 1249 15968 1252
rect 17453 1251 17512 1252
rect 15883 1248 15940 1249
rect 3116 1166 3375 1167
rect 249 1165 1407 1166
rect -310 1158 1407 1165
rect -310 1093 1328 1158
rect 1396 1093 1407 1158
rect 3116 1158 4551 1166
rect 3116 1095 4472 1158
rect -310 1082 1407 1093
rect 3117 1093 4472 1095
rect 4540 1093 4551 1158
rect 3117 1083 4551 1093
rect 6265 1162 7683 1170
rect 6265 1097 7604 1162
rect 7672 1097 7683 1162
rect 6265 1086 7683 1097
rect 9412 1162 10827 1170
rect 9412 1097 10748 1162
rect 10816 1097 10827 1162
rect 9412 1086 10827 1097
rect 12619 1168 12697 1178
rect 12619 1166 12865 1168
rect 15755 1166 15830 1209
rect 18896 1170 18966 3202
rect 20394 2416 20494 2426
rect 20394 2314 20494 2324
rect 19015 1455 19072 1456
rect 19248 1455 19341 1457
rect 19007 1454 20423 1455
rect 19004 1446 20423 1454
rect 19004 1378 19015 1446
rect 19072 1445 20423 1446
rect 19072 1382 19259 1445
rect 19330 1383 20344 1445
rect 20414 1383 20423 1445
rect 19330 1382 20423 1383
rect 19072 1378 20423 1382
rect 19004 1371 20423 1378
rect 19004 1370 19082 1371
rect 19015 1368 19072 1370
rect 19015 1338 19072 1340
rect 19004 1335 19100 1338
rect 19004 1330 20644 1335
rect 19004 1262 19015 1330
rect 19072 1325 20644 1330
rect 19072 1265 20585 1325
rect 19072 1262 20644 1265
rect 19004 1256 20644 1262
rect 19004 1253 19100 1256
rect 20585 1255 20644 1256
rect 19015 1252 19072 1253
rect 22037 1205 22119 3336
rect 31070 3245 31154 3255
rect 31070 3152 31154 3162
rect 30689 2900 33173 2911
rect 30689 2846 33108 2900
rect 33164 2846 33173 2900
rect 30689 2836 33173 2846
rect 30689 2817 30769 2836
rect 30501 2807 30567 2813
rect 30689 2755 30699 2817
rect 30755 2755 30769 2817
rect 30689 2745 30769 2755
rect 23538 2416 23638 2426
rect 23538 2314 23638 2324
rect 29681 1933 29691 2011
rect 29761 1933 29771 2011
rect 22159 1455 22216 1456
rect 22392 1455 22485 1457
rect 22151 1454 23567 1455
rect 22148 1446 23567 1454
rect 22148 1378 22159 1446
rect 22216 1445 23567 1446
rect 22216 1382 22403 1445
rect 22474 1383 23488 1445
rect 23558 1383 23567 1445
rect 22474 1382 23567 1383
rect 22216 1378 23567 1382
rect 22148 1371 23567 1378
rect 30501 1419 30567 2741
rect 31911 1991 31921 2063
rect 31991 1991 32001 2063
rect 22148 1370 22226 1371
rect 22159 1368 22216 1370
rect 30501 1365 30507 1419
rect 30561 1365 30567 1419
rect 22159 1338 22216 1340
rect 22148 1335 22244 1338
rect 22148 1330 23788 1335
rect 22148 1262 22159 1330
rect 22216 1325 23788 1330
rect 22216 1265 23729 1325
rect 22216 1262 23788 1265
rect 22148 1256 23788 1262
rect 22148 1253 22244 1256
rect 23729 1255 23788 1256
rect 22159 1252 22216 1253
rect 22036 1171 22119 1205
rect 31069 1178 31152 1188
rect 22036 1170 22295 1171
rect 12619 1158 14029 1166
rect 12619 1093 13950 1158
rect 14018 1093 14029 1158
rect 15755 1158 17173 1166
rect 15755 1136 17094 1158
rect 3341 1082 4551 1083
rect 12619 1082 14029 1093
rect 15756 1093 17094 1136
rect 17162 1093 17173 1158
rect 15756 1082 17173 1093
rect 18896 1162 20305 1170
rect 18896 1097 20226 1162
rect 20294 1097 20305 1162
rect 22036 1162 23449 1170
rect 22036 1139 23370 1162
rect 18896 1086 20305 1097
rect 22037 1097 23370 1139
rect 23438 1097 23449 1162
rect 22037 1086 23449 1097
rect 18896 1085 18966 1086
rect 22037 1085 22295 1086
rect 31069 1084 31152 1094
rect -310 1079 240 1082
rect 33218 1049 33286 7131
rect 33932 6707 34019 6711
rect 34120 6707 34211 10400
rect 35469 9279 35531 9281
rect 35469 9271 35533 9279
rect 35531 9269 35533 9271
rect 35469 9197 35533 9207
rect 35239 7890 35299 7900
rect 35239 7818 35299 7828
rect 33923 6701 34807 6707
rect 33923 6597 33932 6701
rect 34019 6696 34807 6701
rect 34019 6600 34729 6696
rect 34806 6600 34807 6696
rect 35461 6694 35523 6696
rect 35461 6686 35525 6694
rect 35523 6684 35525 6686
rect 35461 6612 35525 6622
rect 34019 6597 34807 6600
rect 33923 6590 34807 6597
rect 33932 6587 34019 6590
rect 33218 1048 33852 1049
rect 33218 1038 33861 1048
rect 33218 957 33774 1038
rect 33218 947 33861 957
rect 34114 1040 34217 1050
rect 34114 951 34217 961
rect 33218 946 33852 947
rect 30689 832 33173 842
rect 30689 778 33108 832
rect 33164 778 33173 832
rect 30689 767 33173 778
rect 30689 747 30769 767
rect 30503 738 30569 744
rect 30689 687 30703 747
rect 30755 687 30769 747
rect 30689 676 30769 687
rect 1516 168 1592 178
rect 1516 100 1592 110
rect 4660 168 4736 178
rect 4660 100 4736 110
rect 7792 172 7868 182
rect 7792 104 7868 114
rect 10936 172 11012 182
rect 10936 104 11012 114
rect 14138 168 14214 178
rect 14138 100 14214 110
rect 17282 168 17358 178
rect 17282 100 17358 110
rect 20414 172 20490 182
rect 20414 104 20490 114
rect 23558 172 23634 182
rect 23558 104 23634 114
rect 29683 -136 29693 -58
rect 29763 -136 29773 -58
rect -310 -155 -142 -140
rect -550 -314 -446 -307
rect -575 -317 -430 -314
rect -575 -479 -550 -317
rect -446 -380 -430 -317
rect -310 -317 -285 -155
rect -181 -248 -142 -155
rect -181 -317 22136 -248
rect -446 -450 -428 -380
rect -310 -403 22136 -317
rect -310 -404 -142 -403
rect -446 -479 18988 -450
rect -575 -490 18988 -479
rect -813 -604 -663 -592
rect -813 -766 -792 -604
rect -688 -656 -663 -604
rect -575 -613 18986 -490
rect 18871 -647 18986 -613
rect -688 -766 15858 -656
rect -813 -786 15858 -766
rect 1528 -1480 1628 -1470
rect 1528 -1582 1628 -1572
rect 4672 -1480 4772 -1470
rect 4672 -1582 4772 -1572
rect 7804 -1476 7904 -1466
rect 7804 -1578 7904 -1568
rect 10948 -1476 11048 -1466
rect 10948 -1578 11048 -1568
rect 14150 -1480 14250 -1470
rect 14150 -1582 14250 -1572
rect 6425 -2437 6482 -2436
rect 6658 -2437 6751 -2435
rect 9569 -2437 9626 -2436
rect 9802 -2437 9895 -2435
rect 6417 -2438 7833 -2437
rect 9561 -2438 10977 -2437
rect 149 -2441 206 -2440
rect 382 -2441 475 -2439
rect 3293 -2441 3350 -2440
rect 3526 -2441 3619 -2439
rect 141 -2442 1557 -2441
rect 3285 -2442 4701 -2441
rect 138 -2450 1557 -2442
rect 138 -2518 149 -2450
rect 206 -2451 1557 -2450
rect 206 -2514 393 -2451
rect 464 -2513 1478 -2451
rect 1548 -2513 1557 -2451
rect 464 -2514 1557 -2513
rect 206 -2518 1557 -2514
rect 138 -2525 1557 -2518
rect 3282 -2450 4701 -2442
rect 3282 -2518 3293 -2450
rect 3350 -2451 4701 -2450
rect 3350 -2514 3537 -2451
rect 3608 -2513 4622 -2451
rect 4692 -2513 4701 -2451
rect 3608 -2514 4701 -2513
rect 3350 -2518 4701 -2514
rect 3282 -2525 4701 -2518
rect 6414 -2446 7833 -2438
rect 6414 -2514 6425 -2446
rect 6482 -2447 7833 -2446
rect 6482 -2510 6669 -2447
rect 6740 -2509 7754 -2447
rect 7824 -2509 7833 -2447
rect 6740 -2510 7833 -2509
rect 6482 -2514 7833 -2510
rect 6414 -2521 7833 -2514
rect 9558 -2446 10977 -2438
rect 12771 -2441 12828 -2440
rect 13004 -2441 13097 -2439
rect 12763 -2442 14179 -2441
rect 9558 -2514 9569 -2446
rect 9626 -2447 10977 -2446
rect 9626 -2510 9813 -2447
rect 9884 -2509 10898 -2447
rect 10968 -2509 10977 -2447
rect 9884 -2510 10977 -2509
rect 9626 -2514 10977 -2510
rect 9558 -2521 10977 -2514
rect 12760 -2450 14179 -2442
rect 12760 -2518 12771 -2450
rect 12828 -2451 14179 -2450
rect 12828 -2514 13015 -2451
rect 13086 -2513 14100 -2451
rect 14170 -2513 14179 -2451
rect 13086 -2514 14179 -2513
rect 12828 -2518 14179 -2514
rect 6414 -2522 6492 -2521
rect 9558 -2522 9636 -2521
rect 6425 -2524 6482 -2522
rect 9569 -2524 9626 -2522
rect 12760 -2525 14179 -2518
rect 138 -2526 216 -2525
rect 3282 -2526 3360 -2525
rect 12760 -2526 12838 -2525
rect 149 -2528 206 -2526
rect 3293 -2528 3350 -2526
rect 12771 -2528 12828 -2526
rect 6425 -2554 6482 -2552
rect 9569 -2554 9626 -2552
rect 149 -2558 206 -2556
rect 3293 -2558 3350 -2556
rect 6414 -2557 6510 -2554
rect 9558 -2557 9654 -2554
rect 138 -2561 234 -2558
rect 3282 -2561 3378 -2558
rect 138 -2566 1778 -2561
rect 138 -2634 149 -2566
rect 206 -2571 1778 -2566
rect 206 -2631 1719 -2571
rect 206 -2634 1778 -2631
rect 138 -2640 1778 -2634
rect 138 -2643 234 -2640
rect 1719 -2641 1778 -2640
rect 3282 -2566 4922 -2561
rect 3282 -2634 3293 -2566
rect 3350 -2571 4922 -2566
rect 3350 -2631 4863 -2571
rect 3350 -2634 4922 -2631
rect 3282 -2640 4922 -2634
rect 6414 -2562 8054 -2557
rect 6414 -2630 6425 -2562
rect 6482 -2567 8054 -2562
rect 6482 -2627 7995 -2567
rect 6482 -2630 8054 -2627
rect 6414 -2636 8054 -2630
rect 6414 -2639 6510 -2636
rect 7995 -2637 8054 -2636
rect 9558 -2562 11198 -2557
rect 12771 -2558 12828 -2556
rect 9558 -2630 9569 -2562
rect 9626 -2567 11198 -2562
rect 9626 -2627 11139 -2567
rect 9626 -2630 11198 -2627
rect 9558 -2636 11198 -2630
rect 9558 -2639 9654 -2636
rect 11139 -2637 11198 -2636
rect 12760 -2561 12856 -2558
rect 12760 -2566 14400 -2561
rect 12760 -2634 12771 -2566
rect 12828 -2571 14400 -2566
rect 12828 -2631 14341 -2571
rect 12828 -2634 14400 -2631
rect 6425 -2640 6482 -2639
rect 9569 -2640 9626 -2639
rect 12760 -2640 14400 -2634
rect 3282 -2643 3378 -2640
rect 4863 -2641 4922 -2640
rect 12760 -2643 12856 -2640
rect 14341 -2641 14400 -2640
rect 149 -2644 206 -2643
rect 3293 -2644 3350 -2643
rect 12771 -2644 12828 -2643
rect -172 -2718 -63 -2697
rect -172 -2796 -165 -2718
rect -77 -2725 -63 -2718
rect 6309 -2723 6500 -2722
rect 6546 -2723 7715 -2722
rect -77 -2726 265 -2725
rect 3179 -2726 3397 -2724
rect -77 -2734 1439 -2726
rect -77 -2796 1360 -2734
rect -172 -2799 1360 -2796
rect 1428 -2799 1439 -2734
rect -172 -2810 1439 -2799
rect 3179 -2734 4583 -2726
rect 3179 -2798 3188 -2734
rect 3249 -2798 4504 -2734
rect 3179 -2799 4504 -2798
rect 4572 -2799 4583 -2734
rect 3179 -2810 4583 -2799
rect 6309 -2730 7715 -2723
rect 6309 -2737 7636 -2730
rect 6309 -2800 6318 -2737
rect 6401 -2795 7636 -2737
rect 7704 -2795 7715 -2730
rect 6401 -2800 7715 -2795
rect 6309 -2806 7715 -2800
rect 9453 -2730 10859 -2722
rect 12693 -2726 12758 -2720
rect 15745 -2726 15857 -786
rect 17294 -1480 17394 -1470
rect 17294 -1582 17394 -1572
rect 15915 -2441 15972 -2440
rect 16148 -2441 16241 -2439
rect 15907 -2442 17323 -2441
rect 15904 -2450 17323 -2442
rect 15904 -2518 15915 -2450
rect 15972 -2451 17323 -2450
rect 15972 -2514 16159 -2451
rect 16230 -2513 17244 -2451
rect 17314 -2513 17323 -2451
rect 16230 -2514 17323 -2513
rect 15972 -2518 17323 -2514
rect 15904 -2525 17323 -2518
rect 15904 -2526 15982 -2525
rect 15915 -2528 15972 -2526
rect 15915 -2558 15972 -2556
rect 15904 -2561 16000 -2558
rect 15904 -2566 17544 -2561
rect 15904 -2634 15915 -2566
rect 15972 -2571 17544 -2566
rect 15972 -2631 17485 -2571
rect 15972 -2634 17544 -2631
rect 15904 -2640 17544 -2634
rect 15904 -2643 16000 -2640
rect 17485 -2641 17544 -2640
rect 15915 -2644 15972 -2643
rect 18871 -2720 18988 -647
rect 20426 -1476 20526 -1466
rect 20426 -1578 20526 -1568
rect 19047 -2437 19104 -2436
rect 19280 -2437 19373 -2435
rect 19039 -2438 20455 -2437
rect 19036 -2446 20455 -2438
rect 19036 -2514 19047 -2446
rect 19104 -2447 20455 -2446
rect 19104 -2510 19291 -2447
rect 19362 -2509 20376 -2447
rect 20446 -2509 20455 -2447
rect 19362 -2510 20455 -2509
rect 19104 -2514 20455 -2510
rect 19036 -2521 20455 -2514
rect 19036 -2522 19114 -2521
rect 19047 -2524 19104 -2522
rect 19047 -2554 19104 -2552
rect 19036 -2557 19132 -2554
rect 19036 -2562 20676 -2557
rect 19036 -2630 19047 -2562
rect 19104 -2567 20676 -2562
rect 19104 -2627 20617 -2567
rect 19104 -2630 20676 -2627
rect 19036 -2636 20676 -2630
rect 19036 -2639 19132 -2636
rect 20617 -2637 20676 -2636
rect 19047 -2640 19104 -2639
rect 18871 -2722 19156 -2720
rect 22006 -2722 22134 -403
rect 30503 -650 30569 672
rect 31913 -78 31923 -6
rect 31993 -78 32003 -6
rect 30503 -704 30509 -650
rect 30563 -704 30569 -650
rect 31067 -891 31157 -881
rect 31067 -988 31157 -978
rect 33108 -1221 33164 -1220
rect 30688 -1230 33173 -1221
rect 30688 -1284 33108 -1230
rect 33164 -1284 33173 -1230
rect 30688 -1296 33173 -1284
rect 30688 -1318 30769 -1296
rect 30501 -1330 30567 -1324
rect 30688 -1383 30698 -1318
rect 30757 -1383 30769 -1318
rect 30688 -1388 30769 -1383
rect 30698 -1393 30757 -1388
rect 23570 -1476 23670 -1466
rect 23570 -1578 23670 -1568
rect 29681 -2204 29691 -2126
rect 29761 -2204 29771 -2126
rect 22191 -2437 22248 -2436
rect 22424 -2437 22517 -2435
rect 22183 -2438 23599 -2437
rect 22180 -2446 23599 -2438
rect 22180 -2514 22191 -2446
rect 22248 -2447 23599 -2446
rect 22248 -2510 22435 -2447
rect 22506 -2509 23520 -2447
rect 23590 -2509 23599 -2447
rect 22506 -2510 23599 -2509
rect 22248 -2514 23599 -2510
rect 22180 -2521 23599 -2514
rect 22180 -2522 22258 -2521
rect 22191 -2524 22248 -2522
rect 22191 -2554 22248 -2552
rect 22180 -2557 22276 -2554
rect 22180 -2562 23820 -2557
rect 22180 -2630 22191 -2562
rect 22248 -2567 23820 -2562
rect 22248 -2627 23761 -2567
rect 22248 -2630 23820 -2627
rect 22180 -2636 23820 -2630
rect 22180 -2639 22276 -2636
rect 23761 -2637 23820 -2636
rect 22191 -2640 22248 -2639
rect 30501 -2718 30567 -1396
rect 31911 -2146 31921 -2074
rect 31991 -2146 32001 -2074
rect 34250 -2311 34368 6590
rect 35220 4612 35280 4622
rect 35220 4540 35280 4550
rect 35442 3416 35504 3418
rect 35442 3408 35506 3416
rect 35504 3406 35506 3408
rect 35442 3334 35506 3344
rect 35236 1852 35296 1862
rect 35236 1780 35296 1790
rect 35458 656 35520 658
rect 35458 648 35522 656
rect 35520 646 35522 648
rect 35458 574 35522 584
rect 34250 -2397 34260 -2311
rect 34359 -2397 34368 -2311
rect 34250 -2405 34368 -2397
rect 34260 -2407 34359 -2405
rect 9453 -2737 10780 -2730
rect 9453 -2798 9462 -2737
rect 9581 -2795 10780 -2737
rect 10848 -2795 10859 -2730
rect 9581 -2798 10859 -2795
rect 9453 -2806 10859 -2798
rect 12691 -2730 14061 -2726
rect 6309 -2807 6562 -2806
rect 6318 -2810 6401 -2807
rect 9462 -2808 9581 -2806
rect -172 -2811 -63 -2810
rect 12691 -2811 12693 -2730
rect 12758 -2734 14061 -2730
rect 12758 -2799 13982 -2734
rect 14050 -2799 14061 -2734
rect 15745 -2734 17205 -2726
rect 15745 -2780 17126 -2734
rect 12758 -2810 14061 -2799
rect 15746 -2799 17126 -2780
rect 17194 -2799 17205 -2734
rect 15746 -2810 17205 -2799
rect 18871 -2730 20337 -2722
rect 18871 -2795 20258 -2730
rect 20326 -2795 20337 -2730
rect 18871 -2806 20337 -2795
rect 22006 -2730 23481 -2722
rect 22006 -2795 23402 -2730
rect 23470 -2795 23481 -2730
rect 30501 -2772 30507 -2718
rect 30561 -2772 30567 -2718
rect 22006 -2806 23481 -2795
rect 18871 -2807 19156 -2806
rect 12758 -2811 12905 -2810
rect 12693 -2821 12758 -2811
rect 15746 -2812 16043 -2810
rect 36213 -2877 36320 10787
rect 66535 10786 67892 10796
rect 36361 10755 52520 10757
rect 62994 10755 63055 10756
rect 36361 10735 63086 10755
rect 36361 10681 48116 10735
rect 48173 10681 63086 10735
rect 36361 10662 63086 10681
rect 36361 10661 59345 10662
rect 36362 -2199 36480 10661
rect 62994 10535 63086 10662
rect 67590 10624 67652 10626
rect 67590 10616 67654 10624
rect 67652 10614 67654 10616
rect 67590 10542 67654 10552
rect 47257 10421 47410 10431
rect 44775 10367 44928 10377
rect 40708 10333 40861 10343
rect 38226 10279 38379 10289
rect 41855 10333 42008 10343
rect 41120 10238 41176 10248
rect 40708 10194 40861 10204
rect 38226 10140 38379 10150
rect 40995 10172 41120 10234
rect 41176 10172 41177 10234
rect 48404 10421 48557 10431
rect 47669 10326 47725 10336
rect 47257 10282 47410 10292
rect 44775 10228 44928 10238
rect 47544 10260 47669 10322
rect 47725 10260 47726 10322
rect 60536 10421 60689 10431
rect 58054 10367 58207 10377
rect 53911 10353 54064 10363
rect 48404 10282 48557 10292
rect 51429 10299 51582 10309
rect 46539 10211 46605 10214
rect 41855 10194 42008 10204
rect 45613 10204 46605 10211
rect 39990 10123 40056 10126
rect 39064 10116 40056 10123
rect 39064 10050 39990 10116
rect 38497 9087 38507 9240
rect 38636 9087 38646 9240
rect 36997 8652 37164 8653
rect 37504 8652 37620 8653
rect 36997 8642 37620 8652
rect 36997 8625 37503 8642
rect 36997 8519 37009 8625
rect 37121 8536 37503 8625
rect 37615 8536 37620 8642
rect 37121 8519 37620 8536
rect 36997 8510 37620 8519
rect 38240 8629 38393 8639
rect 38240 8490 38393 8500
rect 36996 7531 37161 7541
rect 36996 7530 37164 7531
rect 37786 7530 37904 7533
rect 36996 7523 37904 7530
rect 36996 7513 37786 7523
rect 36996 7407 37008 7513
rect 37120 7511 37786 7513
rect 36996 7405 37014 7407
rect 37126 7405 37786 7511
rect 38511 7437 38521 7590
rect 38650 7437 38660 7590
rect 36996 7398 37904 7405
rect 37002 7396 37904 7398
rect 37039 7395 37904 7396
rect 37273 7151 37388 7161
rect 37273 7044 37388 7054
rect 37783 5744 37899 7395
rect 38235 7025 38388 7035
rect 38235 6886 38388 6896
rect 38833 6267 38896 6273
rect 39064 6267 39132 10050
rect 39990 10040 40056 10050
rect 40995 9511 41055 10172
rect 41120 10162 41176 10172
rect 40917 9510 41055 9511
rect 40655 9500 41055 9510
rect 40655 9403 40656 9500
rect 40755 9403 41055 9500
rect 45613 10138 46539 10204
rect 41812 9489 41877 9490
rect 42907 9489 43121 9499
rect 41811 9480 42945 9489
rect 41811 9426 41812 9480
rect 41877 9426 42945 9480
rect 41811 9415 42945 9426
rect 40655 9395 41055 9403
rect 42907 9414 42945 9415
rect 43090 9414 43121 9489
rect 42907 9401 43121 9414
rect 40655 9391 40964 9395
rect 45046 9175 45056 9328
rect 45185 9175 45195 9328
rect 40055 8932 40208 8942
rect 40055 8793 40208 8803
rect 41197 8930 41350 8940
rect 41197 8791 41350 8801
rect 43546 8740 43713 8741
rect 44053 8740 44169 8741
rect 43546 8730 44169 8740
rect 43546 8713 44052 8730
rect 43546 8607 43558 8713
rect 43670 8624 44052 8713
rect 44164 8624 44169 8730
rect 43670 8607 44169 8624
rect 43546 8598 44169 8607
rect 44789 8717 44942 8727
rect 44789 8578 44942 8588
rect 40053 8286 40206 8296
rect 40053 8147 40206 8157
rect 41951 8286 42104 8296
rect 41951 8147 42104 8157
rect 44335 7618 44453 7621
rect 43543 7611 44453 7618
rect 43543 7493 44335 7611
rect 45060 7525 45070 7678
rect 45199 7525 45209 7678
rect 43543 7483 44453 7493
rect 40694 7315 40772 7325
rect 40694 7219 40772 7229
rect 38828 6263 39132 6267
rect 38828 6211 38833 6263
rect 38896 6211 39132 6263
rect 38828 6205 39132 6211
rect 38833 6201 38896 6205
rect 38506 5833 38516 5986
rect 38645 5833 38655 5986
rect 39999 5889 40152 5899
rect 39999 5750 40152 5760
rect 41897 5889 42050 5899
rect 41897 5750 42050 5760
rect 37783 5734 37900 5744
rect 37783 5628 37788 5734
rect 37783 5618 37900 5628
rect 37783 5617 37899 5618
rect 43543 5299 43709 7483
rect 43822 7239 43937 7249
rect 43822 7132 43937 7142
rect 44332 5832 44448 7483
rect 44784 7113 44937 7123
rect 44784 6974 44937 6984
rect 45382 6355 45445 6361
rect 45613 6355 45681 10138
rect 46539 10128 46605 10138
rect 47544 9599 47604 10260
rect 47669 10250 47725 10260
rect 55058 10353 55211 10363
rect 54323 10258 54379 10268
rect 53911 10214 54064 10224
rect 51429 10160 51582 10170
rect 54198 10192 54323 10254
rect 54379 10192 54380 10254
rect 61683 10421 61836 10431
rect 60948 10326 61004 10336
rect 60536 10282 60689 10292
rect 58054 10228 58207 10238
rect 60823 10260 60948 10322
rect 61004 10260 61005 10322
rect 61683 10282 61836 10292
rect 55058 10214 55211 10224
rect 59818 10211 59884 10214
rect 58892 10204 59884 10211
rect 53193 10143 53259 10146
rect 47466 9598 47604 9599
rect 47204 9588 47604 9598
rect 47204 9491 47205 9588
rect 47304 9491 47604 9588
rect 52267 10136 53259 10143
rect 52267 10070 53193 10136
rect 48361 9577 48426 9578
rect 49456 9577 49524 9587
rect 48360 9568 49456 9577
rect 48360 9514 48361 9568
rect 48426 9514 49456 9568
rect 48360 9503 49456 9514
rect 49456 9492 49524 9502
rect 47204 9483 47604 9491
rect 47204 9479 47513 9483
rect 51700 9107 51710 9260
rect 51839 9107 51849 9260
rect 46604 9020 46757 9030
rect 46604 8881 46757 8891
rect 47746 9018 47899 9028
rect 47746 8879 47899 8889
rect 49525 8672 50469 8675
rect 50707 8672 50823 8673
rect 49525 8662 50823 8672
rect 49525 8556 50706 8662
rect 50818 8556 50823 8662
rect 49525 8530 50823 8556
rect 51443 8649 51596 8659
rect 46602 8374 46755 8384
rect 46602 8235 46755 8245
rect 48500 8374 48653 8384
rect 48500 8235 48653 8245
rect 47243 7403 47321 7413
rect 47243 7307 47321 7317
rect 49525 6890 49645 8530
rect 51443 8510 51596 8520
rect 50199 7551 50364 7561
rect 50199 7550 50367 7551
rect 50989 7550 51107 7553
rect 50199 7543 51107 7550
rect 50199 7533 50989 7543
rect 50199 7427 50211 7533
rect 50323 7531 50989 7533
rect 50199 7425 50217 7427
rect 50329 7425 50989 7531
rect 51714 7457 51724 7610
rect 51853 7457 51863 7610
rect 50199 7418 51107 7425
rect 50205 7416 51107 7418
rect 50242 7415 51107 7416
rect 50476 7171 50591 7181
rect 50476 7064 50591 7074
rect 49525 6791 49645 6801
rect 45377 6351 45681 6355
rect 45377 6299 45382 6351
rect 45445 6299 45681 6351
rect 45377 6293 45681 6299
rect 45382 6289 45445 6293
rect 45055 5921 45065 6074
rect 45194 5921 45204 6074
rect 46548 5977 46701 5987
rect 46548 5838 46701 5848
rect 48446 5977 48599 5987
rect 48446 5838 48599 5848
rect 44332 5822 44449 5832
rect 44332 5716 44337 5822
rect 44332 5706 44449 5716
rect 50986 5764 51102 7415
rect 51438 7045 51591 7055
rect 51438 6906 51591 6916
rect 52036 6287 52099 6293
rect 52267 6287 52335 10070
rect 53193 10060 53259 10070
rect 54198 9531 54258 10192
rect 54323 10182 54379 10192
rect 54120 9530 54258 9531
rect 53858 9520 54258 9530
rect 53858 9423 53859 9520
rect 53958 9423 54258 9520
rect 58892 10138 59818 10204
rect 55015 9509 55080 9510
rect 56079 9509 56176 9519
rect 55014 9500 56079 9509
rect 55014 9446 55015 9500
rect 55080 9446 56079 9500
rect 55014 9435 56079 9446
rect 56176 9435 56177 9509
rect 56079 9425 56176 9435
rect 53858 9415 54258 9423
rect 53858 9411 54167 9415
rect 58325 9175 58335 9328
rect 58464 9175 58474 9328
rect 53258 8952 53411 8962
rect 53258 8813 53411 8823
rect 54400 8950 54553 8960
rect 54400 8811 54553 8821
rect 56825 8740 56992 8741
rect 57332 8740 57448 8741
rect 56825 8730 57448 8740
rect 56825 8713 57331 8730
rect 56825 8607 56837 8713
rect 56949 8624 57331 8713
rect 57443 8624 57448 8730
rect 56949 8607 57448 8624
rect 56825 8598 57448 8607
rect 58068 8717 58221 8727
rect 58068 8578 58221 8588
rect 53256 8306 53409 8316
rect 53256 8167 53409 8177
rect 55154 8306 55307 8316
rect 55154 8167 55307 8177
rect 57614 7618 57732 7621
rect 56851 7611 57732 7618
rect 56851 7493 57614 7611
rect 58339 7525 58349 7678
rect 58478 7525 58488 7678
rect 56851 7484 57732 7493
rect 53897 7335 53975 7345
rect 53897 7239 53975 7249
rect 56632 6824 56728 6834
rect 56632 6714 56728 6724
rect 52031 6283 52335 6287
rect 52031 6231 52036 6283
rect 52099 6231 52335 6283
rect 52031 6225 52335 6231
rect 52036 6221 52099 6225
rect 51709 5853 51719 6006
rect 51848 5853 51858 6006
rect 53202 5909 53355 5919
rect 53202 5770 53355 5780
rect 55100 5909 55253 5919
rect 55100 5770 55253 5780
rect 50986 5754 51103 5764
rect 44332 5705 44448 5706
rect 50986 5648 50991 5754
rect 50986 5638 51103 5648
rect 50986 5637 51102 5638
rect 56152 5520 56294 5530
rect 56152 5377 56294 5386
rect 43543 5153 49457 5299
rect 43632 5148 49457 5153
rect 56852 5277 56962 7484
rect 56993 7483 57732 7484
rect 57101 7239 57216 7249
rect 57101 7132 57216 7142
rect 57611 5832 57727 7483
rect 58063 7113 58216 7123
rect 58063 6974 58216 6984
rect 58661 6355 58724 6361
rect 58892 6355 58960 10138
rect 59818 10128 59884 10138
rect 60823 9599 60883 10260
rect 60948 10250 61004 10260
rect 60745 9598 60883 9599
rect 60483 9588 60883 9598
rect 60483 9491 60484 9588
rect 60583 9491 60883 9588
rect 61640 9577 61705 9578
rect 62618 9577 62686 9587
rect 61639 9568 62618 9577
rect 61639 9514 61640 9568
rect 61705 9514 62618 9568
rect 61639 9503 62618 9514
rect 62618 9492 62686 9502
rect 60483 9483 60883 9491
rect 60483 9479 60792 9483
rect 59883 9020 60036 9030
rect 59883 8881 60036 8891
rect 61025 9018 61178 9028
rect 61025 8879 61178 8889
rect 62994 8725 63085 10535
rect 65935 9838 66146 9848
rect 65935 9671 66146 9681
rect 63762 9657 63822 9667
rect 63762 9585 63822 9595
rect 62994 8714 63493 8725
rect 62994 8633 63411 8714
rect 62994 8624 63493 8633
rect 63411 8623 63493 8624
rect 63984 8461 64046 8463
rect 63984 8453 64048 8461
rect 64046 8451 64048 8453
rect 59881 8374 60034 8384
rect 59881 8235 60034 8245
rect 61779 8374 61932 8384
rect 63984 8379 64048 8389
rect 61779 8235 61932 8245
rect 66015 8077 66168 8087
rect 66015 7938 66168 7948
rect 67370 7729 67430 7739
rect 67370 7657 67430 7667
rect 60522 7403 60600 7413
rect 60522 7307 60600 7317
rect 65223 7157 65290 7162
rect 65216 7152 66932 7157
rect 65216 7089 65223 7152
rect 65290 7147 66932 7152
rect 65290 7091 66879 7147
rect 65290 7089 66932 7091
rect 65216 7081 66932 7089
rect 65223 7079 65290 7081
rect 67003 7044 67076 7054
rect 65223 7035 65290 7036
rect 65483 7035 67003 7044
rect 65215 7034 67003 7035
rect 65215 7026 65483 7034
rect 65215 6963 65223 7026
rect 65290 6966 65483 7026
rect 65538 6966 67003 7034
rect 65290 6963 67003 6966
rect 65215 6956 67003 6963
rect 65216 6955 65305 6956
rect 65223 6953 65290 6955
rect 67003 6945 67076 6955
rect 68233 6807 68333 19076
rect 68767 19071 68873 22120
rect 71202 21971 71286 22120
rect 71319 22119 71404 22147
rect 71486 22119 71571 22147
rect 71200 21960 71286 21971
rect 71200 21889 71212 21960
rect 71275 21889 71286 21960
rect 71200 21878 71286 21889
rect 71202 20875 71286 21878
rect 70231 20725 70241 20825
rect 70333 20725 70343 20825
rect 71202 20805 71212 20875
rect 71274 20805 71286 20875
rect 71202 20796 71286 20805
rect 71322 20634 71401 22119
rect 71487 20993 71571 22119
rect 71487 20925 71495 20993
rect 71560 20925 71571 20993
rect 71487 20914 71571 20925
rect 72475 20729 72485 20805
rect 72543 20729 72553 20805
rect 71322 20575 71332 20634
rect 71392 20575 71402 20634
rect 68767 18992 71287 19071
rect 71319 19060 71404 19071
rect 71486 19060 71571 19071
rect 71317 19003 71327 19060
rect 71395 19003 71405 19060
rect 71485 19003 71495 19060
rect 71563 19003 71573 19060
rect 68767 15939 68873 18992
rect 71202 18948 71287 18992
rect 71319 18975 71404 19003
rect 71486 18975 71571 19003
rect 71202 18827 71286 18948
rect 71200 18816 71286 18827
rect 71200 18745 71212 18816
rect 71275 18745 71286 18816
rect 71200 18734 71286 18745
rect 71202 17731 71286 18734
rect 70231 17581 70241 17681
rect 70333 17581 70343 17681
rect 71202 17661 71212 17731
rect 71274 17661 71286 17731
rect 71202 17652 71286 17661
rect 71322 17490 71401 18975
rect 71487 17849 71571 18975
rect 71487 17781 71495 17849
rect 71560 17781 71571 17849
rect 71487 17770 71571 17781
rect 72475 17585 72485 17661
rect 72543 17585 72553 17661
rect 71322 17431 71332 17490
rect 71392 17431 71402 17490
rect 68767 15860 71282 15939
rect 71315 15928 71400 15939
rect 71482 15928 71567 15939
rect 71313 15871 71323 15928
rect 71391 15871 71401 15928
rect 71481 15871 71491 15928
rect 71559 15871 71569 15928
rect 68767 12877 68873 15860
rect 71198 15695 71282 15860
rect 71315 15843 71400 15871
rect 71482 15843 71567 15871
rect 71196 15684 71282 15695
rect 71196 15613 71208 15684
rect 71271 15613 71282 15684
rect 71196 15602 71282 15613
rect 71198 14599 71282 15602
rect 70227 14449 70237 14549
rect 70329 14449 70339 14549
rect 71198 14529 71208 14599
rect 71270 14529 71282 14599
rect 71198 14520 71282 14529
rect 71318 14358 71397 15843
rect 71483 14717 71567 15843
rect 71483 14649 71491 14717
rect 71556 14649 71567 14717
rect 71483 14638 71567 14649
rect 72471 14453 72481 14529
rect 72539 14453 72549 14529
rect 71318 14299 71328 14358
rect 71388 14299 71398 14358
rect 68478 12865 68873 12877
rect 68478 12784 68502 12865
rect 68646 12797 68873 12865
rect 68646 12784 71283 12797
rect 71315 12784 71400 12795
rect 71483 12788 71567 12798
rect 68478 12774 71283 12784
rect 68478 12773 68728 12774
rect 67716 6806 68333 6807
rect 66537 6796 68333 6806
rect 66599 6705 68333 6796
rect 66537 6695 68333 6705
rect 68115 6694 68333 6695
rect 68767 12717 71283 12774
rect 71313 12727 71323 12784
rect 71391 12727 71401 12784
rect 68767 9593 68873 12717
rect 71197 12682 71283 12717
rect 71315 12699 71400 12727
rect 71198 12551 71282 12682
rect 71196 12540 71282 12551
rect 71196 12469 71208 12540
rect 71271 12469 71282 12540
rect 71196 12458 71282 12469
rect 71198 11455 71282 12458
rect 70227 11305 70237 11405
rect 70329 11305 70339 11405
rect 71198 11385 71208 11455
rect 71270 11385 71282 11455
rect 71198 11376 71282 11385
rect 71318 11214 71397 12699
rect 71483 12691 71494 12788
rect 71557 12691 71567 12788
rect 71483 11573 71567 12691
rect 71483 11505 71491 11573
rect 71556 11505 71567 11573
rect 71483 11494 71567 11505
rect 72471 11309 72481 11385
rect 72539 11309 72549 11385
rect 71318 11155 71328 11214
rect 71388 11155 71398 11214
rect 68767 9515 71286 9593
rect 71319 9582 71404 9593
rect 71486 9582 71571 9593
rect 71317 9525 71327 9582
rect 71395 9525 71405 9582
rect 71485 9525 71495 9582
rect 71563 9525 71573 9582
rect 63762 6624 63822 6634
rect 63762 6552 63822 6562
rect 67592 6533 67654 6535
rect 67592 6525 67656 6533
rect 67654 6523 67656 6525
rect 67592 6451 67656 6461
rect 58656 6351 58960 6355
rect 58656 6299 58661 6351
rect 58724 6299 58960 6351
rect 58656 6293 58960 6299
rect 68767 6449 68873 9515
rect 71202 9349 71286 9515
rect 71319 9497 71404 9525
rect 71486 9497 71571 9525
rect 71200 9338 71286 9349
rect 71200 9267 71212 9338
rect 71275 9267 71286 9338
rect 71200 9256 71286 9267
rect 71202 8253 71286 9256
rect 70231 8103 70241 8203
rect 70333 8103 70343 8203
rect 71202 8183 71212 8253
rect 71274 8183 71286 8253
rect 71202 8174 71286 8183
rect 71322 8012 71401 9497
rect 71487 8371 71571 9497
rect 71487 8303 71495 8371
rect 71560 8303 71571 8371
rect 71487 8292 71571 8303
rect 72475 8107 72485 8183
rect 72543 8107 72553 8183
rect 71322 7953 71332 8012
rect 71392 7953 71402 8012
rect 68767 6371 71287 6449
rect 71319 6438 71404 6449
rect 71486 6441 71572 6452
rect 71317 6381 71327 6438
rect 71395 6381 71405 6438
rect 58661 6289 58724 6293
rect 58334 5921 58344 6074
rect 58473 5921 58483 6074
rect 59827 5977 59980 5987
rect 59827 5838 59980 5848
rect 61725 5977 61878 5987
rect 61725 5838 61878 5848
rect 57611 5822 57728 5832
rect 57611 5716 57616 5822
rect 63516 5814 63605 5823
rect 57611 5706 57728 5716
rect 63000 5813 63605 5814
rect 63000 5726 63516 5813
rect 63000 5722 63605 5726
rect 57611 5705 57727 5706
rect 57261 5520 57403 5530
rect 57261 5376 57403 5386
rect 40700 4553 40853 4563
rect 38218 4499 38371 4509
rect 41847 4553 42000 4563
rect 41112 4458 41168 4468
rect 40700 4414 40853 4424
rect 38218 4360 38371 4370
rect 40987 4392 41112 4454
rect 41168 4392 41169 4454
rect 47251 4551 47404 4561
rect 41847 4414 42000 4424
rect 44769 4497 44922 4507
rect 39982 4343 40048 4346
rect 39056 4336 40048 4343
rect 39056 4270 39982 4336
rect 38489 3307 38499 3460
rect 38628 3307 38638 3460
rect 36989 2872 37156 2873
rect 37496 2872 37612 2873
rect 36989 2862 37612 2872
rect 36989 2845 37495 2862
rect 36989 2739 37001 2845
rect 37113 2756 37495 2845
rect 37607 2756 37612 2862
rect 37113 2739 37612 2756
rect 36989 2730 37612 2739
rect 38232 2849 38385 2859
rect 38232 2710 38385 2720
rect 36885 1761 37119 1766
rect 36885 1756 37153 1761
rect 37119 1751 37153 1756
rect 37119 1750 37156 1751
rect 37778 1750 37896 1753
rect 37119 1743 37896 1750
rect 37119 1625 37778 1743
rect 38503 1657 38513 1810
rect 38642 1657 38652 1810
rect 37119 1619 37896 1625
rect 36885 1615 37896 1619
rect 36885 1609 37119 1615
rect 37265 1371 37380 1381
rect 37265 1264 37380 1274
rect 37775 -36 37891 1615
rect 38227 1245 38380 1255
rect 38227 1106 38380 1116
rect 38825 487 38888 493
rect 39056 487 39124 4270
rect 39982 4260 40048 4270
rect 40987 3731 41047 4392
rect 41112 4382 41168 4392
rect 48398 4551 48551 4561
rect 47663 4456 47719 4466
rect 47251 4412 47404 4422
rect 44769 4358 44922 4368
rect 47538 4390 47663 4452
rect 47719 4390 47720 4452
rect 48398 4412 48551 4422
rect 46533 4341 46599 4344
rect 40909 3730 41047 3731
rect 40647 3720 41047 3730
rect 40647 3623 40648 3720
rect 40747 3623 41047 3720
rect 45607 4334 46599 4341
rect 45607 4268 46533 4334
rect 41804 3709 41869 3710
rect 42899 3709 42967 3719
rect 41803 3700 42899 3709
rect 41803 3646 41804 3700
rect 41869 3646 42899 3700
rect 41803 3635 42899 3646
rect 42899 3624 42967 3634
rect 40647 3615 41047 3623
rect 40647 3611 40956 3615
rect 45040 3305 45050 3458
rect 45179 3305 45189 3458
rect 40047 3152 40200 3162
rect 40047 3013 40200 3023
rect 41189 3150 41342 3160
rect 41189 3011 41342 3021
rect 44047 2870 44163 2871
rect 43786 2867 44163 2870
rect 43540 2860 44163 2867
rect 43540 2843 44046 2860
rect 43540 2737 43552 2843
rect 43664 2754 44046 2843
rect 44158 2754 44163 2860
rect 43664 2737 44163 2754
rect 43540 2728 44163 2737
rect 44783 2847 44936 2857
rect 44783 2708 44936 2718
rect 40045 2506 40198 2516
rect 40045 2367 40198 2377
rect 41943 2506 42096 2516
rect 41943 2367 42096 2377
rect 43520 1749 43743 1759
rect 44329 1748 44447 1751
rect 43743 1741 44447 1748
rect 43743 1623 44329 1741
rect 45054 1655 45064 1808
rect 45193 1655 45203 1808
rect 43743 1613 44447 1623
rect 43520 1603 43743 1613
rect 40686 1535 40764 1545
rect 40686 1439 40764 1449
rect 43816 1369 43931 1379
rect 43816 1262 43931 1272
rect 38820 483 39124 487
rect 38820 431 38825 483
rect 38888 431 39124 483
rect 38820 425 39124 431
rect 38825 421 38888 425
rect 38498 53 38508 206
rect 38637 53 38647 206
rect 39991 109 40144 119
rect 39991 -30 40144 -20
rect 41889 109 42042 119
rect 41889 -30 42042 -20
rect 37775 -46 37892 -36
rect 37775 -152 37780 -46
rect 37775 -162 37892 -152
rect 44326 -38 44442 1613
rect 44778 1243 44931 1253
rect 44778 1104 44931 1114
rect 45376 485 45439 491
rect 45607 485 45675 4268
rect 46533 4258 46599 4268
rect 47538 3729 47598 4390
rect 47663 4380 47719 4390
rect 47460 3728 47598 3729
rect 47198 3718 47598 3728
rect 47198 3621 47199 3718
rect 47298 3621 47598 3718
rect 48355 3707 48420 3708
rect 49323 3707 49453 5148
rect 56852 5145 62761 5277
rect 56852 5144 56956 5145
rect 62632 5121 62761 5145
rect 62632 5032 62762 5121
rect 53906 4552 54059 4562
rect 51424 4498 51577 4508
rect 55053 4552 55206 4562
rect 54318 4457 54374 4467
rect 53906 4413 54059 4423
rect 51424 4359 51577 4369
rect 54193 4391 54318 4453
rect 54374 4391 54375 4453
rect 60528 4553 60681 4563
rect 55053 4413 55206 4423
rect 58046 4499 58199 4509
rect 53188 4342 53254 4345
rect 48354 3698 49453 3707
rect 48354 3644 48355 3698
rect 48420 3644 49453 3698
rect 48354 3633 49453 3644
rect 49323 3630 49453 3633
rect 52262 4335 53254 4342
rect 52262 4269 53188 4335
rect 47198 3613 47598 3621
rect 47198 3609 47507 3613
rect 51695 3306 51705 3459
rect 51834 3306 51844 3459
rect 46598 3150 46751 3160
rect 46598 3011 46751 3021
rect 47740 3148 47893 3158
rect 47740 3009 47893 3019
rect 50128 2872 50294 2874
rect 50128 2871 50362 2872
rect 50702 2871 50818 2872
rect 50128 2861 50818 2871
rect 50128 2849 50701 2861
rect 50128 2736 50140 2849
rect 50344 2755 50701 2849
rect 50813 2755 50818 2861
rect 50128 2735 50292 2736
rect 50344 2735 50818 2755
rect 50128 2729 50818 2735
rect 51438 2848 51591 2858
rect 50128 2728 50352 2729
rect 51438 2709 51591 2719
rect 46596 2504 46749 2514
rect 46596 2365 46749 2375
rect 48494 2504 48647 2514
rect 48494 2365 48647 2375
rect 50194 1750 50359 1760
rect 50194 1749 50362 1750
rect 50984 1749 51102 1752
rect 50194 1742 51102 1749
rect 50194 1734 50984 1742
rect 50194 1622 50201 1734
rect 50345 1624 50984 1734
rect 51709 1656 51719 1809
rect 51848 1656 51858 1809
rect 50345 1622 51102 1624
rect 50194 1617 51102 1622
rect 50200 1615 51102 1617
rect 50201 1614 51102 1615
rect 50201 1612 50345 1614
rect 47237 1533 47315 1543
rect 47237 1437 47315 1447
rect 50471 1370 50586 1380
rect 50471 1263 50586 1273
rect 45371 481 45675 485
rect 45371 429 45376 481
rect 45439 429 45675 481
rect 45371 423 45675 429
rect 45376 419 45439 423
rect 45049 51 45059 204
rect 45188 51 45198 204
rect 46542 107 46695 117
rect 46542 -32 46695 -22
rect 48440 107 48593 117
rect 48440 -32 48593 -22
rect 50981 -37 51097 1614
rect 51433 1244 51586 1254
rect 51433 1105 51586 1115
rect 52031 486 52094 492
rect 52262 486 52330 4269
rect 53188 4259 53254 4269
rect 54193 3730 54253 4391
rect 54318 4381 54374 4391
rect 61675 4553 61828 4563
rect 60940 4458 60996 4468
rect 60528 4414 60681 4424
rect 58046 4360 58199 4370
rect 60815 4392 60940 4454
rect 60996 4392 60997 4454
rect 61675 4414 61828 4424
rect 59810 4343 59876 4346
rect 54115 3729 54253 3730
rect 53853 3719 54253 3729
rect 53853 3622 53854 3719
rect 53953 3622 54253 3719
rect 58884 4336 59876 4343
rect 58884 4270 59810 4336
rect 55010 3708 55075 3709
rect 56105 3708 56173 3718
rect 55009 3699 56105 3708
rect 55009 3645 55010 3699
rect 55075 3645 56105 3699
rect 55009 3634 56105 3645
rect 56105 3623 56173 3633
rect 53853 3614 54253 3622
rect 53853 3610 54162 3614
rect 58317 3307 58327 3460
rect 58456 3307 58466 3460
rect 53253 3151 53406 3161
rect 53253 3012 53406 3022
rect 54395 3149 54548 3159
rect 54395 3010 54548 3020
rect 57324 2872 57440 2873
rect 56817 2862 57440 2872
rect 56817 2845 57323 2862
rect 56817 2739 56829 2845
rect 56941 2756 57323 2845
rect 57435 2756 57440 2862
rect 56941 2739 57440 2756
rect 56817 2730 57440 2739
rect 58060 2849 58213 2859
rect 58060 2710 58213 2720
rect 53251 2505 53404 2515
rect 53251 2366 53404 2376
rect 55149 2505 55302 2515
rect 55149 2366 55302 2376
rect 56816 1751 56981 1761
rect 56816 1750 56984 1751
rect 57606 1750 57724 1753
rect 56816 1743 57724 1750
rect 56816 1733 57606 1743
rect 56816 1627 56828 1733
rect 56940 1731 57606 1733
rect 56816 1625 56834 1627
rect 56946 1625 57606 1731
rect 58331 1657 58341 1810
rect 58470 1657 58480 1810
rect 56816 1618 57724 1625
rect 56822 1616 57724 1618
rect 56859 1615 57724 1616
rect 53892 1534 53970 1544
rect 53892 1438 53970 1448
rect 57093 1371 57208 1381
rect 57093 1264 57208 1274
rect 52026 482 52330 486
rect 52026 430 52031 482
rect 52094 430 52330 482
rect 52026 424 52330 430
rect 52031 420 52094 424
rect 51704 52 51714 205
rect 51843 52 51853 205
rect 53197 108 53350 118
rect 53197 -31 53350 -21
rect 55095 108 55248 118
rect 55095 -31 55248 -21
rect 57603 -36 57719 1615
rect 58055 1245 58208 1255
rect 58055 1106 58208 1116
rect 58653 487 58716 493
rect 58884 487 58952 4270
rect 59810 4260 59876 4270
rect 60815 3731 60875 4392
rect 60940 4382 60996 4392
rect 60737 3730 60875 3731
rect 60475 3720 60875 3730
rect 60475 3623 60476 3720
rect 60575 3623 60875 3720
rect 61632 3709 61697 3710
rect 62632 3709 62763 5032
rect 61631 3700 62763 3709
rect 61631 3646 61632 3700
rect 61697 3646 62763 3700
rect 61631 3635 62763 3646
rect 62632 3633 62763 3635
rect 62727 3632 62763 3633
rect 60475 3615 60875 3623
rect 60475 3611 60784 3615
rect 59875 3152 60028 3162
rect 59875 3013 60028 3023
rect 61017 3150 61170 3160
rect 61017 3011 61170 3021
rect 59873 2506 60026 2516
rect 59873 2367 60026 2377
rect 61771 2506 61924 2516
rect 61771 2367 61924 2377
rect 60514 1535 60592 1545
rect 60514 1439 60592 1449
rect 62787 1023 62919 1033
rect 62787 917 62919 927
rect 58648 483 58952 487
rect 58648 431 58653 483
rect 58716 431 58952 483
rect 63000 564 63097 5722
rect 63516 5716 63605 5722
rect 65937 5747 66148 5757
rect 65937 5580 66148 5590
rect 63984 5428 64046 5430
rect 63984 5420 64048 5428
rect 64046 5418 64048 5420
rect 63984 5346 64048 5356
rect 63833 4704 63893 4714
rect 63833 4632 63893 4642
rect 66015 4582 66168 4592
rect 66015 4443 66168 4453
rect 67370 4234 67430 4244
rect 67370 4162 67430 4172
rect 63568 3692 63654 3702
rect 65216 3669 65309 3673
rect 63568 3581 63654 3591
rect 65186 3663 65323 3669
rect 65186 3586 65216 3663
rect 65309 3662 65323 3663
rect 65309 3652 66932 3662
rect 65309 3596 66879 3652
rect 65309 3586 66932 3596
rect 65186 3579 65323 3586
rect 65216 3576 65309 3579
rect 67003 3549 67076 3559
rect 65223 3540 65290 3541
rect 65483 3540 67003 3549
rect 65215 3539 67003 3540
rect 65215 3531 65483 3539
rect 63340 3518 63425 3528
rect 63340 3448 63425 3458
rect 64055 3508 64117 3510
rect 64055 3500 64119 3508
rect 64117 3498 64119 3500
rect 65215 3468 65223 3531
rect 65290 3471 65483 3531
rect 65538 3471 67003 3539
rect 65290 3468 67003 3471
rect 65215 3461 67003 3468
rect 65216 3460 65305 3461
rect 65223 3458 65290 3460
rect 67003 3450 67076 3460
rect 64055 3426 64119 3436
rect 68767 3318 68873 6371
rect 71202 6331 71287 6371
rect 71319 6353 71404 6381
rect 71486 6368 71495 6441
rect 71565 6368 71572 6441
rect 71202 6205 71286 6331
rect 71200 6194 71286 6205
rect 71200 6123 71212 6194
rect 71275 6123 71286 6194
rect 71200 6112 71286 6123
rect 71202 5109 71286 6112
rect 70231 4959 70241 5059
rect 70333 4959 70343 5059
rect 71202 5039 71212 5109
rect 71274 5039 71286 5109
rect 71202 5030 71286 5039
rect 71322 4868 71401 6353
rect 71486 6335 71572 6368
rect 71487 5227 71571 6335
rect 71487 5159 71495 5227
rect 71560 5159 71571 5227
rect 71487 5148 71571 5159
rect 72475 4963 72485 5039
rect 72543 4963 72553 5039
rect 71322 4809 71332 4868
rect 71392 4809 71402 4868
rect 68767 3317 71267 3318
rect 67830 3311 68312 3312
rect 66537 3301 68312 3311
rect 66599 3300 68312 3301
rect 66599 3210 68186 3300
rect 66537 3209 68186 3210
rect 68296 3209 68312 3300
rect 66537 3200 68312 3209
rect 68767 3239 71282 3317
rect 71315 3306 71400 3317
rect 71482 3306 71567 3317
rect 71313 3249 71323 3306
rect 71391 3249 71401 3306
rect 71481 3249 71491 3306
rect 71559 3249 71569 3306
rect 68186 3199 68296 3200
rect 67592 3038 67654 3040
rect 67592 3030 67656 3038
rect 67654 3028 67656 3030
rect 67592 2956 67656 2966
rect 65937 2252 66148 2262
rect 65937 2085 66148 2095
rect 63830 1634 63890 1644
rect 63830 1562 63890 1572
rect 63170 698 63254 708
rect 63170 599 63254 608
rect 63000 562 63638 564
rect 63000 561 63663 562
rect 63000 551 63670 561
rect 63000 487 63604 551
rect 63000 477 63670 487
rect 64781 534 68317 622
rect 63000 475 63595 477
rect 58648 425 58952 431
rect 64052 438 64114 440
rect 64052 430 64116 438
rect 64114 428 64116 430
rect 58653 421 58716 425
rect 64052 356 64116 366
rect 58326 53 58336 206
rect 58465 53 58475 206
rect 59819 109 59972 119
rect 59819 -30 59972 -20
rect 61717 109 61870 119
rect 61717 -30 61870 -20
rect 44326 -48 44443 -38
rect 44326 -154 44331 -48
rect 50981 -47 51098 -37
rect 37775 -163 37891 -162
rect 44326 -164 44443 -154
rect 50142 -85 50310 -75
rect 44326 -165 44442 -164
rect 50142 -172 50169 -85
rect 50271 -172 50310 -85
rect 50981 -153 50986 -47
rect 50981 -163 51098 -153
rect 57603 -46 57720 -36
rect 57603 -152 57608 -46
rect 57603 -162 57720 -152
rect 57603 -163 57719 -162
rect 50981 -164 51097 -163
rect 50142 -420 50310 -172
rect 64781 -420 64875 534
rect 66015 234 66168 244
rect 66015 95 66168 105
rect 67370 -114 67430 -104
rect 67370 -186 67430 -176
rect 50142 -594 64875 -420
rect 50241 -595 64875 -594
rect 65223 -686 65290 -681
rect 65216 -691 66932 -686
rect 42168 -713 42232 -703
rect 42230 -777 42232 -775
rect 42168 -785 42232 -777
rect 48722 -708 48786 -698
rect 48784 -772 48786 -770
rect 48722 -780 48786 -772
rect 55371 -720 55435 -710
rect 48722 -782 48784 -780
rect 65216 -754 65223 -691
rect 65290 -696 66932 -691
rect 65290 -752 66879 -696
rect 65290 -754 66932 -752
rect 65216 -762 66932 -754
rect 65223 -764 65290 -762
rect 67968 -779 68110 -778
rect 68203 -779 68317 534
rect 68767 173 68873 3239
rect 71198 3073 71282 3239
rect 71315 3221 71400 3249
rect 71482 3221 71567 3249
rect 71196 3062 71282 3073
rect 71196 2991 71208 3062
rect 71271 2991 71282 3062
rect 71196 2980 71282 2991
rect 71198 1977 71282 2980
rect 70227 1827 70237 1927
rect 70329 1827 70339 1927
rect 71198 1907 71208 1977
rect 71270 1907 71282 1977
rect 71198 1898 71282 1907
rect 71318 1736 71397 3221
rect 71483 2095 71567 3221
rect 71483 2027 71491 2095
rect 71556 2027 71567 2095
rect 71483 2016 71567 2027
rect 72471 1831 72481 1907
rect 72539 1831 72549 1907
rect 71318 1677 71328 1736
rect 71388 1677 71398 1736
rect 68767 95 71282 173
rect 71315 162 71400 173
rect 71482 162 71567 172
rect 71313 105 71323 162
rect 71391 105 71401 162
rect 71481 105 71491 162
rect 71559 105 71569 162
rect 71198 -71 71282 95
rect 71315 77 71400 105
rect 71482 77 71567 105
rect 71196 -82 71282 -71
rect 71196 -153 71208 -82
rect 71271 -153 71282 -82
rect 71196 -164 71282 -153
rect 55433 -784 55435 -782
rect 42168 -787 42230 -785
rect 55371 -792 55435 -784
rect 67955 -788 68317 -779
rect 55371 -794 55433 -792
rect 67003 -799 67076 -789
rect 65223 -808 65290 -807
rect 65483 -808 67003 -799
rect 65215 -809 67003 -808
rect 65215 -817 65483 -809
rect 65215 -880 65223 -817
rect 65290 -877 65483 -817
rect 65538 -877 67003 -809
rect 65290 -880 67003 -877
rect 65215 -887 67003 -880
rect 65216 -888 65305 -887
rect 67955 -876 67968 -788
rect 68110 -876 68317 -788
rect 67955 -887 68317 -876
rect 65223 -890 65290 -888
rect 67003 -898 67076 -888
rect 41229 -948 41305 -946
rect 36362 -2268 36374 -2199
rect 36470 -2268 36480 -2199
rect 36362 -2274 36480 -2268
rect 41222 -956 41314 -948
rect 41222 -1042 41229 -956
rect 41305 -1042 41314 -956
rect 36374 -2278 36470 -2274
rect 41222 -2448 41314 -1042
rect 63584 -962 63668 -952
rect 68719 -1036 68845 -1035
rect 67909 -1037 68845 -1036
rect 63584 -1062 63668 -1052
rect 66537 -1047 68845 -1037
rect 41409 -1083 41589 -1073
rect 41409 -1174 41460 -1083
rect 54657 -1092 54726 -1082
rect 41409 -1184 41589 -1174
rect 54649 -1181 54657 -1092
rect 54726 -1181 54727 -1092
rect 66599 -1053 68845 -1047
rect 66599 -1126 68739 -1053
rect 68826 -1126 68845 -1053
rect 66599 -1138 68845 -1126
rect 66537 -1145 68845 -1138
rect 66537 -1148 68726 -1145
rect 41409 -2195 41518 -1184
rect 41946 -1919 42006 -1909
rect 41946 -1991 42006 -1981
rect 48500 -1914 48560 -1904
rect 48500 -1986 48560 -1976
rect 41409 -2269 41414 -2195
rect 41514 -2269 41518 -2195
rect 41409 -2275 41518 -2269
rect 41414 -2279 41514 -2275
rect 41222 -2530 41314 -2520
rect 54649 -2340 54727 -1181
rect 71198 -1167 71282 -164
rect 63837 -1211 63897 -1201
rect 63837 -1283 63897 -1273
rect 67592 -1310 67654 -1308
rect 67592 -1318 67656 -1310
rect 70227 -1317 70237 -1217
rect 70329 -1317 70339 -1217
rect 71198 -1237 71208 -1167
rect 71270 -1237 71282 -1167
rect 71198 -1246 71282 -1237
rect 67654 -1320 67656 -1318
rect 67592 -1392 67656 -1382
rect 71318 -1408 71397 77
rect 71483 -1049 71567 77
rect 71483 -1117 71491 -1049
rect 71556 -1117 71567 -1049
rect 71483 -1128 71567 -1117
rect 72471 -1313 72481 -1237
rect 72539 -1313 72549 -1237
rect 71318 -1467 71328 -1408
rect 71388 -1467 71398 -1408
rect 62999 -1705 63083 -1695
rect 62999 -1805 63083 -1795
rect 55149 -1926 55209 -1916
rect 55149 -1998 55209 -1988
rect 63168 -2021 63252 -2011
rect 63168 -2121 63252 -2111
rect 65937 -2096 66148 -2086
rect 65937 -2263 66148 -2253
rect 54649 -2455 54728 -2340
rect 63481 -2370 63542 -2360
rect 63481 -2455 63542 -2445
rect 64059 -2407 64121 -2405
rect 64059 -2415 64123 -2407
rect 64121 -2417 64123 -2415
rect 54649 -2523 54654 -2455
rect 54723 -2523 54728 -2455
rect 64059 -2489 64123 -2479
rect 54649 -2526 54728 -2523
rect 54654 -2533 54723 -2526
rect 36213 -2931 36220 -2877
rect 36315 -2883 36320 -2877
rect 36315 -2931 36319 -2883
rect 36213 -2942 36319 -2931
rect 31068 -2959 31154 -2949
rect 31068 -3054 31154 -3044
rect 1548 -3724 1624 -3714
rect 1548 -3792 1624 -3782
rect 4692 -3724 4768 -3714
rect 4692 -3792 4768 -3782
rect 7824 -3720 7900 -3710
rect 7824 -3788 7900 -3778
rect 10968 -3720 11044 -3710
rect 10968 -3788 11044 -3778
rect 14170 -3724 14246 -3714
rect 14170 -3792 14246 -3782
rect 17314 -3724 17390 -3714
rect 17314 -3792 17390 -3782
rect 20446 -3720 20522 -3710
rect 20446 -3788 20522 -3778
rect 23590 -3720 23666 -3710
rect 23590 -3788 23666 -3778
<< via2 >>
rect 4272 22240 4372 22268
rect 4272 22180 4280 22240
rect 4280 22180 4360 22240
rect 4360 22180 4372 22240
rect 4272 22176 4372 22180
rect 7416 22240 7516 22268
rect 7416 22180 7424 22240
rect 7424 22180 7504 22240
rect 7504 22180 7516 22240
rect 7416 22176 7516 22180
rect 10548 22236 10648 22264
rect 10548 22176 10556 22236
rect 10556 22176 10636 22236
rect 10636 22176 10648 22236
rect 10548 22172 10648 22176
rect 13692 22236 13792 22264
rect 13692 22176 13700 22236
rect 13700 22176 13780 22236
rect 13780 22176 13792 22236
rect 13692 22172 13792 22176
rect 16894 22240 16994 22268
rect 16894 22180 16902 22240
rect 16902 22180 16982 22240
rect 16982 22180 16994 22240
rect 16894 22176 16994 22180
rect 20038 22240 20138 22268
rect 20038 22180 20046 22240
rect 20046 22180 20126 22240
rect 20126 22180 20138 22240
rect 20038 22176 20138 22180
rect 23170 22236 23270 22264
rect 23170 22176 23178 22236
rect 23178 22176 23258 22236
rect 23258 22176 23270 22236
rect 23170 22172 23270 22176
rect 26314 22236 26414 22264
rect 26314 22176 26322 22236
rect 26322 22176 26402 22236
rect 26402 22176 26414 22236
rect 26314 22172 26414 22176
rect 27948 21443 28042 21444
rect 27948 21386 27952 21443
rect 27952 21386 28039 21443
rect 28039 21386 28042 21443
rect 27948 21381 28042 21386
rect 2735 21234 2840 21242
rect 2735 21167 2748 21234
rect 2748 21167 2827 21234
rect 2827 21167 2840 21234
rect 2735 21152 2840 21167
rect 5683 20935 5762 21024
rect 2744 20814 2837 20890
rect 27738 21113 27794 21169
rect 27948 21009 28044 21013
rect 27948 20947 27957 21009
rect 27957 20947 28037 21009
rect 28037 20947 28044 21009
rect 27948 20939 28044 20947
rect 28530 20865 28598 20867
rect 28530 20813 28535 20865
rect 28535 20813 28595 20865
rect 28595 20813 28598 20865
rect 28530 20811 28598 20813
rect 9146 20672 9210 20731
rect 27951 20663 28043 20667
rect 12290 20509 12346 20578
rect 27951 20611 27956 20663
rect 27956 20611 28038 20663
rect 28038 20611 28043 20663
rect 27951 20610 28043 20611
rect 27946 20521 28046 20522
rect 27946 20466 27949 20521
rect 27949 20466 28039 20521
rect 28039 20466 28046 20521
rect 15509 20359 15571 20427
rect 27941 20392 28050 20395
rect 27941 20339 27945 20392
rect 27945 20339 28046 20392
rect 28046 20339 28050 20392
rect 27941 20336 28050 20339
rect 18687 20222 18746 20279
rect 21813 20096 21872 20162
rect 27940 20150 28050 20154
rect 27940 20098 27945 20150
rect 27945 20098 28045 20150
rect 28045 20098 28050 20150
rect 27940 20094 28050 20098
rect 4276 20022 4352 20024
rect 4276 19970 4280 20022
rect 4280 19970 4346 20022
rect 4346 19970 4352 20022
rect 4276 19966 4352 19970
rect 7420 20022 7496 20024
rect 7420 19970 7424 20022
rect 7424 19970 7490 20022
rect 7490 19970 7496 20022
rect 7420 19966 7496 19970
rect 10552 20018 10628 20020
rect 10552 19966 10556 20018
rect 10556 19966 10622 20018
rect 10622 19966 10628 20018
rect 10552 19962 10628 19966
rect 13696 20018 13772 20020
rect 13696 19966 13700 20018
rect 13700 19966 13766 20018
rect 13766 19966 13772 20018
rect 13696 19962 13772 19966
rect 16898 20022 16974 20024
rect 16898 19970 16902 20022
rect 16902 19970 16968 20022
rect 16968 19970 16974 20022
rect 16898 19966 16974 19970
rect 20042 20022 20118 20024
rect 20042 19970 20046 20022
rect 20046 19970 20112 20022
rect 20112 19970 20118 20022
rect 20042 19966 20118 19970
rect 23174 20018 23250 20020
rect 23174 19966 23178 20018
rect 23178 19966 23244 20018
rect 23244 19966 23250 20018
rect 23174 19962 23250 19966
rect 26318 20018 26394 20020
rect 26318 19966 26322 20018
rect 26322 19966 26388 20018
rect 26388 19966 26394 20018
rect 26318 19962 26394 19966
rect 24932 19801 25005 19882
rect 27943 19929 28047 19933
rect 27943 19875 27945 19929
rect 27945 19875 28043 19929
rect 28043 19875 28047 19929
rect 27943 19872 28047 19875
rect 4622 17027 4712 17048
rect 4622 16975 4638 17027
rect 4638 16975 4690 17027
rect 4690 16975 4712 17027
rect 4622 16957 4712 16975
rect 5790 17027 5880 17048
rect 5790 16975 5806 17027
rect 5806 16975 5858 17027
rect 5858 16975 5880 17027
rect 5790 16957 5880 16975
rect 6958 17027 7048 17048
rect 6958 16975 6974 17027
rect 6974 16975 7026 17027
rect 7026 16975 7048 17027
rect 6958 16957 7048 16975
rect 8126 17027 8216 17048
rect 8126 16975 8142 17027
rect 8142 16975 8194 17027
rect 8194 16975 8216 17027
rect 8126 16957 8216 16975
rect 9300 17025 9390 17046
rect 9300 16973 9316 17025
rect 9316 16973 9368 17025
rect 9368 16973 9390 17025
rect 9300 16955 9390 16973
rect 10468 17025 10558 17046
rect 10468 16973 10484 17025
rect 10484 16973 10536 17025
rect 10536 16973 10558 17025
rect 10468 16955 10558 16973
rect 11636 17025 11726 17046
rect 11636 16973 11652 17025
rect 11652 16973 11704 17025
rect 11704 16973 11726 17025
rect 11636 16955 11726 16973
rect 12804 17025 12894 17046
rect 12804 16973 12820 17025
rect 12820 16973 12872 17025
rect 12872 16973 12894 17025
rect 12804 16955 12894 16973
rect 14498 16777 14558 16839
rect 14830 15901 14915 15902
rect 15946 16777 16006 16839
rect 14830 15813 14915 15901
rect 16288 15884 16349 15897
rect 17444 16775 17504 16837
rect 16288 15830 16292 15884
rect 16292 15830 16346 15884
rect 16346 15830 16349 15884
rect 17788 15878 17848 15888
rect 18892 16775 18952 16837
rect 16288 15818 16349 15830
rect 14830 15812 14915 15813
rect 17788 15824 17789 15878
rect 17789 15824 17843 15878
rect 17843 15824 17848 15878
rect 19238 15884 19298 15895
rect 20412 16777 20472 16839
rect 19238 15830 19241 15884
rect 19241 15830 19295 15884
rect 19295 15830 19298 15884
rect 20750 15884 20817 15897
rect 21860 16777 21920 16839
rect 20750 15830 20757 15884
rect 20757 15830 20811 15884
rect 20811 15830 20817 15884
rect 22202 15879 22266 15891
rect 23358 16775 23418 16837
rect 17788 15820 17848 15824
rect 19238 15820 19298 15830
rect 20750 15819 20817 15830
rect 22202 15825 22205 15879
rect 22205 15825 22259 15879
rect 22259 15825 22266 15879
rect 23692 15881 23768 15899
rect 24806 16775 24866 16837
rect 25630 16122 25701 16181
rect 25346 16021 25415 16085
rect 27800 16801 27858 16802
rect 27800 16747 27801 16801
rect 27801 16747 27857 16801
rect 27857 16747 27858 16801
rect 27800 16746 27858 16747
rect 23692 15826 23703 15881
rect 23703 15826 23757 15881
rect 23757 15826 23768 15881
rect 22202 15817 22266 15825
rect 23692 15812 23768 15826
rect 5087 15703 5177 15721
rect 5087 15651 5109 15703
rect 5109 15651 5161 15703
rect 5161 15651 5177 15703
rect 5087 15630 5177 15651
rect 6255 15703 6345 15721
rect 6255 15651 6277 15703
rect 6277 15651 6329 15703
rect 6329 15651 6345 15703
rect 6255 15630 6345 15651
rect 7423 15703 7513 15721
rect 7423 15651 7445 15703
rect 7445 15651 7497 15703
rect 7497 15651 7513 15703
rect 7423 15630 7513 15651
rect 8591 15703 8681 15721
rect 8591 15651 8613 15703
rect 8613 15651 8665 15703
rect 8665 15651 8681 15703
rect 8591 15630 8681 15651
rect 9765 15701 9855 15719
rect 9765 15649 9787 15701
rect 9787 15649 9839 15701
rect 9839 15649 9855 15701
rect 9765 15628 9855 15649
rect 10933 15701 11023 15719
rect 10933 15649 10955 15701
rect 10955 15649 11007 15701
rect 11007 15649 11023 15701
rect 10933 15628 11023 15649
rect 12101 15701 12191 15719
rect 12101 15649 12123 15701
rect 12123 15649 12175 15701
rect 12175 15649 12191 15701
rect 12101 15628 12191 15649
rect 13269 15701 13359 15719
rect 13269 15649 13291 15701
rect 13291 15649 13343 15701
rect 13343 15649 13359 15701
rect 13269 15628 13359 15649
rect 14272 15575 14274 15633
rect 14274 15575 14336 15633
rect 14272 15571 14336 15575
rect 15720 15575 15722 15633
rect 15722 15575 15784 15633
rect 15720 15571 15784 15575
rect 17218 15573 17220 15631
rect 17220 15573 17282 15631
rect 17218 15569 17282 15573
rect 18666 15573 18668 15631
rect 18668 15573 18730 15631
rect 18666 15569 18730 15573
rect 20186 15575 20188 15633
rect 20188 15575 20250 15633
rect 20186 15571 20250 15575
rect 21634 15575 21636 15633
rect 21636 15575 21698 15633
rect 21634 15571 21698 15575
rect 23132 15573 23134 15631
rect 23134 15573 23196 15631
rect 23132 15569 23196 15573
rect 24580 15573 24582 15631
rect 24582 15573 24644 15631
rect 24580 15569 24644 15573
rect 1770 15102 1870 15130
rect 1770 15042 1778 15102
rect 1778 15042 1858 15102
rect 1858 15042 1870 15102
rect 1770 15038 1870 15042
rect 4914 15102 5014 15130
rect 4914 15042 4922 15102
rect 4922 15042 5002 15102
rect 5002 15042 5014 15102
rect 4914 15038 5014 15042
rect 8046 15098 8146 15126
rect 8046 15038 8054 15098
rect 8054 15038 8134 15098
rect 8134 15038 8146 15098
rect 8046 15034 8146 15038
rect 11190 15098 11290 15126
rect 11190 15038 11198 15098
rect 11198 15038 11278 15098
rect 11278 15038 11290 15098
rect 11190 15034 11290 15038
rect 14392 15102 14492 15130
rect 14392 15042 14400 15102
rect 14400 15042 14480 15102
rect 14480 15042 14492 15102
rect 14392 15038 14492 15042
rect 17536 15102 17636 15130
rect 17536 15042 17544 15102
rect 17544 15042 17624 15102
rect 17624 15042 17636 15102
rect 17536 15038 17636 15042
rect 20668 15098 20768 15126
rect 20668 15038 20676 15098
rect 20676 15038 20756 15098
rect 20756 15038 20768 15098
rect 20668 15034 20768 15038
rect 23812 15098 23912 15126
rect 23812 15038 23820 15098
rect 23820 15038 23900 15098
rect 23900 15038 23912 15098
rect 23812 15034 23912 15038
rect 1774 12884 1850 12886
rect 1774 12832 1778 12884
rect 1778 12832 1844 12884
rect 1844 12832 1850 12884
rect 1774 12828 1850 12832
rect 4918 12884 4994 12886
rect 4918 12832 4922 12884
rect 4922 12832 4988 12884
rect 4988 12832 4994 12884
rect 4918 12828 4994 12832
rect 8050 12880 8126 12882
rect 8050 12828 8054 12880
rect 8054 12828 8120 12880
rect 8120 12828 8126 12880
rect 8050 12824 8126 12828
rect 11194 12880 11270 12882
rect 11194 12828 11198 12880
rect 11198 12828 11264 12880
rect 11264 12828 11270 12880
rect 11194 12824 11270 12828
rect 14396 12884 14472 12886
rect 14396 12832 14400 12884
rect 14400 12832 14466 12884
rect 14466 12832 14472 12884
rect 14396 12828 14472 12832
rect 17540 12884 17616 12886
rect 17540 12832 17544 12884
rect 17544 12832 17610 12884
rect 17610 12832 17616 12884
rect 17540 12828 17616 12832
rect 20672 12880 20748 12882
rect 20672 12828 20676 12880
rect 20676 12828 20742 12880
rect 20742 12828 20748 12880
rect 20672 12824 20748 12828
rect 23816 12880 23892 12882
rect 23816 12828 23820 12880
rect 23820 12828 23886 12880
rect 23886 12828 23892 12880
rect 23816 12824 23892 12828
rect 1770 12368 1870 12396
rect 1770 12308 1778 12368
rect 1778 12308 1858 12368
rect 1858 12308 1870 12368
rect 1770 12304 1870 12308
rect 4914 12368 5014 12396
rect 4914 12308 4922 12368
rect 4922 12308 5002 12368
rect 5002 12308 5014 12368
rect 4914 12304 5014 12308
rect 8046 12364 8146 12392
rect 8046 12304 8054 12364
rect 8054 12304 8134 12364
rect 8134 12304 8146 12364
rect 8046 12300 8146 12304
rect 11190 12364 11290 12392
rect 11190 12304 11198 12364
rect 11198 12304 11278 12364
rect 11278 12304 11290 12364
rect 11190 12300 11290 12304
rect 14392 12368 14492 12396
rect 14392 12308 14400 12368
rect 14400 12308 14480 12368
rect 14480 12308 14492 12368
rect 14392 12304 14492 12308
rect 17536 12368 17636 12396
rect 17536 12308 17544 12368
rect 17544 12308 17624 12368
rect 17624 12308 17636 12368
rect 17536 12304 17636 12308
rect 20668 12364 20768 12392
rect 20668 12304 20676 12364
rect 20676 12304 20756 12364
rect 20756 12304 20768 12364
rect 20668 12300 20768 12304
rect 23812 12364 23912 12392
rect 23812 12304 23820 12364
rect 23820 12304 23900 12364
rect 23900 12304 23912 12364
rect 23812 12300 23912 12304
rect 32913 20306 33097 20318
rect -1727 3217 -1616 3282
rect -791 2757 -659 2840
rect -545 2637 -428 2722
rect 32913 20169 32926 20306
rect 32926 20169 33084 20306
rect 33084 20169 33097 20306
rect 32913 20157 33097 20169
rect 42512 24873 42665 24884
rect 40030 24819 40183 24830
rect 40030 24711 40041 24819
rect 40041 24711 40173 24819
rect 40173 24711 40183 24819
rect 42512 24765 42523 24873
rect 42523 24765 42655 24873
rect 42655 24765 42665 24873
rect 43659 24873 43812 24884
rect 42512 24755 42665 24765
rect 40030 24701 40183 24711
rect 43659 24765 43670 24873
rect 43670 24765 43802 24873
rect 43802 24765 43812 24873
rect 49025 24870 49178 24881
rect 43659 24755 43812 24765
rect 46543 24816 46696 24827
rect 40311 23780 40440 23791
rect 40311 23648 40321 23780
rect 40321 23648 40429 23780
rect 40429 23648 40440 23780
rect 40311 23638 40440 23648
rect 38849 23078 38991 23181
rect 40044 23169 40197 23180
rect 40044 23061 40055 23169
rect 40055 23061 40187 23169
rect 40187 23061 40197 23169
rect 40044 23051 40197 23061
rect 38809 21950 38947 22076
rect 40325 22130 40454 22141
rect 40325 21998 40335 22130
rect 40335 21998 40443 22130
rect 40443 21998 40454 22130
rect 40325 21988 40454 21998
rect 39077 21693 39192 21702
rect 39077 21614 39087 21693
rect 39087 21614 39180 21693
rect 39180 21614 39192 21693
rect 39077 21605 39192 21614
rect 40039 21565 40192 21576
rect 40039 21457 40050 21565
rect 40050 21457 40182 21565
rect 40182 21457 40192 21565
rect 40039 21447 40192 21457
rect 46543 24708 46554 24816
rect 46554 24708 46686 24816
rect 46686 24708 46696 24816
rect 49025 24762 49036 24870
rect 49036 24762 49168 24870
rect 49168 24762 49178 24870
rect 50172 24870 50325 24881
rect 49025 24752 49178 24762
rect 46543 24698 46696 24708
rect 50172 24762 50183 24870
rect 50183 24762 50315 24870
rect 50315 24762 50325 24870
rect 55559 24865 55712 24876
rect 50172 24752 50325 24762
rect 53077 24811 53230 24822
rect 46824 23777 46953 23788
rect 46824 23645 46834 23777
rect 46834 23645 46942 23777
rect 46942 23645 46953 23777
rect 46824 23635 46953 23645
rect 41859 23473 42012 23483
rect 41859 23365 41869 23473
rect 41869 23365 42001 23473
rect 42001 23365 42012 23473
rect 41859 23354 42012 23365
rect 43001 23471 43154 23481
rect 43001 23363 43011 23471
rect 43011 23363 43143 23471
rect 43143 23363 43154 23471
rect 43001 23352 43154 23363
rect 41857 22826 42010 22837
rect 41857 22718 41868 22826
rect 41868 22718 42000 22826
rect 42000 22718 42010 22826
rect 41857 22708 42010 22718
rect 43755 22826 43908 22837
rect 43755 22718 43766 22826
rect 43766 22718 43898 22826
rect 43898 22718 43908 22826
rect 43755 22708 43908 22718
rect 42498 21856 42576 21866
rect 42498 21790 42513 21856
rect 42513 21790 42576 21856
rect 42498 21780 42576 21790
rect 40320 20526 40449 20537
rect 40320 20394 40330 20526
rect 40330 20394 40438 20526
rect 40438 20394 40449 20526
rect 40320 20384 40449 20394
rect 41803 20430 41956 20440
rect 41803 20322 41813 20430
rect 41813 20322 41945 20430
rect 41945 20322 41956 20430
rect 41803 20311 41956 20322
rect 43701 20430 43854 20440
rect 43701 20322 43711 20430
rect 43711 20322 43843 20430
rect 43843 20322 43854 20430
rect 43701 20311 43854 20322
rect 45281 23083 45510 23207
rect 46557 23166 46710 23177
rect 46557 23058 46568 23166
rect 46568 23058 46700 23166
rect 46700 23058 46710 23166
rect 46557 23048 46710 23058
rect 46838 22127 46967 22138
rect 46838 21995 46848 22127
rect 46848 21995 46956 22127
rect 46956 21995 46967 22127
rect 46838 21985 46967 21995
rect 45590 21690 45705 21699
rect 45590 21611 45600 21690
rect 45600 21611 45693 21690
rect 45693 21611 45705 21690
rect 45590 21602 45705 21611
rect 46552 21562 46705 21573
rect 46552 21454 46563 21562
rect 46563 21454 46695 21562
rect 46695 21454 46705 21562
rect 46552 21444 46705 21454
rect 53077 24703 53088 24811
rect 53088 24703 53220 24811
rect 53220 24703 53230 24811
rect 55559 24757 55570 24865
rect 55570 24757 55702 24865
rect 55702 24757 55712 24865
rect 56706 24865 56859 24876
rect 55559 24747 55712 24757
rect 53077 24693 53230 24703
rect 56706 24757 56717 24865
rect 56717 24757 56849 24865
rect 56849 24757 56859 24865
rect 62117 24869 62270 24880
rect 56706 24747 56859 24757
rect 59635 24815 59788 24826
rect 53358 23772 53487 23783
rect 53358 23640 53368 23772
rect 53368 23640 53476 23772
rect 53476 23640 53487 23772
rect 53358 23630 53487 23640
rect 48372 23470 48525 23480
rect 48372 23362 48382 23470
rect 48382 23362 48514 23470
rect 48514 23362 48525 23470
rect 48372 23351 48525 23362
rect 49514 23468 49667 23478
rect 49514 23360 49524 23468
rect 49524 23360 49656 23468
rect 49656 23360 49667 23468
rect 49514 23349 49667 23360
rect 48370 22823 48523 22834
rect 48370 22715 48381 22823
rect 48381 22715 48513 22823
rect 48513 22715 48523 22823
rect 48370 22705 48523 22715
rect 50268 22823 50421 22834
rect 50268 22715 50279 22823
rect 50279 22715 50411 22823
rect 50411 22715 50421 22823
rect 50268 22705 50421 22715
rect 49011 21853 49089 21863
rect 49011 21787 49026 21853
rect 49026 21787 49089 21853
rect 49011 21777 49089 21787
rect 46833 20523 46962 20534
rect 46833 20391 46843 20523
rect 46843 20391 46951 20523
rect 46951 20391 46962 20523
rect 46833 20381 46962 20391
rect 48316 20427 48469 20437
rect 48316 20319 48326 20427
rect 48326 20319 48458 20427
rect 48458 20319 48469 20427
rect 48316 20308 48469 20319
rect 50214 20427 50367 20437
rect 50214 20319 50224 20427
rect 50224 20319 50356 20427
rect 50356 20319 50367 20427
rect 50214 20308 50367 20319
rect 51840 23073 52058 23213
rect 53091 23161 53244 23172
rect 53091 23053 53102 23161
rect 53102 23053 53234 23161
rect 53234 23053 53244 23161
rect 53091 23043 53244 23053
rect 53372 22122 53501 22133
rect 53372 21990 53382 22122
rect 53382 21990 53490 22122
rect 53490 21990 53501 22122
rect 53372 21980 53501 21990
rect 52124 21685 52239 21694
rect 52124 21606 52134 21685
rect 52134 21606 52227 21685
rect 52227 21606 52239 21685
rect 52124 21597 52239 21606
rect 53086 21557 53239 21568
rect 53086 21449 53097 21557
rect 53097 21449 53229 21557
rect 53229 21449 53239 21557
rect 53086 21439 53239 21449
rect 59635 24707 59646 24815
rect 59646 24707 59778 24815
rect 59778 24707 59788 24815
rect 62117 24761 62128 24869
rect 62128 24761 62260 24869
rect 62260 24761 62270 24869
rect 63264 24869 63417 24880
rect 62117 24751 62270 24761
rect 59635 24697 59788 24707
rect 63264 24761 63275 24869
rect 63275 24761 63407 24869
rect 63407 24761 63417 24869
rect 63264 24751 63417 24761
rect 59916 23776 60045 23787
rect 59916 23644 59926 23776
rect 59926 23644 60034 23776
rect 60034 23644 60045 23776
rect 59916 23634 60045 23644
rect 54906 23465 55059 23475
rect 54906 23357 54916 23465
rect 54916 23357 55048 23465
rect 55048 23357 55059 23465
rect 54906 23346 55059 23357
rect 56048 23463 56201 23473
rect 56048 23355 56058 23463
rect 56058 23355 56190 23463
rect 56190 23355 56201 23463
rect 56048 23344 56201 23355
rect 54904 22818 55057 22829
rect 54904 22710 54915 22818
rect 54915 22710 55047 22818
rect 55047 22710 55057 22818
rect 54904 22700 55057 22710
rect 56802 22818 56955 22829
rect 56802 22710 56813 22818
rect 56813 22710 56945 22818
rect 56945 22710 56955 22818
rect 56802 22700 56955 22710
rect 55545 21848 55623 21858
rect 55545 21782 55560 21848
rect 55560 21782 55623 21848
rect 55545 21772 55623 21782
rect 53367 20518 53496 20529
rect 53367 20386 53377 20518
rect 53377 20386 53485 20518
rect 53485 20386 53496 20518
rect 53367 20376 53496 20386
rect 54850 20422 55003 20432
rect 54850 20314 54860 20422
rect 54860 20314 54992 20422
rect 54992 20314 55003 20422
rect 54850 20303 55003 20314
rect 56748 20422 56901 20432
rect 56748 20314 56758 20422
rect 56758 20314 56890 20422
rect 56890 20314 56901 20422
rect 56748 20303 56901 20314
rect 58364 23070 58616 23215
rect 59649 23165 59802 23176
rect 59649 23057 59660 23165
rect 59660 23057 59792 23165
rect 59792 23057 59802 23165
rect 59649 23047 59802 23057
rect 59930 22126 60059 22137
rect 59930 21994 59940 22126
rect 59940 21994 60048 22126
rect 60048 21994 60059 22126
rect 59930 21984 60059 21994
rect 58682 21689 58797 21698
rect 58682 21610 58692 21689
rect 58692 21610 58785 21689
rect 58785 21610 58797 21689
rect 58682 21601 58797 21610
rect 59644 21561 59797 21572
rect 59644 21453 59655 21561
rect 59655 21453 59787 21561
rect 59787 21453 59797 21561
rect 59644 21443 59797 21453
rect 61464 23469 61617 23479
rect 61464 23361 61474 23469
rect 61474 23361 61606 23469
rect 61606 23361 61617 23469
rect 61464 23350 61617 23361
rect 62606 23467 62759 23477
rect 62606 23359 62616 23467
rect 62616 23359 62748 23467
rect 62748 23359 62759 23467
rect 62606 23348 62759 23359
rect 61462 22822 61615 22833
rect 61462 22714 61473 22822
rect 61473 22714 61605 22822
rect 61605 22714 61615 22822
rect 61462 22704 61615 22714
rect 63360 22822 63513 22833
rect 63360 22714 63371 22822
rect 63371 22714 63503 22822
rect 63503 22714 63513 22822
rect 63360 22704 63513 22714
rect 62103 21852 62181 21862
rect 62103 21786 62118 21852
rect 62118 21786 62181 21852
rect 62103 21776 62181 21786
rect 59925 20522 60054 20533
rect 59925 20390 59935 20522
rect 59935 20390 60043 20522
rect 60043 20390 60054 20522
rect 59925 20380 60054 20390
rect 61408 20426 61561 20436
rect 61408 20318 61418 20426
rect 61418 20318 61550 20426
rect 61550 20318 61561 20426
rect 61408 20307 61561 20318
rect 63306 20426 63459 20436
rect 63306 20318 63316 20426
rect 63316 20318 63448 20426
rect 63448 20318 63459 20426
rect 63306 20307 63459 20318
rect 39608 19265 39761 19276
rect 39608 19157 39618 19265
rect 39618 19157 39750 19265
rect 39750 19157 39761 19265
rect 40755 19265 40908 19276
rect 39608 19147 39761 19157
rect 40755 19157 40765 19265
rect 40765 19157 40897 19265
rect 40897 19157 40908 19265
rect 46166 19261 46319 19272
rect 40755 19147 40908 19157
rect 43237 19211 43390 19222
rect 43237 19103 43247 19211
rect 43247 19103 43379 19211
rect 43379 19103 43390 19211
rect 46166 19153 46176 19261
rect 46176 19153 46308 19261
rect 46308 19153 46319 19261
rect 47313 19261 47466 19272
rect 46166 19143 46319 19153
rect 47313 19153 47323 19261
rect 47323 19153 47455 19261
rect 47455 19153 47466 19261
rect 52700 19266 52853 19277
rect 47313 19143 47466 19153
rect 49795 19207 49948 19218
rect 43237 19093 43390 19103
rect 40266 17863 40419 17873
rect 40266 17755 40277 17863
rect 40277 17755 40409 17863
rect 40409 17755 40419 17863
rect 40266 17744 40419 17755
rect 41408 17865 41561 17875
rect 41408 17757 41419 17865
rect 41419 17757 41551 17865
rect 41551 17757 41561 17865
rect 41408 17746 41561 17757
rect 39512 17218 39665 17229
rect 39512 17110 39522 17218
rect 39522 17110 39654 17218
rect 39654 17110 39665 17218
rect 39512 17100 39665 17110
rect 41410 17218 41563 17229
rect 41410 17110 41420 17218
rect 41420 17110 41552 17218
rect 41552 17110 41563 17218
rect 41410 17100 41563 17110
rect 40844 16248 40922 16258
rect 40844 16182 40907 16248
rect 40907 16182 40922 16248
rect 40844 16172 40922 16182
rect 49795 19099 49805 19207
rect 49805 19099 49937 19207
rect 49937 19099 49948 19207
rect 52700 19158 52710 19266
rect 52710 19158 52842 19266
rect 52842 19158 52853 19266
rect 53847 19266 54000 19277
rect 52700 19148 52853 19158
rect 53847 19158 53857 19266
rect 53857 19158 53989 19266
rect 53989 19158 54000 19266
rect 59213 19269 59366 19280
rect 53847 19148 54000 19158
rect 56329 19212 56482 19223
rect 49795 19089 49948 19099
rect 42980 18172 43109 18183
rect 42980 18040 42991 18172
rect 42991 18040 43099 18172
rect 43099 18040 43109 18172
rect 42980 18030 43109 18040
rect 43223 17561 43376 17572
rect 43223 17453 43233 17561
rect 43233 17453 43365 17561
rect 43365 17453 43376 17561
rect 43223 17443 43376 17453
rect 42966 16522 43095 16533
rect 42966 16390 42977 16522
rect 42977 16390 43085 16522
rect 43085 16390 43095 16522
rect 42966 16380 43095 16390
rect 43228 15957 43381 15968
rect 43228 15849 43238 15957
rect 43238 15849 43370 15957
rect 43370 15849 43381 15957
rect 43228 15839 43381 15849
rect 39566 14822 39719 14832
rect 39566 14714 39577 14822
rect 39577 14714 39709 14822
rect 39709 14714 39719 14822
rect 39566 14703 39719 14714
rect 41464 14822 41617 14832
rect 41464 14714 41475 14822
rect 41475 14714 41607 14822
rect 41607 14714 41617 14822
rect 42971 14918 43100 14929
rect 42971 14786 42982 14918
rect 42982 14786 43090 14918
rect 43090 14786 43100 14918
rect 42971 14776 43100 14786
rect 41464 14703 41617 14714
rect 44228 16085 44343 16094
rect 44228 16006 44240 16085
rect 44240 16006 44333 16085
rect 44333 16006 44343 16085
rect 44228 15997 44343 16006
rect 46824 17859 46977 17869
rect 46824 17751 46835 17859
rect 46835 17751 46967 17859
rect 46967 17751 46977 17859
rect 46824 17740 46977 17751
rect 47966 17861 48119 17871
rect 47966 17753 47977 17861
rect 47977 17753 48109 17861
rect 48109 17753 48119 17861
rect 47966 17742 48119 17753
rect 46070 17214 46223 17225
rect 46070 17106 46080 17214
rect 46080 17106 46212 17214
rect 46212 17106 46223 17214
rect 46070 17096 46223 17106
rect 47968 17214 48121 17225
rect 47968 17106 47978 17214
rect 47978 17106 48110 17214
rect 48110 17106 48121 17214
rect 47968 17096 48121 17106
rect 47402 16244 47480 16254
rect 47402 16178 47465 16244
rect 47465 16178 47480 16244
rect 47402 16168 47480 16178
rect 56329 19104 56339 19212
rect 56339 19104 56471 19212
rect 56471 19104 56482 19212
rect 59213 19161 59223 19269
rect 59223 19161 59355 19269
rect 59355 19161 59366 19269
rect 60360 19269 60513 19280
rect 59213 19151 59366 19161
rect 60360 19161 60370 19269
rect 60370 19161 60502 19269
rect 60502 19161 60513 19269
rect 60360 19151 60513 19161
rect 62842 19215 62995 19226
rect 56329 19094 56482 19104
rect 49538 18168 49667 18179
rect 49538 18036 49549 18168
rect 49549 18036 49657 18168
rect 49657 18036 49667 18168
rect 49538 18026 49667 18036
rect 53358 17864 53511 17874
rect 53358 17756 53369 17864
rect 53369 17756 53501 17864
rect 53501 17756 53511 17864
rect 53358 17745 53511 17756
rect 54500 17866 54653 17876
rect 54500 17758 54511 17866
rect 54511 17758 54643 17866
rect 54643 17758 54653 17866
rect 54500 17747 54653 17758
rect 49781 17557 49934 17568
rect 49781 17449 49791 17557
rect 49791 17449 49923 17557
rect 49923 17449 49934 17557
rect 49781 17439 49934 17449
rect 49524 16518 49653 16529
rect 49524 16386 49535 16518
rect 49535 16386 49643 16518
rect 49643 16386 49653 16518
rect 49524 16376 49653 16386
rect 49786 15953 49939 15964
rect 49786 15845 49796 15953
rect 49796 15845 49928 15953
rect 49928 15845 49939 15953
rect 49786 15835 49939 15845
rect 46124 14818 46277 14828
rect 46124 14710 46135 14818
rect 46135 14710 46267 14818
rect 46267 14710 46277 14818
rect 46124 14699 46277 14710
rect 48022 14818 48175 14828
rect 48022 14710 48033 14818
rect 48033 14710 48165 14818
rect 48165 14710 48175 14818
rect 49529 14914 49658 14925
rect 49529 14782 49540 14914
rect 49540 14782 49648 14914
rect 49648 14782 49658 14914
rect 49529 14772 49658 14782
rect 48022 14699 48175 14710
rect 50786 16081 50901 16090
rect 50786 16002 50798 16081
rect 50798 16002 50891 16081
rect 50891 16002 50901 16081
rect 50786 15993 50901 16002
rect 52604 17219 52757 17230
rect 52604 17111 52614 17219
rect 52614 17111 52746 17219
rect 52746 17111 52757 17219
rect 52604 17101 52757 17111
rect 54502 17219 54655 17230
rect 54502 17111 54512 17219
rect 54512 17111 54644 17219
rect 54644 17111 54655 17219
rect 54502 17101 54655 17111
rect 53936 16249 54014 16259
rect 53936 16183 53999 16249
rect 53999 16183 54014 16249
rect 53936 16173 54014 16183
rect 62842 19107 62852 19215
rect 62852 19107 62984 19215
rect 62984 19107 62995 19215
rect 62842 19097 62995 19107
rect 56072 18173 56201 18184
rect 56072 18041 56083 18173
rect 56083 18041 56191 18173
rect 56191 18041 56201 18173
rect 56072 18031 56201 18041
rect 56315 17562 56468 17573
rect 56315 17454 56325 17562
rect 56325 17454 56457 17562
rect 56457 17454 56468 17562
rect 56315 17444 56468 17454
rect 56058 16523 56187 16534
rect 56058 16391 56069 16523
rect 56069 16391 56177 16523
rect 56177 16391 56187 16523
rect 56058 16381 56187 16391
rect 56320 15958 56473 15969
rect 56320 15850 56330 15958
rect 56330 15850 56462 15958
rect 56462 15850 56473 15958
rect 56320 15840 56473 15850
rect 52658 14823 52811 14833
rect 52658 14715 52669 14823
rect 52669 14715 52801 14823
rect 52801 14715 52811 14823
rect 52658 14704 52811 14715
rect 54556 14823 54709 14833
rect 54556 14715 54567 14823
rect 54567 14715 54699 14823
rect 54699 14715 54709 14823
rect 56063 14919 56192 14930
rect 56063 14787 56074 14919
rect 56074 14787 56182 14919
rect 56182 14787 56192 14919
rect 56063 14777 56192 14787
rect 54556 14704 54709 14715
rect 57320 16086 57435 16095
rect 57320 16007 57332 16086
rect 57332 16007 57425 16086
rect 57425 16007 57435 16086
rect 57320 15998 57435 16007
rect 59871 17867 60024 17877
rect 59871 17759 59882 17867
rect 59882 17759 60014 17867
rect 60014 17759 60024 17867
rect 59871 17748 60024 17759
rect 61013 17869 61166 17879
rect 61013 17761 61024 17869
rect 61024 17761 61156 17869
rect 61156 17761 61166 17869
rect 61013 17750 61166 17761
rect 59117 17222 59270 17233
rect 59117 17114 59127 17222
rect 59127 17114 59259 17222
rect 59259 17114 59270 17222
rect 59117 17104 59270 17114
rect 61015 17222 61168 17233
rect 61015 17114 61025 17222
rect 61025 17114 61157 17222
rect 61157 17114 61168 17222
rect 61015 17104 61168 17114
rect 60449 16252 60527 16262
rect 60449 16186 60512 16252
rect 60512 16186 60527 16252
rect 60449 16176 60527 16186
rect 62585 18176 62714 18187
rect 62585 18044 62596 18176
rect 62596 18044 62704 18176
rect 62704 18044 62714 18176
rect 62585 18034 62714 18044
rect 62828 17565 62981 17576
rect 62828 17457 62838 17565
rect 62838 17457 62970 17565
rect 62970 17457 62981 17565
rect 64020 17481 64238 17637
rect 62828 17447 62981 17457
rect 62571 16526 62700 16537
rect 62571 16394 62582 16526
rect 62582 16394 62690 16526
rect 62690 16394 62700 16526
rect 62571 16384 62700 16394
rect 62833 15961 62986 15972
rect 62833 15853 62843 15961
rect 62843 15853 62975 15961
rect 62975 15853 62986 15961
rect 62833 15843 62986 15853
rect 59171 14826 59324 14836
rect 59171 14718 59182 14826
rect 59182 14718 59314 14826
rect 59314 14718 59324 14826
rect 59171 14707 59324 14718
rect 61069 14826 61222 14836
rect 61069 14718 61080 14826
rect 61080 14718 61212 14826
rect 61212 14718 61222 14826
rect 62576 14922 62705 14933
rect 62576 14790 62587 14922
rect 62587 14790 62695 14922
rect 62695 14790 62705 14922
rect 62576 14780 62705 14790
rect 61069 14707 61222 14718
rect 63833 16089 63948 16098
rect 63833 16010 63845 16089
rect 63845 16010 63938 16089
rect 63938 16010 63948 16089
rect 63833 16001 63948 16010
rect 29695 12341 29765 12353
rect 29695 12287 29703 12341
rect 29703 12287 29757 12341
rect 29757 12287 29765 12341
rect 29695 12275 29765 12287
rect 57724 13164 57823 13180
rect 57724 13089 57731 13164
rect 57731 13089 57817 13164
rect 57817 13089 57823 13164
rect 57724 13078 57823 13089
rect 51199 13043 51299 13050
rect 51199 12973 51208 13043
rect 51208 12973 51295 13043
rect 51295 12973 51299 13043
rect 51199 12965 51299 12973
rect 44619 12710 44737 12714
rect 44619 12649 44633 12710
rect 44633 12649 44726 12710
rect 44726 12649 44737 12710
rect 44619 12646 44737 12649
rect 31925 12399 31995 12405
rect 31925 12337 31927 12399
rect 31927 12337 31985 12399
rect 31985 12337 31995 12399
rect 31925 12333 31995 12337
rect 41911 12313 41971 12375
rect 48460 12312 48520 12374
rect 55114 12333 55174 12395
rect 63767 12166 63827 12228
rect 66013 12157 66166 12168
rect 66013 12049 66024 12157
rect 66024 12049 66156 12157
rect 66156 12049 66166 12157
rect 66013 12039 66166 12049
rect 67368 11758 67428 11820
rect 31064 11518 31160 11526
rect 31064 11441 31074 11518
rect 31074 11441 31153 11518
rect 31153 11441 31160 11518
rect 31064 11429 31160 11441
rect 42133 11111 42195 11169
rect 42195 11111 42197 11169
rect 42133 11107 42197 11111
rect 48682 11110 48744 11168
rect 48744 11110 48746 11168
rect 55336 11131 55398 11189
rect 55398 11131 55400 11189
rect 55336 11127 55400 11131
rect 48682 11106 48746 11110
rect 29693 10273 29763 10285
rect 29693 10219 29701 10273
rect 29701 10219 29755 10273
rect 29755 10219 29763 10273
rect 29693 10207 29763 10219
rect 1774 10150 1850 10152
rect 1774 10098 1778 10150
rect 1778 10098 1844 10150
rect 1844 10098 1850 10150
rect 1774 10094 1850 10098
rect 4918 10150 4994 10152
rect 4918 10098 4922 10150
rect 4922 10098 4988 10150
rect 4988 10098 4994 10150
rect 4918 10094 4994 10098
rect 8050 10146 8126 10148
rect 8050 10094 8054 10146
rect 8054 10094 8120 10146
rect 8120 10094 8126 10146
rect 8050 10090 8126 10094
rect 11194 10146 11270 10148
rect 11194 10094 11198 10146
rect 11198 10094 11264 10146
rect 11264 10094 11270 10146
rect 11194 10090 11270 10094
rect 14396 10150 14472 10152
rect 14396 10098 14400 10150
rect 14400 10098 14466 10150
rect 14466 10098 14472 10150
rect 14396 10094 14472 10098
rect 17540 10150 17616 10152
rect 17540 10098 17544 10150
rect 17544 10098 17610 10150
rect 17610 10098 17616 10150
rect 20672 10146 20748 10148
rect 17540 10094 17616 10098
rect 20672 10094 20676 10146
rect 20676 10094 20742 10146
rect 20742 10094 20748 10146
rect 20672 10090 20748 10094
rect 1780 9636 1880 9664
rect 1780 9576 1788 9636
rect 1788 9576 1868 9636
rect 1868 9576 1880 9636
rect 1780 9572 1880 9576
rect 4924 9636 5024 9664
rect 4924 9576 4932 9636
rect 4932 9576 5012 9636
rect 5012 9576 5024 9636
rect 4924 9572 5024 9576
rect 8056 9632 8156 9660
rect 8056 9572 8064 9632
rect 8064 9572 8144 9632
rect 8144 9572 8156 9632
rect 8056 9568 8156 9572
rect 11200 9632 11300 9660
rect 11200 9572 11208 9632
rect 11208 9572 11288 9632
rect 11288 9572 11300 9632
rect 11200 9568 11300 9572
rect 14402 9636 14502 9664
rect 14402 9576 14410 9636
rect 14410 9576 14490 9636
rect 14490 9576 14502 9636
rect 14402 9572 14502 9576
rect 17546 9636 17646 9664
rect 17546 9576 17554 9636
rect 17554 9576 17634 9636
rect 17634 9576 17646 9636
rect 17546 9572 17646 9576
rect 20678 9632 20778 9660
rect 20678 9572 20686 9632
rect 20686 9572 20766 9632
rect 20766 9572 20778 9632
rect 20678 9568 20778 9572
rect 23816 10146 23892 10148
rect 23816 10094 23820 10146
rect 23820 10094 23886 10146
rect 23886 10094 23892 10146
rect 23816 10090 23892 10094
rect 34107 10895 34223 10951
rect 67977 11130 68115 11142
rect 67977 11072 67990 11130
rect 67990 11072 68102 11130
rect 68102 11072 68115 11130
rect 67977 11060 68115 11072
rect 63989 10964 64051 11022
rect 64051 10964 64053 11022
rect 63989 10960 64053 10964
rect 35247 10413 35307 10475
rect 31923 10331 31993 10337
rect 31923 10269 31925 10331
rect 31925 10269 31983 10331
rect 31983 10269 31993 10331
rect 31923 10265 31993 10269
rect 23822 9632 23922 9660
rect 23822 9572 23830 9632
rect 23830 9572 23910 9632
rect 23910 9572 23922 9632
rect 23822 9568 23922 9572
rect 31066 9449 31158 9456
rect 31066 9375 31077 9449
rect 31077 9375 31148 9449
rect 31148 9375 31158 9449
rect 31066 9364 31158 9375
rect 29695 8204 29765 8216
rect 29695 8150 29703 8204
rect 29703 8150 29757 8204
rect 29757 8150 29765 8204
rect 29695 8138 29765 8150
rect 31925 8262 31995 8268
rect 31925 8200 31927 8262
rect 31927 8200 31985 8262
rect 31985 8200 31995 8262
rect 31925 8196 31995 8200
rect 1784 7418 1860 7420
rect 1784 7366 1788 7418
rect 1788 7366 1854 7418
rect 1854 7366 1860 7418
rect 1784 7362 1860 7366
rect 4928 7418 5004 7420
rect 4928 7366 4932 7418
rect 4932 7366 4998 7418
rect 4998 7366 5004 7418
rect 4928 7362 5004 7366
rect 8060 7414 8136 7416
rect 8060 7362 8064 7414
rect 8064 7362 8130 7414
rect 8130 7362 8136 7414
rect 8060 7358 8136 7362
rect 11204 7414 11280 7416
rect 11204 7362 11208 7414
rect 11208 7362 11274 7414
rect 11274 7362 11280 7414
rect 11204 7358 11280 7362
rect 14406 7418 14482 7420
rect 14406 7366 14410 7418
rect 14410 7366 14476 7418
rect 14476 7366 14482 7418
rect 14406 7362 14482 7366
rect 17550 7418 17626 7420
rect 17550 7366 17554 7418
rect 17554 7366 17620 7418
rect 17620 7366 17626 7418
rect 17550 7362 17626 7366
rect 20682 7414 20758 7416
rect 20682 7362 20686 7414
rect 20686 7362 20752 7414
rect 20752 7362 20758 7414
rect 20682 7358 20758 7362
rect 23826 7414 23902 7416
rect 23826 7362 23830 7414
rect 23830 7362 23896 7414
rect 23896 7362 23902 7414
rect 23826 7358 23902 7362
rect 31072 7372 31157 7384
rect 31072 7307 31084 7372
rect 31084 7307 31147 7372
rect 31147 7307 31157 7372
rect 31072 7298 31157 7307
rect 27506 7096 27562 7158
rect 27506 6805 27562 6867
rect 3273 6751 3367 6761
rect 3273 6677 3283 6751
rect 3283 6677 3359 6751
rect 3359 6677 3367 6751
rect 4011 6751 4105 6761
rect 4011 6677 4021 6751
rect 4021 6677 4097 6751
rect 4097 6677 4105 6751
rect 4749 6751 4843 6761
rect 4749 6677 4759 6751
rect 4759 6677 4835 6751
rect 4835 6677 4843 6751
rect 5487 6751 5581 6761
rect 5487 6677 5497 6751
rect 5497 6677 5573 6751
rect 5573 6677 5581 6751
rect 6227 6751 6321 6761
rect 6227 6677 6237 6751
rect 6237 6677 6313 6751
rect 6313 6677 6321 6751
rect 6969 6751 7063 6761
rect 6969 6677 6979 6751
rect 6979 6677 7055 6751
rect 7055 6677 7063 6751
rect 7707 6751 7801 6761
rect 7707 6677 7717 6751
rect 7717 6677 7793 6751
rect 7793 6677 7801 6751
rect 8445 6753 8539 6763
rect 8445 6679 8455 6753
rect 8455 6679 8531 6753
rect 8531 6679 8539 6753
rect 10049 6698 10127 6706
rect 10049 6644 10061 6698
rect 10061 6644 10115 6698
rect 10115 6644 10127 6698
rect 10049 6636 10127 6644
rect 12117 6696 12195 6704
rect 12117 6642 12129 6696
rect 12129 6642 12183 6696
rect 12183 6642 12195 6696
rect 12117 6634 12195 6642
rect 14186 6698 14264 6706
rect 14186 6644 14198 6698
rect 14198 6644 14252 6698
rect 14252 6644 14264 6698
rect 14186 6636 14264 6644
rect 16254 6696 16332 6704
rect 16254 6642 16266 6696
rect 16266 6642 16320 6696
rect 16320 6642 16332 6696
rect 16254 6634 16332 6642
rect 18323 6696 18401 6704
rect 18323 6642 18335 6696
rect 18335 6642 18389 6696
rect 18389 6642 18401 6696
rect 18323 6634 18401 6642
rect 20391 6694 20469 6702
rect 20391 6640 20403 6694
rect 20403 6640 20457 6694
rect 20457 6640 20469 6694
rect 20391 6632 20469 6640
rect 22460 6696 22538 6704
rect 22460 6642 22472 6696
rect 22472 6642 22526 6696
rect 22526 6642 22538 6696
rect 22460 6634 22538 6642
rect 24528 6694 24606 6702
rect 24528 6640 24540 6694
rect 24540 6640 24594 6694
rect 24594 6640 24606 6694
rect 24528 6632 24606 6640
rect 27507 6499 27563 6561
rect 27506 6338 27562 6400
rect 27506 6187 27562 6249
rect 27506 6026 27562 6088
rect 29693 6136 29763 6148
rect 29693 6082 29701 6136
rect 29701 6082 29755 6136
rect 29755 6082 29763 6136
rect 29693 6070 29763 6082
rect 10847 5896 10930 5905
rect 3353 5805 3419 5863
rect 4091 5805 4157 5863
rect 4829 5805 4895 5863
rect 5567 5805 5633 5863
rect 6307 5805 6373 5863
rect 7049 5805 7115 5863
rect 7787 5805 7853 5863
rect 8525 5807 8591 5865
rect 10847 5830 10857 5896
rect 10857 5830 10923 5896
rect 10923 5830 10930 5896
rect 10847 5825 10930 5830
rect 12927 5829 12991 5893
rect 12991 5829 12994 5893
rect 15000 5830 15060 5896
rect 15060 5830 15065 5896
rect 17061 5894 17128 5896
rect 15000 5828 15065 5830
rect 17061 5828 17062 5894
rect 17062 5828 17128 5894
rect 19132 5828 19196 5893
rect 23264 5894 23339 5910
rect 17061 5827 17128 5828
rect 21199 5826 21265 5892
rect 21265 5826 21268 5892
rect 23264 5828 23268 5894
rect 23268 5828 23334 5894
rect 23334 5828 23339 5894
rect 23264 5824 23339 5828
rect 25624 5885 25690 5886
rect 25624 5832 25628 5885
rect 25628 5832 25688 5885
rect 25688 5832 25690 5885
rect 25624 5829 25690 5832
rect 27506 5839 27562 5901
rect 25346 5627 25417 5704
rect 27506 5635 27562 5697
rect 31923 6194 31993 6200
rect 31923 6132 31925 6194
rect 31925 6132 31983 6194
rect 31983 6132 31993 6194
rect 31923 6128 31993 6132
rect 31067 5304 31156 5314
rect 31067 5240 31076 5304
rect 31076 5240 31149 5304
rect 31149 5240 31156 5304
rect 31067 5229 31156 5240
rect 474 4635 569 4640
rect 474 4566 483 4635
rect 483 4566 563 4635
rect 563 4566 569 4635
rect 474 4562 569 4566
rect 248 4483 358 4486
rect 248 4405 257 4483
rect 257 4405 352 4483
rect 352 4405 358 4483
rect 248 4397 358 4405
rect 10107 4474 10179 4476
rect 10107 4416 10111 4474
rect 10111 4416 10173 4474
rect 10173 4416 10179 4474
rect 10107 4406 10179 4416
rect 12175 4472 12247 4474
rect 12175 4414 12179 4472
rect 12179 4414 12241 4472
rect 12241 4414 12247 4472
rect 12175 4404 12247 4414
rect 14244 4474 14316 4476
rect 14244 4416 14248 4474
rect 14248 4416 14310 4474
rect 14310 4416 14316 4474
rect 14244 4406 14316 4416
rect 16312 4472 16384 4474
rect 16312 4414 16316 4472
rect 16316 4414 16378 4472
rect 16378 4414 16384 4472
rect 16312 4404 16384 4414
rect 18381 4472 18453 4474
rect 18381 4414 18385 4472
rect 18385 4414 18447 4472
rect 18447 4414 18453 4472
rect 18381 4404 18453 4414
rect 20449 4470 20521 4472
rect 20449 4412 20453 4470
rect 20453 4412 20515 4470
rect 20515 4412 20521 4470
rect 20449 4402 20521 4412
rect 22518 4472 22590 4474
rect 22518 4414 22522 4472
rect 22522 4414 22584 4472
rect 22584 4414 22590 4472
rect 22518 4404 22590 4414
rect 24586 4470 24658 4472
rect 24586 4412 24590 4470
rect 24590 4412 24652 4470
rect 24652 4412 24658 4470
rect 24586 4402 24658 4412
rect -10 4287 95 4290
rect -10 4213 3 4287
rect 3 4213 84 4287
rect 84 4213 95 4287
rect -10 4206 95 4213
rect 29693 4067 29763 4079
rect 29693 4013 29701 4067
rect 29701 4013 29755 4067
rect 29755 4013 29763 4067
rect 29693 4001 29763 4013
rect 31923 4125 31993 4131
rect 31923 4063 31925 4125
rect 31925 4063 31983 4125
rect 31983 4063 31993 4125
rect 31923 4059 31993 4063
rect 135 3214 214 3277
rect -22 2773 43 2875
rect 130 2627 214 2684
rect 1496 2384 1596 2412
rect 1496 2324 1508 2384
rect 1508 2324 1588 2384
rect 1588 2324 1596 2384
rect 1496 2320 1596 2324
rect 4640 2384 4740 2412
rect 4640 2324 4652 2384
rect 4652 2324 4732 2384
rect 4732 2324 4740 2384
rect 4640 2320 4740 2324
rect 7772 2388 7872 2416
rect 7772 2328 7784 2388
rect 7784 2328 7864 2388
rect 7864 2328 7872 2388
rect 7772 2324 7872 2328
rect 10916 2388 11016 2416
rect 10916 2328 10928 2388
rect 10928 2328 11008 2388
rect 11008 2328 11016 2388
rect 10916 2324 11016 2328
rect 14118 2384 14218 2412
rect 14118 2324 14130 2384
rect 14130 2324 14210 2384
rect 14210 2324 14218 2384
rect 14118 2320 14218 2324
rect 17262 2384 17362 2412
rect 17262 2324 17274 2384
rect 17274 2324 17354 2384
rect 17354 2324 17362 2384
rect 17262 2320 17362 2324
rect 20394 2388 20494 2416
rect 20394 2328 20406 2388
rect 20406 2328 20486 2388
rect 20486 2328 20494 2388
rect 20394 2324 20494 2328
rect 31070 3238 31154 3245
rect 31070 3172 31079 3238
rect 31079 3172 31144 3238
rect 31144 3172 31154 3238
rect 31070 3162 31154 3172
rect 23538 2388 23638 2416
rect 23538 2328 23550 2388
rect 23550 2328 23630 2388
rect 23630 2328 23638 2388
rect 23538 2324 23638 2328
rect 29691 1999 29761 2011
rect 29691 1945 29699 1999
rect 29699 1945 29753 1999
rect 29753 1945 29761 1999
rect 29691 1933 29761 1945
rect 31921 2057 31991 2063
rect 31921 1995 31923 2057
rect 31923 1995 31981 2057
rect 31981 1995 31991 2057
rect 31921 1991 31991 1995
rect 31069 1171 31152 1178
rect 31069 1101 31079 1171
rect 31079 1101 31144 1171
rect 31144 1101 31152 1171
rect 31069 1094 31152 1101
rect 35469 9211 35531 9269
rect 35531 9211 35533 9269
rect 35469 9207 35533 9211
rect 35239 7828 35299 7890
rect 35461 6626 35523 6684
rect 35523 6626 35525 6684
rect 35461 6622 35525 6626
rect 34114 1032 34217 1040
rect 34114 969 34127 1032
rect 34127 969 34208 1032
rect 34208 969 34217 1032
rect 34114 961 34217 969
rect 1516 166 1592 168
rect 1516 114 1522 166
rect 1522 114 1588 166
rect 1588 114 1592 166
rect 1516 110 1592 114
rect 4660 166 4736 168
rect 4660 114 4666 166
rect 4666 114 4732 166
rect 4732 114 4736 166
rect 4660 110 4736 114
rect 7792 170 7868 172
rect 7792 118 7798 170
rect 7798 118 7864 170
rect 7864 118 7868 170
rect 7792 114 7868 118
rect 10936 170 11012 172
rect 10936 118 10942 170
rect 10942 118 11008 170
rect 11008 118 11012 170
rect 10936 114 11012 118
rect 14138 166 14214 168
rect 14138 114 14144 166
rect 14144 114 14210 166
rect 14210 114 14214 166
rect 14138 110 14214 114
rect 17282 166 17358 168
rect 17282 114 17288 166
rect 17288 114 17354 166
rect 17354 114 17358 166
rect 17282 110 17358 114
rect 20414 170 20490 172
rect 20414 118 20420 170
rect 20420 118 20486 170
rect 20486 118 20490 170
rect 20414 114 20490 118
rect 23558 170 23634 172
rect 23558 118 23564 170
rect 23564 118 23630 170
rect 23630 118 23634 170
rect 23558 114 23634 118
rect 29693 -70 29763 -58
rect 29693 -124 29701 -70
rect 29701 -124 29755 -70
rect 29755 -124 29763 -70
rect 29693 -136 29763 -124
rect 1528 -1508 1628 -1480
rect 1528 -1568 1540 -1508
rect 1540 -1568 1620 -1508
rect 1620 -1568 1628 -1508
rect 1528 -1572 1628 -1568
rect 4672 -1508 4772 -1480
rect 4672 -1568 4684 -1508
rect 4684 -1568 4764 -1508
rect 4764 -1568 4772 -1508
rect 4672 -1572 4772 -1568
rect 7804 -1504 7904 -1476
rect 7804 -1564 7816 -1504
rect 7816 -1564 7896 -1504
rect 7896 -1564 7904 -1504
rect 7804 -1568 7904 -1564
rect 10948 -1504 11048 -1476
rect 10948 -1564 10960 -1504
rect 10960 -1564 11040 -1504
rect 11040 -1564 11048 -1504
rect 10948 -1568 11048 -1564
rect 14150 -1508 14250 -1480
rect 14150 -1568 14162 -1508
rect 14162 -1568 14242 -1508
rect 14242 -1568 14250 -1508
rect 14150 -1572 14250 -1568
rect -165 -2796 -77 -2718
rect 3188 -2798 3249 -2734
rect 6318 -2800 6401 -2737
rect 17294 -1508 17394 -1480
rect 17294 -1568 17306 -1508
rect 17306 -1568 17386 -1508
rect 17386 -1568 17394 -1508
rect 17294 -1572 17394 -1568
rect 20426 -1504 20526 -1476
rect 20426 -1564 20438 -1504
rect 20438 -1564 20518 -1504
rect 20518 -1564 20526 -1504
rect 20426 -1568 20526 -1564
rect 31923 -12 31993 -6
rect 31923 -74 31925 -12
rect 31925 -74 31983 -12
rect 31983 -74 31993 -12
rect 31923 -78 31993 -74
rect 31067 -898 31157 -891
rect 31067 -968 31076 -898
rect 31076 -968 31149 -898
rect 31149 -968 31157 -898
rect 31067 -978 31157 -968
rect 23570 -1504 23670 -1476
rect 23570 -1564 23582 -1504
rect 23582 -1564 23662 -1504
rect 23662 -1564 23670 -1504
rect 23570 -1568 23670 -1564
rect 29691 -2138 29761 -2126
rect 29691 -2192 29699 -2138
rect 29699 -2192 29753 -2138
rect 29753 -2192 29761 -2138
rect 29691 -2204 29761 -2192
rect 31921 -2080 31991 -2074
rect 31921 -2142 31923 -2080
rect 31923 -2142 31981 -2080
rect 31981 -2142 31991 -2080
rect 31921 -2146 31991 -2142
rect 35220 4550 35280 4612
rect 35442 3348 35504 3406
rect 35504 3348 35506 3406
rect 35442 3344 35506 3348
rect 35236 1790 35296 1852
rect 35458 588 35520 646
rect 35520 588 35522 646
rect 35458 584 35522 588
rect 9462 -2798 9581 -2737
rect 12693 -2811 12758 -2730
rect 67590 10556 67652 10614
rect 67652 10556 67654 10614
rect 67590 10552 67654 10556
rect 47257 10410 47410 10421
rect 44775 10356 44928 10367
rect 40708 10322 40861 10333
rect 38226 10268 38379 10279
rect 38226 10160 38237 10268
rect 38237 10160 38369 10268
rect 38369 10160 38379 10268
rect 40708 10214 40719 10322
rect 40719 10214 40851 10322
rect 40851 10214 40861 10322
rect 41855 10322 42008 10333
rect 40708 10204 40861 10214
rect 38226 10150 38379 10160
rect 41855 10214 41866 10322
rect 41866 10214 41998 10322
rect 41998 10214 42008 10322
rect 44775 10248 44786 10356
rect 44786 10248 44918 10356
rect 44918 10248 44928 10356
rect 47257 10302 47268 10410
rect 47268 10302 47400 10410
rect 47400 10302 47410 10410
rect 48404 10410 48557 10421
rect 47257 10292 47410 10302
rect 44775 10238 44928 10248
rect 48404 10302 48415 10410
rect 48415 10302 48547 10410
rect 48547 10302 48557 10410
rect 60536 10410 60689 10421
rect 53911 10342 54064 10353
rect 48404 10292 48557 10302
rect 51429 10288 51582 10299
rect 41855 10204 42008 10214
rect 38507 9229 38636 9240
rect 38507 9097 38517 9229
rect 38517 9097 38625 9229
rect 38625 9097 38636 9229
rect 38507 9087 38636 9097
rect 38240 8618 38393 8629
rect 38240 8510 38251 8618
rect 38251 8510 38383 8618
rect 38383 8510 38393 8618
rect 38240 8500 38393 8510
rect 38521 7579 38650 7590
rect 38521 7447 38531 7579
rect 38531 7447 38639 7579
rect 38639 7447 38650 7579
rect 38521 7437 38650 7447
rect 37273 7142 37388 7151
rect 37273 7063 37283 7142
rect 37283 7063 37376 7142
rect 37376 7063 37388 7142
rect 37273 7054 37388 7063
rect 38235 7014 38388 7025
rect 38235 6906 38246 7014
rect 38246 6906 38378 7014
rect 38378 6906 38388 7014
rect 38235 6896 38388 6906
rect 42945 9414 43090 9489
rect 45056 9317 45185 9328
rect 45056 9185 45066 9317
rect 45066 9185 45174 9317
rect 45174 9185 45185 9317
rect 45056 9175 45185 9185
rect 40055 8922 40208 8932
rect 40055 8814 40065 8922
rect 40065 8814 40197 8922
rect 40197 8814 40208 8922
rect 40055 8803 40208 8814
rect 41197 8920 41350 8930
rect 41197 8812 41207 8920
rect 41207 8812 41339 8920
rect 41339 8812 41350 8920
rect 41197 8801 41350 8812
rect 44789 8706 44942 8717
rect 44789 8598 44800 8706
rect 44800 8598 44932 8706
rect 44932 8598 44942 8706
rect 44789 8588 44942 8598
rect 40053 8275 40206 8286
rect 40053 8167 40064 8275
rect 40064 8167 40196 8275
rect 40196 8167 40206 8275
rect 40053 8157 40206 8167
rect 41951 8275 42104 8286
rect 41951 8167 41962 8275
rect 41962 8167 42094 8275
rect 42094 8167 42104 8275
rect 41951 8157 42104 8167
rect 45070 7667 45199 7678
rect 45070 7535 45080 7667
rect 45080 7535 45188 7667
rect 45188 7535 45199 7667
rect 45070 7525 45199 7535
rect 40694 7305 40772 7315
rect 40694 7239 40709 7305
rect 40709 7239 40772 7305
rect 40694 7229 40772 7239
rect 38516 5975 38645 5986
rect 38516 5843 38526 5975
rect 38526 5843 38634 5975
rect 38634 5843 38645 5975
rect 38516 5833 38645 5843
rect 39999 5879 40152 5889
rect 39999 5771 40009 5879
rect 40009 5771 40141 5879
rect 40141 5771 40152 5879
rect 39999 5760 40152 5771
rect 41897 5879 42050 5889
rect 41897 5771 41907 5879
rect 41907 5771 42039 5879
rect 42039 5771 42050 5879
rect 41897 5760 42050 5771
rect 43822 7230 43937 7239
rect 43822 7151 43832 7230
rect 43832 7151 43925 7230
rect 43925 7151 43937 7230
rect 43822 7142 43937 7151
rect 44784 7102 44937 7113
rect 44784 6994 44795 7102
rect 44795 6994 44927 7102
rect 44927 6994 44937 7102
rect 44784 6984 44937 6994
rect 51429 10180 51440 10288
rect 51440 10180 51572 10288
rect 51572 10180 51582 10288
rect 53911 10234 53922 10342
rect 53922 10234 54054 10342
rect 54054 10234 54064 10342
rect 55058 10342 55211 10353
rect 53911 10224 54064 10234
rect 51429 10170 51582 10180
rect 55058 10234 55069 10342
rect 55069 10234 55201 10342
rect 55201 10234 55211 10342
rect 55058 10224 55211 10234
rect 58054 10356 58207 10367
rect 58054 10248 58065 10356
rect 58065 10248 58197 10356
rect 58197 10248 58207 10356
rect 60536 10302 60547 10410
rect 60547 10302 60679 10410
rect 60679 10302 60689 10410
rect 61683 10410 61836 10421
rect 60536 10292 60689 10302
rect 58054 10238 58207 10248
rect 61683 10302 61694 10410
rect 61694 10302 61826 10410
rect 61826 10302 61836 10410
rect 61683 10292 61836 10302
rect 51710 9249 51839 9260
rect 51710 9117 51720 9249
rect 51720 9117 51828 9249
rect 51828 9117 51839 9249
rect 51710 9107 51839 9117
rect 46604 9010 46757 9020
rect 46604 8902 46614 9010
rect 46614 8902 46746 9010
rect 46746 8902 46757 9010
rect 46604 8891 46757 8902
rect 47746 9008 47899 9018
rect 47746 8900 47756 9008
rect 47756 8900 47888 9008
rect 47888 8900 47899 9008
rect 47746 8889 47899 8900
rect 51443 8638 51596 8649
rect 51443 8530 51454 8638
rect 51454 8530 51586 8638
rect 51586 8530 51596 8638
rect 46602 8363 46755 8374
rect 46602 8255 46613 8363
rect 46613 8255 46745 8363
rect 46745 8255 46755 8363
rect 46602 8245 46755 8255
rect 48500 8363 48653 8374
rect 48500 8255 48511 8363
rect 48511 8255 48643 8363
rect 48643 8255 48653 8363
rect 48500 8245 48653 8255
rect 47243 7393 47321 7403
rect 47243 7327 47258 7393
rect 47258 7327 47321 7393
rect 47243 7317 47321 7327
rect 51443 8520 51596 8530
rect 51724 7599 51853 7610
rect 51724 7467 51734 7599
rect 51734 7467 51842 7599
rect 51842 7467 51853 7599
rect 51724 7457 51853 7467
rect 50476 7162 50591 7171
rect 50476 7083 50486 7162
rect 50486 7083 50579 7162
rect 50579 7083 50591 7162
rect 50476 7074 50591 7083
rect 45065 6063 45194 6074
rect 45065 5931 45075 6063
rect 45075 5931 45183 6063
rect 45183 5931 45194 6063
rect 45065 5921 45194 5931
rect 46548 5967 46701 5977
rect 46548 5859 46558 5967
rect 46558 5859 46690 5967
rect 46690 5859 46701 5967
rect 46548 5848 46701 5859
rect 48446 5967 48599 5977
rect 48446 5859 48456 5967
rect 48456 5859 48588 5967
rect 48588 5859 48599 5967
rect 48446 5848 48599 5859
rect 51438 7034 51591 7045
rect 51438 6926 51449 7034
rect 51449 6926 51581 7034
rect 51581 6926 51591 7034
rect 51438 6916 51591 6926
rect 56079 9435 56176 9509
rect 58335 9317 58464 9328
rect 58335 9185 58345 9317
rect 58345 9185 58453 9317
rect 58453 9185 58464 9317
rect 58335 9175 58464 9185
rect 53258 8942 53411 8952
rect 53258 8834 53268 8942
rect 53268 8834 53400 8942
rect 53400 8834 53411 8942
rect 53258 8823 53411 8834
rect 54400 8940 54553 8950
rect 54400 8832 54410 8940
rect 54410 8832 54542 8940
rect 54542 8832 54553 8940
rect 54400 8821 54553 8832
rect 58068 8706 58221 8717
rect 58068 8598 58079 8706
rect 58079 8598 58211 8706
rect 58211 8598 58221 8706
rect 58068 8588 58221 8598
rect 53256 8295 53409 8306
rect 53256 8187 53267 8295
rect 53267 8187 53399 8295
rect 53399 8187 53409 8295
rect 53256 8177 53409 8187
rect 55154 8295 55307 8306
rect 55154 8187 55165 8295
rect 55165 8187 55297 8295
rect 55297 8187 55307 8295
rect 55154 8177 55307 8187
rect 58349 7667 58478 7678
rect 58349 7535 58359 7667
rect 58359 7535 58467 7667
rect 58467 7535 58478 7667
rect 58349 7525 58478 7535
rect 53897 7325 53975 7335
rect 53897 7259 53912 7325
rect 53912 7259 53975 7325
rect 53897 7249 53975 7259
rect 56632 6724 56728 6824
rect 51719 5995 51848 6006
rect 51719 5863 51729 5995
rect 51729 5863 51837 5995
rect 51837 5863 51848 5995
rect 51719 5853 51848 5863
rect 53202 5899 53355 5909
rect 53202 5791 53212 5899
rect 53212 5791 53344 5899
rect 53344 5791 53355 5899
rect 53202 5780 53355 5791
rect 55100 5899 55253 5909
rect 55100 5791 55110 5899
rect 55110 5791 55242 5899
rect 55242 5791 55253 5899
rect 55100 5780 55253 5791
rect 56152 5512 56294 5520
rect 56152 5398 56163 5512
rect 56163 5398 56286 5512
rect 56286 5398 56294 5512
rect 56152 5386 56294 5398
rect 57101 7230 57216 7239
rect 57101 7151 57111 7230
rect 57111 7151 57204 7230
rect 57204 7151 57216 7230
rect 57101 7142 57216 7151
rect 58063 7102 58216 7113
rect 58063 6994 58074 7102
rect 58074 6994 58206 7102
rect 58206 6994 58216 7102
rect 58063 6984 58216 6994
rect 59883 9010 60036 9020
rect 59883 8902 59893 9010
rect 59893 8902 60025 9010
rect 60025 8902 60036 9010
rect 59883 8891 60036 8902
rect 61025 9008 61178 9018
rect 61025 8900 61035 9008
rect 61035 8900 61167 9008
rect 61167 8900 61178 9008
rect 61025 8889 61178 8900
rect 65935 9822 66146 9838
rect 65935 9699 65954 9822
rect 65954 9699 66128 9822
rect 66128 9699 66146 9822
rect 65935 9681 66146 9699
rect 63762 9595 63822 9657
rect 63984 8393 64046 8451
rect 64046 8393 64048 8451
rect 63984 8389 64048 8393
rect 59881 8363 60034 8374
rect 59881 8255 59892 8363
rect 59892 8255 60024 8363
rect 60024 8255 60034 8363
rect 59881 8245 60034 8255
rect 61779 8363 61932 8374
rect 61779 8255 61790 8363
rect 61790 8255 61922 8363
rect 61922 8255 61932 8363
rect 61779 8245 61932 8255
rect 66015 8066 66168 8077
rect 66015 7958 66026 8066
rect 66026 7958 66158 8066
rect 66158 7958 66168 8066
rect 66015 7948 66168 7958
rect 67370 7667 67430 7729
rect 60522 7393 60600 7403
rect 60522 7327 60537 7393
rect 60537 7327 60600 7393
rect 60522 7317 60600 7327
rect 70241 20813 70333 20825
rect 70241 20733 70269 20813
rect 70269 20733 70329 20813
rect 70329 20733 70333 20813
rect 70241 20725 70333 20733
rect 72485 20799 72543 20805
rect 72485 20733 72487 20799
rect 72487 20733 72539 20799
rect 72539 20733 72543 20799
rect 72485 20729 72543 20733
rect 70241 17669 70333 17681
rect 70241 17589 70269 17669
rect 70269 17589 70329 17669
rect 70329 17589 70333 17669
rect 70241 17581 70333 17589
rect 72485 17655 72543 17661
rect 72485 17589 72487 17655
rect 72487 17589 72539 17655
rect 72539 17589 72543 17655
rect 72485 17585 72543 17589
rect 70237 14537 70329 14549
rect 70237 14457 70265 14537
rect 70265 14457 70325 14537
rect 70325 14457 70329 14537
rect 70237 14449 70329 14457
rect 72481 14523 72539 14529
rect 72481 14457 72483 14523
rect 72483 14457 72535 14523
rect 72535 14457 72539 14523
rect 72481 14453 72539 14457
rect 70237 11393 70329 11405
rect 70237 11313 70265 11393
rect 70265 11313 70325 11393
rect 70325 11313 70329 11393
rect 70237 11305 70329 11313
rect 71494 12691 71557 12788
rect 72481 11379 72539 11385
rect 72481 11313 72483 11379
rect 72483 11313 72535 11379
rect 72535 11313 72539 11379
rect 72481 11309 72539 11313
rect 63762 6562 63822 6624
rect 67592 6465 67654 6523
rect 67654 6465 67656 6523
rect 67592 6461 67656 6465
rect 70241 8191 70333 8203
rect 70241 8111 70269 8191
rect 70269 8111 70329 8191
rect 70329 8111 70333 8191
rect 70241 8103 70333 8111
rect 72485 8177 72543 8183
rect 72485 8111 72487 8177
rect 72487 8111 72539 8177
rect 72539 8111 72543 8177
rect 72485 8107 72543 8111
rect 58344 6063 58473 6074
rect 58344 5931 58354 6063
rect 58354 5931 58462 6063
rect 58462 5931 58473 6063
rect 58344 5921 58473 5931
rect 59827 5967 59980 5977
rect 59827 5859 59837 5967
rect 59837 5859 59969 5967
rect 59969 5859 59980 5967
rect 59827 5848 59980 5859
rect 61725 5967 61878 5977
rect 61725 5859 61735 5967
rect 61735 5859 61867 5967
rect 61867 5859 61878 5967
rect 61725 5848 61878 5859
rect 57261 5512 57403 5520
rect 57261 5398 57272 5512
rect 57272 5398 57395 5512
rect 57395 5398 57403 5512
rect 57261 5386 57403 5398
rect 40700 4542 40853 4553
rect 38218 4488 38371 4499
rect 38218 4380 38229 4488
rect 38229 4380 38361 4488
rect 38361 4380 38371 4488
rect 40700 4434 40711 4542
rect 40711 4434 40843 4542
rect 40843 4434 40853 4542
rect 41847 4542 42000 4553
rect 40700 4424 40853 4434
rect 38218 4370 38371 4380
rect 41847 4434 41858 4542
rect 41858 4434 41990 4542
rect 41990 4434 42000 4542
rect 47251 4540 47404 4551
rect 41847 4424 42000 4434
rect 44769 4486 44922 4497
rect 38499 3449 38628 3460
rect 38499 3317 38509 3449
rect 38509 3317 38617 3449
rect 38617 3317 38628 3449
rect 38499 3307 38628 3317
rect 38232 2838 38385 2849
rect 38232 2730 38243 2838
rect 38243 2730 38375 2838
rect 38375 2730 38385 2838
rect 38232 2720 38385 2730
rect 36885 1619 37119 1756
rect 38513 1799 38642 1810
rect 38513 1667 38523 1799
rect 38523 1667 38631 1799
rect 38631 1667 38642 1799
rect 38513 1657 38642 1667
rect 37265 1362 37380 1371
rect 37265 1283 37275 1362
rect 37275 1283 37368 1362
rect 37368 1283 37380 1362
rect 37265 1274 37380 1283
rect 38227 1234 38380 1245
rect 38227 1126 38238 1234
rect 38238 1126 38370 1234
rect 38370 1126 38380 1234
rect 38227 1116 38380 1126
rect 44769 4378 44780 4486
rect 44780 4378 44912 4486
rect 44912 4378 44922 4486
rect 47251 4432 47262 4540
rect 47262 4432 47394 4540
rect 47394 4432 47404 4540
rect 48398 4540 48551 4551
rect 47251 4422 47404 4432
rect 44769 4368 44922 4378
rect 48398 4432 48409 4540
rect 48409 4432 48541 4540
rect 48541 4432 48551 4540
rect 48398 4422 48551 4432
rect 45050 3447 45179 3458
rect 45050 3315 45060 3447
rect 45060 3315 45168 3447
rect 45168 3315 45179 3447
rect 45050 3305 45179 3315
rect 40047 3142 40200 3152
rect 40047 3034 40057 3142
rect 40057 3034 40189 3142
rect 40189 3034 40200 3142
rect 40047 3023 40200 3034
rect 41189 3140 41342 3150
rect 41189 3032 41199 3140
rect 41199 3032 41331 3140
rect 41331 3032 41342 3140
rect 41189 3021 41342 3032
rect 44783 2836 44936 2847
rect 44783 2728 44794 2836
rect 44794 2728 44926 2836
rect 44926 2728 44936 2836
rect 44783 2718 44936 2728
rect 40045 2495 40198 2506
rect 40045 2387 40056 2495
rect 40056 2387 40188 2495
rect 40188 2387 40198 2495
rect 40045 2377 40198 2387
rect 41943 2495 42096 2506
rect 41943 2387 41954 2495
rect 41954 2387 42086 2495
rect 42086 2387 42096 2495
rect 41943 2377 42096 2387
rect 43520 1613 43743 1749
rect 45064 1797 45193 1808
rect 45064 1665 45074 1797
rect 45074 1665 45182 1797
rect 45182 1665 45193 1797
rect 45064 1655 45193 1665
rect 40686 1525 40764 1535
rect 40686 1459 40701 1525
rect 40701 1459 40764 1525
rect 40686 1449 40764 1459
rect 43816 1360 43931 1369
rect 43816 1281 43826 1360
rect 43826 1281 43919 1360
rect 43919 1281 43931 1360
rect 43816 1272 43931 1281
rect 38508 195 38637 206
rect 38508 63 38518 195
rect 38518 63 38626 195
rect 38626 63 38637 195
rect 38508 53 38637 63
rect 39991 99 40144 109
rect 39991 -9 40001 99
rect 40001 -9 40133 99
rect 40133 -9 40144 99
rect 39991 -20 40144 -9
rect 41889 99 42042 109
rect 41889 -9 41899 99
rect 41899 -9 42031 99
rect 42031 -9 42042 99
rect 41889 -20 42042 -9
rect 44778 1232 44931 1243
rect 44778 1124 44789 1232
rect 44789 1124 44921 1232
rect 44921 1124 44931 1232
rect 44778 1114 44931 1124
rect 53906 4541 54059 4552
rect 51424 4487 51577 4498
rect 51424 4379 51435 4487
rect 51435 4379 51567 4487
rect 51567 4379 51577 4487
rect 53906 4433 53917 4541
rect 53917 4433 54049 4541
rect 54049 4433 54059 4541
rect 55053 4541 55206 4552
rect 53906 4423 54059 4433
rect 51424 4369 51577 4379
rect 55053 4433 55064 4541
rect 55064 4433 55196 4541
rect 55196 4433 55206 4541
rect 60528 4542 60681 4553
rect 55053 4423 55206 4433
rect 58046 4488 58199 4499
rect 51705 3448 51834 3459
rect 51705 3316 51715 3448
rect 51715 3316 51823 3448
rect 51823 3316 51834 3448
rect 51705 3306 51834 3316
rect 46598 3140 46751 3150
rect 46598 3032 46608 3140
rect 46608 3032 46740 3140
rect 46740 3032 46751 3140
rect 46598 3021 46751 3032
rect 47740 3138 47893 3148
rect 47740 3030 47750 3138
rect 47750 3030 47882 3138
rect 47882 3030 47893 3138
rect 47740 3019 47893 3030
rect 51438 2837 51591 2848
rect 51438 2729 51449 2837
rect 51449 2729 51581 2837
rect 51581 2729 51591 2837
rect 51438 2719 51591 2729
rect 46596 2493 46749 2504
rect 46596 2385 46607 2493
rect 46607 2385 46739 2493
rect 46739 2385 46749 2493
rect 46596 2375 46749 2385
rect 48494 2493 48647 2504
rect 48494 2385 48505 2493
rect 48505 2385 48637 2493
rect 48637 2385 48647 2493
rect 48494 2375 48647 2385
rect 50201 1622 50345 1734
rect 51719 1798 51848 1809
rect 51719 1666 51729 1798
rect 51729 1666 51837 1798
rect 51837 1666 51848 1798
rect 51719 1656 51848 1666
rect 47237 1523 47315 1533
rect 47237 1457 47252 1523
rect 47252 1457 47315 1523
rect 47237 1447 47315 1457
rect 50471 1361 50586 1370
rect 50471 1282 50481 1361
rect 50481 1282 50574 1361
rect 50574 1282 50586 1361
rect 50471 1273 50586 1282
rect 45059 193 45188 204
rect 45059 61 45069 193
rect 45069 61 45177 193
rect 45177 61 45188 193
rect 45059 51 45188 61
rect 46542 97 46695 107
rect 46542 -11 46552 97
rect 46552 -11 46684 97
rect 46684 -11 46695 97
rect 46542 -22 46695 -11
rect 48440 97 48593 107
rect 48440 -11 48450 97
rect 48450 -11 48582 97
rect 48582 -11 48593 97
rect 48440 -22 48593 -11
rect 51433 1233 51586 1244
rect 51433 1125 51444 1233
rect 51444 1125 51576 1233
rect 51576 1125 51586 1233
rect 51433 1115 51586 1125
rect 58046 4380 58057 4488
rect 58057 4380 58189 4488
rect 58189 4380 58199 4488
rect 60528 4434 60539 4542
rect 60539 4434 60671 4542
rect 60671 4434 60681 4542
rect 61675 4542 61828 4553
rect 60528 4424 60681 4434
rect 58046 4370 58199 4380
rect 61675 4434 61686 4542
rect 61686 4434 61818 4542
rect 61818 4434 61828 4542
rect 61675 4424 61828 4434
rect 58327 3449 58456 3460
rect 58327 3317 58337 3449
rect 58337 3317 58445 3449
rect 58445 3317 58456 3449
rect 58327 3307 58456 3317
rect 53253 3141 53406 3151
rect 53253 3033 53263 3141
rect 53263 3033 53395 3141
rect 53395 3033 53406 3141
rect 53253 3022 53406 3033
rect 54395 3139 54548 3149
rect 54395 3031 54405 3139
rect 54405 3031 54537 3139
rect 54537 3031 54548 3139
rect 54395 3020 54548 3031
rect 58060 2838 58213 2849
rect 58060 2730 58071 2838
rect 58071 2730 58203 2838
rect 58203 2730 58213 2838
rect 58060 2720 58213 2730
rect 53251 2494 53404 2505
rect 53251 2386 53262 2494
rect 53262 2386 53394 2494
rect 53394 2386 53404 2494
rect 53251 2376 53404 2386
rect 55149 2494 55302 2505
rect 55149 2386 55160 2494
rect 55160 2386 55292 2494
rect 55292 2386 55302 2494
rect 55149 2376 55302 2386
rect 58341 1799 58470 1810
rect 58341 1667 58351 1799
rect 58351 1667 58459 1799
rect 58459 1667 58470 1799
rect 58341 1657 58470 1667
rect 53892 1524 53970 1534
rect 53892 1458 53907 1524
rect 53907 1458 53970 1524
rect 53892 1448 53970 1458
rect 57093 1362 57208 1371
rect 57093 1283 57103 1362
rect 57103 1283 57196 1362
rect 57196 1283 57208 1362
rect 57093 1274 57208 1283
rect 51714 194 51843 205
rect 51714 62 51724 194
rect 51724 62 51832 194
rect 51832 62 51843 194
rect 51714 52 51843 62
rect 53197 98 53350 108
rect 53197 -10 53207 98
rect 53207 -10 53339 98
rect 53339 -10 53350 98
rect 53197 -21 53350 -10
rect 55095 98 55248 108
rect 55095 -10 55105 98
rect 55105 -10 55237 98
rect 55237 -10 55248 98
rect 55095 -21 55248 -10
rect 58055 1234 58208 1245
rect 58055 1126 58066 1234
rect 58066 1126 58198 1234
rect 58198 1126 58208 1234
rect 58055 1116 58208 1126
rect 59875 3142 60028 3152
rect 59875 3034 59885 3142
rect 59885 3034 60017 3142
rect 60017 3034 60028 3142
rect 59875 3023 60028 3034
rect 61017 3140 61170 3150
rect 61017 3032 61027 3140
rect 61027 3032 61159 3140
rect 61159 3032 61170 3140
rect 61017 3021 61170 3032
rect 59873 2495 60026 2506
rect 59873 2387 59884 2495
rect 59884 2387 60016 2495
rect 60016 2387 60026 2495
rect 59873 2377 60026 2387
rect 61771 2495 61924 2506
rect 61771 2387 61782 2495
rect 61782 2387 61914 2495
rect 61914 2387 61924 2495
rect 61771 2377 61924 2387
rect 60514 1525 60592 1535
rect 60514 1459 60529 1525
rect 60529 1459 60592 1525
rect 60514 1449 60592 1459
rect 62787 1017 62919 1023
rect 62787 936 62795 1017
rect 62795 936 62912 1017
rect 62912 936 62919 1017
rect 62787 927 62919 936
rect 65937 5731 66148 5747
rect 65937 5608 65956 5731
rect 65956 5608 66130 5731
rect 66130 5608 66148 5731
rect 65937 5590 66148 5608
rect 63984 5360 64046 5418
rect 64046 5360 64048 5418
rect 63984 5356 64048 5360
rect 63833 4642 63893 4704
rect 66015 4571 66168 4582
rect 66015 4463 66026 4571
rect 66026 4463 66158 4571
rect 66158 4463 66168 4571
rect 66015 4453 66168 4463
rect 67370 4172 67430 4234
rect 63568 3591 63654 3692
rect 65216 3586 65309 3663
rect 63340 3458 63425 3518
rect 64055 3440 64117 3498
rect 64117 3440 64119 3498
rect 64055 3436 64119 3440
rect 71495 6368 71565 6441
rect 70241 5047 70333 5059
rect 70241 4967 70269 5047
rect 70269 4967 70329 5047
rect 70329 4967 70333 5047
rect 70241 4959 70333 4967
rect 72485 5033 72543 5039
rect 72485 4967 72487 5033
rect 72487 4967 72539 5033
rect 72539 4967 72543 5033
rect 72485 4963 72543 4967
rect 67592 2970 67654 3028
rect 67654 2970 67656 3028
rect 67592 2966 67656 2970
rect 65937 2236 66148 2252
rect 65937 2113 65956 2236
rect 65956 2113 66130 2236
rect 66130 2113 66148 2236
rect 65937 2095 66148 2113
rect 63830 1572 63890 1634
rect 63170 608 63254 698
rect 63604 487 63670 551
rect 64052 370 64114 428
rect 64114 370 64116 428
rect 64052 366 64116 370
rect 58336 195 58465 206
rect 58336 63 58346 195
rect 58346 63 58454 195
rect 58454 63 58465 195
rect 58336 53 58465 63
rect 59819 99 59972 109
rect 59819 -9 59829 99
rect 59829 -9 59961 99
rect 59961 -9 59972 99
rect 59819 -20 59972 -9
rect 61717 99 61870 109
rect 61717 -9 61727 99
rect 61727 -9 61859 99
rect 61859 -9 61870 99
rect 61717 -20 61870 -9
rect 66015 223 66168 234
rect 66015 115 66026 223
rect 66026 115 66158 223
rect 66158 115 66168 223
rect 66015 105 66168 115
rect 67370 -176 67430 -114
rect 42168 -717 42232 -713
rect 42168 -775 42230 -717
rect 42230 -775 42232 -717
rect 48722 -712 48786 -708
rect 48722 -770 48784 -712
rect 48784 -770 48786 -712
rect 55371 -724 55435 -720
rect 55371 -782 55433 -724
rect 55433 -782 55435 -724
rect 70237 1915 70329 1927
rect 70237 1835 70265 1915
rect 70265 1835 70325 1915
rect 70325 1835 70329 1915
rect 70237 1827 70329 1835
rect 72481 1901 72539 1907
rect 72481 1835 72483 1901
rect 72483 1835 72535 1901
rect 72535 1835 72539 1901
rect 72481 1831 72539 1835
rect 63584 -1052 63668 -962
rect 68739 -1126 68826 -1053
rect 41946 -1981 42006 -1919
rect 48500 -1976 48560 -1914
rect 63837 -1273 63897 -1211
rect 70237 -1229 70329 -1217
rect 70237 -1309 70265 -1229
rect 70265 -1309 70325 -1229
rect 70325 -1309 70329 -1229
rect 70237 -1317 70329 -1309
rect 67592 -1378 67654 -1320
rect 67654 -1378 67656 -1320
rect 67592 -1382 67656 -1378
rect 72481 -1243 72539 -1237
rect 72481 -1309 72483 -1243
rect 72483 -1309 72535 -1243
rect 72535 -1309 72539 -1243
rect 72481 -1313 72539 -1309
rect 63001 -1795 63083 -1705
rect 55149 -1988 55209 -1926
rect 63168 -2111 63252 -2021
rect 65937 -2112 66148 -2096
rect 65937 -2235 65956 -2112
rect 65956 -2235 66130 -2112
rect 66130 -2235 66148 -2112
rect 65937 -2253 66148 -2235
rect 63481 -2445 63542 -2370
rect 64059 -2475 64121 -2417
rect 64121 -2475 64123 -2417
rect 64059 -2479 64123 -2475
rect 31068 -2968 31154 -2959
rect 31068 -3033 31078 -2968
rect 31078 -3033 31142 -2968
rect 31142 -3033 31154 -2968
rect 31068 -3044 31154 -3033
rect 1548 -3726 1624 -3724
rect 1548 -3778 1554 -3726
rect 1554 -3778 1620 -3726
rect 1620 -3778 1624 -3726
rect 1548 -3782 1624 -3778
rect 4692 -3726 4768 -3724
rect 4692 -3778 4698 -3726
rect 4698 -3778 4764 -3726
rect 4764 -3778 4768 -3726
rect 4692 -3782 4768 -3778
rect 7824 -3722 7900 -3720
rect 7824 -3774 7830 -3722
rect 7830 -3774 7896 -3722
rect 7896 -3774 7900 -3722
rect 7824 -3778 7900 -3774
rect 10968 -3722 11044 -3720
rect 10968 -3774 10974 -3722
rect 10974 -3774 11040 -3722
rect 11040 -3774 11044 -3722
rect 10968 -3778 11044 -3774
rect 14170 -3726 14246 -3724
rect 14170 -3778 14176 -3726
rect 14176 -3778 14242 -3726
rect 14242 -3778 14246 -3726
rect 14170 -3782 14246 -3778
rect 17314 -3726 17390 -3724
rect 17314 -3778 17320 -3726
rect 17320 -3778 17386 -3726
rect 17386 -3778 17390 -3726
rect 17314 -3782 17390 -3778
rect 20446 -3722 20522 -3720
rect 20446 -3774 20452 -3722
rect 20452 -3774 20518 -3722
rect 20518 -3774 20522 -3722
rect 20446 -3778 20522 -3774
rect 23590 -3722 23666 -3720
rect 23590 -3774 23596 -3722
rect 23596 -3774 23662 -3722
rect 23662 -3774 23666 -3722
rect 23590 -3778 23666 -3774
<< metal3 >>
rect 39998 24682 40008 24861
rect 40207 24682 40217 24861
rect 42480 24736 42490 24915
rect 42689 24736 42699 24915
rect 43627 24736 43637 24915
rect 43836 24736 43846 24915
rect 46511 24679 46521 24858
rect 46720 24679 46730 24858
rect 48993 24733 49003 24912
rect 49202 24733 49212 24912
rect 50140 24733 50150 24912
rect 50349 24733 50359 24912
rect 53045 24674 53055 24853
rect 53254 24674 53264 24853
rect 55527 24728 55537 24907
rect 55736 24728 55746 24907
rect 56674 24728 56684 24907
rect 56883 24728 56893 24907
rect 59603 24678 59613 24857
rect 59812 24678 59822 24857
rect 62085 24732 62095 24911
rect 62294 24732 62304 24911
rect 63232 24732 63242 24911
rect 63441 24732 63451 24911
rect 40292 23813 40471 23823
rect 40292 23605 40471 23614
rect 46805 23810 46984 23820
rect 46805 23602 46984 23611
rect 53339 23805 53518 23815
rect 53339 23597 53518 23606
rect 59897 23809 60076 23819
rect 59897 23601 60076 23610
rect 41826 23323 41835 23502
rect 42034 23323 42044 23502
rect 42968 23321 42977 23500
rect 43176 23321 43186 23500
rect 48339 23320 48348 23499
rect 48547 23320 48557 23499
rect 49481 23318 49490 23497
rect 49689 23318 49699 23497
rect 54873 23315 54882 23494
rect 55081 23315 55091 23494
rect 56015 23313 56024 23492
rect 56223 23313 56233 23492
rect 61431 23319 61440 23498
rect 61639 23319 61649 23498
rect 62573 23317 62582 23496
rect 62781 23317 62791 23496
rect 45151 23228 45534 23229
rect 32099 23181 39025 23204
rect 32099 23078 38849 23181
rect 38991 23078 39025 23181
rect 32099 23061 39025 23078
rect 4262 22268 4382 22273
rect 4262 22174 4272 22268
rect 4372 22174 4382 22268
rect 4262 22171 4382 22174
rect 7406 22268 7526 22273
rect 7406 22174 7416 22268
rect 7516 22174 7526 22268
rect 7406 22171 7526 22174
rect 10538 22264 10658 22269
rect 10538 22170 10548 22264
rect 10648 22170 10658 22264
rect 10538 22167 10658 22170
rect 13682 22264 13802 22269
rect 13682 22170 13692 22264
rect 13792 22170 13802 22264
rect 16884 22268 17004 22273
rect 16884 22174 16894 22268
rect 16994 22174 17004 22268
rect 16884 22171 17004 22174
rect 20028 22268 20148 22273
rect 20028 22174 20038 22268
rect 20138 22174 20148 22268
rect 20028 22171 20148 22174
rect 23160 22264 23280 22269
rect 13682 22167 13802 22170
rect 23160 22170 23170 22264
rect 23270 22170 23280 22264
rect 23160 22167 23280 22170
rect 26304 22264 26424 22269
rect 26304 22170 26314 22264
rect 26414 22170 26424 22264
rect 26304 22167 26424 22170
rect 27938 21446 28052 21449
rect 27936 21445 28138 21446
rect 27936 21444 29062 21445
rect 27936 21381 27948 21444
rect 28042 21381 29062 21444
rect 27938 21376 28052 21381
rect 1121 21254 2852 21256
rect 1072 21242 2852 21254
rect 1072 21152 2735 21242
rect 2840 21152 2852 21242
rect 1072 21138 2852 21152
rect 27717 21183 27814 21184
rect 1072 17992 1202 21138
rect 27717 21100 27727 21183
rect 27804 21100 27814 21183
rect 27717 21081 27814 21100
rect 5663 20925 5673 21034
rect 5773 20925 5783 21034
rect 27938 21013 28054 21018
rect 27938 20939 27948 21013
rect 28044 20998 28054 21013
rect 28044 20939 28917 20998
rect 27938 20934 28917 20939
rect 27944 20932 28917 20934
rect -1500 17991 -1397 17992
rect -527 17991 1202 17992
rect -1500 17878 1202 17991
rect 1264 20890 2858 20901
rect 1264 20814 2744 20890
rect 2837 20814 2858 20890
rect 1264 20800 2858 20814
rect 28520 20867 28774 20872
rect 28520 20811 28530 20867
rect 28598 20811 28774 20867
rect 28520 20806 28774 20811
rect -1500 17875 1096 17878
rect -1500 15335 -1397 17875
rect -1326 17727 -386 17728
rect 1264 17727 1399 20800
rect -1326 17611 1399 17727
rect 1476 20737 1583 20738
rect 1476 20736 1823 20737
rect 1476 20731 9220 20736
rect 1476 20672 9146 20731
rect 9210 20672 9220 20731
rect 1476 20667 9220 20672
rect 27936 20667 28635 20679
rect 1476 20666 2828 20667
rect 1476 20663 1823 20666
rect -1326 17610 1338 17611
rect -1325 15460 -1222 17610
rect 1476 17470 1583 20663
rect 27936 20610 27951 20667
rect 28043 20619 28635 20667
rect 28043 20610 28634 20619
rect 27936 20589 28634 20610
rect 27936 20588 28082 20589
rect 12280 20578 12356 20583
rect 28562 20582 28634 20589
rect 1645 20571 1713 20573
rect 12280 20572 12290 20578
rect 1785 20571 12290 20572
rect 1645 20524 12290 20571
rect -1151 17467 -461 17468
rect -120 17467 1583 17470
rect -1151 17353 1583 17467
rect -1151 17350 1095 17353
rect 1476 17350 1583 17353
rect 1644 20509 12290 20524
rect 12346 20509 12356 20578
rect 1644 20504 12356 20509
rect 27936 20523 28056 20527
rect 27936 20522 28486 20523
rect 1644 20503 2828 20504
rect -1151 17349 -461 17350
rect -1151 15611 -1048 17349
rect -527 17191 1096 17192
rect -971 17190 1096 17191
rect 1644 17190 1774 20503
rect 27936 20466 27946 20522
rect 28046 20466 28487 20522
rect 27936 20461 28487 20466
rect 27937 20460 28487 20461
rect 28415 20458 28487 20460
rect 15499 20427 15581 20432
rect 15499 20426 15509 20427
rect -971 17076 1774 17190
rect 1850 20359 15509 20426
rect 15571 20359 15581 20427
rect 1850 20358 15581 20359
rect 1850 20357 2828 20358
rect -971 17075 1668 17076
rect -971 15763 -868 17075
rect 45 17073 1668 17075
rect -785 16923 -424 16925
rect 1850 16923 1969 20357
rect 15499 20354 15581 20358
rect 27931 20397 28060 20400
rect 27931 20396 28348 20397
rect 27931 20395 28349 20396
rect 27931 20336 27941 20395
rect 28050 20336 28349 20395
rect 27931 20334 28349 20336
rect 27931 20331 28060 20334
rect -785 16808 1969 16923
rect 2043 20284 18701 20286
rect 2043 20279 18756 20284
rect 2043 20222 18687 20279
rect 18746 20222 18756 20279
rect 2043 20218 18756 20222
rect 2043 20217 2828 20218
rect 18677 20217 18756 20218
rect -785 16806 1958 16808
rect -785 16805 -424 16806
rect -785 15865 -682 16805
rect -616 16645 -439 16646
rect 2043 16645 2164 20217
rect 21803 20162 21882 20167
rect 3900 20153 4136 20158
rect 21803 20153 21813 20162
rect 3900 20151 21813 20153
rect 2227 20096 21813 20151
rect 21872 20096 21882 20162
rect 2227 20092 21882 20096
rect 2227 20084 4136 20092
rect 21803 20091 21882 20092
rect 27930 20156 28060 20159
rect 27930 20154 28213 20156
rect 27930 20094 27940 20154
rect 28050 20094 28213 20154
rect 27930 20091 28213 20094
rect 27930 20089 28060 20091
rect 2227 20083 2828 20084
rect -616 16528 2164 16645
rect 2228 16621 2365 20083
rect 4226 20024 4392 20032
rect 4226 19956 4274 20024
rect 4358 19956 4392 20024
rect 4226 19952 4392 19956
rect 7370 20024 7536 20032
rect 7370 19956 7418 20024
rect 7502 19956 7536 20024
rect 7370 19952 7536 19956
rect 10502 20020 10668 20028
rect 10502 19952 10550 20020
rect 10634 19952 10668 20020
rect 10502 19948 10668 19952
rect 13646 20020 13812 20028
rect 13646 19952 13694 20020
rect 13778 19952 13812 20020
rect 16848 20024 17014 20032
rect 16848 19956 16896 20024
rect 16980 19956 17014 20024
rect 16848 19952 17014 19956
rect 19992 20024 20158 20032
rect 19992 19956 20040 20024
rect 20124 19956 20158 20024
rect 19992 19952 20158 19956
rect 23124 20020 23290 20028
rect 23124 19952 23172 20020
rect 23256 19952 23290 20020
rect 13646 19948 13812 19952
rect 23124 19948 23290 19952
rect 26268 20020 26434 20028
rect 26268 19952 26316 20020
rect 26400 19952 26434 20020
rect 26268 19948 26434 19952
rect 27933 19933 28057 19938
rect 2516 19883 2683 19884
rect -616 16526 -439 16528
rect -616 16107 -513 16526
rect 2226 16507 2365 16621
rect 2457 19882 2683 19883
rect 24922 19882 25015 19887
rect 2457 19802 24932 19882
rect 2457 16538 2576 19802
rect 24922 19801 24932 19802
rect 25005 19801 25015 19882
rect 27933 19872 27943 19933
rect 28047 19872 28057 19933
rect 27933 19867 28057 19872
rect 24922 19796 25015 19801
rect 27936 19859 28054 19867
rect 4598 17048 4740 17062
rect 4598 16957 4622 17048
rect 4712 16957 4740 17048
rect 4598 16942 4740 16957
rect 5766 17048 5908 17062
rect 5766 16957 5790 17048
rect 5880 16957 5908 17048
rect 5766 16942 5908 16957
rect 6934 17048 7076 17062
rect 6934 16957 6958 17048
rect 7048 16957 7076 17048
rect 6934 16942 7076 16957
rect 8102 17048 8244 17062
rect 8102 16957 8126 17048
rect 8216 16957 8244 17048
rect 8102 16942 8244 16957
rect 9276 17046 9418 17060
rect 9276 16955 9300 17046
rect 9390 16955 9418 17046
rect 9276 16940 9418 16955
rect 10444 17046 10586 17060
rect 10444 16955 10468 17046
rect 10558 16955 10586 17046
rect 10444 16940 10586 16955
rect 11612 17046 11754 17060
rect 11612 16955 11636 17046
rect 11726 16955 11754 17046
rect 11612 16940 11754 16955
rect 12780 16940 12790 17060
rect 12912 16940 12922 17060
rect 14476 16843 14574 16861
rect 14476 16771 14494 16843
rect 14564 16771 14574 16843
rect 14476 16763 14574 16771
rect 15924 16843 16022 16861
rect 15924 16771 15942 16843
rect 16012 16771 16022 16843
rect 15924 16763 16022 16771
rect 17422 16841 17520 16859
rect 17422 16769 17440 16841
rect 17510 16769 17520 16841
rect 17422 16761 17520 16769
rect 18870 16841 18968 16859
rect 18870 16769 18888 16841
rect 18958 16769 18968 16841
rect 18870 16761 18968 16769
rect 20390 16843 20488 16861
rect 20390 16771 20408 16843
rect 20478 16771 20488 16843
rect 20390 16763 20488 16771
rect 21838 16843 21936 16861
rect 21838 16771 21856 16843
rect 21926 16771 21936 16843
rect 21838 16763 21936 16771
rect 23336 16841 23434 16859
rect 23336 16769 23354 16841
rect 23424 16769 23434 16841
rect 23336 16761 23434 16769
rect 24784 16841 24882 16859
rect 24784 16769 24802 16841
rect 24872 16769 24882 16841
rect 27790 16805 27868 16807
rect 24784 16761 24882 16769
rect 27318 16802 27868 16805
rect 27318 16759 27800 16802
rect 27314 16746 27800 16759
rect 27858 16746 27868 16802
rect 27314 16743 27868 16746
rect 2226 16416 2364 16507
rect -438 16300 2364 16416
rect -438 16299 2277 16300
rect -1500 5292 -1399 15335
rect -1323 5292 -1222 15460
rect -1150 5292 -1049 15611
rect -971 5292 -870 15763
rect -784 5292 -683 15865
rect -614 5292 -513 16107
rect -437 5292 -336 16299
rect 521 16090 2144 16091
rect 2457 16090 2579 16538
rect 25629 16186 25701 16191
rect 25620 16181 25711 16186
rect 25620 16122 25630 16181
rect 25701 16122 25711 16181
rect 25620 16117 25711 16122
rect -237 15974 2579 16090
rect 25336 16085 25425 16090
rect 25336 16021 25346 16085
rect 25415 16021 25425 16085
rect 25336 16016 25425 16021
rect -237 15973 2531 15974
rect -237 15859 -130 15973
rect 14820 15902 14925 15907
rect 15498 15903 16359 15905
rect 11472 15894 11557 15895
rect 14820 15894 14830 15902
rect -237 5292 -131 15859
rect 11472 15817 14830 15894
rect 5067 15620 5077 15731
rect 5187 15620 5197 15731
rect 6235 15620 6245 15731
rect 6355 15620 6365 15731
rect 7403 15620 7413 15731
rect 7523 15620 7533 15731
rect 8571 15620 8581 15731
rect 8691 15620 8701 15731
rect 9745 15618 9755 15729
rect 9865 15618 9875 15729
rect 10913 15618 10923 15729
rect 11033 15618 11043 15729
rect 11472 15385 11557 15817
rect 14820 15812 14830 15817
rect 14915 15812 14925 15902
rect 14820 15807 14925 15812
rect 15443 15897 16359 15903
rect 15443 15818 16288 15897
rect 16349 15818 16359 15897
rect 18992 15900 19058 15901
rect 18992 15895 19308 15900
rect 15443 15813 16359 15818
rect 16763 15893 17781 15894
rect 16763 15888 17858 15893
rect 16763 15820 17788 15888
rect 17848 15820 17858 15888
rect 16763 15816 17858 15820
rect 12081 15618 12091 15729
rect 12201 15618 12211 15729
rect 13249 15618 13259 15729
rect 13369 15618 13379 15729
rect 14574 15667 15010 15668
rect 15443 15667 15506 15813
rect 14254 15639 14356 15655
rect 14254 15571 14268 15639
rect 14342 15571 14356 15639
rect 14254 15557 14356 15571
rect 14574 15582 15506 15667
rect 15702 15639 15804 15655
rect 14574 15476 14635 15582
rect 15702 15571 15716 15639
rect 15790 15571 15804 15639
rect 15702 15557 15804 15571
rect 10968 15380 11557 15385
rect 13324 15416 14635 15476
rect 15010 15460 15076 15462
rect 16763 15460 16845 15816
rect 17778 15815 17858 15816
rect 18992 15820 19238 15895
rect 19298 15820 19308 15895
rect 18992 15816 19308 15820
rect 17200 15637 17302 15653
rect 17200 15569 17214 15637
rect 17288 15569 17302 15637
rect 17200 15555 17302 15569
rect 18648 15637 18750 15653
rect 18648 15569 18662 15637
rect 18736 15569 18750 15637
rect 18648 15555 18750 15569
rect 10968 15315 11556 15380
rect 1760 15130 1880 15135
rect 1760 15036 1770 15130
rect 1870 15036 1880 15130
rect 1760 15033 1880 15036
rect 4904 15130 5024 15135
rect 4904 15036 4914 15130
rect 5014 15036 5024 15130
rect 4904 15033 5024 15036
rect 8036 15126 8156 15131
rect 8036 15032 8046 15126
rect 8146 15032 8156 15126
rect 8036 15029 8156 15032
rect 1724 12886 1890 12894
rect 1724 12818 1772 12886
rect 1856 12818 1890 12886
rect 1724 12814 1890 12818
rect 4868 12886 5034 12894
rect 4868 12818 4916 12886
rect 5000 12818 5034 12886
rect 4868 12814 5034 12818
rect 8000 12882 8166 12890
rect 8000 12814 8048 12882
rect 8132 12814 8166 12882
rect 8000 12810 8166 12814
rect 1760 12396 1880 12401
rect 1760 12302 1770 12396
rect 1870 12302 1880 12396
rect 1760 12299 1880 12302
rect 4904 12396 5024 12401
rect 4904 12302 4914 12396
rect 5014 12302 5024 12396
rect 4904 12299 5024 12302
rect 8036 12392 8156 12397
rect 8036 12298 8046 12392
rect 8146 12298 8156 12392
rect 8036 12295 8156 12298
rect 1724 10152 1890 10160
rect 1724 10084 1772 10152
rect 1856 10084 1890 10152
rect 1724 10080 1890 10084
rect 4868 10152 5034 10160
rect 4868 10084 4916 10152
rect 5000 10084 5034 10152
rect 4868 10080 5034 10084
rect 8000 10148 8166 10156
rect 8000 10080 8048 10148
rect 8132 10080 8166 10148
rect 8000 10076 8166 10080
rect 1770 9664 1890 9669
rect 1770 9570 1780 9664
rect 1880 9570 1890 9664
rect 1770 9567 1890 9570
rect 4914 9664 5034 9669
rect 4914 9570 4924 9664
rect 5024 9570 5034 9664
rect 4914 9567 5034 9570
rect 8046 9660 8166 9665
rect 8046 9566 8056 9660
rect 8156 9566 8166 9660
rect 8046 9563 8166 9566
rect 1734 7420 1900 7428
rect 1734 7352 1782 7420
rect 1866 7352 1900 7420
rect 1734 7348 1900 7352
rect 4878 7420 5044 7428
rect 4878 7352 4926 7420
rect 5010 7352 5044 7420
rect 4878 7348 5044 7352
rect 8010 7416 8176 7424
rect 8010 7348 8058 7416
rect 8142 7348 8176 7416
rect 8010 7344 8176 7348
rect 3129 6775 3523 6781
rect 3129 6667 3265 6775
rect 3375 6667 3523 6775
rect 3129 6631 3523 6667
rect 3867 6775 4261 6781
rect 3867 6667 4003 6775
rect 4113 6667 4261 6775
rect 3867 6631 4261 6667
rect 4605 6775 4999 6781
rect 4605 6667 4741 6775
rect 4851 6667 4999 6775
rect 4605 6631 4999 6667
rect 5343 6775 5737 6781
rect 5343 6667 5479 6775
rect 5589 6667 5737 6775
rect 5343 6631 5737 6667
rect 6083 6775 6477 6781
rect 6083 6667 6219 6775
rect 6329 6667 6477 6775
rect 6083 6631 6477 6667
rect 6825 6775 7219 6781
rect 6825 6667 6961 6775
rect 7071 6667 7219 6775
rect 6825 6631 7219 6667
rect 7563 6775 7957 6781
rect 7563 6667 7699 6775
rect 7809 6667 7957 6775
rect 7563 6631 7957 6667
rect 8301 6777 8695 6783
rect 8301 6669 8437 6777
rect 8547 6669 8695 6777
rect 8301 6633 8695 6669
rect 9983 6708 10197 6712
rect 9983 6706 10051 6708
rect 9983 6636 10049 6706
rect 10127 6636 10197 6708
rect 9983 6634 10197 6636
rect 10039 6631 10137 6634
rect 10970 5910 11041 15315
rect 11180 15126 11300 15131
rect 11180 15032 11190 15126
rect 11290 15032 11300 15126
rect 11180 15029 11300 15032
rect 11144 12882 11310 12890
rect 11144 12814 11192 12882
rect 11276 12814 11310 12882
rect 11144 12810 11310 12814
rect 11180 12392 11300 12397
rect 11180 12298 11190 12392
rect 11290 12298 11300 12392
rect 11180 12295 11300 12298
rect 11144 10148 11310 10156
rect 11144 10080 11192 10148
rect 11276 10080 11310 10148
rect 11144 10076 11310 10080
rect 11190 9660 11310 9665
rect 11190 9566 11200 9660
rect 11300 9566 11310 9660
rect 11190 9563 11310 9566
rect 11154 7416 11320 7424
rect 11154 7348 11202 7416
rect 11286 7348 11320 7416
rect 11154 7344 11320 7348
rect 12051 6706 12265 6710
rect 12051 6704 12119 6706
rect 12051 6634 12117 6704
rect 12195 6634 12265 6706
rect 12051 6632 12265 6634
rect 12107 6629 12205 6632
rect 10837 5905 11041 5910
rect 8477 5885 8637 5887
rect 3305 5883 3465 5885
rect 3305 5783 3333 5883
rect 3435 5873 3465 5883
rect 4043 5883 4203 5885
rect 3435 5791 3467 5873
rect 3435 5783 3465 5791
rect 3305 5777 3465 5783
rect 4043 5783 4071 5883
rect 4173 5873 4203 5883
rect 4781 5883 4941 5885
rect 4173 5791 4205 5873
rect 4173 5783 4203 5791
rect 4043 5777 4203 5783
rect 4781 5783 4809 5883
rect 4911 5873 4941 5883
rect 5519 5883 5679 5885
rect 4911 5791 4943 5873
rect 4911 5783 4941 5791
rect 4781 5777 4941 5783
rect 5519 5783 5547 5883
rect 5649 5873 5679 5883
rect 6259 5883 6419 5885
rect 5649 5791 5681 5873
rect 5649 5783 5679 5791
rect 5519 5777 5679 5783
rect 6259 5783 6287 5883
rect 6389 5873 6419 5883
rect 7001 5883 7161 5885
rect 6389 5791 6421 5873
rect 6389 5783 6419 5791
rect 6259 5777 6419 5783
rect 7001 5783 7029 5883
rect 7131 5873 7161 5883
rect 7739 5883 7899 5885
rect 7131 5791 7163 5873
rect 7131 5783 7161 5791
rect 7001 5777 7161 5783
rect 7739 5783 7767 5883
rect 7869 5873 7899 5883
rect 7869 5791 7901 5873
rect 7869 5783 7899 5791
rect 7739 5777 7899 5783
rect 8477 5785 8505 5885
rect 8607 5875 8637 5885
rect 8607 5793 8639 5875
rect 10837 5825 10847 5905
rect 10930 5825 11041 5905
rect 13324 5899 13389 15416
rect 15006 15371 16845 15460
rect 14382 15130 14502 15135
rect 14382 15036 14392 15130
rect 14492 15036 14502 15130
rect 14382 15033 14502 15036
rect 14346 12886 14512 12894
rect 14346 12818 14394 12886
rect 14478 12818 14512 12886
rect 14346 12814 14512 12818
rect 14382 12396 14502 12401
rect 14382 12302 14392 12396
rect 14492 12302 14502 12396
rect 14382 12299 14502 12302
rect 14346 10152 14512 10160
rect 14346 10084 14394 10152
rect 14478 10084 14512 10152
rect 14346 10080 14512 10084
rect 14392 9664 14512 9669
rect 14392 9570 14402 9664
rect 14502 9570 14512 9664
rect 14392 9567 14512 9570
rect 14356 7420 14522 7428
rect 14356 7352 14404 7420
rect 14488 7352 14522 7420
rect 14356 7348 14522 7352
rect 14120 6708 14334 6712
rect 14120 6706 14188 6708
rect 14120 6636 14186 6706
rect 14264 6636 14334 6708
rect 14120 6634 14334 6636
rect 14176 6631 14274 6634
rect 15010 5901 15076 15371
rect 16763 15369 16845 15371
rect 17063 15451 17137 15452
rect 18992 15451 19058 15816
rect 19228 15815 19308 15816
rect 20740 15897 20827 15902
rect 20740 15819 20750 15897
rect 20817 15819 20827 15897
rect 20740 15682 20827 15819
rect 21214 15891 22279 15902
rect 21214 15817 22202 15891
rect 22266 15817 22279 15891
rect 21214 15811 22279 15817
rect 23292 15899 23778 15911
rect 23292 15812 23692 15899
rect 23768 15812 23778 15899
rect 20168 15639 20270 15655
rect 20168 15571 20182 15639
rect 20256 15571 20270 15639
rect 20168 15557 20270 15571
rect 20740 15481 20826 15682
rect 17063 15376 19058 15451
rect 16188 6706 16402 6710
rect 16188 6704 16256 6706
rect 16188 6634 16254 6704
rect 16332 6634 16402 6706
rect 16188 6632 16402 6634
rect 16244 6629 16342 6632
rect 17063 5901 17137 15376
rect 18992 15375 19058 15376
rect 19140 15409 20826 15481
rect 17526 15130 17646 15135
rect 17526 15036 17536 15130
rect 17636 15036 17646 15130
rect 17526 15033 17646 15036
rect 17490 12886 17656 12894
rect 17490 12818 17538 12886
rect 17622 12818 17656 12886
rect 17490 12814 17656 12818
rect 17526 12396 17646 12401
rect 17526 12302 17536 12396
rect 17636 12302 17646 12396
rect 17526 12299 17646 12302
rect 17490 10152 17656 10160
rect 17490 10084 17538 10152
rect 17622 10084 17656 10152
rect 17490 10080 17656 10084
rect 17536 9664 17656 9669
rect 17536 9570 17546 9664
rect 17646 9570 17656 9664
rect 17536 9567 17656 9570
rect 17500 7420 17666 7428
rect 17500 7352 17548 7420
rect 17632 7352 17666 7420
rect 17500 7348 17666 7352
rect 18257 6706 18471 6710
rect 18257 6704 18325 6706
rect 18257 6634 18323 6704
rect 18401 6634 18471 6706
rect 18257 6632 18471 6634
rect 18313 6629 18411 6632
rect 12969 5898 13389 5899
rect 10837 5812 11041 5825
rect 12917 5893 13389 5898
rect 12917 5829 12927 5893
rect 12994 5829 13389 5893
rect 12917 5825 13389 5829
rect 12917 5824 13104 5825
rect 13324 5824 13389 5825
rect 14990 5896 15076 5901
rect 14990 5828 15000 5896
rect 15065 5828 15076 5896
rect 14990 5823 15076 5828
rect 15010 5814 15076 5823
rect 17051 5896 17138 5901
rect 19140 5898 19207 15409
rect 20658 15126 20778 15131
rect 20658 15032 20668 15126
rect 20768 15032 20778 15126
rect 20658 15029 20778 15032
rect 20622 12882 20788 12890
rect 20622 12814 20670 12882
rect 20754 12814 20788 12882
rect 20622 12810 20788 12814
rect 20658 12392 20778 12397
rect 20658 12298 20668 12392
rect 20768 12298 20778 12392
rect 20658 12295 20778 12298
rect 20622 10148 20788 10156
rect 20622 10080 20670 10148
rect 20754 10080 20788 10148
rect 20622 10076 20788 10080
rect 20668 9660 20788 9665
rect 20668 9566 20678 9660
rect 20778 9566 20788 9660
rect 20668 9563 20788 9566
rect 20632 7416 20798 7424
rect 20632 7348 20680 7416
rect 20764 7348 20798 7416
rect 20632 7344 20798 7348
rect 20325 6704 20539 6708
rect 20325 6702 20393 6704
rect 20325 6632 20391 6702
rect 20469 6632 20539 6704
rect 20325 6630 20539 6632
rect 20381 6627 20479 6630
rect 17051 5827 17061 5896
rect 17128 5827 17138 5896
rect 17051 5822 17138 5827
rect 19122 5893 19207 5898
rect 21214 5897 21278 15811
rect 23292 15806 23778 15812
rect 21616 15639 21718 15655
rect 21616 15571 21630 15639
rect 21704 15571 21718 15639
rect 21616 15557 21718 15571
rect 23114 15637 23216 15653
rect 23114 15569 23128 15637
rect 23202 15569 23216 15637
rect 23114 15555 23216 15569
rect 22394 6706 22608 6710
rect 22394 6704 22462 6706
rect 22394 6634 22460 6704
rect 22538 6634 22608 6706
rect 22394 6632 22608 6634
rect 22450 6629 22548 6632
rect 23292 5915 23357 15806
rect 24562 15637 24664 15653
rect 24562 15569 24576 15637
rect 24650 15569 24664 15637
rect 24562 15555 24664 15569
rect 23802 15126 23922 15131
rect 23802 15032 23812 15126
rect 23912 15032 23922 15126
rect 23802 15029 23922 15032
rect 23766 12882 23932 12890
rect 23766 12814 23814 12882
rect 23898 12814 23932 12882
rect 23766 12810 23932 12814
rect 23802 12392 23922 12397
rect 23802 12298 23812 12392
rect 23912 12298 23922 12392
rect 23802 12295 23922 12298
rect 23766 10148 23932 10156
rect 23766 10080 23814 10148
rect 23898 10080 23932 10148
rect 23766 10076 23932 10080
rect 23812 9660 23932 9665
rect 23812 9566 23822 9660
rect 23922 9566 23932 9660
rect 23812 9563 23932 9566
rect 23776 7416 23942 7424
rect 23776 7348 23824 7416
rect 23908 7348 23942 7416
rect 23776 7344 23942 7348
rect 24462 6704 24676 6708
rect 24462 6702 24530 6704
rect 24462 6632 24528 6702
rect 24606 6632 24676 6704
rect 24462 6630 24676 6632
rect 24518 6627 24616 6630
rect 19122 5828 19132 5893
rect 19196 5828 19207 5893
rect 19122 5823 19207 5828
rect 17063 5810 17137 5822
rect 19140 5815 19207 5823
rect 21189 5892 21278 5897
rect 21189 5826 21199 5892
rect 21268 5826 21278 5892
rect 21189 5821 21278 5826
rect 21214 5814 21278 5821
rect 23254 5910 23357 5915
rect 23254 5824 23264 5910
rect 23339 5824 23357 5910
rect 23254 5819 23357 5824
rect 23292 5805 23357 5819
rect 8607 5785 8637 5793
rect 8477 5779 8637 5785
rect 25345 5749 25417 16016
rect 25629 15509 25701 16117
rect 27314 15509 27400 16743
rect 27790 16741 27868 16743
rect 25629 15464 27400 15509
rect 25629 15447 27395 15464
rect 25629 5891 25701 15447
rect 27936 7293 28007 19859
rect 28142 7293 28213 20091
rect 28278 7293 28349 20334
rect 28416 20253 28487 20458
rect 28416 20097 28488 20253
rect 28417 19935 28488 20097
rect 28417 19859 28489 19935
rect 28418 7293 28489 19859
rect 28563 7293 28634 20582
rect 28701 19902 28774 20806
rect 28703 7293 28774 19902
rect 28844 20755 28917 20932
rect 28988 20811 29062 21381
rect 28844 19841 28916 20755
rect 28988 19849 29060 20811
rect 28844 7293 28915 19841
rect 28988 7293 29059 19849
rect 31911 12443 32009 12445
rect 29689 12363 29767 12423
rect 31909 12415 32019 12443
rect 29689 12353 29770 12363
rect 29689 12277 29693 12353
rect 29689 12275 29695 12277
rect 29765 12275 29770 12353
rect 31909 12321 31915 12415
rect 32003 12321 32019 12415
rect 31909 12291 32019 12321
rect 29689 12265 29770 12275
rect 29689 12209 29767 12265
rect 32099 11533 32191 23061
rect 40012 23032 40022 23211
rect 40221 23032 40231 23211
rect 45149 23207 45534 23228
rect 51655 23213 52090 23232
rect 45149 23083 45281 23207
rect 45510 23083 45534 23207
rect 45149 23058 45534 23083
rect 45149 22985 45316 23058
rect 46525 23029 46535 23208
rect 46734 23029 46744 23208
rect 51655 23074 51840 23213
rect 51657 23073 51840 23074
rect 52058 23073 52090 23213
rect 58234 23215 58642 23235
rect 51657 23050 52090 23073
rect 41825 22689 41835 22868
rect 42034 22689 42044 22868
rect 43723 22689 43733 22868
rect 43932 22689 43942 22868
rect 40306 22163 40485 22173
rect 34395 22081 38951 22084
rect 34395 22076 38957 22081
rect 34395 21950 38809 22076
rect 38947 21950 38957 22076
rect 40306 21955 40485 21964
rect 34395 21945 38957 21950
rect 34395 21941 38951 21945
rect 32903 20321 33107 20323
rect 34395 20321 34499 21941
rect 39088 21870 39180 21871
rect 42486 21870 42590 21872
rect 39088 21866 42590 21870
rect 39088 21780 42498 21866
rect 42576 21780 42590 21866
rect 39088 21767 42590 21780
rect 39088 21707 39180 21767
rect 39067 21702 39202 21707
rect 39067 21605 39077 21702
rect 39192 21605 39202 21702
rect 39067 21600 39202 21605
rect 40007 21428 40017 21607
rect 40216 21428 40226 21607
rect 40301 20559 40480 20569
rect 40301 20351 40480 20360
rect 32903 20318 34499 20321
rect 32903 20157 32913 20318
rect 33097 20157 34499 20318
rect 41769 20280 41779 20459
rect 41978 20280 41988 20459
rect 43667 20280 43677 20459
rect 43876 20280 43886 20459
rect 32903 20153 34499 20157
rect 32903 20152 33107 20153
rect 45149 19998 45315 22985
rect 48338 22686 48348 22865
rect 48547 22686 48557 22865
rect 50236 22686 50246 22865
rect 50445 22686 50455 22865
rect 46819 22160 46998 22170
rect 46819 21952 46998 21961
rect 45601 21867 45693 21868
rect 48999 21867 49103 21869
rect 45601 21863 49103 21867
rect 45601 21777 49011 21863
rect 49089 21777 49103 21863
rect 45601 21764 49103 21777
rect 45601 21704 45693 21764
rect 45580 21699 45715 21704
rect 45580 21602 45590 21699
rect 45705 21602 45715 21699
rect 45580 21597 45715 21602
rect 46520 21425 46530 21604
rect 46729 21425 46739 21604
rect 46814 20556 46993 20566
rect 46814 20348 46993 20357
rect 48282 20277 48292 20456
rect 48491 20277 48501 20456
rect 50180 20277 50190 20456
rect 50389 20277 50399 20456
rect 31054 11526 32191 11533
rect 31054 11429 31064 11526
rect 31160 11429 32191 11526
rect 31054 11414 32191 11429
rect 32099 11413 32191 11414
rect 32263 19889 45315 19998
rect 31909 10375 32007 10377
rect 29687 10295 29765 10355
rect 31907 10347 32017 10375
rect 29687 10285 29768 10295
rect 29687 10209 29691 10285
rect 29687 10207 29693 10209
rect 29763 10207 29768 10285
rect 31907 10253 31913 10347
rect 32001 10253 32017 10347
rect 31907 10223 32017 10253
rect 29687 10197 29768 10207
rect 29687 10141 29765 10197
rect 32263 9461 32343 19889
rect 51657 19819 51818 23050
rect 53059 23024 53069 23203
rect 53268 23024 53278 23203
rect 58234 23070 58364 23215
rect 58616 23070 58642 23215
rect 58234 23057 58642 23070
rect 54872 22681 54882 22860
rect 55081 22681 55091 22860
rect 56770 22681 56780 22860
rect 56979 22681 56989 22860
rect 53353 22155 53532 22165
rect 53353 21947 53532 21956
rect 52135 21862 52227 21863
rect 55533 21862 55637 21864
rect 52135 21858 55637 21862
rect 52135 21772 55545 21858
rect 55623 21772 55637 21858
rect 52135 21759 55637 21772
rect 52135 21699 52227 21759
rect 52114 21694 52249 21699
rect 52114 21597 52124 21694
rect 52239 21597 52249 21694
rect 52114 21592 52249 21597
rect 53054 21420 53064 21599
rect 53263 21420 53273 21599
rect 53348 20551 53527 20561
rect 53348 20343 53527 20352
rect 54816 20272 54826 20451
rect 55025 20272 55035 20451
rect 56714 20272 56724 20451
rect 56923 20272 56933 20451
rect 31056 9456 32343 9461
rect 31056 9364 31066 9456
rect 31158 9364 32343 9456
rect 31056 9359 32343 9364
rect 32407 19705 51818 19819
rect 32407 19704 32486 19705
rect 31911 8306 32009 8308
rect 29689 8226 29767 8286
rect 31909 8278 32019 8306
rect 29689 8216 29770 8226
rect 29689 8140 29693 8216
rect 29689 8138 29695 8140
rect 29765 8138 29770 8216
rect 31909 8184 31915 8278
rect 32003 8184 32019 8278
rect 31909 8154 32019 8184
rect 29689 8128 29770 8138
rect 29689 8072 29767 8128
rect 32407 7392 32483 19704
rect 58234 19645 58404 23057
rect 59617 23028 59627 23207
rect 59826 23028 59836 23207
rect 61430 22685 61440 22864
rect 61639 22685 61649 22864
rect 63328 22685 63338 22864
rect 63537 22685 63547 22864
rect 59911 22159 60090 22169
rect 59911 21951 60090 21960
rect 58693 21866 58785 21867
rect 62091 21866 62195 21868
rect 58693 21862 62195 21866
rect 58693 21776 62103 21862
rect 62181 21776 62195 21862
rect 58693 21763 62195 21776
rect 58693 21703 58785 21763
rect 58672 21698 58807 21703
rect 58672 21601 58682 21698
rect 58797 21601 58807 21698
rect 58672 21596 58807 21601
rect 59612 21424 59622 21603
rect 59821 21424 59831 21603
rect 70236 20825 70338 20835
rect 70236 20725 70241 20825
rect 70335 20725 70338 20825
rect 70236 20715 70338 20725
rect 72477 20811 72557 20845
rect 72477 20727 72485 20811
rect 72553 20727 72557 20811
rect 72477 20679 72557 20727
rect 59906 20555 60085 20565
rect 59906 20347 60085 20356
rect 61374 20276 61384 20455
rect 61583 20276 61593 20455
rect 63272 20276 63282 20455
rect 63481 20276 63491 20455
rect 27935 7170 28007 7293
rect 27493 7158 28007 7170
rect 27493 7096 27506 7158
rect 27562 7096 28007 7158
rect 27493 7081 28007 7096
rect 28141 7091 28213 7293
rect 28277 7091 28349 7293
rect 28417 7091 28489 7293
rect 28141 6878 28212 7091
rect 27492 6867 28212 6878
rect 27492 6805 27506 6867
rect 27562 6805 28212 6867
rect 27492 6793 28212 6805
rect 27492 6792 28208 6793
rect 28277 6572 28348 7091
rect 27495 6561 28348 6572
rect 27495 6499 27507 6561
rect 27563 6499 28348 6561
rect 27495 6486 28348 6499
rect 28277 6485 28348 6486
rect 28417 6410 28488 7091
rect 27493 6400 28488 6410
rect 27493 6338 27506 6400
rect 27562 6338 28488 6400
rect 27493 6327 28488 6338
rect 28562 7089 28634 7293
rect 28702 7090 28774 7293
rect 28843 7090 28915 7293
rect 27493 6323 28482 6327
rect 28562 6262 28633 7089
rect 27491 6249 28633 6262
rect 27491 6187 27506 6249
rect 27562 6187 28633 6249
rect 27491 6175 28633 6187
rect 28702 6103 28773 7090
rect 27491 6088 28773 6103
rect 27491 6026 27506 6088
rect 27562 6026 28773 6088
rect 27491 6013 28773 6026
rect 28843 5914 28914 7090
rect 25614 5886 25701 5891
rect 25614 5829 25624 5886
rect 25690 5829 25701 5886
rect 25614 5824 25701 5829
rect 27493 5901 28914 5914
rect 27493 5839 27506 5901
rect 27562 5839 28914 5901
rect 27493 5826 28914 5839
rect 28843 5825 28914 5826
rect 28987 7085 29059 7293
rect 31062 7384 32483 7392
rect 31062 7298 31072 7384
rect 31157 7298 32483 7384
rect 31062 7280 32483 7298
rect 32407 7277 32483 7280
rect 32543 19535 58405 19645
rect 25629 5815 25701 5824
rect 25327 5704 25437 5749
rect 28987 5709 29058 7085
rect 31909 6238 32007 6240
rect 29687 6158 29765 6218
rect 31907 6210 32017 6238
rect 29687 6148 29768 6158
rect 29687 6072 29691 6148
rect 29687 6070 29693 6072
rect 29763 6070 29768 6148
rect 31907 6116 31913 6210
rect 32001 6116 32017 6210
rect 31907 6086 32017 6116
rect 29687 6060 29768 6070
rect 29687 6004 29765 6060
rect 25327 5627 25346 5704
rect 25417 5627 25437 5704
rect 25327 5607 25437 5627
rect 27493 5697 29058 5709
rect 27493 5635 27506 5697
rect 27562 5635 29058 5697
rect 27493 5620 29058 5635
rect 32543 5327 32622 19535
rect 33918 19534 34130 19535
rect 39574 19128 39584 19307
rect 39783 19128 39793 19307
rect 40721 19128 40731 19307
rect 40930 19128 40940 19307
rect 43203 19074 43213 19253
rect 43412 19074 43422 19253
rect 46132 19124 46142 19303
rect 46341 19124 46351 19303
rect 47279 19124 47289 19303
rect 47488 19124 47498 19303
rect 49761 19070 49771 19249
rect 49970 19070 49980 19249
rect 52666 19129 52676 19308
rect 52875 19129 52885 19308
rect 53813 19129 53823 19308
rect 54022 19129 54032 19308
rect 56295 19075 56305 19254
rect 56504 19075 56514 19254
rect 59179 19132 59189 19311
rect 59388 19132 59398 19311
rect 60326 19132 60336 19311
rect 60535 19132 60545 19311
rect 62808 19078 62818 19257
rect 63017 19078 63027 19257
rect 42949 18205 43128 18215
rect 42949 17997 43128 18006
rect 49507 18201 49686 18211
rect 49507 17993 49686 18002
rect 56041 18206 56220 18216
rect 56041 17998 56220 18007
rect 62554 18209 62733 18219
rect 62554 18001 62733 18010
rect 40234 17713 40244 17892
rect 40443 17713 40452 17892
rect 41376 17715 41386 17894
rect 41585 17715 41594 17894
rect 46792 17709 46802 17888
rect 47001 17709 47010 17888
rect 47934 17711 47944 17890
rect 48143 17711 48152 17890
rect 53326 17714 53336 17893
rect 53535 17714 53544 17893
rect 54468 17716 54478 17895
rect 54677 17716 54686 17895
rect 59839 17717 59849 17896
rect 60048 17717 60057 17896
rect 60981 17719 60991 17898
rect 61190 17719 61199 17898
rect 70236 17681 70338 17691
rect 64005 17637 64407 17659
rect 43189 17424 43199 17603
rect 43398 17424 43408 17603
rect 49747 17420 49757 17599
rect 49956 17420 49966 17599
rect 56281 17425 56291 17604
rect 56490 17425 56500 17604
rect 62794 17428 62804 17607
rect 63003 17428 63013 17607
rect 64005 17481 64020 17637
rect 64238 17481 64407 17637
rect 70236 17581 70241 17681
rect 70335 17581 70338 17681
rect 70236 17571 70338 17581
rect 72477 17667 72557 17701
rect 72477 17583 72485 17667
rect 72553 17583 72557 17667
rect 72477 17535 72557 17583
rect 64005 17456 64407 17481
rect 39478 17081 39488 17260
rect 39687 17081 39697 17260
rect 41376 17081 41386 17260
rect 41585 17081 41595 17260
rect 46036 17077 46046 17256
rect 46245 17077 46255 17256
rect 47934 17077 47944 17256
rect 48143 17077 48153 17256
rect 52570 17082 52580 17261
rect 52779 17082 52789 17261
rect 54468 17082 54478 17261
rect 54677 17082 54687 17261
rect 59083 17085 59093 17264
rect 59292 17085 59302 17264
rect 60981 17085 60991 17264
rect 61190 17085 61200 17264
rect 42935 16555 43114 16565
rect 42935 16347 43114 16356
rect 49493 16551 49672 16561
rect 49493 16343 49672 16352
rect 56027 16556 56206 16566
rect 56027 16348 56206 16357
rect 62540 16559 62719 16569
rect 62540 16351 62719 16360
rect 60435 16266 60539 16268
rect 63845 16266 63937 16267
rect 40830 16262 40934 16264
rect 53922 16263 54026 16265
rect 57332 16263 57424 16264
rect 44240 16262 44332 16263
rect 40830 16258 44332 16262
rect 40830 16172 40844 16258
rect 40922 16172 44332 16258
rect 40830 16159 44332 16172
rect 44240 16099 44332 16159
rect 47388 16258 47492 16260
rect 53922 16259 57424 16263
rect 50798 16258 50890 16259
rect 47388 16254 50890 16258
rect 47388 16168 47402 16254
rect 47480 16168 50890 16254
rect 47388 16155 50890 16168
rect 53922 16173 53936 16259
rect 54014 16173 57424 16259
rect 53922 16160 57424 16173
rect 60435 16262 63937 16266
rect 60435 16176 60449 16262
rect 60527 16176 63937 16262
rect 60435 16163 63937 16176
rect 44218 16094 44353 16099
rect 50798 16095 50890 16155
rect 57332 16100 57424 16160
rect 63845 16103 63937 16163
rect 57310 16095 57445 16100
rect 43194 15820 43204 15999
rect 43403 15820 43413 15999
rect 44218 15997 44228 16094
rect 44343 15997 44353 16094
rect 44218 15992 44353 15997
rect 50776 16090 50911 16095
rect 49752 15816 49762 15995
rect 49961 15816 49971 15995
rect 50776 15993 50786 16090
rect 50901 15993 50911 16090
rect 50776 15988 50911 15993
rect 56286 15821 56296 16000
rect 56495 15821 56505 16000
rect 57310 15998 57320 16095
rect 57435 15998 57445 16095
rect 63823 16098 63958 16103
rect 57310 15993 57445 15998
rect 62799 15824 62809 16003
rect 63008 15824 63018 16003
rect 63823 16001 63833 16098
rect 63948 16001 63958 16098
rect 63823 15996 63958 16001
rect 42940 14951 43119 14961
rect 39534 14672 39544 14851
rect 39743 14672 39753 14851
rect 41432 14672 41442 14851
rect 41641 14672 41651 14851
rect 49498 14947 49677 14957
rect 42940 14743 43119 14752
rect 46092 14668 46102 14847
rect 46301 14668 46311 14847
rect 47990 14668 48000 14847
rect 48199 14668 48209 14847
rect 56032 14952 56211 14962
rect 49498 14739 49677 14748
rect 52626 14673 52636 14852
rect 52835 14673 52845 14852
rect 54524 14673 54534 14852
rect 54733 14673 54743 14852
rect 62545 14955 62724 14965
rect 56032 14744 56211 14753
rect 59139 14676 59149 14855
rect 59348 14676 59358 14855
rect 61037 14676 61047 14855
rect 61246 14676 61256 14855
rect 62545 14747 62724 14756
rect 32738 13515 32870 13516
rect 64226 13515 64407 17456
rect 70232 14549 70334 14559
rect 70232 14449 70237 14549
rect 70331 14449 70334 14549
rect 70232 14439 70334 14449
rect 72473 14535 72553 14569
rect 72473 14451 72481 14535
rect 72549 14451 72553 14535
rect 72473 14403 72553 14451
rect 31056 5314 32622 5327
rect -1500 4136 -1396 5292
rect -1323 4262 -1219 5292
rect -1150 4389 -1046 5292
rect -971 4555 -867 5292
rect -784 4705 -680 5292
rect -614 4872 -510 5292
rect -437 5046 -333 5292
rect -237 5211 -128 5292
rect 31056 5229 31067 5314
rect 31156 5229 32622 5314
rect 31056 5218 32622 5229
rect 32683 13398 64407 13515
rect -1497 3566 -1396 4136
rect -1320 3711 -1219 4262
rect -1147 3903 -1046 4389
rect -968 3960 -867 4555
rect -781 4077 -680 4705
rect -611 4302 -510 4872
rect -434 4506 -333 5046
rect -234 4645 -128 5211
rect -234 4644 585 4645
rect -234 4640 589 4644
rect -234 4562 474 4640
rect 569 4562 589 4640
rect -234 4557 589 4562
rect 452 4555 589 4557
rect -437 4496 -332 4506
rect -437 4486 368 4496
rect -437 4397 248 4486
rect 358 4397 368 4486
rect -437 4390 368 4397
rect 199 4387 368 4390
rect 10065 4490 10217 4492
rect 14202 4490 14354 4492
rect 10065 4486 10219 4490
rect 10065 4398 10095 4486
rect 10189 4398 10219 4486
rect 10065 4392 10219 4398
rect 12133 4488 12285 4490
rect 12133 4484 12287 4488
rect 12133 4396 12163 4484
rect 12257 4396 12287 4484
rect 10065 4382 10217 4392
rect 12133 4390 12287 4396
rect 14202 4486 14356 4490
rect 14202 4398 14232 4486
rect 14326 4398 14356 4486
rect 14202 4392 14356 4398
rect 16270 4488 16422 4490
rect 18339 4488 18491 4490
rect 22476 4488 22628 4490
rect 16270 4484 16424 4488
rect 16270 4396 16300 4484
rect 16394 4396 16424 4484
rect 12133 4380 12285 4390
rect 14202 4382 14354 4392
rect 16270 4390 16424 4396
rect 18339 4484 18493 4488
rect 18339 4396 18369 4484
rect 18463 4396 18493 4484
rect 18339 4390 18493 4396
rect 20407 4486 20559 4488
rect 20407 4482 20561 4486
rect 20407 4394 20437 4482
rect 20531 4394 20561 4482
rect 16270 4380 16422 4390
rect 18339 4380 18491 4390
rect 20407 4388 20561 4394
rect 22476 4484 22630 4488
rect 22476 4396 22506 4484
rect 22600 4396 22630 4484
rect 22476 4390 22630 4396
rect 24544 4486 24696 4488
rect 24544 4482 24698 4486
rect 24544 4394 24574 4482
rect 24668 4394 24698 4482
rect 20407 4378 20559 4388
rect 22476 4380 22628 4390
rect 24544 4388 24698 4394
rect 24544 4378 24696 4388
rect -24 4302 105 4304
rect -611 4290 105 4302
rect -611 4257 -10 4290
rect -612 4206 -10 4257
rect 95 4206 105 4290
rect -612 4196 105 4206
rect -589 4194 105 4196
rect -24 4191 105 4194
rect 31909 4169 32007 4171
rect 29687 4089 29765 4149
rect 31907 4141 32017 4169
rect 29687 4079 29768 4089
rect -781 4017 15756 4077
rect -969 3956 -866 3960
rect -1147 3835 -1047 3903
rect -969 3896 12620 3956
rect 12527 3862 12620 3896
rect -1147 3776 9384 3835
rect -1129 3774 9384 3776
rect 9270 3747 9384 3774
rect -1321 3627 6208 3711
rect -1497 3480 3113 3566
rect -1483 3478 3113 3480
rect -1745 3282 232 3287
rect -1745 3217 -1727 3282
rect -1616 3277 232 3282
rect -1616 3217 135 3277
rect -1745 3214 135 3217
rect 214 3214 232 3277
rect -1745 3199 232 3214
rect -804 2875 54 2891
rect -804 2840 -22 2875
rect -804 2765 -791 2840
rect -801 2757 -791 2765
rect -659 2798 -22 2840
rect -659 2765 -640 2798
rect -52 2773 -22 2798
rect 43 2773 54 2875
rect -52 2765 54 2773
rect -659 2757 -649 2765
rect -801 2752 -649 2757
rect -572 2722 -402 2735
rect -572 2637 -545 2722
rect -428 2699 -402 2722
rect -428 2684 227 2699
rect -428 2637 130 2684
rect -572 2627 130 2637
rect 214 2627 227 2684
rect -572 2616 227 2627
rect -572 2614 -402 2616
rect 1486 2412 1606 2417
rect 1486 2318 1496 2412
rect 1596 2318 1606 2412
rect 1486 2315 1606 2318
rect 1476 168 1642 176
rect 1476 100 1510 168
rect 1594 100 1642 168
rect 1476 96 1642 100
rect 2990 -870 3110 3478
rect 4630 2412 4750 2417
rect 4630 2318 4640 2412
rect 4740 2318 4750 2412
rect 4630 2315 4750 2318
rect 4620 168 4786 176
rect 4620 100 4654 168
rect 4738 100 4786 168
rect 4620 96 4786 100
rect -173 -981 3110 -870
rect 3178 -867 3260 -864
rect 6095 -867 6205 3627
rect 7762 2416 7882 2421
rect 7762 2322 7772 2416
rect 7872 2322 7882 2416
rect 7762 2319 7882 2322
rect 7752 172 7918 180
rect 7752 104 7786 172
rect 7870 104 7918 172
rect 7752 100 7918 104
rect 3178 -981 6205 -867
rect 9270 -870 9385 3747
rect 10906 2416 11026 2421
rect 10906 2322 10916 2416
rect 11016 2322 11026 2416
rect 10906 2319 11026 2322
rect 10896 172 11062 180
rect 10896 104 10930 172
rect 11014 104 11062 172
rect 10896 100 11062 104
rect 12527 -862 12624 3862
rect 14108 2412 14228 2417
rect 14108 2318 14118 2412
rect 14218 2318 14228 2412
rect 14108 2315 14228 2318
rect 14098 168 14264 176
rect 14098 100 14132 168
rect 14216 100 14264 168
rect 14098 96 14264 100
rect 15635 -862 15756 4017
rect 29687 4003 29691 4079
rect 29687 4001 29693 4003
rect 29763 4001 29768 4079
rect 31907 4047 31913 4141
rect 32001 4047 32017 4141
rect 31907 4017 32017 4047
rect 29687 3991 29768 4001
rect 29687 3935 29765 3991
rect 32683 3255 32762 13398
rect 57714 13336 57833 13338
rect 31056 3245 32762 3255
rect 31056 3162 31070 3245
rect 31154 3162 32762 3245
rect 31056 3152 32762 3162
rect 32827 13244 57833 13336
rect 32646 3151 32724 3152
rect 17252 2412 17372 2417
rect 17252 2318 17262 2412
rect 17362 2318 17372 2412
rect 20384 2416 20504 2421
rect 20384 2322 20394 2416
rect 20494 2322 20504 2416
rect 20384 2319 20504 2322
rect 23528 2416 23648 2421
rect 23528 2322 23538 2416
rect 23638 2322 23648 2416
rect 23528 2319 23648 2322
rect 17252 2315 17372 2318
rect 31907 2101 32005 2103
rect 29685 2021 29763 2081
rect 31905 2073 32015 2101
rect 29685 2011 29766 2021
rect 29685 1935 29689 2011
rect 29685 1933 29691 1935
rect 29761 1933 29766 2011
rect 31905 1979 31911 2073
rect 31999 1979 32015 2073
rect 31905 1949 32015 1979
rect 29685 1923 29766 1933
rect 29685 1867 29763 1923
rect 32827 1188 32900 13244
rect 51189 13181 51309 13182
rect 31059 1178 32900 1188
rect 31059 1094 31069 1178
rect 31152 1094 32900 1178
rect 31059 1084 32900 1094
rect 32960 13081 51310 13181
rect 57714 13180 57833 13244
rect 17242 168 17408 176
rect 17242 100 17276 168
rect 17360 100 17408 168
rect 20374 172 20540 180
rect 20374 104 20408 172
rect 20492 104 20540 172
rect 20374 100 20540 104
rect 23518 172 23684 180
rect 23518 104 23552 172
rect 23636 104 23684 172
rect 23518 100 23684 104
rect 17242 96 17408 100
rect 31909 32 32007 34
rect 29687 -48 29765 12
rect 31907 4 32017 32
rect 29687 -58 29768 -48
rect 29687 -134 29691 -58
rect 29687 -136 29693 -134
rect 29763 -136 29768 -58
rect 31907 -90 31913 4
rect 32001 -90 32017 4
rect 31907 -120 32017 -90
rect 29687 -146 29768 -136
rect 29687 -202 29765 -146
rect -173 -982 3064 -981
rect -172 -2713 -63 -982
rect 1518 -1480 1638 -1475
rect 1518 -1574 1528 -1480
rect 1628 -1574 1638 -1480
rect 1518 -1577 1638 -1574
rect -175 -2718 -63 -2713
rect -175 -2796 -165 -2718
rect -77 -2796 -63 -2718
rect -175 -2801 -63 -2796
rect -172 -2810 -63 -2801
rect 3178 -2734 3260 -981
rect 6095 -988 6205 -981
rect 6309 -995 9391 -870
rect 4662 -1480 4782 -1475
rect 4662 -1574 4672 -1480
rect 4772 -1574 4782 -1480
rect 4662 -1577 4782 -1574
rect 6309 -2689 6413 -995
rect 9453 -1006 12624 -862
rect 12694 -1005 15756 -862
rect 32960 -882 33035 13081
rect 51189 13050 51309 13081
rect 57714 13078 57724 13180
rect 57823 13078 57833 13180
rect 57714 13069 57833 13078
rect 33096 12918 44744 13019
rect 51189 12965 51199 13050
rect 51299 12965 51309 13050
rect 51189 12954 51309 12965
rect 33096 12844 33172 12918
rect 31057 -891 33035 -882
rect 31057 -978 31067 -891
rect 31157 -978 33035 -891
rect 31057 -989 33035 -978
rect 12694 -1006 12841 -1005
rect 7794 -1476 7914 -1471
rect 7794 -1570 7804 -1476
rect 7904 -1570 7914 -1476
rect 7794 -1573 7914 -1570
rect 3178 -2798 3188 -2734
rect 3249 -2798 3260 -2734
rect 3178 -2808 3260 -2798
rect 6308 -2737 6413 -2689
rect 9453 -2732 9596 -1006
rect 10938 -1476 11058 -1471
rect 10938 -1570 10948 -1476
rect 11048 -1570 11058 -1476
rect 10938 -1573 11058 -1570
rect 12694 -2667 12797 -1006
rect 14140 -1480 14260 -1475
rect 14140 -1574 14150 -1480
rect 14250 -1574 14260 -1480
rect 14140 -1577 14260 -1574
rect 17284 -1480 17404 -1475
rect 17284 -1574 17294 -1480
rect 17394 -1574 17404 -1480
rect 20416 -1476 20536 -1471
rect 20416 -1570 20426 -1476
rect 20526 -1570 20536 -1476
rect 20416 -1573 20536 -1570
rect 23560 -1476 23680 -1471
rect 23560 -1570 23570 -1476
rect 23670 -1570 23680 -1476
rect 23560 -1573 23680 -1570
rect 17284 -1577 17404 -1574
rect 31907 -2036 32005 -2034
rect 29685 -2116 29763 -2056
rect 31905 -2064 32015 -2036
rect 29685 -2126 29766 -2116
rect 29685 -2202 29689 -2126
rect 29685 -2204 29691 -2202
rect 29761 -2204 29766 -2126
rect 31905 -2158 31911 -2064
rect 31999 -2158 32015 -2064
rect 31905 -2188 32015 -2158
rect 29685 -2214 29766 -2204
rect 29685 -2270 29763 -2214
rect 12693 -2725 12797 -2667
rect 6308 -2800 6318 -2737
rect 6401 -2800 6413 -2737
rect 6308 -2808 6413 -2800
rect 9452 -2737 9596 -2732
rect 9452 -2798 9462 -2737
rect 9581 -2798 9596 -2737
rect 9452 -2803 9596 -2798
rect 9453 -2805 9596 -2803
rect 12683 -2730 12797 -2725
rect 12683 -2811 12693 -2730
rect 12758 -2811 12797 -2730
rect 12683 -2816 12797 -2811
rect 12733 -2822 12797 -2816
rect 33097 -2943 33172 12844
rect 44612 12719 44744 12918
rect 68718 12895 71566 12898
rect 68717 12799 71566 12895
rect 44609 12714 44747 12719
rect 44609 12646 44619 12714
rect 44737 12646 44747 12714
rect 44609 12641 44747 12646
rect 44612 12636 44744 12641
rect 55098 12399 55196 12417
rect 41895 12379 41993 12397
rect 41895 12307 41905 12379
rect 41975 12307 41993 12379
rect 41895 12299 41993 12307
rect 48444 12378 48542 12396
rect 48444 12306 48454 12378
rect 48524 12306 48542 12378
rect 55098 12327 55108 12399
rect 55178 12327 55196 12399
rect 55098 12319 55196 12327
rect 48444 12298 48542 12306
rect 63751 12232 63849 12250
rect 63751 12160 63761 12232
rect 63831 12160 63849 12232
rect 63751 12152 63849 12160
rect 65981 12020 65991 12199
rect 66190 12020 66200 12199
rect 68717 12019 68844 12799
rect 71434 12798 71566 12799
rect 71483 12793 71566 12798
rect 71483 12788 71567 12793
rect 71483 12691 71494 12788
rect 71557 12691 71567 12788
rect 71483 12686 71567 12691
rect 71483 12682 71566 12686
rect 68717 11918 68845 12019
rect 67352 11824 67450 11842
rect 67352 11752 67362 11824
rect 67432 11752 67450 11824
rect 67352 11744 67450 11752
rect 55316 11195 55418 11211
rect 42113 11175 42215 11191
rect 42113 11107 42127 11175
rect 42201 11107 42215 11175
rect 42113 11093 42215 11107
rect 48662 11174 48764 11190
rect 48662 11106 48676 11174
rect 48750 11106 48764 11174
rect 55316 11127 55330 11195
rect 55404 11127 55418 11195
rect 55316 11113 55418 11127
rect 67967 11150 68326 11151
rect 67967 11142 68422 11150
rect 48662 11092 48764 11106
rect 67967 11060 67977 11142
rect 68115 11060 68422 11142
rect 67967 11051 68422 11060
rect 63969 11028 64071 11044
rect 63969 10960 63983 11028
rect 64057 10960 64071 11028
rect 34097 10951 34233 10956
rect 34097 10895 34107 10951
rect 34223 10895 34233 10951
rect 63969 10946 64071 10960
rect 34097 10890 34233 10895
rect 34104 1040 34227 10890
rect 68248 10721 68422 11051
rect 67447 10530 67457 10646
rect 67795 10530 67805 10646
rect 35231 10479 35329 10497
rect 35231 10407 35241 10479
rect 35311 10407 35329 10479
rect 35231 10399 35329 10407
rect 38194 10131 38204 10310
rect 38403 10131 38413 10310
rect 40676 10185 40686 10364
rect 40885 10185 40895 10364
rect 41823 10185 41833 10364
rect 42032 10185 42042 10364
rect 44743 10219 44753 10398
rect 44952 10219 44962 10398
rect 47225 10273 47235 10452
rect 47434 10273 47444 10452
rect 48372 10273 48382 10452
rect 48581 10273 48591 10452
rect 51397 10151 51407 10330
rect 51606 10151 51616 10330
rect 53879 10205 53889 10384
rect 54088 10205 54098 10384
rect 55026 10205 55036 10384
rect 55235 10205 55245 10384
rect 58022 10219 58032 10398
rect 58231 10219 58241 10398
rect 60504 10273 60514 10452
rect 60713 10273 60723 10452
rect 61651 10273 61661 10452
rect 61860 10273 61870 10452
rect 63746 9661 63844 9679
rect 63746 9589 63756 9661
rect 63826 9589 63844 9661
rect 65902 9659 65912 9854
rect 66178 9659 66188 9854
rect 63746 9581 63844 9589
rect 56277 9514 56534 9515
rect 56069 9509 56534 9514
rect 42935 9491 43100 9494
rect 42935 9489 43299 9491
rect 42935 9414 42945 9489
rect 43090 9414 43299 9489
rect 56069 9435 56079 9509
rect 56176 9435 56534 9509
rect 56069 9430 56534 9435
rect 42935 9409 43299 9414
rect 35449 9275 35551 9291
rect 35449 9207 35463 9275
rect 35537 9207 35551 9275
rect 35449 9193 35551 9207
rect 38488 9262 38667 9272
rect 38488 9054 38667 9063
rect 40022 8772 40031 8951
rect 40230 8772 40240 8951
rect 41164 8770 41173 8949
rect 41372 8770 41382 8949
rect 38208 8481 38218 8660
rect 38417 8481 38427 8660
rect 40021 8138 40031 8317
rect 40230 8138 40240 8317
rect 41919 8138 41929 8317
rect 42128 8138 42138 8317
rect 35223 7894 35321 7912
rect 35223 7822 35233 7894
rect 35303 7822 35321 7894
rect 35223 7814 35321 7822
rect 38502 7612 38681 7622
rect 38502 7404 38681 7413
rect 37284 7319 37376 7320
rect 40682 7319 40786 7321
rect 37284 7315 40786 7319
rect 37284 7229 40694 7315
rect 40772 7229 40786 7315
rect 37284 7216 40786 7229
rect 37284 7156 37376 7216
rect 37263 7151 37398 7156
rect 37263 7054 37273 7151
rect 37388 7054 37398 7151
rect 37263 7049 37398 7054
rect 38203 6877 38213 7056
rect 38412 6877 38422 7056
rect 35441 6690 35543 6706
rect 35441 6622 35455 6690
rect 35529 6622 35543 6690
rect 35441 6608 35543 6622
rect 38497 6008 38676 6018
rect 38497 5800 38676 5809
rect 39965 5729 39975 5908
rect 40174 5729 40184 5908
rect 41863 5729 41873 5908
rect 42072 5729 42082 5908
rect 36521 5006 36722 5007
rect 43155 5006 43299 9409
rect 45037 9350 45216 9360
rect 45037 9142 45216 9151
rect 51691 9282 51870 9292
rect 51691 9074 51870 9083
rect 46571 8860 46580 9039
rect 46779 8860 46789 9039
rect 47713 8858 47722 9037
rect 47921 8858 47931 9037
rect 53225 8792 53234 8971
rect 53433 8792 53443 8971
rect 54367 8790 54376 8969
rect 54575 8790 54585 8969
rect 44757 8569 44767 8748
rect 44966 8569 44976 8748
rect 51411 8501 51421 8680
rect 51620 8501 51630 8680
rect 46570 8226 46580 8405
rect 46779 8226 46789 8405
rect 48468 8226 48478 8405
rect 48677 8226 48687 8405
rect 53224 8158 53234 8337
rect 53433 8158 53443 8337
rect 55122 8158 55132 8337
rect 55331 8158 55341 8337
rect 45051 7700 45230 7710
rect 45051 7492 45230 7501
rect 51705 7632 51884 7642
rect 51705 7424 51884 7433
rect 43833 7407 43925 7408
rect 47231 7407 47335 7409
rect 43833 7403 47335 7407
rect 43833 7317 47243 7403
rect 47321 7317 47335 7403
rect 43833 7304 47335 7317
rect 50487 7339 50579 7340
rect 53885 7339 53989 7341
rect 50487 7335 53989 7339
rect 43833 7244 43925 7304
rect 50487 7249 53897 7335
rect 53975 7249 53989 7335
rect 43812 7239 43947 7244
rect 43812 7142 43822 7239
rect 43937 7142 43947 7239
rect 50487 7236 53989 7249
rect 50487 7176 50579 7236
rect 50466 7171 50601 7176
rect 43812 7137 43947 7142
rect 44752 6965 44762 7144
rect 44961 6965 44971 7144
rect 50466 7074 50476 7171
rect 50591 7074 50601 7171
rect 50466 7069 50601 7074
rect 51406 6897 51416 7076
rect 51615 6897 51625 7076
rect 45046 6096 45225 6106
rect 51700 6028 51879 6038
rect 45046 5888 45225 5897
rect 46514 5817 46524 5996
rect 46723 5817 46733 5996
rect 48412 5817 48422 5996
rect 48621 5817 48631 5996
rect 51700 5820 51879 5829
rect 53168 5749 53178 5928
rect 53377 5749 53387 5928
rect 55066 5749 55076 5928
rect 55275 5749 55285 5928
rect 56141 5520 56308 5530
rect 56141 5386 56152 5520
rect 56294 5386 56308 5520
rect 56141 5260 56308 5386
rect 44408 5259 56308 5260
rect 36521 4834 43299 5006
rect 43520 5088 56308 5259
rect 43520 5087 55419 5088
rect 35204 4616 35302 4634
rect 35204 4544 35214 4616
rect 35284 4544 35302 4616
rect 35204 4536 35302 4544
rect 35422 3412 35524 3428
rect 35422 3344 35436 3412
rect 35510 3344 35524 3412
rect 35422 3330 35524 3344
rect 35220 1856 35318 1874
rect 35220 1784 35230 1856
rect 35300 1784 35318 1856
rect 35220 1776 35318 1784
rect 36521 1761 36722 4834
rect 38186 4351 38196 4530
rect 38395 4351 38405 4530
rect 40668 4405 40678 4584
rect 40877 4405 40887 4584
rect 41815 4405 41825 4584
rect 42024 4405 42034 4584
rect 38480 3482 38659 3492
rect 38480 3274 38659 3283
rect 40014 2992 40023 3171
rect 40222 2992 40232 3171
rect 41156 2990 41165 3169
rect 41364 2990 41374 3169
rect 38200 2701 38210 2880
rect 38409 2701 38419 2880
rect 40013 2358 40023 2537
rect 40222 2358 40232 2537
rect 41911 2358 41921 2537
rect 42120 2358 42130 2537
rect 43520 1928 43706 5087
rect 56385 5006 56534 9430
rect 58316 9350 58495 9360
rect 58316 9142 58495 9151
rect 59850 8860 59859 9039
rect 60058 8860 60068 9039
rect 60992 8858 61001 9037
rect 61200 8858 61210 9037
rect 58036 8569 58046 8748
rect 58245 8569 58255 8748
rect 63964 8457 64066 8473
rect 59849 8226 59859 8405
rect 60058 8226 60068 8405
rect 61747 8226 61757 8405
rect 61956 8226 61966 8405
rect 63964 8389 63978 8457
rect 64052 8389 64066 8457
rect 63964 8375 64066 8389
rect 65983 7929 65993 8108
rect 66192 7929 66202 8108
rect 67354 7733 67452 7751
rect 58330 7700 58509 7710
rect 67354 7661 67364 7733
rect 67434 7661 67452 7733
rect 67354 7653 67452 7661
rect 58330 7492 58509 7501
rect 57112 7407 57204 7408
rect 60510 7407 60614 7409
rect 57112 7403 60614 7407
rect 57112 7317 60522 7403
rect 60600 7317 60614 7403
rect 57112 7304 60614 7317
rect 57112 7244 57204 7304
rect 57091 7239 57226 7244
rect 57091 7142 57101 7239
rect 57216 7142 57226 7239
rect 57091 7137 57226 7142
rect 58031 6965 58041 7144
rect 58240 6965 58250 7144
rect 56622 6824 56964 6829
rect 56622 6724 56632 6824
rect 56728 6724 56964 6824
rect 56622 6719 56964 6724
rect 56623 6716 56964 6719
rect 49925 4819 56534 5006
rect 56814 5010 56964 6716
rect 63746 6628 63844 6646
rect 63746 6556 63756 6628
rect 63826 6556 63844 6628
rect 63746 6548 63844 6556
rect 67449 6439 67459 6555
rect 67797 6439 67807 6555
rect 58325 6096 58504 6106
rect 58325 5888 58504 5897
rect 59793 5817 59803 5996
rect 60002 5817 60012 5996
rect 61691 5817 61701 5996
rect 61900 5817 61910 5996
rect 65904 5568 65914 5763
rect 66180 5568 66190 5763
rect 57250 5520 57417 5530
rect 57250 5386 57261 5520
rect 57403 5386 57417 5520
rect 57250 5258 57417 5386
rect 63964 5424 64066 5440
rect 63964 5356 63978 5424
rect 64052 5356 64066 5424
rect 63964 5342 64066 5356
rect 68248 5258 68421 10721
rect 57250 5172 68421 5258
rect 57251 5088 68421 5172
rect 68248 5085 68421 5088
rect 64963 5010 65082 5012
rect 44737 4349 44747 4528
rect 44946 4349 44956 4528
rect 47219 4403 47229 4582
rect 47428 4403 47438 4582
rect 48366 4403 48376 4582
rect 48575 4403 48585 4582
rect 45031 3480 45210 3490
rect 45031 3272 45210 3281
rect 46565 2990 46574 3169
rect 46773 2990 46783 3169
rect 47707 2988 47716 3167
rect 47915 2988 47925 3167
rect 44751 2699 44761 2878
rect 44960 2699 44970 2878
rect 46564 2356 46574 2535
rect 46773 2356 46783 2535
rect 48462 2356 48472 2535
rect 48671 2356 48681 2535
rect 38494 1832 38673 1842
rect 36520 1756 37132 1761
rect 36520 1619 36885 1756
rect 37119 1619 37132 1756
rect 43519 1803 43707 1928
rect 45045 1830 45224 1840
rect 43509 1749 43753 1803
rect 43509 1708 43520 1749
rect 38494 1624 38673 1633
rect 36520 1615 37132 1619
rect 36875 1614 37129 1615
rect 43510 1613 43520 1708
rect 43743 1613 43753 1749
rect 49925 1765 50126 4819
rect 56814 4815 65082 5010
rect 63817 4708 63915 4726
rect 63817 4636 63827 4708
rect 63897 4636 63915 4708
rect 63817 4628 63915 4636
rect 51392 4350 51402 4529
rect 51601 4350 51611 4529
rect 53874 4404 53884 4583
rect 54083 4404 54093 4583
rect 55021 4404 55031 4583
rect 55230 4404 55240 4583
rect 58014 4351 58024 4530
rect 58223 4351 58233 4530
rect 60496 4405 60506 4584
rect 60705 4405 60715 4584
rect 61643 4405 61653 4584
rect 61852 4405 61862 4584
rect 62996 3695 63664 3697
rect 62995 3692 63664 3695
rect 62995 3591 63568 3692
rect 63654 3591 63664 3692
rect 62995 3586 63664 3591
rect 64963 3668 65082 4815
rect 65983 4434 65993 4613
rect 66192 4434 66202 4613
rect 67354 4238 67452 4256
rect 67354 4166 67364 4238
rect 67434 4166 67452 4238
rect 67354 4158 67452 4166
rect 64963 3663 65319 3668
rect 64963 3586 65216 3663
rect 65309 3586 65319 3663
rect 51686 3481 51865 3491
rect 51686 3273 51865 3282
rect 58308 3482 58487 3492
rect 58308 3274 58487 3283
rect 53220 2991 53229 3170
rect 53428 2991 53438 3170
rect 54362 2989 54371 3168
rect 54570 2989 54580 3168
rect 59842 2992 59851 3171
rect 60050 2992 60060 3171
rect 60984 2990 60993 3169
rect 61192 2990 61202 3169
rect 51406 2700 51416 2879
rect 51615 2700 51625 2879
rect 58028 2701 58038 2880
rect 58237 2701 58247 2880
rect 53219 2357 53229 2536
rect 53428 2357 53438 2536
rect 55117 2357 55127 2536
rect 55326 2357 55336 2536
rect 59841 2358 59851 2537
rect 60050 2358 60060 2537
rect 61739 2358 61749 2537
rect 61948 2358 61958 2537
rect 51700 1831 51879 1841
rect 49925 1734 50373 1765
rect 49925 1712 50201 1734
rect 45045 1622 45224 1631
rect 49926 1622 50201 1712
rect 50345 1622 50373 1734
rect 51700 1623 51879 1632
rect 58322 1832 58501 1842
rect 58322 1624 58501 1633
rect 43510 1608 43753 1613
rect 49926 1604 50373 1622
rect 37276 1539 37368 1540
rect 40674 1539 40778 1541
rect 37276 1535 40778 1539
rect 37276 1449 40686 1535
rect 40764 1449 40778 1535
rect 37276 1436 40778 1449
rect 43827 1537 43919 1538
rect 47225 1537 47329 1539
rect 43827 1533 47329 1537
rect 43827 1447 47237 1533
rect 47315 1447 47329 1533
rect 37276 1376 37368 1436
rect 43827 1434 47329 1447
rect 50482 1538 50574 1539
rect 53880 1538 53984 1540
rect 50482 1534 53984 1538
rect 50482 1448 53892 1534
rect 53970 1448 53984 1534
rect 50482 1435 53984 1448
rect 57104 1539 57196 1540
rect 60502 1539 60606 1541
rect 57104 1535 60606 1539
rect 57104 1449 60514 1535
rect 60592 1449 60606 1535
rect 57104 1436 60606 1449
rect 37255 1371 37390 1376
rect 43827 1374 43919 1434
rect 50482 1375 50574 1435
rect 57104 1376 57196 1436
rect 37255 1274 37265 1371
rect 37380 1274 37390 1371
rect 43806 1369 43941 1374
rect 37255 1269 37390 1274
rect 38195 1097 38205 1276
rect 38404 1097 38414 1276
rect 43806 1272 43816 1369
rect 43931 1272 43941 1369
rect 50461 1370 50596 1375
rect 43806 1267 43941 1272
rect 44746 1095 44756 1274
rect 44955 1095 44965 1274
rect 50461 1273 50471 1370
rect 50586 1273 50596 1370
rect 57083 1371 57218 1376
rect 50461 1268 50596 1273
rect 51401 1096 51411 1275
rect 51610 1096 51620 1275
rect 57083 1274 57093 1371
rect 57208 1274 57218 1371
rect 57083 1269 57218 1274
rect 58023 1097 58033 1276
rect 58232 1097 58242 1276
rect 34104 961 34114 1040
rect 34217 961 34227 1040
rect 34104 956 34227 961
rect 62774 1023 62934 1029
rect 62774 927 62787 1023
rect 62919 927 62934 1023
rect 35438 652 35540 668
rect 35438 584 35452 652
rect 35526 584 35540 652
rect 35438 570 35540 584
rect 38489 228 38668 238
rect 45040 226 45219 236
rect 38489 20 38668 29
rect 39957 -51 39967 128
rect 40166 -51 40176 128
rect 41855 -51 41865 128
rect 42064 -51 42074 128
rect 51695 227 51874 237
rect 45040 18 45219 27
rect 46508 -53 46518 126
rect 46717 -53 46727 126
rect 48406 -53 48416 126
rect 48615 -53 48625 126
rect 58317 228 58496 238
rect 51695 19 51874 28
rect 53163 -52 53173 127
rect 53372 -52 53382 127
rect 55061 -52 55071 127
rect 55270 -52 55280 127
rect 58317 20 58496 29
rect 59785 -51 59795 128
rect 59994 -51 60004 128
rect 61683 -51 61693 128
rect 61892 -51 61902 128
rect 42148 -713 42250 -699
rect 42148 -781 42162 -713
rect 42236 -781 42250 -713
rect 42148 -797 42250 -781
rect 48702 -708 48804 -694
rect 48702 -776 48716 -708
rect 48790 -776 48804 -708
rect 48702 -792 48804 -776
rect 55351 -720 55453 -706
rect 55351 -788 55365 -720
rect 55439 -788 55453 -720
rect 55351 -804 55453 -788
rect 41930 -1913 42028 -1905
rect 41930 -1985 41940 -1913
rect 42010 -1985 42028 -1913
rect 41930 -2003 42028 -1985
rect 48484 -1908 48582 -1900
rect 48484 -1980 48494 -1908
rect 48564 -1980 48582 -1908
rect 48484 -1998 48582 -1980
rect 55133 -1920 55231 -1912
rect 55133 -1992 55143 -1920
rect 55213 -1992 55231 -1920
rect 55133 -2010 55231 -1992
rect 62774 -2579 62934 927
rect 62995 919 63095 3586
rect 64963 3581 65319 3586
rect 64963 3579 65282 3581
rect 63330 3518 63435 3523
rect 63330 3458 63340 3518
rect 63425 3458 63435 3518
rect 63330 3421 63435 3458
rect 64035 3504 64137 3520
rect 64035 3436 64049 3504
rect 64123 3436 64137 3504
rect 64035 3422 64137 3436
rect 62995 -1705 63096 919
rect 63164 703 63266 712
rect 63160 698 63266 703
rect 63160 608 63170 698
rect 63254 608 63266 698
rect 63160 603 63266 608
rect 62995 -1795 63001 -1705
rect 63083 -1795 63096 -1705
rect 62995 -1805 63096 -1795
rect 63164 601 63266 603
rect 63164 -2016 63264 601
rect 63158 -2021 63264 -2016
rect 63158 -2111 63168 -2021
rect 63252 -2111 63264 -2021
rect 63158 -2116 63264 -2111
rect 63164 -2118 63264 -2116
rect 63341 -2365 63418 3421
rect 67449 2944 67459 3060
rect 67797 2944 67807 3060
rect 65904 2073 65914 2268
rect 66180 2073 66190 2268
rect 63814 1638 63912 1656
rect 63814 1566 63824 1638
rect 63894 1566 63912 1638
rect 63814 1558 63912 1566
rect 63594 551 63680 556
rect 63594 487 63604 551
rect 63670 487 63680 551
rect 63594 -947 63680 487
rect 64032 434 64134 450
rect 64032 366 64046 434
rect 64120 366 64134 434
rect 64032 352 64134 366
rect 65983 86 65993 265
rect 66192 86 66202 265
rect 67354 -110 67452 -92
rect 67354 -182 67364 -110
rect 67434 -182 67452 -110
rect 67354 -190 67452 -182
rect 63579 -962 63680 -947
rect 63579 -1052 63584 -962
rect 63668 -1052 63680 -962
rect 63579 -1061 63680 -1052
rect 68719 -1053 68845 11918
rect 70232 11405 70334 11415
rect 70232 11305 70237 11405
rect 70331 11305 70334 11405
rect 70232 11295 70334 11305
rect 72473 11391 72553 11425
rect 72473 11307 72481 11391
rect 72549 11307 72553 11391
rect 72473 11259 72553 11307
rect 70236 8203 70338 8213
rect 70236 8103 70241 8203
rect 70335 8103 70338 8203
rect 70236 8093 70338 8103
rect 72477 8189 72557 8223
rect 72477 8105 72485 8189
rect 72553 8105 72557 8189
rect 72477 8057 72557 8105
rect 68719 -1126 68739 -1053
rect 68826 -1126 68845 -1053
rect 68719 -1145 68845 -1126
rect 69014 6458 71576 6575
rect 63821 -1207 63919 -1189
rect 63821 -1279 63831 -1207
rect 63901 -1279 63919 -1207
rect 63821 -1287 63919 -1279
rect 67449 -1404 67459 -1288
rect 67797 -1404 67807 -1288
rect 65904 -2275 65914 -2080
rect 66180 -2275 66190 -2080
rect 63341 -2370 63552 -2365
rect 63341 -2445 63481 -2370
rect 63542 -2445 63552 -2370
rect 63341 -2450 63552 -2445
rect 64039 -2411 64141 -2395
rect 64039 -2479 64053 -2411
rect 64127 -2479 64141 -2411
rect 64039 -2493 64141 -2479
rect 62773 -2710 62934 -2579
rect 69014 -2710 69118 6458
rect 71484 6441 71576 6458
rect 71484 6373 71495 6441
rect 71485 6368 71495 6373
rect 71565 6373 71576 6441
rect 71565 6368 71575 6373
rect 71485 6363 71575 6368
rect 70236 5059 70338 5069
rect 70236 4959 70241 5059
rect 70335 4959 70338 5059
rect 70236 4949 70338 4959
rect 72477 5045 72557 5079
rect 72477 4961 72485 5045
rect 72553 4961 72557 5045
rect 72477 4913 72557 4961
rect 70232 1927 70334 1937
rect 70232 1827 70237 1927
rect 70331 1827 70334 1927
rect 70232 1817 70334 1827
rect 72473 1913 72553 1947
rect 72473 1829 72481 1913
rect 72549 1829 72553 1913
rect 72473 1781 72553 1829
rect 70232 -1217 70334 -1207
rect 70232 -1317 70237 -1217
rect 70331 -1317 70334 -1217
rect 70232 -1327 70334 -1317
rect 72473 -1231 72553 -1197
rect 72473 -1315 72481 -1231
rect 72549 -1315 72553 -1231
rect 72473 -1363 72553 -1315
rect 62773 -2814 69118 -2710
rect 32438 -2945 33172 -2943
rect 31058 -2959 33172 -2945
rect 31058 -3044 31068 -2959
rect 31154 -3044 33172 -2959
rect 31058 -3059 33172 -3044
rect 32294 -3060 33172 -3059
rect 1508 -3724 1674 -3716
rect 1508 -3792 1542 -3724
rect 1626 -3792 1674 -3724
rect 1508 -3796 1674 -3792
rect 4652 -3724 4818 -3716
rect 4652 -3792 4686 -3724
rect 4770 -3792 4818 -3724
rect 7784 -3720 7950 -3712
rect 7784 -3788 7818 -3720
rect 7902 -3788 7950 -3720
rect 7784 -3792 7950 -3788
rect 10928 -3720 11094 -3712
rect 10928 -3788 10962 -3720
rect 11046 -3788 11094 -3720
rect 10928 -3792 11094 -3788
rect 14130 -3724 14296 -3716
rect 14130 -3792 14164 -3724
rect 14248 -3792 14296 -3724
rect 4652 -3796 4818 -3792
rect 14130 -3796 14296 -3792
rect 17274 -3724 17440 -3716
rect 17274 -3792 17308 -3724
rect 17392 -3792 17440 -3724
rect 20406 -3720 20572 -3712
rect 20406 -3788 20440 -3720
rect 20524 -3788 20572 -3720
rect 20406 -3792 20572 -3788
rect 23550 -3720 23716 -3712
rect 23550 -3788 23584 -3720
rect 23668 -3788 23716 -3720
rect 23550 -3792 23716 -3788
rect 17274 -3796 17440 -3792
<< via3 >>
rect 40008 24830 40207 24861
rect 40008 24701 40030 24830
rect 40030 24701 40183 24830
rect 40183 24701 40207 24830
rect 40008 24682 40207 24701
rect 42490 24884 42689 24915
rect 42490 24755 42512 24884
rect 42512 24755 42665 24884
rect 42665 24755 42689 24884
rect 42490 24736 42689 24755
rect 43637 24884 43836 24915
rect 43637 24755 43659 24884
rect 43659 24755 43812 24884
rect 43812 24755 43836 24884
rect 43637 24736 43836 24755
rect 46521 24827 46720 24858
rect 46521 24698 46543 24827
rect 46543 24698 46696 24827
rect 46696 24698 46720 24827
rect 46521 24679 46720 24698
rect 49003 24881 49202 24912
rect 49003 24752 49025 24881
rect 49025 24752 49178 24881
rect 49178 24752 49202 24881
rect 49003 24733 49202 24752
rect 50150 24881 50349 24912
rect 50150 24752 50172 24881
rect 50172 24752 50325 24881
rect 50325 24752 50349 24881
rect 50150 24733 50349 24752
rect 53055 24822 53254 24853
rect 53055 24693 53077 24822
rect 53077 24693 53230 24822
rect 53230 24693 53254 24822
rect 53055 24674 53254 24693
rect 55537 24876 55736 24907
rect 55537 24747 55559 24876
rect 55559 24747 55712 24876
rect 55712 24747 55736 24876
rect 55537 24728 55736 24747
rect 56684 24876 56883 24907
rect 56684 24747 56706 24876
rect 56706 24747 56859 24876
rect 56859 24747 56883 24876
rect 56684 24728 56883 24747
rect 59613 24826 59812 24857
rect 59613 24697 59635 24826
rect 59635 24697 59788 24826
rect 59788 24697 59812 24826
rect 59613 24678 59812 24697
rect 62095 24880 62294 24911
rect 62095 24751 62117 24880
rect 62117 24751 62270 24880
rect 62270 24751 62294 24880
rect 62095 24732 62294 24751
rect 63242 24880 63441 24911
rect 63242 24751 63264 24880
rect 63264 24751 63417 24880
rect 63417 24751 63441 24880
rect 63242 24732 63441 24751
rect 40292 23791 40471 23813
rect 40292 23638 40311 23791
rect 40311 23638 40440 23791
rect 40440 23638 40471 23791
rect 40292 23614 40471 23638
rect 46805 23788 46984 23810
rect 46805 23635 46824 23788
rect 46824 23635 46953 23788
rect 46953 23635 46984 23788
rect 46805 23611 46984 23635
rect 53339 23783 53518 23805
rect 53339 23630 53358 23783
rect 53358 23630 53487 23783
rect 53487 23630 53518 23783
rect 53339 23606 53518 23630
rect 59897 23787 60076 23809
rect 59897 23634 59916 23787
rect 59916 23634 60045 23787
rect 60045 23634 60076 23787
rect 59897 23610 60076 23634
rect 41835 23483 42034 23502
rect 41835 23354 41859 23483
rect 41859 23354 42012 23483
rect 42012 23354 42034 23483
rect 41835 23323 42034 23354
rect 42977 23481 43176 23500
rect 42977 23352 43001 23481
rect 43001 23352 43154 23481
rect 43154 23352 43176 23481
rect 42977 23321 43176 23352
rect 48348 23480 48547 23499
rect 48348 23351 48372 23480
rect 48372 23351 48525 23480
rect 48525 23351 48547 23480
rect 48348 23320 48547 23351
rect 49490 23478 49689 23497
rect 49490 23349 49514 23478
rect 49514 23349 49667 23478
rect 49667 23349 49689 23478
rect 49490 23318 49689 23349
rect 54882 23475 55081 23494
rect 54882 23346 54906 23475
rect 54906 23346 55059 23475
rect 55059 23346 55081 23475
rect 54882 23315 55081 23346
rect 56024 23473 56223 23492
rect 56024 23344 56048 23473
rect 56048 23344 56201 23473
rect 56201 23344 56223 23473
rect 56024 23313 56223 23344
rect 61440 23479 61639 23498
rect 61440 23350 61464 23479
rect 61464 23350 61617 23479
rect 61617 23350 61639 23479
rect 61440 23319 61639 23350
rect 62582 23477 62781 23496
rect 62582 23348 62606 23477
rect 62606 23348 62759 23477
rect 62759 23348 62781 23477
rect 62582 23317 62781 23348
rect 4272 22176 4372 22266
rect 4272 22174 4372 22176
rect 7416 22176 7516 22266
rect 7416 22174 7516 22176
rect 10548 22172 10648 22262
rect 10548 22170 10648 22172
rect 13692 22172 13792 22262
rect 13692 22170 13792 22172
rect 16894 22176 16994 22266
rect 16894 22174 16994 22176
rect 20038 22176 20138 22266
rect 20038 22174 20138 22176
rect 23170 22172 23270 22262
rect 23170 22170 23270 22172
rect 26314 22172 26414 22262
rect 26314 22170 26414 22172
rect 27727 21169 27804 21183
rect 27727 21113 27738 21169
rect 27738 21113 27794 21169
rect 27794 21113 27804 21169
rect 27727 21100 27804 21113
rect 5673 21024 5773 21034
rect 5673 20935 5683 21024
rect 5683 20935 5762 21024
rect 5762 20935 5773 21024
rect 5673 20925 5773 20935
rect 4274 19966 4276 20024
rect 4276 19966 4352 20024
rect 4352 19966 4358 20024
rect 4274 19956 4358 19966
rect 7418 19966 7420 20024
rect 7420 19966 7496 20024
rect 7496 19966 7502 20024
rect 7418 19956 7502 19966
rect 10550 19962 10552 20020
rect 10552 19962 10628 20020
rect 10628 19962 10634 20020
rect 10550 19952 10634 19962
rect 13694 19962 13696 20020
rect 13696 19962 13772 20020
rect 13772 19962 13778 20020
rect 13694 19952 13778 19962
rect 16896 19966 16898 20024
rect 16898 19966 16974 20024
rect 16974 19966 16980 20024
rect 16896 19956 16980 19966
rect 20040 19966 20042 20024
rect 20042 19966 20118 20024
rect 20118 19966 20124 20024
rect 20040 19956 20124 19966
rect 23172 19962 23174 20020
rect 23174 19962 23250 20020
rect 23250 19962 23256 20020
rect 23172 19952 23256 19962
rect 26316 19962 26318 20020
rect 26318 19962 26394 20020
rect 26394 19962 26400 20020
rect 26316 19952 26400 19962
rect 4632 16970 4696 17034
rect 5800 16970 5864 17034
rect 6968 16968 7032 17032
rect 8136 16970 8200 17034
rect 9308 16970 9372 17034
rect 10478 16968 10542 17032
rect 11646 16968 11710 17032
rect 12790 17046 12912 17060
rect 12790 16955 12804 17046
rect 12804 16955 12894 17046
rect 12894 16955 12912 17046
rect 12790 16940 12912 16955
rect 14494 16839 14564 16843
rect 14494 16777 14498 16839
rect 14498 16777 14558 16839
rect 14558 16777 14564 16839
rect 14494 16771 14564 16777
rect 15942 16839 16012 16843
rect 15942 16777 15946 16839
rect 15946 16777 16006 16839
rect 16006 16777 16012 16839
rect 15942 16771 16012 16777
rect 17440 16837 17510 16841
rect 17440 16775 17444 16837
rect 17444 16775 17504 16837
rect 17504 16775 17510 16837
rect 17440 16769 17510 16775
rect 18888 16837 18958 16841
rect 18888 16775 18892 16837
rect 18892 16775 18952 16837
rect 18952 16775 18958 16837
rect 18888 16769 18958 16775
rect 20408 16839 20478 16843
rect 20408 16777 20412 16839
rect 20412 16777 20472 16839
rect 20472 16777 20478 16839
rect 20408 16771 20478 16777
rect 21856 16839 21926 16843
rect 21856 16777 21860 16839
rect 21860 16777 21920 16839
rect 21920 16777 21926 16839
rect 21856 16771 21926 16777
rect 23354 16837 23424 16841
rect 23354 16775 23358 16837
rect 23358 16775 23418 16837
rect 23418 16775 23424 16837
rect 23354 16769 23424 16775
rect 24802 16837 24872 16841
rect 24802 16775 24806 16837
rect 24806 16775 24866 16837
rect 24866 16775 24872 16837
rect 24802 16769 24872 16775
rect 5077 15721 5187 15731
rect 5077 15630 5087 15721
rect 5087 15630 5177 15721
rect 5177 15630 5187 15721
rect 5077 15620 5187 15630
rect 6245 15721 6355 15731
rect 6245 15630 6255 15721
rect 6255 15630 6345 15721
rect 6345 15630 6355 15721
rect 6245 15620 6355 15630
rect 7413 15721 7523 15731
rect 7413 15630 7423 15721
rect 7423 15630 7513 15721
rect 7513 15630 7523 15721
rect 7413 15620 7523 15630
rect 8581 15721 8691 15731
rect 8581 15630 8591 15721
rect 8591 15630 8681 15721
rect 8681 15630 8691 15721
rect 8581 15620 8691 15630
rect 9755 15719 9865 15729
rect 9755 15628 9765 15719
rect 9765 15628 9855 15719
rect 9855 15628 9865 15719
rect 9755 15618 9865 15628
rect 10923 15719 11033 15729
rect 10923 15628 10933 15719
rect 10933 15628 11023 15719
rect 11023 15628 11033 15719
rect 10923 15618 11033 15628
rect 12091 15719 12201 15729
rect 12091 15628 12101 15719
rect 12101 15628 12191 15719
rect 12191 15628 12201 15719
rect 12091 15618 12201 15628
rect 13259 15719 13369 15729
rect 13259 15628 13269 15719
rect 13269 15628 13359 15719
rect 13359 15628 13369 15719
rect 13259 15618 13369 15628
rect 14268 15633 14342 15639
rect 14268 15571 14272 15633
rect 14272 15571 14336 15633
rect 14336 15571 14342 15633
rect 15716 15633 15790 15639
rect 15716 15571 15720 15633
rect 15720 15571 15784 15633
rect 15784 15571 15790 15633
rect 17214 15631 17288 15637
rect 17214 15569 17218 15631
rect 17218 15569 17282 15631
rect 17282 15569 17288 15631
rect 18662 15631 18736 15637
rect 18662 15569 18666 15631
rect 18666 15569 18730 15631
rect 18730 15569 18736 15631
rect 1770 15038 1870 15128
rect 1770 15036 1870 15038
rect 4914 15038 5014 15128
rect 4914 15036 5014 15038
rect 8046 15034 8146 15124
rect 8046 15032 8146 15034
rect 1772 12828 1774 12886
rect 1774 12828 1850 12886
rect 1850 12828 1856 12886
rect 1772 12818 1856 12828
rect 4916 12828 4918 12886
rect 4918 12828 4994 12886
rect 4994 12828 5000 12886
rect 4916 12818 5000 12828
rect 8048 12824 8050 12882
rect 8050 12824 8126 12882
rect 8126 12824 8132 12882
rect 8048 12814 8132 12824
rect 1770 12304 1870 12394
rect 1770 12302 1870 12304
rect 4914 12304 5014 12394
rect 4914 12302 5014 12304
rect 8046 12300 8146 12390
rect 8046 12298 8146 12300
rect 1772 10094 1774 10152
rect 1774 10094 1850 10152
rect 1850 10094 1856 10152
rect 1772 10084 1856 10094
rect 4916 10094 4918 10152
rect 4918 10094 4994 10152
rect 4994 10094 5000 10152
rect 4916 10084 5000 10094
rect 8048 10090 8050 10148
rect 8050 10090 8126 10148
rect 8126 10090 8132 10148
rect 8048 10080 8132 10090
rect 1780 9572 1880 9662
rect 1780 9570 1880 9572
rect 4924 9572 5024 9662
rect 4924 9570 5024 9572
rect 8056 9568 8156 9658
rect 8056 9566 8156 9568
rect 1782 7362 1784 7420
rect 1784 7362 1860 7420
rect 1860 7362 1866 7420
rect 1782 7352 1866 7362
rect 4926 7362 4928 7420
rect 4928 7362 5004 7420
rect 5004 7362 5010 7420
rect 4926 7352 5010 7362
rect 8058 7358 8060 7416
rect 8060 7358 8136 7416
rect 8136 7358 8142 7416
rect 8058 7348 8142 7358
rect 3265 6761 3375 6775
rect 3265 6677 3273 6761
rect 3273 6677 3367 6761
rect 3367 6677 3375 6761
rect 3265 6667 3375 6677
rect 4003 6761 4113 6775
rect 4003 6677 4011 6761
rect 4011 6677 4105 6761
rect 4105 6677 4113 6761
rect 4003 6667 4113 6677
rect 4741 6761 4851 6775
rect 4741 6677 4749 6761
rect 4749 6677 4843 6761
rect 4843 6677 4851 6761
rect 4741 6667 4851 6677
rect 5479 6761 5589 6775
rect 5479 6677 5487 6761
rect 5487 6677 5581 6761
rect 5581 6677 5589 6761
rect 5479 6667 5589 6677
rect 6219 6761 6329 6775
rect 6219 6677 6227 6761
rect 6227 6677 6321 6761
rect 6321 6677 6329 6761
rect 6219 6667 6329 6677
rect 6961 6761 7071 6775
rect 6961 6677 6969 6761
rect 6969 6677 7063 6761
rect 7063 6677 7071 6761
rect 6961 6667 7071 6677
rect 7699 6761 7809 6775
rect 7699 6677 7707 6761
rect 7707 6677 7801 6761
rect 7801 6677 7809 6761
rect 7699 6667 7809 6677
rect 8437 6763 8547 6777
rect 8437 6679 8445 6763
rect 8445 6679 8539 6763
rect 8539 6679 8547 6763
rect 8437 6669 8547 6679
rect 10051 6706 10127 6708
rect 10051 6642 10127 6706
rect 11190 15034 11290 15124
rect 11190 15032 11290 15034
rect 11192 12824 11194 12882
rect 11194 12824 11270 12882
rect 11270 12824 11276 12882
rect 11192 12814 11276 12824
rect 11190 12300 11290 12390
rect 11190 12298 11290 12300
rect 11192 10090 11194 10148
rect 11194 10090 11270 10148
rect 11270 10090 11276 10148
rect 11192 10080 11276 10090
rect 11200 9568 11300 9658
rect 11200 9566 11300 9568
rect 11202 7358 11204 7416
rect 11204 7358 11280 7416
rect 11280 7358 11286 7416
rect 11202 7348 11286 7358
rect 12119 6704 12195 6706
rect 12119 6640 12195 6704
rect 3333 5863 3435 5883
rect 3333 5805 3353 5863
rect 3353 5805 3419 5863
rect 3419 5805 3435 5863
rect 3333 5783 3435 5805
rect 4071 5863 4173 5883
rect 4071 5805 4091 5863
rect 4091 5805 4157 5863
rect 4157 5805 4173 5863
rect 4071 5783 4173 5805
rect 4809 5863 4911 5883
rect 4809 5805 4829 5863
rect 4829 5805 4895 5863
rect 4895 5805 4911 5863
rect 4809 5783 4911 5805
rect 5547 5863 5649 5883
rect 5547 5805 5567 5863
rect 5567 5805 5633 5863
rect 5633 5805 5649 5863
rect 5547 5783 5649 5805
rect 6287 5863 6389 5883
rect 6287 5805 6307 5863
rect 6307 5805 6373 5863
rect 6373 5805 6389 5863
rect 6287 5783 6389 5805
rect 7029 5863 7131 5883
rect 7029 5805 7049 5863
rect 7049 5805 7115 5863
rect 7115 5805 7131 5863
rect 7029 5783 7131 5805
rect 7767 5863 7869 5883
rect 7767 5805 7787 5863
rect 7787 5805 7853 5863
rect 7853 5805 7869 5863
rect 7767 5783 7869 5805
rect 8505 5865 8607 5885
rect 8505 5807 8525 5865
rect 8525 5807 8591 5865
rect 8591 5807 8607 5865
rect 8505 5785 8607 5807
rect 14392 15038 14492 15128
rect 14392 15036 14492 15038
rect 14394 12828 14396 12886
rect 14396 12828 14472 12886
rect 14472 12828 14478 12886
rect 14394 12818 14478 12828
rect 14392 12304 14492 12394
rect 14392 12302 14492 12304
rect 14394 10094 14396 10152
rect 14396 10094 14472 10152
rect 14472 10094 14478 10152
rect 14394 10084 14478 10094
rect 14402 9572 14502 9662
rect 14402 9570 14502 9572
rect 14404 7362 14406 7420
rect 14406 7362 14482 7420
rect 14482 7362 14488 7420
rect 14404 7352 14488 7362
rect 14188 6706 14264 6708
rect 14188 6642 14264 6706
rect 20182 15633 20256 15639
rect 20182 15571 20186 15633
rect 20186 15571 20250 15633
rect 20250 15571 20256 15633
rect 16256 6704 16332 6706
rect 16256 6640 16332 6704
rect 17536 15038 17636 15128
rect 17536 15036 17636 15038
rect 17538 12828 17540 12886
rect 17540 12828 17616 12886
rect 17616 12828 17622 12886
rect 17538 12818 17622 12828
rect 17536 12304 17636 12394
rect 17536 12302 17636 12304
rect 17538 10094 17540 10152
rect 17540 10094 17616 10152
rect 17616 10094 17622 10152
rect 17538 10084 17622 10094
rect 17546 9572 17646 9662
rect 17546 9570 17646 9572
rect 17548 7362 17550 7420
rect 17550 7362 17626 7420
rect 17626 7362 17632 7420
rect 17548 7352 17632 7362
rect 18325 6704 18401 6706
rect 18325 6640 18401 6704
rect 20668 15034 20768 15124
rect 20668 15032 20768 15034
rect 20670 12824 20672 12882
rect 20672 12824 20748 12882
rect 20748 12824 20754 12882
rect 20670 12814 20754 12824
rect 20668 12300 20768 12390
rect 20668 12298 20768 12300
rect 20670 10090 20672 10148
rect 20672 10090 20748 10148
rect 20748 10090 20754 10148
rect 20670 10080 20754 10090
rect 20678 9568 20778 9658
rect 20678 9566 20778 9568
rect 20680 7358 20682 7416
rect 20682 7358 20758 7416
rect 20758 7358 20764 7416
rect 20680 7348 20764 7358
rect 20393 6702 20469 6704
rect 20393 6638 20469 6702
rect 21630 15633 21704 15639
rect 21630 15571 21634 15633
rect 21634 15571 21698 15633
rect 21698 15571 21704 15633
rect 23128 15631 23202 15637
rect 23128 15569 23132 15631
rect 23132 15569 23196 15631
rect 23196 15569 23202 15631
rect 22462 6704 22538 6706
rect 22462 6640 22538 6704
rect 24576 15631 24650 15637
rect 24576 15569 24580 15631
rect 24580 15569 24644 15631
rect 24644 15569 24650 15631
rect 23812 15034 23912 15124
rect 23812 15032 23912 15034
rect 23814 12824 23816 12882
rect 23816 12824 23892 12882
rect 23892 12824 23898 12882
rect 23814 12814 23898 12824
rect 23812 12300 23912 12390
rect 23812 12298 23912 12300
rect 23814 10090 23816 10148
rect 23816 10090 23892 10148
rect 23892 10090 23898 10148
rect 23814 10080 23898 10090
rect 23822 9568 23922 9658
rect 23822 9566 23922 9568
rect 23824 7358 23826 7416
rect 23826 7358 23902 7416
rect 23902 7358 23908 7416
rect 23824 7348 23908 7358
rect 24530 6702 24606 6704
rect 24530 6638 24606 6702
rect 29693 12277 29695 12353
rect 29695 12277 29759 12353
rect 31915 12405 32003 12415
rect 31915 12333 31925 12405
rect 31925 12333 31995 12405
rect 31995 12333 32003 12405
rect 31915 12321 32003 12333
rect 40022 23180 40221 23211
rect 40022 23051 40044 23180
rect 40044 23051 40197 23180
rect 40197 23051 40221 23180
rect 40022 23032 40221 23051
rect 46535 23177 46734 23208
rect 46535 23048 46557 23177
rect 46557 23048 46710 23177
rect 46710 23048 46734 23177
rect 46535 23029 46734 23048
rect 41835 22837 42034 22868
rect 41835 22708 41857 22837
rect 41857 22708 42010 22837
rect 42010 22708 42034 22837
rect 41835 22689 42034 22708
rect 43733 22837 43932 22868
rect 43733 22708 43755 22837
rect 43755 22708 43908 22837
rect 43908 22708 43932 22837
rect 43733 22689 43932 22708
rect 40306 22141 40485 22163
rect 40306 21988 40325 22141
rect 40325 21988 40454 22141
rect 40454 21988 40485 22141
rect 40306 21964 40485 21988
rect 40017 21576 40216 21607
rect 40017 21447 40039 21576
rect 40039 21447 40192 21576
rect 40192 21447 40216 21576
rect 40017 21428 40216 21447
rect 40301 20537 40480 20559
rect 40301 20384 40320 20537
rect 40320 20384 40449 20537
rect 40449 20384 40480 20537
rect 40301 20360 40480 20384
rect 41779 20440 41978 20459
rect 41779 20311 41803 20440
rect 41803 20311 41956 20440
rect 41956 20311 41978 20440
rect 41779 20280 41978 20311
rect 43677 20440 43876 20459
rect 43677 20311 43701 20440
rect 43701 20311 43854 20440
rect 43854 20311 43876 20440
rect 43677 20280 43876 20311
rect 48348 22834 48547 22865
rect 48348 22705 48370 22834
rect 48370 22705 48523 22834
rect 48523 22705 48547 22834
rect 48348 22686 48547 22705
rect 50246 22834 50445 22865
rect 50246 22705 50268 22834
rect 50268 22705 50421 22834
rect 50421 22705 50445 22834
rect 50246 22686 50445 22705
rect 46819 22138 46998 22160
rect 46819 21985 46838 22138
rect 46838 21985 46967 22138
rect 46967 21985 46998 22138
rect 46819 21961 46998 21985
rect 46530 21573 46729 21604
rect 46530 21444 46552 21573
rect 46552 21444 46705 21573
rect 46705 21444 46729 21573
rect 46530 21425 46729 21444
rect 46814 20534 46993 20556
rect 46814 20381 46833 20534
rect 46833 20381 46962 20534
rect 46962 20381 46993 20534
rect 46814 20357 46993 20381
rect 48292 20437 48491 20456
rect 48292 20308 48316 20437
rect 48316 20308 48469 20437
rect 48469 20308 48491 20437
rect 48292 20277 48491 20308
rect 50190 20437 50389 20456
rect 50190 20308 50214 20437
rect 50214 20308 50367 20437
rect 50367 20308 50389 20437
rect 50190 20277 50389 20308
rect 29691 10209 29693 10285
rect 29693 10209 29757 10285
rect 31913 10337 32001 10347
rect 31913 10265 31923 10337
rect 31923 10265 31993 10337
rect 31993 10265 32001 10337
rect 31913 10253 32001 10265
rect 53069 23172 53268 23203
rect 53069 23043 53091 23172
rect 53091 23043 53244 23172
rect 53244 23043 53268 23172
rect 53069 23024 53268 23043
rect 54882 22829 55081 22860
rect 54882 22700 54904 22829
rect 54904 22700 55057 22829
rect 55057 22700 55081 22829
rect 54882 22681 55081 22700
rect 56780 22829 56979 22860
rect 56780 22700 56802 22829
rect 56802 22700 56955 22829
rect 56955 22700 56979 22829
rect 56780 22681 56979 22700
rect 53353 22133 53532 22155
rect 53353 21980 53372 22133
rect 53372 21980 53501 22133
rect 53501 21980 53532 22133
rect 53353 21956 53532 21980
rect 53064 21568 53263 21599
rect 53064 21439 53086 21568
rect 53086 21439 53239 21568
rect 53239 21439 53263 21568
rect 53064 21420 53263 21439
rect 53348 20529 53527 20551
rect 53348 20376 53367 20529
rect 53367 20376 53496 20529
rect 53496 20376 53527 20529
rect 53348 20352 53527 20376
rect 54826 20432 55025 20451
rect 54826 20303 54850 20432
rect 54850 20303 55003 20432
rect 55003 20303 55025 20432
rect 54826 20272 55025 20303
rect 56724 20432 56923 20451
rect 56724 20303 56748 20432
rect 56748 20303 56901 20432
rect 56901 20303 56923 20432
rect 56724 20272 56923 20303
rect 29693 8140 29695 8216
rect 29695 8140 29759 8216
rect 31915 8268 32003 8278
rect 31915 8196 31925 8268
rect 31925 8196 31995 8268
rect 31995 8196 32003 8268
rect 31915 8184 32003 8196
rect 59627 23176 59826 23207
rect 59627 23047 59649 23176
rect 59649 23047 59802 23176
rect 59802 23047 59826 23176
rect 59627 23028 59826 23047
rect 61440 22833 61639 22864
rect 61440 22704 61462 22833
rect 61462 22704 61615 22833
rect 61615 22704 61639 22833
rect 61440 22685 61639 22704
rect 63338 22833 63537 22864
rect 63338 22704 63360 22833
rect 63360 22704 63513 22833
rect 63513 22704 63537 22833
rect 63338 22685 63537 22704
rect 59911 22137 60090 22159
rect 59911 21984 59930 22137
rect 59930 21984 60059 22137
rect 60059 21984 60090 22137
rect 59911 21960 60090 21984
rect 59622 21572 59821 21603
rect 59622 21443 59644 21572
rect 59644 21443 59797 21572
rect 59797 21443 59821 21572
rect 59622 21424 59821 21443
rect 70243 20725 70333 20825
rect 70333 20725 70335 20825
rect 72485 20805 72553 20811
rect 72485 20729 72543 20805
rect 72543 20729 72553 20805
rect 72485 20727 72553 20729
rect 59906 20533 60085 20555
rect 59906 20380 59925 20533
rect 59925 20380 60054 20533
rect 60054 20380 60085 20533
rect 59906 20356 60085 20380
rect 61384 20436 61583 20455
rect 61384 20307 61408 20436
rect 61408 20307 61561 20436
rect 61561 20307 61583 20436
rect 61384 20276 61583 20307
rect 63282 20436 63481 20455
rect 63282 20307 63306 20436
rect 63306 20307 63459 20436
rect 63459 20307 63481 20436
rect 63282 20276 63481 20307
rect 29691 6072 29693 6148
rect 29693 6072 29757 6148
rect 31913 6200 32001 6210
rect 31913 6128 31923 6200
rect 31923 6128 31993 6200
rect 31993 6128 32001 6200
rect 31913 6116 32001 6128
rect 39584 19276 39783 19307
rect 39584 19147 39608 19276
rect 39608 19147 39761 19276
rect 39761 19147 39783 19276
rect 39584 19128 39783 19147
rect 40731 19276 40930 19307
rect 40731 19147 40755 19276
rect 40755 19147 40908 19276
rect 40908 19147 40930 19276
rect 40731 19128 40930 19147
rect 43213 19222 43412 19253
rect 43213 19093 43237 19222
rect 43237 19093 43390 19222
rect 43390 19093 43412 19222
rect 43213 19074 43412 19093
rect 46142 19272 46341 19303
rect 46142 19143 46166 19272
rect 46166 19143 46319 19272
rect 46319 19143 46341 19272
rect 46142 19124 46341 19143
rect 47289 19272 47488 19303
rect 47289 19143 47313 19272
rect 47313 19143 47466 19272
rect 47466 19143 47488 19272
rect 47289 19124 47488 19143
rect 49771 19218 49970 19249
rect 49771 19089 49795 19218
rect 49795 19089 49948 19218
rect 49948 19089 49970 19218
rect 49771 19070 49970 19089
rect 52676 19277 52875 19308
rect 52676 19148 52700 19277
rect 52700 19148 52853 19277
rect 52853 19148 52875 19277
rect 52676 19129 52875 19148
rect 53823 19277 54022 19308
rect 53823 19148 53847 19277
rect 53847 19148 54000 19277
rect 54000 19148 54022 19277
rect 53823 19129 54022 19148
rect 56305 19223 56504 19254
rect 56305 19094 56329 19223
rect 56329 19094 56482 19223
rect 56482 19094 56504 19223
rect 56305 19075 56504 19094
rect 59189 19280 59388 19311
rect 59189 19151 59213 19280
rect 59213 19151 59366 19280
rect 59366 19151 59388 19280
rect 59189 19132 59388 19151
rect 60336 19280 60535 19311
rect 60336 19151 60360 19280
rect 60360 19151 60513 19280
rect 60513 19151 60535 19280
rect 60336 19132 60535 19151
rect 62818 19226 63017 19257
rect 62818 19097 62842 19226
rect 62842 19097 62995 19226
rect 62995 19097 63017 19226
rect 62818 19078 63017 19097
rect 42949 18183 43128 18205
rect 42949 18030 42980 18183
rect 42980 18030 43109 18183
rect 43109 18030 43128 18183
rect 42949 18006 43128 18030
rect 49507 18179 49686 18201
rect 49507 18026 49538 18179
rect 49538 18026 49667 18179
rect 49667 18026 49686 18179
rect 49507 18002 49686 18026
rect 56041 18184 56220 18206
rect 56041 18031 56072 18184
rect 56072 18031 56201 18184
rect 56201 18031 56220 18184
rect 56041 18007 56220 18031
rect 62554 18187 62733 18209
rect 62554 18034 62585 18187
rect 62585 18034 62714 18187
rect 62714 18034 62733 18187
rect 62554 18010 62733 18034
rect 40244 17873 40443 17892
rect 40244 17744 40266 17873
rect 40266 17744 40419 17873
rect 40419 17744 40443 17873
rect 40244 17713 40443 17744
rect 41386 17875 41585 17894
rect 41386 17746 41408 17875
rect 41408 17746 41561 17875
rect 41561 17746 41585 17875
rect 41386 17715 41585 17746
rect 46802 17869 47001 17888
rect 46802 17740 46824 17869
rect 46824 17740 46977 17869
rect 46977 17740 47001 17869
rect 46802 17709 47001 17740
rect 47944 17871 48143 17890
rect 47944 17742 47966 17871
rect 47966 17742 48119 17871
rect 48119 17742 48143 17871
rect 47944 17711 48143 17742
rect 53336 17874 53535 17893
rect 53336 17745 53358 17874
rect 53358 17745 53511 17874
rect 53511 17745 53535 17874
rect 53336 17714 53535 17745
rect 54478 17876 54677 17895
rect 54478 17747 54500 17876
rect 54500 17747 54653 17876
rect 54653 17747 54677 17876
rect 54478 17716 54677 17747
rect 59849 17877 60048 17896
rect 59849 17748 59871 17877
rect 59871 17748 60024 17877
rect 60024 17748 60048 17877
rect 59849 17717 60048 17748
rect 60991 17879 61190 17898
rect 60991 17750 61013 17879
rect 61013 17750 61166 17879
rect 61166 17750 61190 17879
rect 60991 17719 61190 17750
rect 43199 17572 43398 17603
rect 43199 17443 43223 17572
rect 43223 17443 43376 17572
rect 43376 17443 43398 17572
rect 43199 17424 43398 17443
rect 49757 17568 49956 17599
rect 49757 17439 49781 17568
rect 49781 17439 49934 17568
rect 49934 17439 49956 17568
rect 49757 17420 49956 17439
rect 56291 17573 56490 17604
rect 56291 17444 56315 17573
rect 56315 17444 56468 17573
rect 56468 17444 56490 17573
rect 56291 17425 56490 17444
rect 62804 17576 63003 17607
rect 62804 17447 62828 17576
rect 62828 17447 62981 17576
rect 62981 17447 63003 17576
rect 62804 17428 63003 17447
rect 70243 17581 70333 17681
rect 70333 17581 70335 17681
rect 72485 17661 72553 17667
rect 72485 17585 72543 17661
rect 72543 17585 72553 17661
rect 72485 17583 72553 17585
rect 39488 17229 39687 17260
rect 39488 17100 39512 17229
rect 39512 17100 39665 17229
rect 39665 17100 39687 17229
rect 39488 17081 39687 17100
rect 41386 17229 41585 17260
rect 41386 17100 41410 17229
rect 41410 17100 41563 17229
rect 41563 17100 41585 17229
rect 41386 17081 41585 17100
rect 46046 17225 46245 17256
rect 46046 17096 46070 17225
rect 46070 17096 46223 17225
rect 46223 17096 46245 17225
rect 46046 17077 46245 17096
rect 47944 17225 48143 17256
rect 47944 17096 47968 17225
rect 47968 17096 48121 17225
rect 48121 17096 48143 17225
rect 47944 17077 48143 17096
rect 52580 17230 52779 17261
rect 52580 17101 52604 17230
rect 52604 17101 52757 17230
rect 52757 17101 52779 17230
rect 52580 17082 52779 17101
rect 54478 17230 54677 17261
rect 54478 17101 54502 17230
rect 54502 17101 54655 17230
rect 54655 17101 54677 17230
rect 54478 17082 54677 17101
rect 59093 17233 59292 17264
rect 59093 17104 59117 17233
rect 59117 17104 59270 17233
rect 59270 17104 59292 17233
rect 59093 17085 59292 17104
rect 60991 17233 61190 17264
rect 60991 17104 61015 17233
rect 61015 17104 61168 17233
rect 61168 17104 61190 17233
rect 60991 17085 61190 17104
rect 42935 16533 43114 16555
rect 42935 16380 42966 16533
rect 42966 16380 43095 16533
rect 43095 16380 43114 16533
rect 42935 16356 43114 16380
rect 49493 16529 49672 16551
rect 49493 16376 49524 16529
rect 49524 16376 49653 16529
rect 49653 16376 49672 16529
rect 49493 16352 49672 16376
rect 56027 16534 56206 16556
rect 56027 16381 56058 16534
rect 56058 16381 56187 16534
rect 56187 16381 56206 16534
rect 56027 16357 56206 16381
rect 62540 16537 62719 16559
rect 62540 16384 62571 16537
rect 62571 16384 62700 16537
rect 62700 16384 62719 16537
rect 62540 16360 62719 16384
rect 43204 15968 43403 15999
rect 43204 15839 43228 15968
rect 43228 15839 43381 15968
rect 43381 15839 43403 15968
rect 43204 15820 43403 15839
rect 49762 15964 49961 15995
rect 49762 15835 49786 15964
rect 49786 15835 49939 15964
rect 49939 15835 49961 15964
rect 49762 15816 49961 15835
rect 56296 15969 56495 16000
rect 56296 15840 56320 15969
rect 56320 15840 56473 15969
rect 56473 15840 56495 15969
rect 56296 15821 56495 15840
rect 62809 15972 63008 16003
rect 62809 15843 62833 15972
rect 62833 15843 62986 15972
rect 62986 15843 63008 15972
rect 62809 15824 63008 15843
rect 42940 14929 43119 14951
rect 39544 14832 39743 14851
rect 39544 14703 39566 14832
rect 39566 14703 39719 14832
rect 39719 14703 39743 14832
rect 39544 14672 39743 14703
rect 41442 14832 41641 14851
rect 41442 14703 41464 14832
rect 41464 14703 41617 14832
rect 41617 14703 41641 14832
rect 41442 14672 41641 14703
rect 42940 14776 42971 14929
rect 42971 14776 43100 14929
rect 43100 14776 43119 14929
rect 49498 14925 49677 14947
rect 42940 14752 43119 14776
rect 46102 14828 46301 14847
rect 46102 14699 46124 14828
rect 46124 14699 46277 14828
rect 46277 14699 46301 14828
rect 46102 14668 46301 14699
rect 48000 14828 48199 14847
rect 48000 14699 48022 14828
rect 48022 14699 48175 14828
rect 48175 14699 48199 14828
rect 48000 14668 48199 14699
rect 49498 14772 49529 14925
rect 49529 14772 49658 14925
rect 49658 14772 49677 14925
rect 56032 14930 56211 14952
rect 49498 14748 49677 14772
rect 52636 14833 52835 14852
rect 52636 14704 52658 14833
rect 52658 14704 52811 14833
rect 52811 14704 52835 14833
rect 52636 14673 52835 14704
rect 54534 14833 54733 14852
rect 54534 14704 54556 14833
rect 54556 14704 54709 14833
rect 54709 14704 54733 14833
rect 54534 14673 54733 14704
rect 56032 14777 56063 14930
rect 56063 14777 56192 14930
rect 56192 14777 56211 14930
rect 62545 14933 62724 14955
rect 56032 14753 56211 14777
rect 59149 14836 59348 14855
rect 59149 14707 59171 14836
rect 59171 14707 59324 14836
rect 59324 14707 59348 14836
rect 59149 14676 59348 14707
rect 61047 14836 61246 14855
rect 61047 14707 61069 14836
rect 61069 14707 61222 14836
rect 61222 14707 61246 14836
rect 61047 14676 61246 14707
rect 62545 14780 62576 14933
rect 62576 14780 62705 14933
rect 62705 14780 62724 14933
rect 62545 14756 62724 14780
rect 70239 14449 70329 14549
rect 70329 14449 70331 14549
rect 72481 14529 72549 14535
rect 72481 14453 72539 14529
rect 72539 14453 72549 14529
rect 72481 14451 72549 14453
rect 10095 4476 10189 4486
rect 10095 4406 10107 4476
rect 10107 4406 10179 4476
rect 10179 4406 10189 4476
rect 10095 4398 10189 4406
rect 12163 4474 12257 4484
rect 12163 4404 12175 4474
rect 12175 4404 12247 4474
rect 12247 4404 12257 4474
rect 12163 4396 12257 4404
rect 14232 4476 14326 4486
rect 14232 4406 14244 4476
rect 14244 4406 14316 4476
rect 14316 4406 14326 4476
rect 14232 4398 14326 4406
rect 16300 4474 16394 4484
rect 16300 4404 16312 4474
rect 16312 4404 16384 4474
rect 16384 4404 16394 4474
rect 16300 4396 16394 4404
rect 18369 4474 18463 4484
rect 18369 4404 18381 4474
rect 18381 4404 18453 4474
rect 18453 4404 18463 4474
rect 18369 4396 18463 4404
rect 20437 4472 20531 4482
rect 20437 4402 20449 4472
rect 20449 4402 20521 4472
rect 20521 4402 20531 4472
rect 20437 4394 20531 4402
rect 22506 4474 22600 4484
rect 22506 4404 22518 4474
rect 22518 4404 22590 4474
rect 22590 4404 22600 4474
rect 22506 4396 22600 4404
rect 24574 4472 24668 4482
rect 24574 4402 24586 4472
rect 24586 4402 24658 4472
rect 24658 4402 24668 4472
rect 24574 4394 24668 4402
rect 1496 2320 1596 2410
rect 1496 2318 1596 2320
rect 1510 110 1516 168
rect 1516 110 1592 168
rect 1592 110 1594 168
rect 1510 100 1594 110
rect 4640 2320 4740 2410
rect 4640 2318 4740 2320
rect 4654 110 4660 168
rect 4660 110 4736 168
rect 4736 110 4738 168
rect 4654 100 4738 110
rect 7772 2324 7872 2414
rect 7772 2322 7872 2324
rect 7786 114 7792 172
rect 7792 114 7868 172
rect 7868 114 7870 172
rect 7786 104 7870 114
rect 10916 2324 11016 2414
rect 10916 2322 11016 2324
rect 10930 114 10936 172
rect 10936 114 11012 172
rect 11012 114 11014 172
rect 10930 104 11014 114
rect 14118 2320 14218 2410
rect 14118 2318 14218 2320
rect 14132 110 14138 168
rect 14138 110 14214 168
rect 14214 110 14216 168
rect 14132 100 14216 110
rect 29691 4003 29693 4079
rect 29693 4003 29757 4079
rect 31913 4131 32001 4141
rect 31913 4059 31923 4131
rect 31923 4059 31993 4131
rect 31993 4059 32001 4131
rect 31913 4047 32001 4059
rect 17262 2320 17362 2410
rect 17262 2318 17362 2320
rect 20394 2324 20494 2414
rect 20394 2322 20494 2324
rect 23538 2324 23638 2414
rect 23538 2322 23638 2324
rect 29689 1935 29691 2011
rect 29691 1935 29755 2011
rect 31911 2063 31999 2073
rect 31911 1991 31921 2063
rect 31921 1991 31991 2063
rect 31991 1991 31999 2063
rect 31911 1979 31999 1991
rect 17276 110 17282 168
rect 17282 110 17358 168
rect 17358 110 17360 168
rect 17276 100 17360 110
rect 20408 114 20414 172
rect 20414 114 20490 172
rect 20490 114 20492 172
rect 20408 104 20492 114
rect 23552 114 23558 172
rect 23558 114 23634 172
rect 23634 114 23636 172
rect 23552 104 23636 114
rect 29691 -134 29693 -58
rect 29693 -134 29757 -58
rect 31913 -6 32001 4
rect 31913 -78 31923 -6
rect 31923 -78 31993 -6
rect 31993 -78 32001 -6
rect 31913 -90 32001 -78
rect 1528 -1572 1628 -1482
rect 1528 -1574 1628 -1572
rect 4672 -1572 4772 -1482
rect 4672 -1574 4772 -1572
rect 7804 -1568 7904 -1478
rect 7804 -1570 7904 -1568
rect 10948 -1568 11048 -1478
rect 10948 -1570 11048 -1568
rect 14150 -1572 14250 -1482
rect 14150 -1574 14250 -1572
rect 17294 -1572 17394 -1482
rect 17294 -1574 17394 -1572
rect 20426 -1568 20526 -1478
rect 20426 -1570 20526 -1568
rect 23570 -1568 23670 -1478
rect 23570 -1570 23670 -1568
rect 29689 -2202 29691 -2126
rect 29691 -2202 29755 -2126
rect 31911 -2074 31999 -2064
rect 31911 -2146 31921 -2074
rect 31921 -2146 31991 -2074
rect 31991 -2146 31999 -2074
rect 31911 -2158 31999 -2146
rect 41905 12375 41975 12379
rect 41905 12313 41911 12375
rect 41911 12313 41971 12375
rect 41971 12313 41975 12375
rect 41905 12307 41975 12313
rect 48454 12374 48524 12378
rect 48454 12312 48460 12374
rect 48460 12312 48520 12374
rect 48520 12312 48524 12374
rect 48454 12306 48524 12312
rect 55108 12395 55178 12399
rect 55108 12333 55114 12395
rect 55114 12333 55174 12395
rect 55174 12333 55178 12395
rect 55108 12327 55178 12333
rect 63761 12228 63831 12232
rect 63761 12166 63767 12228
rect 63767 12166 63827 12228
rect 63827 12166 63831 12228
rect 63761 12160 63831 12166
rect 65991 12168 66190 12199
rect 65991 12039 66013 12168
rect 66013 12039 66166 12168
rect 66166 12039 66190 12168
rect 65991 12020 66190 12039
rect 67362 11820 67432 11824
rect 67362 11758 67368 11820
rect 67368 11758 67428 11820
rect 67428 11758 67432 11820
rect 67362 11752 67432 11758
rect 42127 11169 42201 11175
rect 42127 11107 42133 11169
rect 42133 11107 42197 11169
rect 42197 11107 42201 11169
rect 48676 11168 48750 11174
rect 48676 11106 48682 11168
rect 48682 11106 48746 11168
rect 48746 11106 48750 11168
rect 55330 11189 55404 11195
rect 55330 11127 55336 11189
rect 55336 11127 55400 11189
rect 55400 11127 55404 11189
rect 63983 11022 64057 11028
rect 63983 10960 63989 11022
rect 63989 10960 64053 11022
rect 64053 10960 64057 11022
rect 67457 10614 67795 10646
rect 67457 10552 67590 10614
rect 67590 10552 67654 10614
rect 67654 10552 67795 10614
rect 67457 10530 67795 10552
rect 35241 10475 35311 10479
rect 35241 10413 35247 10475
rect 35247 10413 35307 10475
rect 35307 10413 35311 10475
rect 35241 10407 35311 10413
rect 38204 10279 38403 10310
rect 38204 10150 38226 10279
rect 38226 10150 38379 10279
rect 38379 10150 38403 10279
rect 38204 10131 38403 10150
rect 40686 10333 40885 10364
rect 40686 10204 40708 10333
rect 40708 10204 40861 10333
rect 40861 10204 40885 10333
rect 40686 10185 40885 10204
rect 41833 10333 42032 10364
rect 41833 10204 41855 10333
rect 41855 10204 42008 10333
rect 42008 10204 42032 10333
rect 41833 10185 42032 10204
rect 44753 10367 44952 10398
rect 44753 10238 44775 10367
rect 44775 10238 44928 10367
rect 44928 10238 44952 10367
rect 44753 10219 44952 10238
rect 47235 10421 47434 10452
rect 47235 10292 47257 10421
rect 47257 10292 47410 10421
rect 47410 10292 47434 10421
rect 47235 10273 47434 10292
rect 48382 10421 48581 10452
rect 48382 10292 48404 10421
rect 48404 10292 48557 10421
rect 48557 10292 48581 10421
rect 48382 10273 48581 10292
rect 51407 10299 51606 10330
rect 51407 10170 51429 10299
rect 51429 10170 51582 10299
rect 51582 10170 51606 10299
rect 51407 10151 51606 10170
rect 53889 10353 54088 10384
rect 53889 10224 53911 10353
rect 53911 10224 54064 10353
rect 54064 10224 54088 10353
rect 53889 10205 54088 10224
rect 55036 10353 55235 10384
rect 55036 10224 55058 10353
rect 55058 10224 55211 10353
rect 55211 10224 55235 10353
rect 55036 10205 55235 10224
rect 58032 10367 58231 10398
rect 58032 10238 58054 10367
rect 58054 10238 58207 10367
rect 58207 10238 58231 10367
rect 58032 10219 58231 10238
rect 60514 10421 60713 10452
rect 60514 10292 60536 10421
rect 60536 10292 60689 10421
rect 60689 10292 60713 10421
rect 60514 10273 60713 10292
rect 61661 10421 61860 10452
rect 61661 10292 61683 10421
rect 61683 10292 61836 10421
rect 61836 10292 61860 10421
rect 61661 10273 61860 10292
rect 63756 9657 63826 9661
rect 63756 9595 63762 9657
rect 63762 9595 63822 9657
rect 63822 9595 63826 9657
rect 63756 9589 63826 9595
rect 65912 9838 66178 9854
rect 65912 9681 65935 9838
rect 65935 9681 66146 9838
rect 66146 9681 66178 9838
rect 65912 9659 66178 9681
rect 35463 9269 35537 9275
rect 35463 9207 35469 9269
rect 35469 9207 35533 9269
rect 35533 9207 35537 9269
rect 38488 9240 38667 9262
rect 38488 9087 38507 9240
rect 38507 9087 38636 9240
rect 38636 9087 38667 9240
rect 38488 9063 38667 9087
rect 40031 8932 40230 8951
rect 40031 8803 40055 8932
rect 40055 8803 40208 8932
rect 40208 8803 40230 8932
rect 40031 8772 40230 8803
rect 41173 8930 41372 8949
rect 41173 8801 41197 8930
rect 41197 8801 41350 8930
rect 41350 8801 41372 8930
rect 41173 8770 41372 8801
rect 38218 8629 38417 8660
rect 38218 8500 38240 8629
rect 38240 8500 38393 8629
rect 38393 8500 38417 8629
rect 38218 8481 38417 8500
rect 40031 8286 40230 8317
rect 40031 8157 40053 8286
rect 40053 8157 40206 8286
rect 40206 8157 40230 8286
rect 40031 8138 40230 8157
rect 41929 8286 42128 8317
rect 41929 8157 41951 8286
rect 41951 8157 42104 8286
rect 42104 8157 42128 8286
rect 41929 8138 42128 8157
rect 35233 7890 35303 7894
rect 35233 7828 35239 7890
rect 35239 7828 35299 7890
rect 35299 7828 35303 7890
rect 35233 7822 35303 7828
rect 38502 7590 38681 7612
rect 38502 7437 38521 7590
rect 38521 7437 38650 7590
rect 38650 7437 38681 7590
rect 38502 7413 38681 7437
rect 38213 7025 38412 7056
rect 38213 6896 38235 7025
rect 38235 6896 38388 7025
rect 38388 6896 38412 7025
rect 38213 6877 38412 6896
rect 35455 6684 35529 6690
rect 35455 6622 35461 6684
rect 35461 6622 35525 6684
rect 35525 6622 35529 6684
rect 38497 5986 38676 6008
rect 38497 5833 38516 5986
rect 38516 5833 38645 5986
rect 38645 5833 38676 5986
rect 38497 5809 38676 5833
rect 39975 5889 40174 5908
rect 39975 5760 39999 5889
rect 39999 5760 40152 5889
rect 40152 5760 40174 5889
rect 39975 5729 40174 5760
rect 41873 5889 42072 5908
rect 41873 5760 41897 5889
rect 41897 5760 42050 5889
rect 42050 5760 42072 5889
rect 41873 5729 42072 5760
rect 45037 9328 45216 9350
rect 45037 9175 45056 9328
rect 45056 9175 45185 9328
rect 45185 9175 45216 9328
rect 45037 9151 45216 9175
rect 51691 9260 51870 9282
rect 51691 9107 51710 9260
rect 51710 9107 51839 9260
rect 51839 9107 51870 9260
rect 51691 9083 51870 9107
rect 46580 9020 46779 9039
rect 46580 8891 46604 9020
rect 46604 8891 46757 9020
rect 46757 8891 46779 9020
rect 46580 8860 46779 8891
rect 47722 9018 47921 9037
rect 47722 8889 47746 9018
rect 47746 8889 47899 9018
rect 47899 8889 47921 9018
rect 47722 8858 47921 8889
rect 53234 8952 53433 8971
rect 53234 8823 53258 8952
rect 53258 8823 53411 8952
rect 53411 8823 53433 8952
rect 53234 8792 53433 8823
rect 54376 8950 54575 8969
rect 54376 8821 54400 8950
rect 54400 8821 54553 8950
rect 54553 8821 54575 8950
rect 54376 8790 54575 8821
rect 44767 8717 44966 8748
rect 44767 8588 44789 8717
rect 44789 8588 44942 8717
rect 44942 8588 44966 8717
rect 44767 8569 44966 8588
rect 51421 8649 51620 8680
rect 51421 8520 51443 8649
rect 51443 8520 51596 8649
rect 51596 8520 51620 8649
rect 51421 8501 51620 8520
rect 46580 8374 46779 8405
rect 46580 8245 46602 8374
rect 46602 8245 46755 8374
rect 46755 8245 46779 8374
rect 46580 8226 46779 8245
rect 48478 8374 48677 8405
rect 48478 8245 48500 8374
rect 48500 8245 48653 8374
rect 48653 8245 48677 8374
rect 48478 8226 48677 8245
rect 53234 8306 53433 8337
rect 53234 8177 53256 8306
rect 53256 8177 53409 8306
rect 53409 8177 53433 8306
rect 53234 8158 53433 8177
rect 55132 8306 55331 8337
rect 55132 8177 55154 8306
rect 55154 8177 55307 8306
rect 55307 8177 55331 8306
rect 55132 8158 55331 8177
rect 45051 7678 45230 7700
rect 45051 7525 45070 7678
rect 45070 7525 45199 7678
rect 45199 7525 45230 7678
rect 45051 7501 45230 7525
rect 51705 7610 51884 7632
rect 51705 7457 51724 7610
rect 51724 7457 51853 7610
rect 51853 7457 51884 7610
rect 51705 7433 51884 7457
rect 44762 7113 44961 7144
rect 44762 6984 44784 7113
rect 44784 6984 44937 7113
rect 44937 6984 44961 7113
rect 44762 6965 44961 6984
rect 51416 7045 51615 7076
rect 51416 6916 51438 7045
rect 51438 6916 51591 7045
rect 51591 6916 51615 7045
rect 51416 6897 51615 6916
rect 45046 6074 45225 6096
rect 45046 5921 45065 6074
rect 45065 5921 45194 6074
rect 45194 5921 45225 6074
rect 51700 6006 51879 6028
rect 45046 5897 45225 5921
rect 46524 5977 46723 5996
rect 46524 5848 46548 5977
rect 46548 5848 46701 5977
rect 46701 5848 46723 5977
rect 46524 5817 46723 5848
rect 48422 5977 48621 5996
rect 48422 5848 48446 5977
rect 48446 5848 48599 5977
rect 48599 5848 48621 5977
rect 48422 5817 48621 5848
rect 51700 5853 51719 6006
rect 51719 5853 51848 6006
rect 51848 5853 51879 6006
rect 51700 5829 51879 5853
rect 53178 5909 53377 5928
rect 53178 5780 53202 5909
rect 53202 5780 53355 5909
rect 53355 5780 53377 5909
rect 53178 5749 53377 5780
rect 55076 5909 55275 5928
rect 55076 5780 55100 5909
rect 55100 5780 55253 5909
rect 55253 5780 55275 5909
rect 55076 5749 55275 5780
rect 35214 4612 35284 4616
rect 35214 4550 35220 4612
rect 35220 4550 35280 4612
rect 35280 4550 35284 4612
rect 35214 4544 35284 4550
rect 35436 3406 35510 3412
rect 35436 3344 35442 3406
rect 35442 3344 35506 3406
rect 35506 3344 35510 3406
rect 35230 1852 35300 1856
rect 35230 1790 35236 1852
rect 35236 1790 35296 1852
rect 35296 1790 35300 1852
rect 35230 1784 35300 1790
rect 38196 4499 38395 4530
rect 38196 4370 38218 4499
rect 38218 4370 38371 4499
rect 38371 4370 38395 4499
rect 38196 4351 38395 4370
rect 40678 4553 40877 4584
rect 40678 4424 40700 4553
rect 40700 4424 40853 4553
rect 40853 4424 40877 4553
rect 40678 4405 40877 4424
rect 41825 4553 42024 4584
rect 41825 4424 41847 4553
rect 41847 4424 42000 4553
rect 42000 4424 42024 4553
rect 41825 4405 42024 4424
rect 38480 3460 38659 3482
rect 38480 3307 38499 3460
rect 38499 3307 38628 3460
rect 38628 3307 38659 3460
rect 38480 3283 38659 3307
rect 40023 3152 40222 3171
rect 40023 3023 40047 3152
rect 40047 3023 40200 3152
rect 40200 3023 40222 3152
rect 40023 2992 40222 3023
rect 41165 3150 41364 3169
rect 41165 3021 41189 3150
rect 41189 3021 41342 3150
rect 41342 3021 41364 3150
rect 41165 2990 41364 3021
rect 38210 2849 38409 2880
rect 38210 2720 38232 2849
rect 38232 2720 38385 2849
rect 38385 2720 38409 2849
rect 38210 2701 38409 2720
rect 40023 2506 40222 2537
rect 40023 2377 40045 2506
rect 40045 2377 40198 2506
rect 40198 2377 40222 2506
rect 40023 2358 40222 2377
rect 41921 2506 42120 2537
rect 41921 2377 41943 2506
rect 41943 2377 42096 2506
rect 42096 2377 42120 2506
rect 41921 2358 42120 2377
rect 58316 9328 58495 9350
rect 58316 9175 58335 9328
rect 58335 9175 58464 9328
rect 58464 9175 58495 9328
rect 58316 9151 58495 9175
rect 59859 9020 60058 9039
rect 59859 8891 59883 9020
rect 59883 8891 60036 9020
rect 60036 8891 60058 9020
rect 59859 8860 60058 8891
rect 61001 9018 61200 9037
rect 61001 8889 61025 9018
rect 61025 8889 61178 9018
rect 61178 8889 61200 9018
rect 61001 8858 61200 8889
rect 58046 8717 58245 8748
rect 58046 8588 58068 8717
rect 58068 8588 58221 8717
rect 58221 8588 58245 8717
rect 58046 8569 58245 8588
rect 59859 8374 60058 8405
rect 59859 8245 59881 8374
rect 59881 8245 60034 8374
rect 60034 8245 60058 8374
rect 59859 8226 60058 8245
rect 61757 8374 61956 8405
rect 61757 8245 61779 8374
rect 61779 8245 61932 8374
rect 61932 8245 61956 8374
rect 61757 8226 61956 8245
rect 63978 8451 64052 8457
rect 63978 8389 63984 8451
rect 63984 8389 64048 8451
rect 64048 8389 64052 8451
rect 65993 8077 66192 8108
rect 65993 7948 66015 8077
rect 66015 7948 66168 8077
rect 66168 7948 66192 8077
rect 65993 7929 66192 7948
rect 58330 7678 58509 7700
rect 58330 7525 58349 7678
rect 58349 7525 58478 7678
rect 58478 7525 58509 7678
rect 67364 7729 67434 7733
rect 67364 7667 67370 7729
rect 67370 7667 67430 7729
rect 67430 7667 67434 7729
rect 67364 7661 67434 7667
rect 58330 7501 58509 7525
rect 58041 7113 58240 7144
rect 58041 6984 58063 7113
rect 58063 6984 58216 7113
rect 58216 6984 58240 7113
rect 58041 6965 58240 6984
rect 63756 6624 63826 6628
rect 63756 6562 63762 6624
rect 63762 6562 63822 6624
rect 63822 6562 63826 6624
rect 63756 6556 63826 6562
rect 67459 6523 67797 6555
rect 67459 6461 67592 6523
rect 67592 6461 67656 6523
rect 67656 6461 67797 6523
rect 67459 6439 67797 6461
rect 58325 6074 58504 6096
rect 58325 5921 58344 6074
rect 58344 5921 58473 6074
rect 58473 5921 58504 6074
rect 58325 5897 58504 5921
rect 59803 5977 60002 5996
rect 59803 5848 59827 5977
rect 59827 5848 59980 5977
rect 59980 5848 60002 5977
rect 59803 5817 60002 5848
rect 61701 5977 61900 5996
rect 61701 5848 61725 5977
rect 61725 5848 61878 5977
rect 61878 5848 61900 5977
rect 61701 5817 61900 5848
rect 65914 5747 66180 5763
rect 65914 5590 65937 5747
rect 65937 5590 66148 5747
rect 66148 5590 66180 5747
rect 65914 5568 66180 5590
rect 63978 5418 64052 5424
rect 63978 5356 63984 5418
rect 63984 5356 64048 5418
rect 64048 5356 64052 5418
rect 44747 4497 44946 4528
rect 44747 4368 44769 4497
rect 44769 4368 44922 4497
rect 44922 4368 44946 4497
rect 44747 4349 44946 4368
rect 47229 4551 47428 4582
rect 47229 4422 47251 4551
rect 47251 4422 47404 4551
rect 47404 4422 47428 4551
rect 47229 4403 47428 4422
rect 48376 4551 48575 4582
rect 48376 4422 48398 4551
rect 48398 4422 48551 4551
rect 48551 4422 48575 4551
rect 48376 4403 48575 4422
rect 45031 3458 45210 3480
rect 45031 3305 45050 3458
rect 45050 3305 45179 3458
rect 45179 3305 45210 3458
rect 45031 3281 45210 3305
rect 46574 3150 46773 3169
rect 46574 3021 46598 3150
rect 46598 3021 46751 3150
rect 46751 3021 46773 3150
rect 46574 2990 46773 3021
rect 47716 3148 47915 3167
rect 47716 3019 47740 3148
rect 47740 3019 47893 3148
rect 47893 3019 47915 3148
rect 47716 2988 47915 3019
rect 44761 2847 44960 2878
rect 44761 2718 44783 2847
rect 44783 2718 44936 2847
rect 44936 2718 44960 2847
rect 44761 2699 44960 2718
rect 46574 2504 46773 2535
rect 46574 2375 46596 2504
rect 46596 2375 46749 2504
rect 46749 2375 46773 2504
rect 46574 2356 46773 2375
rect 48472 2504 48671 2535
rect 48472 2375 48494 2504
rect 48494 2375 48647 2504
rect 48647 2375 48671 2504
rect 48472 2356 48671 2375
rect 38494 1810 38673 1832
rect 38494 1657 38513 1810
rect 38513 1657 38642 1810
rect 38642 1657 38673 1810
rect 45045 1808 45224 1830
rect 38494 1633 38673 1657
rect 45045 1655 45064 1808
rect 45064 1655 45193 1808
rect 45193 1655 45224 1808
rect 63827 4704 63897 4708
rect 63827 4642 63833 4704
rect 63833 4642 63893 4704
rect 63893 4642 63897 4704
rect 63827 4636 63897 4642
rect 51402 4498 51601 4529
rect 51402 4369 51424 4498
rect 51424 4369 51577 4498
rect 51577 4369 51601 4498
rect 51402 4350 51601 4369
rect 53884 4552 54083 4583
rect 53884 4423 53906 4552
rect 53906 4423 54059 4552
rect 54059 4423 54083 4552
rect 53884 4404 54083 4423
rect 55031 4552 55230 4583
rect 55031 4423 55053 4552
rect 55053 4423 55206 4552
rect 55206 4423 55230 4552
rect 55031 4404 55230 4423
rect 58024 4499 58223 4530
rect 58024 4370 58046 4499
rect 58046 4370 58199 4499
rect 58199 4370 58223 4499
rect 58024 4351 58223 4370
rect 60506 4553 60705 4584
rect 60506 4424 60528 4553
rect 60528 4424 60681 4553
rect 60681 4424 60705 4553
rect 60506 4405 60705 4424
rect 61653 4553 61852 4584
rect 61653 4424 61675 4553
rect 61675 4424 61828 4553
rect 61828 4424 61852 4553
rect 61653 4405 61852 4424
rect 65993 4582 66192 4613
rect 65993 4453 66015 4582
rect 66015 4453 66168 4582
rect 66168 4453 66192 4582
rect 65993 4434 66192 4453
rect 67364 4234 67434 4238
rect 67364 4172 67370 4234
rect 67370 4172 67430 4234
rect 67430 4172 67434 4234
rect 67364 4166 67434 4172
rect 51686 3459 51865 3481
rect 51686 3306 51705 3459
rect 51705 3306 51834 3459
rect 51834 3306 51865 3459
rect 51686 3282 51865 3306
rect 58308 3460 58487 3482
rect 58308 3307 58327 3460
rect 58327 3307 58456 3460
rect 58456 3307 58487 3460
rect 58308 3283 58487 3307
rect 53229 3151 53428 3170
rect 53229 3022 53253 3151
rect 53253 3022 53406 3151
rect 53406 3022 53428 3151
rect 53229 2991 53428 3022
rect 54371 3149 54570 3168
rect 54371 3020 54395 3149
rect 54395 3020 54548 3149
rect 54548 3020 54570 3149
rect 54371 2989 54570 3020
rect 59851 3152 60050 3171
rect 59851 3023 59875 3152
rect 59875 3023 60028 3152
rect 60028 3023 60050 3152
rect 59851 2992 60050 3023
rect 60993 3150 61192 3169
rect 60993 3021 61017 3150
rect 61017 3021 61170 3150
rect 61170 3021 61192 3150
rect 60993 2990 61192 3021
rect 51416 2848 51615 2879
rect 51416 2719 51438 2848
rect 51438 2719 51591 2848
rect 51591 2719 51615 2848
rect 51416 2700 51615 2719
rect 58038 2849 58237 2880
rect 58038 2720 58060 2849
rect 58060 2720 58213 2849
rect 58213 2720 58237 2849
rect 58038 2701 58237 2720
rect 53229 2505 53428 2536
rect 53229 2376 53251 2505
rect 53251 2376 53404 2505
rect 53404 2376 53428 2505
rect 53229 2357 53428 2376
rect 55127 2505 55326 2536
rect 55127 2376 55149 2505
rect 55149 2376 55302 2505
rect 55302 2376 55326 2505
rect 55127 2357 55326 2376
rect 59851 2506 60050 2537
rect 59851 2377 59873 2506
rect 59873 2377 60026 2506
rect 60026 2377 60050 2506
rect 59851 2358 60050 2377
rect 61749 2506 61948 2537
rect 61749 2377 61771 2506
rect 61771 2377 61924 2506
rect 61924 2377 61948 2506
rect 61749 2358 61948 2377
rect 51700 1809 51879 1831
rect 45045 1631 45224 1655
rect 51700 1656 51719 1809
rect 51719 1656 51848 1809
rect 51848 1656 51879 1809
rect 51700 1632 51879 1656
rect 58322 1810 58501 1832
rect 58322 1657 58341 1810
rect 58341 1657 58470 1810
rect 58470 1657 58501 1810
rect 58322 1633 58501 1657
rect 38205 1245 38404 1276
rect 38205 1116 38227 1245
rect 38227 1116 38380 1245
rect 38380 1116 38404 1245
rect 38205 1097 38404 1116
rect 44756 1243 44955 1274
rect 44756 1114 44778 1243
rect 44778 1114 44931 1243
rect 44931 1114 44955 1243
rect 44756 1095 44955 1114
rect 51411 1244 51610 1275
rect 51411 1115 51433 1244
rect 51433 1115 51586 1244
rect 51586 1115 51610 1244
rect 51411 1096 51610 1115
rect 58033 1245 58232 1276
rect 58033 1116 58055 1245
rect 58055 1116 58208 1245
rect 58208 1116 58232 1245
rect 58033 1097 58232 1116
rect 35452 646 35526 652
rect 35452 584 35458 646
rect 35458 584 35522 646
rect 35522 584 35526 646
rect 38489 206 38668 228
rect 38489 53 38508 206
rect 38508 53 38637 206
rect 38637 53 38668 206
rect 45040 204 45219 226
rect 38489 29 38668 53
rect 39967 109 40166 128
rect 39967 -20 39991 109
rect 39991 -20 40144 109
rect 40144 -20 40166 109
rect 39967 -51 40166 -20
rect 41865 109 42064 128
rect 41865 -20 41889 109
rect 41889 -20 42042 109
rect 42042 -20 42064 109
rect 41865 -51 42064 -20
rect 45040 51 45059 204
rect 45059 51 45188 204
rect 45188 51 45219 204
rect 51695 205 51874 227
rect 45040 27 45219 51
rect 46518 107 46717 126
rect 46518 -22 46542 107
rect 46542 -22 46695 107
rect 46695 -22 46717 107
rect 46518 -53 46717 -22
rect 48416 107 48615 126
rect 48416 -22 48440 107
rect 48440 -22 48593 107
rect 48593 -22 48615 107
rect 48416 -53 48615 -22
rect 51695 52 51714 205
rect 51714 52 51843 205
rect 51843 52 51874 205
rect 58317 206 58496 228
rect 51695 28 51874 52
rect 53173 108 53372 127
rect 53173 -21 53197 108
rect 53197 -21 53350 108
rect 53350 -21 53372 108
rect 53173 -52 53372 -21
rect 55071 108 55270 127
rect 55071 -21 55095 108
rect 55095 -21 55248 108
rect 55248 -21 55270 108
rect 55071 -52 55270 -21
rect 58317 53 58336 206
rect 58336 53 58465 206
rect 58465 53 58496 206
rect 58317 29 58496 53
rect 59795 109 59994 128
rect 59795 -20 59819 109
rect 59819 -20 59972 109
rect 59972 -20 59994 109
rect 59795 -51 59994 -20
rect 61693 109 61892 128
rect 61693 -20 61717 109
rect 61717 -20 61870 109
rect 61870 -20 61892 109
rect 61693 -51 61892 -20
rect 42162 -775 42168 -713
rect 42168 -775 42232 -713
rect 42232 -775 42236 -713
rect 42162 -781 42236 -775
rect 48716 -770 48722 -708
rect 48722 -770 48786 -708
rect 48786 -770 48790 -708
rect 48716 -776 48790 -770
rect 55365 -782 55371 -720
rect 55371 -782 55435 -720
rect 55435 -782 55439 -720
rect 55365 -788 55439 -782
rect 41940 -1919 42010 -1913
rect 41940 -1981 41946 -1919
rect 41946 -1981 42006 -1919
rect 42006 -1981 42010 -1919
rect 41940 -1985 42010 -1981
rect 48494 -1914 48564 -1908
rect 48494 -1976 48500 -1914
rect 48500 -1976 48560 -1914
rect 48560 -1976 48564 -1914
rect 48494 -1980 48564 -1976
rect 55143 -1926 55213 -1920
rect 55143 -1988 55149 -1926
rect 55149 -1988 55209 -1926
rect 55209 -1988 55213 -1926
rect 55143 -1992 55213 -1988
rect 64049 3498 64123 3504
rect 64049 3436 64055 3498
rect 64055 3436 64119 3498
rect 64119 3436 64123 3498
rect 67459 3028 67797 3060
rect 67459 2966 67592 3028
rect 67592 2966 67656 3028
rect 67656 2966 67797 3028
rect 67459 2944 67797 2966
rect 65914 2252 66180 2268
rect 65914 2095 65937 2252
rect 65937 2095 66148 2252
rect 66148 2095 66180 2252
rect 65914 2073 66180 2095
rect 63824 1634 63894 1638
rect 63824 1572 63830 1634
rect 63830 1572 63890 1634
rect 63890 1572 63894 1634
rect 63824 1566 63894 1572
rect 64046 428 64120 434
rect 64046 366 64052 428
rect 64052 366 64116 428
rect 64116 366 64120 428
rect 65993 234 66192 265
rect 65993 105 66015 234
rect 66015 105 66168 234
rect 66168 105 66192 234
rect 65993 86 66192 105
rect 67364 -114 67434 -110
rect 67364 -176 67370 -114
rect 67370 -176 67430 -114
rect 67430 -176 67434 -114
rect 67364 -182 67434 -176
rect 70239 11305 70329 11405
rect 70329 11305 70331 11405
rect 72481 11385 72549 11391
rect 72481 11309 72539 11385
rect 72539 11309 72549 11385
rect 72481 11307 72549 11309
rect 70243 8103 70333 8203
rect 70333 8103 70335 8203
rect 72485 8183 72553 8189
rect 72485 8107 72543 8183
rect 72543 8107 72553 8183
rect 72485 8105 72553 8107
rect 63831 -1211 63901 -1207
rect 63831 -1273 63837 -1211
rect 63837 -1273 63897 -1211
rect 63897 -1273 63901 -1211
rect 63831 -1279 63901 -1273
rect 67459 -1320 67797 -1288
rect 67459 -1382 67592 -1320
rect 67592 -1382 67656 -1320
rect 67656 -1382 67797 -1320
rect 67459 -1404 67797 -1382
rect 65914 -2096 66180 -2080
rect 65914 -2253 65937 -2096
rect 65937 -2253 66148 -2096
rect 66148 -2253 66180 -2096
rect 65914 -2275 66180 -2253
rect 64053 -2417 64127 -2411
rect 64053 -2479 64059 -2417
rect 64059 -2479 64123 -2417
rect 64123 -2479 64127 -2417
rect 70243 4959 70333 5059
rect 70333 4959 70335 5059
rect 72485 5039 72553 5045
rect 72485 4963 72543 5039
rect 72543 4963 72553 5039
rect 72485 4961 72553 4963
rect 70239 1827 70329 1927
rect 70329 1827 70331 1927
rect 72481 1907 72549 1913
rect 72481 1831 72539 1907
rect 72539 1831 72549 1907
rect 72481 1829 72549 1831
rect 70239 -1317 70329 -1217
rect 70329 -1317 70331 -1217
rect 72481 -1237 72549 -1231
rect 72481 -1313 72539 -1237
rect 72539 -1313 72549 -1237
rect 72481 -1315 72549 -1313
rect 1542 -3782 1548 -3724
rect 1548 -3782 1624 -3724
rect 1624 -3782 1626 -3724
rect 1542 -3792 1626 -3782
rect 4686 -3782 4692 -3724
rect 4692 -3782 4768 -3724
rect 4768 -3782 4770 -3724
rect 4686 -3792 4770 -3782
rect 7818 -3778 7824 -3720
rect 7824 -3778 7900 -3720
rect 7900 -3778 7902 -3720
rect 7818 -3788 7902 -3778
rect 10962 -3778 10968 -3720
rect 10968 -3778 11044 -3720
rect 11044 -3778 11046 -3720
rect 10962 -3788 11046 -3778
rect 14164 -3782 14170 -3724
rect 14170 -3782 14246 -3724
rect 14246 -3782 14248 -3724
rect 14164 -3792 14248 -3782
rect 17308 -3782 17314 -3724
rect 17314 -3782 17390 -3724
rect 17390 -3782 17392 -3724
rect 17308 -3792 17392 -3782
rect 20440 -3778 20446 -3720
rect 20446 -3778 20522 -3720
rect 20522 -3778 20524 -3720
rect 20440 -3788 20524 -3778
rect 23584 -3778 23590 -3720
rect 23590 -3778 23666 -3720
rect 23666 -3778 23668 -3720
rect 23584 -3788 23668 -3778
<< metal4 >>
rect 1700 25190 70358 26422
rect 1700 25052 70369 25190
rect 24031 24915 70369 25052
rect 24031 24861 42490 24915
rect 24031 24682 40008 24861
rect 40207 24736 42490 24861
rect 42689 24736 43637 24915
rect 43836 24912 70369 24915
rect 43836 24858 49003 24912
rect 43836 24736 46521 24858
rect 40207 24682 46521 24736
rect 24031 24679 46521 24682
rect 46720 24733 49003 24858
rect 49202 24733 50150 24912
rect 50349 24911 70369 24912
rect 50349 24907 62095 24911
rect 50349 24853 55537 24907
rect 50349 24733 53055 24853
rect 46720 24679 53055 24733
rect 24031 24674 53055 24679
rect 53254 24728 55537 24853
rect 55736 24728 56684 24907
rect 56883 24857 62095 24907
rect 56883 24728 59613 24857
rect 53254 24678 59613 24728
rect 59812 24732 62095 24857
rect 62294 24732 63242 24911
rect 63441 24732 70369 24911
rect 59812 24678 70369 24732
rect 53254 24674 70369 24678
rect 24031 24477 70369 24674
rect 24031 24476 38546 24477
rect 24031 24458 38298 24476
rect 39142 24472 70369 24477
rect 24031 22372 27295 24458
rect 28199 24453 29654 24458
rect 3340 22266 27295 22372
rect 3340 22174 4272 22266
rect 4372 22174 7416 22266
rect 7516 22262 16894 22266
rect 7516 22174 10548 22262
rect 3340 22170 10548 22174
rect 10648 22170 13692 22262
rect 13792 22174 16894 22262
rect 16994 22174 20038 22266
rect 20138 22262 27295 22266
rect 20138 22174 23170 22262
rect 13792 22170 23170 22174
rect 23270 22170 26314 22262
rect 26414 22170 27295 22262
rect 3340 22138 27295 22170
rect 24031 22120 27295 22138
rect 27726 21183 27814 21184
rect 27726 21100 27727 21183
rect 27804 21100 27814 21183
rect 5662 21034 5783 21035
rect 5662 20925 5673 21034
rect 5773 20925 5783 21034
rect 3916 19852 3962 20032
rect 5662 20032 5783 20925
rect 4736 19852 7095 20032
rect 7869 19852 10151 20032
rect 10925 19852 13267 20032
rect 14041 19852 16526 20032
rect 17300 19852 19675 20032
rect 20449 19852 22797 20032
rect 23571 19852 25990 20032
rect 26764 20031 27290 20032
rect 27726 20031 27814 21100
rect 26764 19852 27814 20031
rect 4500 17060 14277 17126
rect 4500 17034 12790 17060
rect 4500 16970 4632 17034
rect 4696 16970 5800 17034
rect 5864 17032 8136 17034
rect 5864 16970 6968 17032
rect 4500 16968 6968 16970
rect 7032 16970 8136 17032
rect 8200 16970 9308 17034
rect 9372 17032 12790 17034
rect 9372 16970 10478 17032
rect 7032 16968 10478 16970
rect 10542 16968 11646 17032
rect 11710 16968 12790 17032
rect 4500 16940 12790 16968
rect 12912 16940 14277 17060
rect 4500 16930 14277 16940
rect 13421 16899 14277 16930
rect 28853 16929 29654 24453
rect 25064 16899 29654 16929
rect 13421 16843 29654 16899
rect 13421 16771 14494 16843
rect 14564 16771 15942 16843
rect 16012 16841 20408 16843
rect 16012 16771 17440 16841
rect 13421 16769 17440 16771
rect 17510 16769 18888 16841
rect 18958 16771 20408 16841
rect 20478 16771 21856 16843
rect 21926 16841 29654 16843
rect 21926 16771 23354 16841
rect 18958 16769 23354 16771
rect 23424 16769 24802 16841
rect 24872 16769 29654 16841
rect 13421 16742 29654 16769
rect 14094 16741 29654 16742
rect 25017 16363 29654 16741
rect 36128 19573 37642 24458
rect 39142 23425 39994 24472
rect 39142 23211 40362 23425
rect 39142 23032 40022 23211
rect 40221 23043 40362 23211
rect 40221 23038 40707 23043
rect 42585 23038 42932 23041
rect 43799 23038 44415 24472
rect 40221 23032 44415 23038
rect 39142 22868 44415 23032
rect 39142 22689 41835 22868
rect 42034 22689 43733 22868
rect 43932 22689 44415 22868
rect 39142 22533 44415 22689
rect 39142 21803 39994 22533
rect 43799 22528 44415 22533
rect 45980 23208 46875 23422
rect 45980 23029 46535 23208
rect 46734 23040 46875 23208
rect 46734 23035 47220 23040
rect 49098 23035 49445 23038
rect 50312 23035 50928 24472
rect 53034 24468 57462 24472
rect 46734 23029 50928 23035
rect 45980 22865 50928 23029
rect 45980 22686 48348 22865
rect 48547 22686 50246 22865
rect 50445 22686 50928 22865
rect 45980 22530 50928 22686
rect 39142 21607 40735 21803
rect 39142 21428 40017 21607
rect 40216 21428 40735 21607
rect 39142 21159 40735 21428
rect 45980 21800 46150 22530
rect 50312 22525 50928 22530
rect 52514 23203 53409 23417
rect 52514 23024 53069 23203
rect 53268 23035 53409 23203
rect 53268 23030 53754 23035
rect 55632 23030 55979 23033
rect 56846 23030 57462 24468
rect 53268 23024 57462 23030
rect 52514 22860 57462 23024
rect 52514 22681 54882 22860
rect 55081 22681 56780 22860
rect 56979 22681 57462 22860
rect 52514 22525 57462 22681
rect 45980 21604 47248 21800
rect 45980 21425 46530 21604
rect 46729 21425 47248 21604
rect 39142 19872 39994 21159
rect 45980 21156 47248 21425
rect 52514 21795 52684 22525
rect 56846 22520 57462 22525
rect 59072 23207 59967 23421
rect 59072 23028 59627 23207
rect 59826 23039 59967 23207
rect 59826 23034 60312 23039
rect 62190 23034 62537 23037
rect 63404 23034 70369 24472
rect 59826 23028 70369 23034
rect 59072 22948 70369 23028
rect 59072 22864 64020 22948
rect 59072 22685 61440 22864
rect 61639 22685 63338 22864
rect 63537 22685 64020 22864
rect 59072 22529 64020 22685
rect 59072 21799 59242 22529
rect 63404 22524 64020 22529
rect 52514 21599 53782 21795
rect 52514 21420 53064 21599
rect 53263 21420 53782 21599
rect 52514 21151 53782 21420
rect 59072 21603 60340 21799
rect 68378 21681 70369 22948
rect 59072 21424 59622 21603
rect 59821 21424 60340 21603
rect 59072 21155 60340 21424
rect 68370 21520 70369 21681
rect 68370 20825 70367 21520
rect 68370 20725 70243 20825
rect 70335 20725 70367 20825
rect 41755 20459 42000 20462
rect 41755 20441 41779 20459
rect 41978 20441 42000 20459
rect 43653 20459 43898 20462
rect 43653 20441 43677 20459
rect 43876 20441 43898 20459
rect 41651 20137 41675 20374
rect 42185 20137 43521 20323
rect 48268 20456 48513 20459
rect 48268 20438 48292 20456
rect 48491 20438 48513 20456
rect 50166 20456 50411 20459
rect 50166 20438 50190 20456
rect 50389 20438 50411 20456
rect 41651 20132 44018 20137
rect 48164 20134 48188 20371
rect 48698 20134 50034 20320
rect 54802 20451 55047 20454
rect 54802 20433 54826 20451
rect 55025 20433 55047 20451
rect 56700 20451 56945 20454
rect 56700 20433 56724 20451
rect 56923 20433 56945 20451
rect 42039 20130 43710 20132
rect 48164 20129 50531 20134
rect 54698 20129 54722 20366
rect 55232 20129 56568 20315
rect 61360 20455 61605 20458
rect 61360 20437 61384 20455
rect 61583 20437 61605 20455
rect 63258 20455 63503 20458
rect 63258 20437 63282 20455
rect 63481 20437 63503 20455
rect 61256 20133 61280 20370
rect 61790 20133 63126 20319
rect 48552 20127 50223 20129
rect 54698 20124 57065 20129
rect 61256 20128 63623 20133
rect 61644 20126 63315 20128
rect 55086 20122 56757 20124
rect 39138 19578 39995 19872
rect 63031 19603 63883 19608
rect 68370 19603 70367 20725
rect 72473 20552 72653 20585
rect 63031 19596 70367 19603
rect 42195 19578 70367 19596
rect 39134 19573 70367 19578
rect 36128 19311 70367 19573
rect 36128 19308 59189 19311
rect 36128 19307 52676 19308
rect 36128 19128 39584 19307
rect 39783 19128 40731 19307
rect 40930 19303 52676 19307
rect 40930 19253 46142 19303
rect 40930 19128 43213 19253
rect 36128 19074 43213 19128
rect 43412 19124 46142 19253
rect 46341 19124 47289 19303
rect 47488 19249 52676 19303
rect 47488 19124 49771 19249
rect 43412 19074 49771 19124
rect 36128 19070 49771 19074
rect 49970 19129 52676 19249
rect 52875 19129 53823 19308
rect 54022 19254 59189 19308
rect 54022 19129 56305 19254
rect 49970 19075 56305 19129
rect 56504 19132 59189 19254
rect 59388 19132 60336 19311
rect 60535 19257 70367 19311
rect 60535 19132 62818 19257
rect 56504 19078 62818 19132
rect 63017 19078 70367 19257
rect 56504 19075 70367 19078
rect 49970 19070 70367 19075
rect 36128 18868 70367 19070
rect 36128 18858 39621 18868
rect 36128 16363 37642 18858
rect 39134 17430 39621 18858
rect 42195 18856 70367 18868
rect 42677 18276 43187 18283
rect 43058 17603 43953 17817
rect 43058 17435 43199 17603
rect 40488 17430 40835 17433
rect 42713 17430 43199 17435
rect 39134 17424 43199 17430
rect 43398 17424 43953 17603
rect 39134 17260 43953 17424
rect 39134 17081 39488 17260
rect 39687 17081 41386 17260
rect 41585 17081 43953 17260
rect 39134 16925 43953 17081
rect 39134 16920 39621 16925
rect 838 15231 24768 15234
rect 25017 15231 37642 16363
rect 43783 16195 43953 16925
rect 45563 17426 46179 18856
rect 49616 17599 50511 17813
rect 49616 17431 49757 17599
rect 47046 17426 47393 17429
rect 49271 17426 49757 17431
rect 45563 17420 49757 17426
rect 49956 17420 50511 17599
rect 45563 17256 50511 17420
rect 45563 17077 46046 17256
rect 46245 17077 47944 17256
rect 48143 17077 50511 17256
rect 45563 16921 50511 17077
rect 52097 17431 52713 18856
rect 56150 17604 57045 17818
rect 56150 17436 56291 17604
rect 53580 17431 53927 17434
rect 55805 17431 56291 17436
rect 52097 17425 56291 17431
rect 56490 17425 57045 17604
rect 52097 17261 57045 17425
rect 52097 17082 52580 17261
rect 52779 17082 54478 17261
rect 54677 17082 57045 17261
rect 52097 16926 57045 17082
rect 52097 16921 52713 16926
rect 45563 16916 46179 16921
rect 42685 15999 43953 16195
rect 50341 16191 50511 16921
rect 56875 16196 57045 16926
rect 58610 17434 59226 18856
rect 63031 18823 70367 18856
rect 63806 18821 70367 18823
rect 62663 17607 63558 17821
rect 62663 17439 62804 17607
rect 60093 17434 60440 17437
rect 62318 17434 62804 17439
rect 58610 17428 62804 17434
rect 63003 17428 63558 17607
rect 58610 17264 63558 17428
rect 58610 17085 59093 17264
rect 59292 17085 60991 17264
rect 61190 17085 63558 17264
rect 58610 16929 63558 17085
rect 58610 16924 59226 16929
rect 63388 16199 63558 16929
rect 42685 15820 43204 15999
rect 43403 15820 43953 15999
rect 42685 15551 43953 15820
rect 49243 15995 50511 16191
rect 49243 15816 49762 15995
rect 49961 15816 50511 15995
rect 49243 15547 50511 15816
rect 55777 16000 57045 16196
rect 55777 15821 56296 16000
rect 56495 15821 57045 16000
rect 55777 15552 57045 15821
rect 62290 16003 63558 16199
rect 62290 15824 62809 16003
rect 63008 15824 63558 16003
rect 62290 15555 63558 15824
rect 68370 17681 70367 18821
rect 72473 17758 72653 17821
rect 68370 17581 70243 17681
rect 70335 17581 70367 17681
rect 838 15128 37642 15231
rect 838 15036 1770 15128
rect 1870 15036 4914 15128
rect 5014 15124 14392 15128
rect 5014 15036 8046 15124
rect 838 15032 8046 15036
rect 8146 15032 11190 15124
rect 11290 15036 14392 15124
rect 14492 15036 17536 15128
rect 17636 15124 37642 15128
rect 17636 15036 20668 15124
rect 11290 15032 20668 15036
rect 20768 15032 23812 15124
rect 23912 15032 37642 15124
rect 838 15000 37642 15032
rect 24657 14998 37642 15000
rect 25058 13888 37642 14998
rect 39522 14851 39767 14854
rect 39522 14833 39544 14851
rect 39743 14833 39767 14851
rect 41420 14851 41665 14854
rect 41420 14833 41442 14851
rect 41641 14833 41665 14851
rect 39899 14529 41235 14715
rect 41745 14529 41769 14766
rect 46080 14847 46325 14850
rect 46080 14829 46102 14847
rect 46301 14829 46325 14847
rect 47978 14847 48223 14850
rect 47978 14829 48000 14847
rect 48199 14829 48223 14847
rect 39402 14524 41769 14529
rect 46457 14525 47793 14711
rect 48303 14525 48327 14762
rect 52614 14852 52859 14855
rect 52614 14834 52636 14852
rect 52835 14834 52859 14852
rect 54512 14852 54757 14855
rect 54512 14834 54534 14852
rect 54733 14834 54757 14852
rect 52991 14530 54327 14716
rect 54837 14530 54861 14767
rect 59127 14855 59372 14858
rect 59127 14837 59149 14855
rect 59348 14837 59372 14855
rect 61025 14855 61270 14858
rect 61025 14837 61047 14855
rect 61246 14837 61270 14855
rect 59504 14533 60840 14719
rect 61350 14533 61374 14770
rect 52494 14525 54861 14530
rect 59007 14528 61374 14533
rect 68370 14549 70367 17581
rect 72473 17372 72653 17427
rect 72473 14625 72653 14688
rect 59315 14526 60986 14528
rect 39710 14522 41381 14524
rect 45960 14520 48327 14525
rect 52802 14523 54473 14525
rect 46268 14518 47939 14520
rect 25058 13036 30031 13888
rect 838 12498 24768 12500
rect 25058 12498 29801 13036
rect 838 12394 29801 12498
rect 838 12302 1770 12394
rect 1870 12302 4914 12394
rect 5014 12390 14392 12394
rect 5014 12302 8046 12390
rect 838 12298 8046 12302
rect 8146 12298 11190 12390
rect 11290 12302 14392 12390
rect 14492 12302 17536 12394
rect 17636 12390 29801 12394
rect 17636 12302 20668 12390
rect 11290 12298 20668 12302
rect 20768 12298 23812 12390
rect 23912 12353 29801 12390
rect 23912 12298 29693 12353
rect 838 12277 29693 12298
rect 29759 12277 29801 12353
rect 838 12266 29801 12277
rect 24547 12263 29801 12266
rect 25058 10285 29801 12263
rect 36128 12560 37642 13888
rect 68370 14449 70239 14549
rect 70331 14449 70367 14549
rect 68370 12568 70367 14449
rect 72473 14284 72653 14294
rect 66442 12567 70367 12568
rect 63039 12566 70367 12567
rect 36121 12559 41773 12560
rect 48172 12559 70367 12566
rect 36121 12399 70367 12559
rect 36121 12379 55108 12399
rect 36121 12307 41905 12379
rect 41975 12378 55108 12379
rect 41975 12307 48454 12378
rect 36121 12306 48454 12307
rect 48524 12327 55108 12378
rect 55178 12327 70367 12399
rect 48524 12306 70367 12327
rect 36121 12268 70367 12306
rect 36121 12261 56673 12268
rect 36121 12260 41773 12261
rect 31909 12158 32099 12194
rect 36121 10639 36527 12260
rect 62826 12232 70367 12268
rect 62826 12160 63761 12232
rect 63831 12199 70367 12232
rect 63831 12160 65991 12199
rect 62826 12108 65991 12160
rect 42439 11074 42440 11282
rect 48471 11258 48981 11259
rect 48471 11077 48472 11258
rect 55138 11066 55139 11242
rect 42434 10640 45991 10672
rect 48747 10645 52304 10672
rect 55582 10645 59139 10672
rect 62826 10652 63293 12108
rect 65849 12105 65991 12108
rect 65969 12020 65991 12105
rect 66190 12106 70367 12199
rect 66190 12105 66318 12106
rect 66190 12020 66214 12105
rect 65969 12017 66214 12020
rect 67202 11824 67588 12106
rect 67202 11783 67362 11824
rect 67204 11752 67362 11783
rect 67432 11783 67588 11824
rect 67432 11752 67586 11783
rect 67204 11730 67586 11752
rect 67931 11405 70367 12106
rect 67931 11305 70239 11405
rect 70331 11305 70367 11405
rect 64200 10898 64201 11069
rect 62201 10645 63293 10652
rect 67456 10647 67512 10648
rect 48747 10640 63293 10645
rect 35005 10635 39162 10639
rect 42434 10635 63293 10640
rect 31907 10502 32099 10508
rect 25058 10209 29691 10285
rect 29757 10209 29801 10285
rect 25058 9775 29801 10209
rect 35005 10479 63293 10635
rect 35005 10407 35241 10479
rect 35311 10452 63293 10479
rect 35311 10407 47235 10452
rect 35005 10398 47235 10407
rect 35005 10385 44753 10398
rect 36126 10364 44753 10385
rect 36126 10310 40686 10364
rect 36126 10131 38204 10310
rect 38403 10185 40686 10310
rect 40885 10185 41833 10364
rect 42032 10219 44753 10364
rect 44952 10273 47235 10398
rect 47434 10273 48382 10452
rect 48581 10398 60514 10452
rect 48581 10384 58032 10398
rect 48581 10330 53889 10384
rect 48581 10273 51407 10330
rect 44952 10219 51407 10273
rect 42032 10185 51407 10219
rect 38403 10151 51407 10185
rect 51606 10205 53889 10330
rect 54088 10205 55036 10384
rect 55235 10219 58032 10384
rect 58231 10273 60514 10398
rect 60713 10273 61661 10452
rect 61860 10273 63293 10452
rect 67452 10646 67512 10647
rect 67749 10647 67788 10648
rect 67749 10646 67803 10647
rect 67452 10530 67457 10646
rect 67795 10530 67803 10646
rect 67452 10389 67512 10530
rect 58231 10219 63293 10273
rect 67749 10389 67803 10530
rect 55235 10205 63293 10219
rect 51606 10151 63293 10205
rect 38403 10131 63293 10151
rect 31907 10018 32099 10100
rect 24583 9768 29801 9775
rect 848 9662 29801 9768
rect 848 9570 1780 9662
rect 1880 9570 4924 9662
rect 5024 9658 14402 9662
rect 5024 9570 8056 9658
rect 848 9566 8056 9570
rect 8156 9566 11200 9658
rect 11300 9570 14402 9658
rect 14502 9570 17546 9662
rect 17646 9658 29801 9662
rect 17646 9570 20678 9658
rect 11300 9566 20678 9570
rect 20778 9566 23822 9658
rect 23922 9566 29801 9658
rect 848 9540 29801 9566
rect 848 9534 24778 9540
rect 25058 8216 29801 9540
rect 36126 10013 63293 10131
rect 36126 10012 45991 10013
rect 48544 10012 59139 10013
rect 36126 9925 42611 10012
rect 36126 9910 40020 9925
rect 31909 8434 32099 8466
rect 25058 8140 29693 8216
rect 29759 8140 29801 8216
rect 8674 6851 9432 6852
rect 3077 6840 9432 6851
rect 25058 6840 29801 8140
rect 36126 8041 36804 9910
rect 31909 8001 32099 8032
rect 34992 7894 36804 8041
rect 34992 7822 35233 7894
rect 35303 7822 36804 7894
rect 34992 7800 36804 7822
rect 3077 6777 29801 6840
rect 3077 6775 8437 6777
rect 3077 6667 3265 6775
rect 3375 6667 4003 6775
rect 4113 6667 4741 6775
rect 4851 6667 5479 6775
rect 5589 6667 6219 6775
rect 6329 6667 6961 6775
rect 7071 6667 7699 6775
rect 7809 6669 8437 6775
rect 8547 6708 29801 6777
rect 8547 6669 10051 6708
rect 7809 6667 10051 6669
rect 3077 6661 10051 6667
rect 8674 6642 10051 6661
rect 10127 6706 14188 6708
rect 10127 6642 12119 6706
rect 8674 6640 12119 6642
rect 12195 6642 14188 6706
rect 14264 6706 29801 6708
rect 14264 6642 16256 6706
rect 12195 6640 16256 6642
rect 16332 6640 18325 6706
rect 18401 6704 22462 6706
rect 18401 6640 20393 6704
rect 8674 6638 20393 6640
rect 20469 6640 22462 6704
rect 22538 6704 29801 6706
rect 22538 6640 24530 6704
rect 20469 6638 24530 6640
rect 24606 6648 29801 6704
rect 24606 6638 25450 6648
rect 8674 6596 25450 6638
rect 8674 6594 9432 6596
rect 25058 6587 25346 6596
rect 28853 6148 29801 6648
rect 31907 6371 32099 6485
rect 28853 6072 29691 6148
rect 29757 6072 29801 6148
rect 3261 5751 3274 5941
rect 3510 5751 3523 5941
rect 3999 5751 4001 5941
rect 4237 5751 4260 5941
rect 4736 5751 4747 5941
rect 4983 5751 4997 5941
rect 5473 5751 5486 5941
rect 5722 5751 5735 5941
rect 6214 5751 6217 5941
rect 6453 5751 6475 5941
rect 6957 5751 6958 5941
rect 7194 5751 7217 5941
rect 7693 5751 7706 5941
rect 7942 5751 7955 5941
rect 8433 5751 8440 5941
rect 8676 5751 8694 5941
rect 10011 4298 10020 4492
rect 10256 4298 10266 4492
rect 12080 4298 12093 4490
rect 12329 4298 12334 4490
rect 14148 4298 14156 4492
rect 14392 4298 14404 4492
rect 16218 4298 16220 4490
rect 16456 4298 16471 4490
rect 18285 4298 18293 4490
rect 18529 4298 18539 4490
rect 20353 4298 20361 4488
rect 20597 4298 20608 4488
rect 22424 4298 22434 4490
rect 22670 4298 22676 4490
rect 24491 4298 24501 4488
rect 24737 4298 24743 4488
rect 28853 4079 29801 6072
rect 31907 5923 32099 5969
rect 36126 4786 36804 7800
rect 37663 8660 38558 8874
rect 37663 8481 38218 8660
rect 38417 8492 38558 8660
rect 38417 8487 38903 8492
rect 40781 8487 41128 8490
rect 41995 8487 42611 9925
rect 38417 8481 42611 8487
rect 37663 8317 42611 8481
rect 37663 8138 40031 8317
rect 40230 8138 41929 8317
rect 42128 8138 42611 8317
rect 37663 7982 42611 8138
rect 37663 7252 37833 7982
rect 41995 7977 42611 7982
rect 44212 8748 45107 8962
rect 44212 8569 44767 8748
rect 44966 8580 45107 8748
rect 44966 8575 45452 8580
rect 47330 8575 47677 8578
rect 48544 8575 49160 10012
rect 51386 9945 55814 10012
rect 44966 8569 49160 8575
rect 44212 8405 49160 8569
rect 44212 8226 46580 8405
rect 46779 8226 48478 8405
rect 48677 8226 49160 8405
rect 44212 8070 49160 8226
rect 44212 7340 44382 8070
rect 48544 8065 49160 8070
rect 50866 8680 51761 8894
rect 50866 8501 51421 8680
rect 51620 8512 51761 8680
rect 51620 8507 52106 8512
rect 53984 8507 54331 8510
rect 55198 8507 55814 9945
rect 61823 9990 63293 10013
rect 51620 8501 55814 8507
rect 50866 8337 55814 8501
rect 50866 8158 53234 8337
rect 53433 8158 55132 8337
rect 55331 8158 55814 8337
rect 50866 8002 55814 8158
rect 37663 7056 38931 7252
rect 37663 6877 38213 7056
rect 38412 6877 38931 7056
rect 37663 6608 38931 6877
rect 44212 7144 45480 7340
rect 44212 6965 44762 7144
rect 44961 6965 45480 7144
rect 44212 6696 45480 6965
rect 50866 7272 51036 8002
rect 55198 7997 55814 8002
rect 57491 8748 58386 8962
rect 57491 8569 58046 8748
rect 58245 8580 58386 8748
rect 58245 8575 58731 8580
rect 60609 8575 60956 8578
rect 61823 8575 62439 9990
rect 58245 8569 62439 8575
rect 57491 8405 62439 8569
rect 57491 8226 59859 8405
rect 60058 8226 61757 8405
rect 61956 8226 62439 8405
rect 57491 8070 62439 8226
rect 57491 7340 57661 8070
rect 61823 8065 62439 8070
rect 62826 9759 63293 9990
rect 62826 9661 64308 9759
rect 62826 9589 63756 9661
rect 63826 9589 64308 9661
rect 62826 9521 64308 9589
rect 50866 7076 52134 7272
rect 50866 6897 51416 7076
rect 51615 6897 52134 7076
rect 50866 6628 52134 6897
rect 57491 7144 58759 7340
rect 57491 6965 58041 7144
rect 58240 6965 58759 7144
rect 57491 6696 58759 6965
rect 62826 6743 63293 9521
rect 63846 8506 64205 8508
rect 65734 8273 67087 8284
rect 67931 8273 70367 11305
rect 72473 11156 72653 11176
rect 72473 8316 72653 8349
rect 65734 8203 70367 8273
rect 65734 8108 70243 8203
rect 65734 8014 65993 8108
rect 65971 7929 65993 8014
rect 66192 8103 70243 8108
rect 70335 8103 70367 8203
rect 66192 8014 70367 8103
rect 66192 7929 66216 8014
rect 66889 8012 70367 8014
rect 65971 7926 66216 7929
rect 67204 7733 67590 8012
rect 67204 7692 67364 7733
rect 67206 7661 67364 7692
rect 67434 7692 67590 7733
rect 67434 7661 67588 7692
rect 67206 7639 67588 7661
rect 62826 6628 64311 6743
rect 62826 6556 63756 6628
rect 63826 6556 64311 6628
rect 67458 6556 67514 6557
rect 62826 6505 64311 6556
rect 67454 6555 67514 6556
rect 67751 6556 67790 6557
rect 67751 6555 67805 6556
rect 39951 5908 40196 5911
rect 39951 5890 39975 5908
rect 40174 5890 40196 5908
rect 41849 5908 42094 5911
rect 41849 5890 41873 5908
rect 42072 5890 42094 5908
rect 46500 5996 46745 5999
rect 46500 5978 46524 5996
rect 46723 5978 46745 5996
rect 48398 5996 48643 5999
rect 48398 5978 48422 5996
rect 48621 5978 48643 5996
rect 39847 5586 39871 5823
rect 40381 5586 41717 5772
rect 46396 5674 46420 5911
rect 46930 5674 48266 5860
rect 53154 5928 53399 5931
rect 53154 5910 53178 5928
rect 53377 5910 53399 5928
rect 55052 5928 55297 5931
rect 55052 5910 55076 5928
rect 55275 5910 55297 5928
rect 46396 5669 48763 5674
rect 46784 5667 48455 5669
rect 53050 5606 53074 5843
rect 53584 5606 54920 5792
rect 59779 5996 60024 5999
rect 59779 5978 59803 5996
rect 60002 5978 60024 5996
rect 61677 5996 61922 5999
rect 61677 5978 61701 5996
rect 61900 5978 61922 5996
rect 59675 5674 59699 5911
rect 60209 5674 61545 5860
rect 59675 5669 62042 5674
rect 60063 5667 61734 5669
rect 53050 5601 55417 5606
rect 53438 5599 55109 5601
rect 39847 5581 42214 5586
rect 40235 5579 41906 5581
rect 62826 5048 63293 6505
rect 67454 6439 67459 6555
rect 67797 6439 67805 6555
rect 67454 6298 67514 6439
rect 67751 6298 67805 6439
rect 63847 5468 64208 5470
rect 63846 5313 63847 5468
rect 64207 5310 64208 5468
rect 67931 5059 70367 8012
rect 72473 7980 72653 7985
rect 72473 5150 72653 5168
rect 67931 5051 70243 5059
rect 67112 5048 70243 5051
rect 62826 4959 70243 5048
rect 70335 4959 70367 5059
rect 44725 4786 49158 4792
rect 51380 4786 55813 4800
rect 58002 4786 62435 4802
rect 62826 4786 70367 4959
rect 36126 4745 70367 4786
rect 34985 4708 70367 4745
rect 34985 4636 63827 4708
rect 63897 4636 70367 4708
rect 34985 4616 70367 4636
rect 34985 4544 35214 4616
rect 35284 4613 70367 4616
rect 35284 4584 65993 4613
rect 35284 4544 40678 4584
rect 34985 4530 40678 4544
rect 34985 4504 38196 4530
rect 36126 4351 38196 4504
rect 38395 4405 40678 4530
rect 40877 4405 41825 4584
rect 42024 4583 60506 4584
rect 42024 4582 53884 4583
rect 42024 4528 47229 4582
rect 42024 4405 44747 4528
rect 38395 4351 44747 4405
rect 36126 4349 44747 4351
rect 44946 4403 47229 4528
rect 47428 4403 48376 4582
rect 48575 4529 53884 4582
rect 48575 4403 51402 4529
rect 44946 4350 51402 4403
rect 51601 4404 53884 4529
rect 54083 4404 55031 4583
rect 55230 4530 60506 4583
rect 55230 4404 58024 4530
rect 51601 4351 58024 4404
rect 58223 4405 60506 4530
rect 60705 4405 61653 4584
rect 61852 4511 65993 4584
rect 61852 4405 63293 4511
rect 65971 4434 65993 4511
rect 66192 4511 70367 4613
rect 66192 4434 66216 4511
rect 67112 4506 70367 4511
rect 65971 4431 66216 4434
rect 58223 4351 63293 4405
rect 51601 4350 63293 4351
rect 44946 4349 63293 4350
rect 31907 4272 32099 4324
rect 28853 4003 29691 4079
rect 29757 4003 29801 4079
rect 28853 2945 29801 4003
rect 36126 4123 63293 4349
rect 67204 4238 67590 4506
rect 67204 4197 67364 4238
rect 67206 4166 67364 4197
rect 67434 4197 67590 4238
rect 67434 4166 67588 4197
rect 67206 4144 67588 4166
rect 31907 3819 32099 3870
rect 708 2520 29801 2945
rect 640 2414 29801 2520
rect 640 2410 7772 2414
rect 640 2318 1496 2410
rect 1596 2318 4640 2410
rect 4740 2322 7772 2410
rect 7872 2322 10916 2414
rect 11016 2410 20394 2414
rect 11016 2322 14118 2410
rect 4740 2318 14118 2322
rect 14218 2318 17262 2410
rect 17362 2322 20394 2410
rect 20494 2322 23538 2414
rect 23638 2322 29801 2414
rect 17362 2318 29801 2322
rect 640 2286 29801 2318
rect 21341 2232 29801 2286
rect 28853 2011 29801 2232
rect 31905 2209 32099 2297
rect 28853 1935 29689 2011
rect 29755 1935 29801 2011
rect 1130 0 1239 180
rect 1875 0 1940 180
rect 4315 0 4439 180
rect 5075 0 5090 180
rect 7465 0 7565 180
rect 10566 0 10640 180
rect 11276 0 11396 180
rect 13771 0 13830 180
rect 14466 0 14581 180
rect 16956 0 17055 180
rect 17691 0 17796 180
rect 20171 0 20176 180
rect 20812 0 20842 180
rect 23217 0 23263 180
rect 23899 0 23994 180
rect 28853 -58 29801 1935
rect 36126 1988 36804 4123
rect 34979 1856 36804 1988
rect 31905 1683 32099 1807
rect 34979 1784 35230 1856
rect 35300 1784 36804 1856
rect 34979 1747 36804 1784
rect 31907 167 32099 198
rect 28853 -134 29691 -58
rect 29757 -134 29801 -58
rect 708 -847 23929 -824
rect 28853 -847 29801 -134
rect 31907 -369 32099 -235
rect 708 -1372 29801 -847
rect 672 -1478 29801 -1372
rect 672 -1482 7804 -1478
rect 672 -1574 1528 -1482
rect 1628 -1574 4672 -1482
rect 4772 -1570 7804 -1482
rect 7904 -1570 10948 -1478
rect 11048 -1482 20426 -1478
rect 11048 -1570 14150 -1482
rect 4772 -1574 14150 -1570
rect 14250 -1574 17294 -1482
rect 17394 -1570 20426 -1482
rect 20526 -1570 23570 -1478
rect 23670 -1570 29801 -1478
rect 17394 -1574 29801 -1570
rect 672 -1606 29801 -1574
rect 22590 -1672 29801 -1606
rect 28853 -2126 29801 -1672
rect 36126 -1868 36804 1747
rect 37655 2880 38550 3094
rect 37655 2701 38210 2880
rect 38409 2712 38550 2880
rect 38409 2707 38895 2712
rect 40773 2707 41120 2710
rect 41987 2707 42603 4123
rect 38409 2701 42603 2707
rect 37655 2537 42603 2701
rect 37655 2358 40023 2537
rect 40222 2358 41921 2537
rect 42120 2358 42603 2537
rect 37655 2202 42603 2358
rect 37655 1472 37825 2202
rect 41987 2197 42603 2202
rect 44206 2878 45101 3092
rect 44206 2699 44761 2878
rect 44960 2710 45101 2878
rect 44960 2705 45446 2710
rect 47324 2705 47671 2708
rect 48538 2705 49154 4123
rect 44960 2699 49154 2705
rect 44206 2535 49154 2699
rect 44206 2356 46574 2535
rect 46773 2356 48472 2535
rect 48671 2356 49154 2535
rect 44206 2200 49154 2356
rect 37655 1276 38923 1472
rect 37655 1097 38205 1276
rect 38404 1097 38923 1276
rect 37655 828 38923 1097
rect 44206 1470 44376 2200
rect 48538 2195 49154 2200
rect 50861 2879 51756 3093
rect 50861 2700 51416 2879
rect 51615 2711 51756 2879
rect 51615 2706 52101 2711
rect 53979 2706 54326 2709
rect 55193 2706 55809 4123
rect 51615 2700 55809 2706
rect 50861 2536 55809 2700
rect 50861 2357 53229 2536
rect 53428 2357 55127 2536
rect 55326 2357 55809 2536
rect 50861 2201 55809 2357
rect 50861 1471 51031 2201
rect 55193 2196 55809 2201
rect 57483 2880 58378 3094
rect 57483 2701 58038 2880
rect 58237 2712 58378 2880
rect 58237 2707 58723 2712
rect 60601 2707 60948 2710
rect 61815 2707 62431 4123
rect 58237 2701 62431 2707
rect 57483 2537 62431 2701
rect 57483 2358 59851 2537
rect 60050 2358 61749 2537
rect 61948 2358 62431 2537
rect 57483 2202 62431 2358
rect 57483 1472 57653 2202
rect 61815 2197 62431 2202
rect 62826 1731 63293 4123
rect 63907 3547 64270 3548
rect 64267 3387 64270 3547
rect 67458 3061 67514 3062
rect 67454 3060 67514 3061
rect 67751 3061 67790 3062
rect 67751 3060 67805 3061
rect 67454 2944 67459 3060
rect 67797 2944 67805 3060
rect 67454 2803 67514 2944
rect 67751 2803 67805 2944
rect 65851 1931 66224 2001
rect 67931 1927 70367 4506
rect 72473 2007 72653 2050
rect 67931 1827 70239 1927
rect 70331 1827 70367 1927
rect 62826 1638 64311 1731
rect 62826 1566 63824 1638
rect 63894 1566 64311 1638
rect 62826 1493 64311 1566
rect 44206 1274 45474 1470
rect 44206 1095 44756 1274
rect 44955 1095 45474 1274
rect 44206 826 45474 1095
rect 50861 1275 52129 1471
rect 50861 1096 51411 1275
rect 51610 1096 52129 1275
rect 50861 827 52129 1096
rect 57483 1276 58751 1472
rect 57483 1097 58033 1276
rect 58232 1097 58751 1276
rect 57483 828 58751 1097
rect 39943 128 40188 131
rect 39943 110 39967 128
rect 40166 110 40188 128
rect 41841 128 42086 131
rect 41841 110 41865 128
rect 42064 110 42086 128
rect 39839 -194 39863 43
rect 40373 -194 41709 -8
rect 46494 126 46739 129
rect 46494 108 46518 126
rect 46717 108 46739 126
rect 48392 126 48637 129
rect 48392 108 48416 126
rect 48615 108 48637 126
rect 39839 -199 42206 -194
rect 46390 -196 46414 41
rect 46924 -196 48260 -10
rect 53149 127 53394 130
rect 53149 109 53173 127
rect 53372 109 53394 127
rect 55047 127 55292 130
rect 55047 109 55071 127
rect 55270 109 55292 127
rect 53045 -195 53069 42
rect 53579 -195 54915 -9
rect 59771 128 60016 131
rect 59771 110 59795 128
rect 59994 110 60016 128
rect 61669 128 61914 131
rect 61669 110 61693 128
rect 61892 110 61914 128
rect 59667 -194 59691 43
rect 60201 -194 61537 -8
rect 40227 -201 41898 -199
rect 46390 -201 48757 -196
rect 53045 -200 55412 -195
rect 59667 -199 62034 -194
rect 46778 -203 48449 -201
rect 53433 -202 55104 -200
rect 60055 -201 61726 -199
rect 62826 -1081 63293 1493
rect 63902 479 64264 480
rect 63902 305 63903 479
rect 64263 305 64264 479
rect 66260 414 67398 416
rect 67931 414 70367 1827
rect 72473 1669 72653 1676
rect 66260 413 70367 414
rect 65786 265 70367 413
rect 65786 167 65993 265
rect 65971 86 65993 167
rect 66192 172 70367 265
rect 66192 167 66643 172
rect 67204 170 70367 172
rect 66192 86 66216 167
rect 65971 83 66216 86
rect 67204 -110 67590 170
rect 68370 161 70367 170
rect 67204 -151 67364 -110
rect 67206 -182 67364 -151
rect 67434 -151 67590 -110
rect 67434 -182 67588 -151
rect 67206 -204 67588 -182
rect 62826 -1207 64305 -1081
rect 62826 -1279 63831 -1207
rect 63901 -1279 64305 -1207
rect 70133 -1217 70367 161
rect 72473 -1111 72653 -1083
rect 62826 -1319 64305 -1279
rect 67458 -1287 67514 -1286
rect 67454 -1288 67514 -1287
rect 67751 -1287 67790 -1286
rect 67751 -1288 67805 -1287
rect 62826 -1868 63293 -1319
rect 67454 -1404 67459 -1288
rect 67797 -1404 67805 -1288
rect 67454 -1545 67514 -1404
rect 67751 -1545 67805 -1404
rect 70133 -1317 70239 -1217
rect 70331 -1317 70367 -1217
rect 31905 -1922 32099 -1886
rect 36121 -1908 63295 -1868
rect 36121 -1913 48494 -1908
rect 28853 -2202 29689 -2126
rect 29755 -2202 29801 -2126
rect 28853 -3018 29801 -2202
rect 36121 -1985 41940 -1913
rect 42010 -1980 48494 -1913
rect 48564 -1920 63295 -1908
rect 48564 -1980 55143 -1920
rect 42010 -1985 55143 -1980
rect 36121 -1992 55143 -1985
rect 55213 -1992 63295 -1920
rect 36121 -2122 63295 -1992
rect 70133 -2249 70367 -1317
rect 63912 -2532 63913 -2374
rect 64273 -2532 64274 -2374
rect 29557 -3041 29801 -3018
rect 1217 -3892 1240 -3712
rect 4191 -3892 4448 -3712
rect 5087 -3892 5128 -3712
rect 7474 -3892 7568 -3712
rect 8207 -3892 8256 -3712
rect 10602 -3892 10632 -3712
rect 11271 -3892 11467 -3712
rect 13813 -3892 13834 -3712
rect 14473 -3892 14627 -3712
rect 16973 -3892 17011 -3712
rect 17650 -3892 17755 -3712
rect 20101 -3892 20163 -3712
rect 20802 -3892 20894 -3712
rect 23240 -3892 23319 -3712
rect 23958 -3892 24026 -3712
<< via4 >>
rect 3962 20024 4736 20067
rect 3962 19956 4274 20024
rect 4274 19956 4358 20024
rect 4358 19956 4736 20024
rect 3962 19755 4736 19956
rect 7095 20024 7869 20073
rect 7095 19956 7418 20024
rect 7418 19956 7502 20024
rect 7502 19956 7869 20024
rect 7095 19761 7869 19956
rect 10151 20020 10925 20089
rect 10151 19952 10550 20020
rect 10550 19952 10634 20020
rect 10634 19952 10925 20020
rect 10151 19777 10925 19952
rect 13267 20020 14041 20106
rect 13267 19952 13694 20020
rect 13694 19952 13778 20020
rect 13778 19952 14041 20020
rect 13267 19794 14041 19952
rect 16526 20024 17300 20095
rect 16526 19956 16896 20024
rect 16896 19956 16980 20024
rect 16980 19956 17300 20024
rect 16526 19783 17300 19956
rect 19675 20024 20449 20073
rect 19675 19956 20040 20024
rect 20040 19956 20124 20024
rect 20124 19956 20449 20024
rect 19675 19761 20449 19956
rect 22797 20020 23571 20067
rect 22797 19952 23172 20020
rect 23172 19952 23256 20020
rect 23256 19952 23571 20020
rect 22797 19755 23571 19952
rect 25990 20020 26764 20084
rect 25990 19952 26316 20020
rect 26316 19952 26400 20020
rect 26400 19952 26764 20020
rect 25990 19772 26764 19952
rect 40233 23813 40743 23891
rect 40233 23614 40292 23813
rect 40292 23614 40471 23813
rect 40471 23614 40743 23813
rect 40233 23587 40743 23614
rect 41801 23502 42105 23653
rect 41801 23323 41835 23502
rect 41835 23323 42034 23502
rect 42034 23323 42105 23502
rect 41801 23143 42105 23323
rect 42935 23500 43239 23663
rect 42935 23321 42977 23500
rect 42977 23321 43176 23500
rect 43176 23321 43239 23500
rect 42935 23153 43239 23321
rect 46746 23810 47256 23888
rect 46746 23611 46805 23810
rect 46805 23611 46984 23810
rect 46984 23611 47256 23810
rect 46746 23584 47256 23611
rect 48314 23499 48618 23650
rect 48314 23320 48348 23499
rect 48348 23320 48547 23499
rect 48547 23320 48618 23499
rect 48314 23140 48618 23320
rect 49448 23497 49752 23660
rect 49448 23318 49490 23497
rect 49490 23318 49689 23497
rect 49689 23318 49752 23497
rect 49448 23150 49752 23318
rect 53280 23805 53790 23883
rect 53280 23606 53339 23805
rect 53339 23606 53518 23805
rect 53518 23606 53790 23805
rect 53280 23579 53790 23606
rect 54848 23494 55152 23645
rect 40227 22163 40737 22231
rect 40227 21964 40306 22163
rect 40306 21964 40485 22163
rect 40485 21964 40737 22163
rect 40227 21927 40737 21964
rect 54848 23315 54882 23494
rect 54882 23315 55081 23494
rect 55081 23315 55152 23494
rect 54848 23135 55152 23315
rect 55982 23492 56286 23655
rect 55982 23313 56024 23492
rect 56024 23313 56223 23492
rect 56223 23313 56286 23492
rect 55982 23145 56286 23313
rect 59838 23809 60348 23887
rect 59838 23610 59897 23809
rect 59897 23610 60076 23809
rect 60076 23610 60348 23809
rect 59838 23583 60348 23610
rect 61406 23498 61710 23649
rect 46740 22160 47250 22228
rect 46740 21961 46819 22160
rect 46819 21961 46998 22160
rect 46998 21961 47250 22160
rect 46740 21924 47250 21961
rect 61406 23319 61440 23498
rect 61440 23319 61639 23498
rect 61639 23319 61710 23498
rect 61406 23139 61710 23319
rect 62540 23496 62844 23659
rect 62540 23317 62582 23496
rect 62582 23317 62781 23496
rect 62781 23317 62844 23496
rect 62540 23149 62844 23317
rect 53274 22155 53784 22223
rect 53274 21956 53353 22155
rect 53353 21956 53532 22155
rect 53532 21956 53784 22155
rect 53274 21919 53784 21956
rect 59832 22159 60342 22227
rect 59832 21960 59911 22159
rect 59911 21960 60090 22159
rect 60090 21960 60342 22159
rect 59832 21923 60342 21960
rect 40226 20559 40736 20626
rect 40226 20360 40301 20559
rect 40301 20360 40480 20559
rect 40480 20360 40736 20559
rect 46739 20556 47249 20623
rect 40226 20322 40736 20360
rect 41675 20280 41779 20441
rect 41779 20280 41978 20441
rect 41978 20280 42185 20441
rect 41675 20137 42185 20280
rect 43521 20280 43677 20441
rect 43677 20280 43876 20441
rect 43876 20280 44031 20441
rect 46739 20357 46814 20556
rect 46814 20357 46993 20556
rect 46993 20357 47249 20556
rect 53273 20551 53783 20618
rect 46739 20319 47249 20357
rect 43521 20137 44031 20280
rect 48188 20277 48292 20438
rect 48292 20277 48491 20438
rect 48491 20277 48698 20438
rect 48188 20134 48698 20277
rect 50034 20277 50190 20438
rect 50190 20277 50389 20438
rect 50389 20277 50544 20438
rect 53273 20352 53348 20551
rect 53348 20352 53527 20551
rect 53527 20352 53783 20551
rect 59831 20555 60341 20622
rect 53273 20314 53783 20352
rect 50034 20134 50544 20277
rect 54722 20272 54826 20433
rect 54826 20272 55025 20433
rect 55025 20272 55232 20433
rect 54722 20129 55232 20272
rect 56568 20272 56724 20433
rect 56724 20272 56923 20433
rect 56923 20272 57078 20433
rect 59831 20356 59906 20555
rect 59906 20356 60085 20555
rect 60085 20356 60341 20555
rect 59831 20318 60341 20356
rect 56568 20129 57078 20272
rect 61280 20276 61384 20437
rect 61384 20276 61583 20437
rect 61583 20276 61790 20437
rect 61280 20133 61790 20276
rect 63126 20276 63282 20437
rect 63282 20276 63481 20437
rect 63481 20276 63636 20437
rect 63126 20133 63636 20276
rect 72463 20811 72707 20916
rect 72463 20727 72485 20811
rect 72485 20727 72553 20811
rect 72553 20727 72707 20811
rect 72463 20585 72707 20727
rect 42677 18205 43187 18276
rect 40181 17892 40485 18055
rect 40181 17713 40244 17892
rect 40244 17713 40443 17892
rect 40443 17713 40485 17892
rect 40181 17545 40485 17713
rect 41315 17894 41619 18045
rect 42677 18006 42949 18205
rect 42949 18006 43128 18205
rect 43128 18006 43187 18205
rect 42677 17979 43187 18006
rect 41315 17715 41386 17894
rect 41386 17715 41585 17894
rect 41585 17715 41619 17894
rect 41315 17535 41619 17715
rect 5010 15731 5246 15748
rect 5010 15620 5077 15731
rect 5077 15620 5187 15731
rect 5187 15620 5246 15731
rect 5010 15512 5246 15620
rect 6175 15731 6411 15764
rect 6175 15620 6245 15731
rect 6245 15620 6355 15731
rect 6355 15620 6411 15731
rect 6175 15528 6411 15620
rect 7353 15731 7589 15752
rect 7353 15620 7413 15731
rect 7413 15620 7523 15731
rect 7523 15620 7589 15731
rect 7353 15516 7589 15620
rect 8522 15731 8758 15786
rect 8522 15620 8581 15731
rect 8581 15620 8691 15731
rect 8691 15620 8758 15731
rect 8522 15550 8758 15620
rect 9692 15729 9928 15788
rect 9692 15618 9755 15729
rect 9755 15618 9865 15729
rect 9865 15618 9928 15729
rect 9692 15552 9928 15618
rect 10856 15729 11092 15746
rect 10856 15618 10923 15729
rect 10923 15618 11033 15729
rect 11033 15618 11092 15729
rect 10856 15510 11092 15618
rect 12030 15729 12266 15759
rect 12030 15618 12091 15729
rect 12091 15618 12201 15729
rect 12201 15618 12266 15729
rect 12030 15523 12266 15618
rect 13202 15729 13438 15746
rect 13202 15618 13259 15729
rect 13259 15618 13369 15729
rect 13369 15618 13438 15729
rect 13202 15510 13438 15618
rect 14189 15639 14425 15724
rect 14189 15571 14268 15639
rect 14268 15571 14342 15639
rect 14342 15571 14425 15639
rect 14189 15488 14425 15571
rect 15638 15639 15874 15730
rect 15638 15571 15716 15639
rect 15716 15571 15790 15639
rect 15790 15571 15874 15639
rect 15638 15494 15874 15571
rect 17133 15637 17369 15715
rect 17133 15569 17214 15637
rect 17214 15569 17288 15637
rect 17288 15569 17369 15637
rect 17133 15479 17369 15569
rect 18581 15637 18817 15719
rect 18581 15569 18662 15637
rect 18662 15569 18736 15637
rect 18736 15569 18817 15637
rect 18581 15483 18817 15569
rect 20100 15639 20336 15719
rect 20100 15571 20182 15639
rect 20182 15571 20256 15639
rect 20256 15571 20336 15639
rect 20100 15483 20336 15571
rect 21549 15639 21785 15724
rect 21549 15571 21630 15639
rect 21630 15571 21704 15639
rect 21704 15571 21785 15639
rect 21549 15488 21785 15571
rect 23044 15637 23280 15715
rect 23044 15569 23128 15637
rect 23128 15569 23202 15637
rect 23202 15569 23280 15637
rect 23044 15479 23280 15569
rect 24493 15637 24729 15730
rect 24493 15569 24576 15637
rect 24576 15569 24650 15637
rect 24650 15569 24729 15637
rect 24493 15494 24729 15569
rect 42683 16555 43193 16623
rect 42683 16356 42935 16555
rect 42935 16356 43114 16555
rect 43114 16356 43193 16555
rect 42683 16319 43193 16356
rect 49235 18201 49745 18279
rect 46739 17888 47043 18051
rect 46739 17709 46802 17888
rect 46802 17709 47001 17888
rect 47001 17709 47043 17888
rect 46739 17541 47043 17709
rect 47873 17890 48177 18041
rect 49235 18002 49507 18201
rect 49507 18002 49686 18201
rect 49686 18002 49745 18201
rect 49235 17975 49745 18002
rect 47873 17711 47944 17890
rect 47944 17711 48143 17890
rect 48143 17711 48177 17890
rect 47873 17531 48177 17711
rect 55769 18206 56279 18284
rect 53273 17893 53577 18056
rect 53273 17714 53336 17893
rect 53336 17714 53535 17893
rect 53535 17714 53577 17893
rect 53273 17546 53577 17714
rect 54407 17895 54711 18046
rect 55769 18007 56041 18206
rect 56041 18007 56220 18206
rect 56220 18007 56279 18206
rect 55769 17980 56279 18007
rect 54407 17716 54478 17895
rect 54478 17716 54677 17895
rect 54677 17716 54711 17895
rect 54407 17536 54711 17716
rect 49241 16551 49751 16619
rect 49241 16352 49493 16551
rect 49493 16352 49672 16551
rect 49672 16352 49751 16551
rect 49241 16315 49751 16352
rect 55775 16556 56285 16624
rect 55775 16357 56027 16556
rect 56027 16357 56206 16556
rect 56206 16357 56285 16556
rect 55775 16320 56285 16357
rect 62282 18209 62792 18287
rect 59786 17896 60090 18059
rect 59786 17717 59849 17896
rect 59849 17717 60048 17896
rect 60048 17717 60090 17896
rect 59786 17549 60090 17717
rect 60920 17898 61224 18049
rect 62282 18010 62554 18209
rect 62554 18010 62733 18209
rect 62733 18010 62792 18209
rect 62282 17983 62792 18010
rect 60920 17719 60991 17898
rect 60991 17719 61190 17898
rect 61190 17719 61224 17898
rect 60920 17539 61224 17719
rect 62288 16559 62798 16627
rect 62288 16360 62540 16559
rect 62540 16360 62719 16559
rect 62719 16360 62798 16559
rect 62288 16323 62798 16360
rect 42684 14951 43194 15018
rect 39389 14672 39544 14833
rect 39544 14672 39743 14833
rect 39743 14672 39899 14833
rect 39389 14529 39899 14672
rect 41235 14672 41442 14833
rect 41442 14672 41641 14833
rect 41641 14672 41745 14833
rect 41235 14529 41745 14672
rect 42684 14752 42940 14951
rect 42940 14752 43119 14951
rect 43119 14752 43194 14951
rect 49242 14947 49752 15014
rect 42684 14714 43194 14752
rect 45947 14668 46102 14829
rect 46102 14668 46301 14829
rect 46301 14668 46457 14829
rect 45947 14525 46457 14668
rect 47793 14668 48000 14829
rect 48000 14668 48199 14829
rect 48199 14668 48303 14829
rect 47793 14525 48303 14668
rect 49242 14748 49498 14947
rect 49498 14748 49677 14947
rect 49677 14748 49752 14947
rect 55776 14952 56286 15019
rect 49242 14710 49752 14748
rect 52481 14673 52636 14834
rect 52636 14673 52835 14834
rect 52835 14673 52991 14834
rect 52481 14530 52991 14673
rect 54327 14673 54534 14834
rect 54534 14673 54733 14834
rect 54733 14673 54837 14834
rect 54327 14530 54837 14673
rect 55776 14753 56032 14952
rect 56032 14753 56211 14952
rect 56211 14753 56286 14952
rect 62289 14955 62799 15022
rect 55776 14715 56286 14753
rect 58994 14676 59149 14837
rect 59149 14676 59348 14837
rect 59348 14676 59504 14837
rect 58994 14533 59504 14676
rect 60840 14676 61047 14837
rect 61047 14676 61246 14837
rect 61246 14676 61350 14837
rect 60840 14533 61350 14676
rect 62289 14756 62545 14955
rect 62545 14756 62724 14955
rect 62724 14756 62799 14955
rect 62289 14718 62799 14756
rect 72465 17667 72709 17758
rect 72465 17583 72485 17667
rect 72485 17583 72553 17667
rect 72553 17583 72709 17667
rect 72465 17427 72709 17583
rect 1701 12886 1937 12908
rect 1701 12818 1772 12886
rect 1772 12818 1856 12886
rect 1856 12818 1937 12886
rect 1701 12672 1937 12818
rect 4856 12886 5092 12935
rect 4856 12818 4916 12886
rect 4916 12818 5000 12886
rect 5000 12818 5092 12886
rect 4856 12699 5092 12818
rect 7974 12882 8210 12926
rect 7974 12814 8048 12882
rect 8048 12814 8132 12882
rect 8132 12814 8210 12882
rect 7974 12690 8210 12814
rect 11120 12882 11356 12930
rect 11120 12814 11192 12882
rect 11192 12814 11276 12882
rect 11276 12814 11356 12882
rect 11120 12694 11356 12814
rect 14310 12886 14546 12917
rect 14310 12818 14394 12886
rect 14394 12818 14478 12886
rect 14478 12818 14546 12886
rect 14310 12681 14546 12818
rect 17461 12886 17697 12926
rect 17461 12818 17538 12886
rect 17538 12818 17622 12886
rect 17622 12818 17697 12886
rect 17461 12690 17697 12818
rect 20597 12882 20833 12908
rect 20597 12814 20670 12882
rect 20670 12814 20754 12882
rect 20754 12814 20833 12882
rect 20597 12672 20833 12814
rect 23734 12882 23970 12922
rect 23734 12814 23814 12882
rect 23814 12814 23898 12882
rect 23898 12814 23970 12882
rect 23734 12686 23970 12814
rect 31880 12415 32303 12596
rect 72463 14535 72707 14625
rect 72463 14451 72481 14535
rect 72481 14451 72549 14535
rect 72549 14451 72707 14535
rect 72463 14294 72707 14451
rect 31880 12321 31915 12415
rect 31915 12321 32003 12415
rect 32003 12321 32303 12415
rect 31880 12194 32303 12321
rect 41930 11175 42439 11283
rect 41930 11107 42127 11175
rect 42127 11107 42201 11175
rect 42201 11107 42439 11175
rect 41930 10975 42439 11107
rect 48472 11174 48981 11258
rect 48472 11106 48676 11174
rect 48676 11106 48750 11174
rect 48750 11106 48981 11174
rect 48472 10950 48981 11106
rect 55139 11195 55648 11243
rect 55139 11127 55330 11195
rect 55330 11127 55404 11195
rect 55404 11127 55648 11195
rect 55139 10936 55648 11127
rect 63840 11028 64200 11069
rect 63840 10960 63983 11028
rect 63983 10960 64057 11028
rect 64057 10960 64200 11028
rect 63840 10796 64200 10960
rect 1710 10152 1946 10185
rect 1710 10084 1772 10152
rect 1772 10084 1856 10152
rect 1856 10084 1946 10152
rect 1710 9949 1946 10084
rect 4842 10152 5078 10194
rect 4842 10084 4916 10152
rect 4916 10084 5000 10152
rect 5000 10084 5078 10152
rect 4842 9958 5078 10084
rect 7975 10148 8211 10185
rect 7975 10080 8048 10148
rect 8048 10080 8132 10148
rect 8132 10080 8211 10148
rect 7975 9949 8211 10080
rect 11108 10148 11344 10185
rect 11108 10080 11192 10148
rect 11192 10080 11276 10148
rect 11276 10080 11344 10148
rect 11108 9949 11344 10080
rect 14305 10152 14541 10189
rect 14305 10084 14394 10152
rect 14394 10084 14478 10152
rect 14478 10084 14541 10152
rect 14305 9953 14541 10084
rect 17461 10152 17697 10185
rect 17461 10084 17538 10152
rect 17538 10084 17622 10152
rect 17622 10084 17697 10152
rect 17461 9949 17697 10084
rect 20583 10148 20819 10193
rect 20583 10080 20670 10148
rect 20670 10080 20754 10148
rect 20754 10080 20819 10148
rect 20583 9957 20819 10080
rect 23723 10148 23959 10207
rect 23723 10080 23814 10148
rect 23814 10080 23898 10148
rect 23898 10080 23959 10148
rect 23723 9971 23959 10080
rect 31875 10347 32298 10502
rect 31875 10253 31913 10347
rect 31913 10253 32001 10347
rect 32001 10253 32298 10347
rect 31875 10100 32298 10253
rect 67512 10646 67749 10705
rect 67512 10530 67749 10646
rect 67512 10248 67749 10530
rect 35267 9275 35775 9345
rect 35267 9207 35463 9275
rect 35463 9207 35537 9275
rect 35537 9207 35775 9275
rect 35267 9037 35775 9207
rect 1706 7420 1942 7465
rect 1706 7352 1782 7420
rect 1782 7352 1866 7420
rect 1866 7352 1942 7420
rect 1706 7229 1942 7352
rect 4846 7420 5082 7447
rect 4846 7352 4926 7420
rect 4926 7352 5010 7420
rect 5010 7352 5082 7420
rect 4846 7211 5082 7352
rect 7981 7416 8217 7461
rect 7981 7348 8058 7416
rect 8058 7348 8142 7416
rect 8142 7348 8217 7416
rect 7981 7225 8217 7348
rect 11122 7416 11358 7442
rect 11122 7348 11202 7416
rect 11202 7348 11286 7416
rect 11286 7348 11358 7416
rect 11122 7206 11358 7348
rect 14331 7420 14567 7447
rect 14331 7352 14404 7420
rect 14404 7352 14488 7420
rect 14488 7352 14567 7420
rect 14331 7211 14567 7352
rect 17462 7420 17698 7447
rect 17462 7352 17548 7420
rect 17548 7352 17632 7420
rect 17632 7352 17698 7420
rect 17462 7211 17698 7352
rect 20593 7416 20829 7447
rect 20593 7348 20680 7416
rect 20680 7348 20764 7416
rect 20764 7348 20829 7416
rect 20593 7211 20829 7348
rect 23747 7416 23983 7456
rect 23747 7348 23824 7416
rect 23824 7348 23908 7416
rect 23908 7348 23983 7416
rect 23747 7220 23983 7348
rect 31865 8278 32288 8434
rect 31865 8184 31915 8278
rect 31915 8184 32003 8278
rect 32003 8184 32288 8278
rect 31865 8032 32288 8184
rect 38429 9262 38939 9340
rect 38429 9063 38488 9262
rect 38488 9063 38667 9262
rect 38667 9063 38939 9262
rect 38429 9036 38939 9063
rect 39997 8951 40301 9102
rect 35242 6690 35750 6763
rect 35242 6622 35455 6690
rect 35455 6622 35529 6690
rect 35529 6622 35750 6690
rect 35242 6455 35750 6622
rect 3274 5883 3510 5958
rect 3274 5783 3333 5883
rect 3333 5783 3435 5883
rect 3435 5783 3510 5883
rect 3274 5722 3510 5783
rect 4001 5883 4237 5960
rect 4001 5783 4071 5883
rect 4071 5783 4173 5883
rect 4173 5783 4237 5883
rect 4001 5724 4237 5783
rect 4747 5883 4983 5962
rect 4747 5783 4809 5883
rect 4809 5783 4911 5883
rect 4911 5783 4983 5883
rect 4747 5726 4983 5783
rect 5486 5883 5722 5962
rect 5486 5783 5547 5883
rect 5547 5783 5649 5883
rect 5649 5783 5722 5883
rect 5486 5726 5722 5783
rect 6217 5883 6453 5951
rect 6217 5783 6287 5883
rect 6287 5783 6389 5883
rect 6389 5783 6453 5883
rect 6217 5715 6453 5783
rect 6958 5883 7194 5956
rect 6958 5783 7029 5883
rect 7029 5783 7131 5883
rect 7131 5783 7194 5883
rect 6958 5720 7194 5783
rect 7706 5883 7942 5958
rect 7706 5783 7767 5883
rect 7767 5783 7869 5883
rect 7869 5783 7942 5883
rect 7706 5722 7942 5783
rect 8440 5885 8676 5960
rect 8440 5785 8505 5885
rect 8505 5785 8607 5885
rect 8607 5785 8676 5885
rect 8440 5724 8676 5785
rect 10020 4486 10256 4531
rect 10020 4398 10095 4486
rect 10095 4398 10189 4486
rect 10189 4398 10256 4486
rect 10020 4295 10256 4398
rect 12093 4484 12329 4519
rect 12093 4396 12163 4484
rect 12163 4396 12257 4484
rect 12257 4396 12329 4484
rect 12093 4283 12329 4396
rect 14156 4486 14392 4519
rect 14156 4398 14232 4486
rect 14232 4398 14326 4486
rect 14326 4398 14392 4486
rect 14156 4283 14392 4398
rect 16220 4484 16456 4515
rect 16220 4396 16300 4484
rect 16300 4396 16394 4484
rect 16394 4396 16456 4484
rect 16220 4279 16456 4396
rect 18293 4484 18529 4522
rect 18293 4396 18369 4484
rect 18369 4396 18463 4484
rect 18463 4396 18529 4484
rect 18293 4286 18529 4396
rect 20361 4482 20597 4529
rect 20361 4394 20437 4482
rect 20437 4394 20531 4482
rect 20531 4394 20597 4482
rect 20361 4293 20597 4394
rect 22434 4484 22670 4524
rect 22434 4396 22506 4484
rect 22506 4396 22600 4484
rect 22600 4396 22670 4484
rect 22434 4288 22670 4396
rect 24501 4482 24737 4515
rect 24501 4394 24574 4482
rect 24574 4394 24668 4482
rect 24668 4394 24737 4482
rect 24501 4279 24737 4394
rect 31891 6210 32314 6371
rect 31891 6116 31913 6210
rect 31913 6116 32001 6210
rect 32001 6116 32314 6210
rect 31891 5969 32314 6116
rect 39997 8772 40031 8951
rect 40031 8772 40230 8951
rect 40230 8772 40301 8951
rect 39997 8592 40301 8772
rect 41131 8949 41435 9112
rect 41131 8770 41173 8949
rect 41173 8770 41372 8949
rect 41372 8770 41435 8949
rect 41131 8602 41435 8770
rect 44978 9350 45488 9428
rect 44978 9151 45037 9350
rect 45037 9151 45216 9350
rect 45216 9151 45488 9350
rect 44978 9124 45488 9151
rect 46546 9039 46850 9190
rect 46546 8860 46580 9039
rect 46580 8860 46779 9039
rect 46779 8860 46850 9039
rect 46546 8680 46850 8860
rect 47680 9037 47984 9200
rect 47680 8858 47722 9037
rect 47722 8858 47921 9037
rect 47921 8858 47984 9037
rect 47680 8690 47984 8858
rect 51632 9282 52142 9360
rect 51632 9083 51691 9282
rect 51691 9083 51870 9282
rect 51870 9083 52142 9282
rect 51632 9056 52142 9083
rect 53200 8971 53504 9122
rect 38423 7612 38933 7680
rect 38423 7413 38502 7612
rect 38502 7413 38681 7612
rect 38681 7413 38933 7612
rect 38423 7376 38933 7413
rect 53200 8792 53234 8971
rect 53234 8792 53433 8971
rect 53433 8792 53504 8971
rect 53200 8612 53504 8792
rect 54334 8969 54638 9132
rect 54334 8790 54376 8969
rect 54376 8790 54575 8969
rect 54575 8790 54638 8969
rect 54334 8622 54638 8790
rect 58257 9350 58767 9428
rect 58257 9151 58316 9350
rect 58316 9151 58495 9350
rect 58495 9151 58767 9350
rect 58257 9124 58767 9151
rect 59825 9039 60129 9190
rect 44972 7700 45482 7768
rect 44972 7501 45051 7700
rect 45051 7501 45230 7700
rect 45230 7501 45482 7700
rect 44972 7464 45482 7501
rect 59825 8860 59859 9039
rect 59859 8860 60058 9039
rect 60058 8860 60129 9039
rect 59825 8680 60129 8860
rect 60959 9037 61263 9200
rect 60959 8858 61001 9037
rect 61001 8858 61200 9037
rect 61200 8858 61263 9037
rect 60959 8690 61263 8858
rect 51626 7632 52136 7700
rect 51626 7433 51705 7632
rect 51705 7433 51884 7632
rect 51884 7433 52136 7632
rect 51626 7396 52136 7433
rect 65849 9854 66222 9856
rect 65849 9659 65912 9854
rect 65912 9659 66178 9854
rect 66178 9659 66222 9854
rect 58251 7700 58761 7768
rect 58251 7501 58330 7700
rect 58330 7501 58509 7700
rect 58509 7501 58761 7700
rect 58251 7464 58761 7501
rect 65849 9517 66222 9659
rect 63846 8457 64206 8506
rect 63846 8389 63978 8457
rect 63978 8389 64052 8457
rect 64052 8389 64206 8457
rect 63846 8233 64206 8389
rect 72465 11391 72709 11507
rect 72465 11307 72481 11391
rect 72481 11307 72549 11391
rect 72549 11307 72709 11391
rect 72465 11176 72709 11307
rect 67514 6555 67751 6614
rect 44971 6096 45481 6163
rect 38422 6008 38932 6075
rect 38422 5809 38497 6008
rect 38497 5809 38676 6008
rect 38676 5809 38932 6008
rect 44971 5897 45046 6096
rect 45046 5897 45225 6096
rect 45225 5897 45481 6096
rect 58250 6096 58760 6163
rect 51625 6028 52135 6095
rect 38422 5771 38932 5809
rect 39871 5729 39975 5890
rect 39975 5729 40174 5890
rect 40174 5729 40381 5890
rect 39871 5586 40381 5729
rect 41717 5729 41873 5890
rect 41873 5729 42072 5890
rect 42072 5729 42227 5890
rect 44971 5859 45481 5897
rect 41717 5586 42227 5729
rect 46420 5817 46524 5978
rect 46524 5817 46723 5978
rect 46723 5817 46930 5978
rect 46420 5674 46930 5817
rect 48266 5817 48422 5978
rect 48422 5817 48621 5978
rect 48621 5817 48776 5978
rect 48266 5674 48776 5817
rect 51625 5829 51700 6028
rect 51700 5829 51879 6028
rect 51879 5829 52135 6028
rect 51625 5791 52135 5829
rect 53074 5749 53178 5910
rect 53178 5749 53377 5910
rect 53377 5749 53584 5910
rect 53074 5606 53584 5749
rect 54920 5749 55076 5910
rect 55076 5749 55275 5910
rect 55275 5749 55430 5910
rect 58250 5897 58325 6096
rect 58325 5897 58504 6096
rect 58504 5897 58760 6096
rect 58250 5859 58760 5897
rect 54920 5606 55430 5749
rect 59699 5817 59803 5978
rect 59803 5817 60002 5978
rect 60002 5817 60209 5978
rect 59699 5674 60209 5817
rect 61545 5817 61701 5978
rect 61701 5817 61900 5978
rect 61900 5817 62055 5978
rect 61545 5674 62055 5817
rect 67514 6439 67751 6555
rect 67514 6157 67751 6439
rect 65851 5763 66224 5765
rect 65851 5568 65914 5763
rect 65914 5568 66180 5763
rect 66180 5568 66224 5763
rect 63847 5424 64207 5468
rect 63847 5356 63978 5424
rect 63978 5356 64052 5424
rect 64052 5356 64207 5424
rect 63847 5195 64207 5356
rect 65851 5426 66224 5568
rect 72465 8189 72709 8316
rect 72465 8105 72485 8189
rect 72485 8105 72553 8189
rect 72553 8105 72709 8189
rect 72465 7985 72709 8105
rect 72465 5045 72709 5150
rect 72465 4961 72485 5045
rect 72485 4961 72553 5045
rect 72553 4961 72709 5045
rect 72465 4819 72709 4961
rect 31875 4141 32298 4272
rect 31875 4047 31913 4141
rect 31913 4047 32001 4141
rect 32001 4047 32298 4141
rect 31875 3870 32298 4047
rect 35218 3412 35726 3458
rect 35218 3344 35436 3412
rect 35436 3344 35510 3412
rect 35510 3344 35726 3412
rect 35218 3150 35726 3344
rect 1239 168 1875 226
rect 1239 100 1510 168
rect 1510 100 1594 168
rect 1594 100 1875 168
rect 1239 -197 1875 100
rect 4439 168 5075 226
rect 4439 100 4654 168
rect 4654 100 4738 168
rect 4738 100 5075 168
rect 4439 -197 5075 100
rect 7565 172 8201 231
rect 7565 104 7786 172
rect 7786 104 7870 172
rect 7870 104 8201 172
rect 7565 -192 8201 104
rect 10640 172 11276 231
rect 10640 104 10930 172
rect 10930 104 11014 172
rect 11014 104 11276 172
rect 10640 -192 11276 104
rect 13830 168 14466 231
rect 13830 100 14132 168
rect 14132 100 14216 168
rect 14216 100 14466 168
rect 13830 -192 14466 100
rect 17055 168 17691 226
rect 17055 100 17276 168
rect 17276 100 17360 168
rect 17360 100 17691 168
rect 17055 -197 17691 100
rect 20176 172 20812 226
rect 20176 104 20408 172
rect 20408 104 20492 172
rect 20492 104 20812 172
rect 20176 -197 20812 104
rect 23263 172 23899 224
rect 23263 104 23552 172
rect 23552 104 23636 172
rect 23636 104 23899 172
rect 23263 -199 23899 104
rect 31880 2073 32303 2209
rect 31880 1979 31911 2073
rect 31911 1979 31999 2073
rect 31999 1979 32303 2073
rect 38421 3482 38931 3560
rect 38421 3283 38480 3482
rect 38480 3283 38659 3482
rect 38659 3283 38931 3482
rect 38421 3256 38931 3283
rect 39989 3171 40293 3322
rect 31880 1807 32303 1979
rect 35193 652 35701 694
rect 35193 584 35452 652
rect 35452 584 35526 652
rect 35526 584 35701 652
rect 35193 386 35701 584
rect 31885 4 32308 167
rect 31885 -90 31913 4
rect 31913 -90 32001 4
rect 32001 -90 32308 4
rect 31885 -235 32308 -90
rect 39989 2992 40023 3171
rect 40023 2992 40222 3171
rect 40222 2992 40293 3171
rect 39989 2812 40293 2992
rect 41123 3169 41427 3332
rect 41123 2990 41165 3169
rect 41165 2990 41364 3169
rect 41364 2990 41427 3169
rect 41123 2822 41427 2990
rect 44972 3480 45482 3558
rect 44972 3281 45031 3480
rect 45031 3281 45210 3480
rect 45210 3281 45482 3480
rect 44972 3254 45482 3281
rect 46540 3169 46844 3320
rect 46540 2990 46574 3169
rect 46574 2990 46773 3169
rect 46773 2990 46844 3169
rect 46540 2810 46844 2990
rect 47674 3167 47978 3330
rect 47674 2988 47716 3167
rect 47716 2988 47915 3167
rect 47915 2988 47978 3167
rect 47674 2820 47978 2988
rect 51627 3481 52137 3559
rect 51627 3282 51686 3481
rect 51686 3282 51865 3481
rect 51865 3282 52137 3481
rect 51627 3255 52137 3282
rect 53195 3170 53499 3321
rect 38415 1832 38925 1900
rect 38415 1633 38494 1832
rect 38494 1633 38673 1832
rect 38673 1633 38925 1832
rect 38415 1596 38925 1633
rect 53195 2991 53229 3170
rect 53229 2991 53428 3170
rect 53428 2991 53499 3170
rect 53195 2811 53499 2991
rect 54329 3168 54633 3331
rect 54329 2989 54371 3168
rect 54371 2989 54570 3168
rect 54570 2989 54633 3168
rect 54329 2821 54633 2989
rect 58249 3482 58759 3560
rect 58249 3283 58308 3482
rect 58308 3283 58487 3482
rect 58487 3283 58759 3482
rect 58249 3256 58759 3283
rect 59817 3171 60121 3322
rect 44966 1830 45476 1898
rect 44966 1631 45045 1830
rect 45045 1631 45224 1830
rect 45224 1631 45476 1830
rect 44966 1594 45476 1631
rect 59817 2992 59851 3171
rect 59851 2992 60050 3171
rect 60050 2992 60121 3171
rect 59817 2812 60121 2992
rect 60951 3169 61255 3332
rect 60951 2990 60993 3169
rect 60993 2990 61192 3169
rect 61192 2990 61255 3169
rect 60951 2822 61255 2990
rect 51621 1831 52131 1899
rect 51621 1632 51700 1831
rect 51700 1632 51879 1831
rect 51879 1632 52131 1831
rect 51621 1595 52131 1632
rect 58243 1832 58753 1900
rect 58243 1633 58322 1832
rect 58322 1633 58501 1832
rect 58501 1633 58753 1832
rect 58243 1596 58753 1633
rect 63907 3504 64267 3547
rect 63907 3436 64049 3504
rect 64049 3436 64123 3504
rect 64123 3436 64267 3504
rect 63907 3274 64267 3436
rect 67514 3060 67751 3119
rect 67514 2944 67751 3060
rect 67514 2662 67751 2944
rect 65851 2268 66224 2270
rect 65851 2073 65914 2268
rect 65914 2073 66180 2268
rect 66180 2073 66224 2268
rect 65851 2001 66224 2073
rect 38414 228 38924 295
rect 38414 29 38489 228
rect 38489 29 38668 228
rect 38668 29 38924 228
rect 44965 226 45475 293
rect 38414 -9 38924 29
rect 39863 -51 39967 110
rect 39967 -51 40166 110
rect 40166 -51 40373 110
rect 39863 -194 40373 -51
rect 41709 -51 41865 110
rect 41865 -51 42064 110
rect 42064 -51 42219 110
rect 44965 27 45040 226
rect 45040 27 45219 226
rect 45219 27 45475 226
rect 51620 227 52130 294
rect 44965 -11 45475 27
rect 41709 -194 42219 -51
rect 46414 -53 46518 108
rect 46518 -53 46717 108
rect 46717 -53 46924 108
rect 46414 -196 46924 -53
rect 48260 -53 48416 108
rect 48416 -53 48615 108
rect 48615 -53 48770 108
rect 51620 28 51695 227
rect 51695 28 51874 227
rect 51874 28 52130 227
rect 58242 228 58752 295
rect 51620 -10 52130 28
rect 48260 -196 48770 -53
rect 53069 -52 53173 109
rect 53173 -52 53372 109
rect 53372 -52 53579 109
rect 53069 -195 53579 -52
rect 54915 -52 55071 109
rect 55071 -52 55270 109
rect 55270 -52 55425 109
rect 58242 29 58317 228
rect 58317 29 58496 228
rect 58496 29 58752 228
rect 58242 -9 58752 29
rect 54915 -195 55425 -52
rect 59691 -51 59795 110
rect 59795 -51 59994 110
rect 59994 -51 60201 110
rect 59691 -194 60201 -51
rect 61537 -51 61693 110
rect 61693 -51 61892 110
rect 61892 -51 62047 110
rect 61537 -194 62047 -51
rect 41892 -713 42400 -523
rect 41892 -781 42162 -713
rect 42162 -781 42236 -713
rect 42236 -781 42400 -713
rect 41892 -831 42400 -781
rect 48431 -708 48939 -542
rect 48431 -776 48716 -708
rect 48716 -776 48790 -708
rect 48790 -776 48939 -708
rect 48431 -850 48939 -776
rect 55137 -720 55645 -567
rect 55137 -788 55365 -720
rect 55365 -788 55439 -720
rect 55439 -788 55645 -720
rect 55137 -875 55645 -788
rect 63903 434 64263 479
rect 63903 366 64046 434
rect 64046 366 64120 434
rect 64120 366 64263 434
rect 63903 206 64263 366
rect 72463 1913 72707 2007
rect 72463 1829 72481 1913
rect 72481 1829 72549 1913
rect 72549 1829 72707 1913
rect 72463 1676 72707 1829
rect 67514 -1288 67751 -1229
rect 67514 -1404 67751 -1288
rect 67514 -1686 67751 -1404
rect 31885 -2064 32308 -1922
rect 31885 -2158 31911 -2064
rect 31911 -2158 31999 -2064
rect 31999 -2158 32308 -2064
rect 65851 -2080 66224 -2078
rect 31885 -2324 32308 -2158
rect 65851 -2275 65914 -2080
rect 65914 -2275 66180 -2080
rect 66180 -2275 66224 -2080
rect 72465 -1231 72709 -1111
rect 72465 -1315 72481 -1231
rect 72481 -1315 72549 -1231
rect 72549 -1315 72709 -1231
rect 72465 -1442 72709 -1315
rect 63913 -2411 64273 -2374
rect 63913 -2479 64053 -2411
rect 64053 -2479 64127 -2411
rect 64127 -2479 64273 -2411
rect 63913 -2647 64273 -2479
rect 65851 -2417 66224 -2275
rect 1240 -3724 1879 -3653
rect 1240 -3792 1542 -3724
rect 1542 -3792 1626 -3724
rect 1626 -3792 1879 -3724
rect 1240 -4061 1879 -3792
rect 4448 -3724 5087 -3653
rect 4448 -3792 4686 -3724
rect 4686 -3792 4770 -3724
rect 4770 -3792 5087 -3724
rect 4448 -4061 5087 -3792
rect 7568 -3720 8207 -3642
rect 7568 -3788 7818 -3720
rect 7818 -3788 7902 -3720
rect 7902 -3788 8207 -3720
rect 7568 -4050 8207 -3788
rect 10632 -3720 11271 -3673
rect 10632 -3788 10962 -3720
rect 10962 -3788 11046 -3720
rect 11046 -3788 11271 -3720
rect 10632 -4081 11271 -3788
rect 13834 -3724 14473 -3663
rect 13834 -3792 14164 -3724
rect 14164 -3792 14248 -3724
rect 14248 -3792 14473 -3724
rect 13834 -4071 14473 -3792
rect 17011 -3724 17650 -3673
rect 17011 -3792 17308 -3724
rect 17308 -3792 17392 -3724
rect 17392 -3792 17650 -3724
rect 17011 -4081 17650 -3792
rect 20163 -3720 20802 -3673
rect 20163 -3788 20440 -3720
rect 20440 -3788 20524 -3720
rect 20524 -3788 20802 -3720
rect 20163 -4081 20802 -3788
rect 23319 -3720 23958 -3673
rect 23319 -3788 23584 -3720
rect 23584 -3788 23668 -3720
rect 23668 -3788 23958 -3720
rect 23319 -4081 23958 -3788
<< metal5 >>
rect -753 23891 73229 24297
rect -753 23587 40233 23891
rect 40743 23888 73229 23891
rect 40743 23663 46746 23888
rect 40743 23653 42935 23663
rect 40743 23587 41801 23653
rect -753 23143 41801 23587
rect 42105 23153 42935 23653
rect 43239 23584 46746 23663
rect 47256 23887 73229 23888
rect 47256 23883 59838 23887
rect 47256 23660 53280 23883
rect 47256 23650 49448 23660
rect 47256 23584 48314 23650
rect 43239 23153 48314 23584
rect 42105 23143 48314 23153
rect -753 23140 48314 23143
rect 48618 23150 49448 23650
rect 49752 23579 53280 23660
rect 53790 23655 59838 23883
rect 53790 23645 55982 23655
rect 53790 23579 54848 23645
rect 49752 23150 54848 23579
rect 48618 23140 54848 23150
rect -753 23135 54848 23140
rect 55152 23145 55982 23645
rect 56286 23583 59838 23655
rect 60348 23659 73229 23887
rect 60348 23649 62540 23659
rect 60348 23583 61406 23649
rect 56286 23145 61406 23583
rect 55152 23139 61406 23145
rect 61710 23149 62540 23649
rect 62844 23149 73229 23659
rect 61710 23139 73229 23149
rect 55152 23135 73229 23139
rect -753 22231 73229 23135
rect -753 21927 40227 22231
rect 40737 22228 73229 22231
rect 40737 21927 46740 22228
rect -753 21924 46740 21927
rect 47250 22227 73229 22228
rect 47250 22223 59832 22227
rect 47250 21924 53274 22223
rect -753 21919 53274 21924
rect 53784 21923 59832 22223
rect 60342 21923 73229 22227
rect 53784 21919 73229 21923
rect -753 20916 73229 21919
rect -753 20626 72463 20916
rect -753 20322 40226 20626
rect 40736 20623 72463 20626
rect 40736 20441 46739 20623
rect 40736 20322 41675 20441
rect -753 20137 41675 20322
rect 42185 20137 43521 20441
rect 44031 20319 46739 20441
rect 47249 20622 72463 20623
rect 47249 20618 59831 20622
rect 47249 20438 53273 20618
rect 47249 20319 48188 20438
rect 44031 20137 48188 20319
rect -753 20134 48188 20137
rect 48698 20134 50034 20438
rect 50544 20314 53273 20438
rect 53783 20433 59831 20618
rect 53783 20314 54722 20433
rect 50544 20134 54722 20314
rect -753 20129 54722 20134
rect 55232 20129 56568 20433
rect 57078 20318 59831 20433
rect 60341 20585 72463 20622
rect 72707 20585 73229 20916
rect 60341 20437 73229 20585
rect 60341 20318 61280 20437
rect 57078 20133 61280 20318
rect 61790 20133 63126 20437
rect 63636 20133 73229 20437
rect 57078 20129 73229 20133
rect -753 20106 73229 20129
rect -753 20089 13267 20106
rect -753 20073 10151 20089
rect -753 20067 7095 20073
rect -753 19755 3962 20067
rect 4736 19761 7095 20067
rect 7869 19777 10151 20073
rect 10925 19794 13267 20089
rect 14041 20095 73229 20106
rect 14041 19794 16526 20095
rect 10925 19783 16526 19794
rect 17300 20084 73229 20095
rect 17300 20073 25990 20084
rect 17300 19783 19675 20073
rect 10925 19777 19675 19783
rect 7869 19761 19675 19777
rect 20449 20067 25990 20073
rect 20449 19761 22797 20067
rect 4736 19755 22797 19761
rect 23571 19772 25990 20067
rect 26764 19772 73229 20084
rect 23571 19755 73229 19772
rect -753 18287 73229 19755
rect -753 18284 62282 18287
rect -753 18279 55769 18284
rect -753 18276 49235 18279
rect -753 18055 42677 18276
rect -753 17545 40181 18055
rect 40485 18045 42677 18055
rect 40485 17545 41315 18045
rect -753 17535 41315 17545
rect 41619 17979 42677 18045
rect 43187 18051 49235 18276
rect 43187 17979 46739 18051
rect 41619 17541 46739 17979
rect 47043 18041 49235 18051
rect 47043 17541 47873 18041
rect 41619 17535 47873 17541
rect -753 17531 47873 17535
rect 48177 17975 49235 18041
rect 49745 18056 55769 18279
rect 49745 17975 53273 18056
rect 48177 17546 53273 17975
rect 53577 18046 55769 18056
rect 53577 17546 54407 18046
rect 48177 17536 54407 17546
rect 54711 17980 55769 18046
rect 56279 18059 62282 18284
rect 56279 17980 59786 18059
rect 54711 17549 59786 17980
rect 60090 18049 62282 18059
rect 60090 17549 60920 18049
rect 54711 17539 60920 17549
rect 61224 17983 62282 18049
rect 62792 17983 73229 18287
rect 61224 17758 73229 17983
rect 61224 17539 72465 17758
rect 54711 17536 72465 17539
rect 48177 17531 72465 17536
rect -753 17427 72465 17531
rect 72709 17427 73229 17758
rect -753 16627 73229 17427
rect -753 16624 62288 16627
rect -753 16623 55775 16624
rect -753 16319 42683 16623
rect 43193 16619 55775 16623
rect 43193 16319 49241 16619
rect -753 16315 49241 16319
rect 49751 16320 55775 16619
rect 56285 16323 62288 16624
rect 62798 16323 73229 16627
rect 56285 16320 73229 16323
rect 49751 16315 73229 16320
rect -753 15788 73229 16315
rect -753 15786 9692 15788
rect -753 15764 8522 15786
rect -753 15748 6175 15764
rect -753 15512 5010 15748
rect 5246 15528 6175 15748
rect 6411 15752 8522 15764
rect 6411 15528 7353 15752
rect 5246 15516 7353 15528
rect 7589 15550 8522 15752
rect 8758 15552 9692 15786
rect 9928 15759 73229 15788
rect 9928 15746 12030 15759
rect 9928 15552 10856 15746
rect 8758 15550 10856 15552
rect 7589 15516 10856 15550
rect 5246 15512 10856 15516
rect -753 15510 10856 15512
rect 11092 15523 12030 15746
rect 12266 15746 73229 15759
rect 12266 15523 13202 15746
rect 11092 15510 13202 15523
rect 13438 15730 73229 15746
rect 13438 15724 15638 15730
rect 13438 15510 14189 15724
rect -753 15488 14189 15510
rect 14425 15494 15638 15724
rect 15874 15724 24493 15730
rect 15874 15719 21549 15724
rect 15874 15715 18581 15719
rect 15874 15494 17133 15715
rect 14425 15488 17133 15494
rect -753 15479 17133 15488
rect 17369 15483 18581 15715
rect 18817 15483 20100 15719
rect 20336 15488 21549 15719
rect 21785 15715 24493 15724
rect 21785 15488 23044 15715
rect 20336 15483 23044 15488
rect 17369 15479 23044 15483
rect 23280 15494 24493 15715
rect 24729 15494 73229 15730
rect 23280 15479 73229 15494
rect -753 15022 73229 15479
rect -753 15019 62289 15022
rect -753 15018 55776 15019
rect -753 14833 42684 15018
rect -753 14529 39389 14833
rect 39899 14529 41235 14833
rect 41745 14714 42684 14833
rect 43194 15014 55776 15018
rect 43194 14829 49242 15014
rect 43194 14714 45947 14829
rect 41745 14529 45947 14714
rect -753 14525 45947 14529
rect 46457 14525 47793 14829
rect 48303 14710 49242 14829
rect 49752 14834 55776 15014
rect 49752 14710 52481 14834
rect 48303 14530 52481 14710
rect 52991 14530 54327 14834
rect 54837 14715 55776 14834
rect 56286 14837 62289 15019
rect 56286 14715 58994 14837
rect 54837 14533 58994 14715
rect 59504 14533 60840 14837
rect 61350 14718 62289 14837
rect 62799 14718 73229 15022
rect 61350 14625 73229 14718
rect 61350 14533 72463 14625
rect 54837 14530 72463 14533
rect 48303 14525 72463 14530
rect -753 14294 72463 14525
rect 72707 14294 73229 14625
rect -753 12935 73229 14294
rect -753 12908 4856 12935
rect -753 12672 1701 12908
rect 1937 12699 4856 12908
rect 5092 12930 73229 12935
rect 5092 12926 11120 12930
rect 5092 12699 7974 12926
rect 1937 12690 7974 12699
rect 8210 12694 11120 12926
rect 11356 12926 73229 12930
rect 11356 12917 17461 12926
rect 11356 12694 14310 12917
rect 8210 12690 14310 12694
rect 1937 12681 14310 12690
rect 14546 12690 17461 12917
rect 17697 12922 73229 12926
rect 17697 12908 23734 12922
rect 17697 12690 20597 12908
rect 14546 12681 20597 12690
rect 1937 12672 20597 12681
rect 20833 12686 23734 12908
rect 23970 12686 73229 12922
rect 20833 12672 73229 12686
rect -753 12596 73229 12672
rect -753 12194 31880 12596
rect 32303 12194 73229 12596
rect -753 11507 73229 12194
rect -753 11283 72465 11507
rect -753 10975 41930 11283
rect 42439 11258 72465 11283
rect 42439 10975 48472 11258
rect -753 10950 48472 10975
rect 48981 11243 72465 11258
rect 48981 10950 55139 11243
rect -753 10936 55139 10950
rect 55648 11176 72465 11243
rect 72709 11176 73229 11507
rect 55648 11069 73229 11176
rect 55648 10936 63840 11069
rect -753 10796 63840 10936
rect 64200 10796 73229 11069
rect -753 10705 73229 10796
rect -753 10502 67512 10705
rect -753 10207 31875 10502
rect -753 10194 23723 10207
rect -753 10185 4842 10194
rect -753 9949 1710 10185
rect 1946 9958 4842 10185
rect 5078 10193 23723 10194
rect 5078 10189 20583 10193
rect 5078 10185 14305 10189
rect 5078 9958 7975 10185
rect 1946 9949 7975 9958
rect 8211 9949 11108 10185
rect 11344 9953 14305 10185
rect 14541 10185 20583 10189
rect 14541 9953 17461 10185
rect 11344 9949 17461 9953
rect 17697 9957 20583 10185
rect 20819 9971 23723 10193
rect 23959 10100 31875 10207
rect 32298 10248 67512 10502
rect 67749 10248 73229 10705
rect 32298 10100 73229 10248
rect 23959 9971 73229 10100
rect 20819 9957 73229 9971
rect 17697 9949 73229 9957
rect -753 9856 73229 9949
rect -753 9517 65849 9856
rect 66222 9517 73229 9856
rect -753 9428 73229 9517
rect -753 9345 44978 9428
rect -753 9037 35267 9345
rect 35775 9340 44978 9345
rect 35775 9037 38429 9340
rect -753 9036 38429 9037
rect 38939 9124 44978 9340
rect 45488 9360 58257 9428
rect 45488 9200 51632 9360
rect 45488 9190 47680 9200
rect 45488 9124 46546 9190
rect 38939 9112 46546 9124
rect 38939 9102 41131 9112
rect 38939 9036 39997 9102
rect -753 8592 39997 9036
rect 40301 8602 41131 9102
rect 41435 8680 46546 9112
rect 46850 8690 47680 9190
rect 47984 9056 51632 9200
rect 52142 9132 58257 9360
rect 52142 9122 54334 9132
rect 52142 9056 53200 9122
rect 47984 8690 53200 9056
rect 46850 8680 53200 8690
rect 41435 8612 53200 8680
rect 53504 8622 54334 9122
rect 54638 9124 58257 9132
rect 58767 9200 73229 9428
rect 58767 9190 60959 9200
rect 58767 9124 59825 9190
rect 54638 8680 59825 9124
rect 60129 8690 60959 9190
rect 61263 8690 73229 9200
rect 60129 8680 73229 8690
rect 54638 8622 73229 8680
rect 53504 8612 73229 8622
rect 41435 8602 73229 8612
rect 40301 8592 73229 8602
rect -753 8506 73229 8592
rect -753 8434 63846 8506
rect -753 8032 31865 8434
rect 32288 8233 63846 8434
rect 64206 8316 73229 8506
rect 64206 8233 72465 8316
rect 32288 8032 72465 8233
rect -753 7985 72465 8032
rect 72709 7985 73229 8316
rect -753 7768 73229 7985
rect -753 7680 44972 7768
rect -753 7465 38423 7680
rect -753 7229 1706 7465
rect 1942 7461 38423 7465
rect 1942 7447 7981 7461
rect 1942 7229 4846 7447
rect -753 7211 4846 7229
rect 5082 7225 7981 7447
rect 8217 7456 38423 7461
rect 8217 7447 23747 7456
rect 8217 7442 14331 7447
rect 8217 7225 11122 7442
rect 5082 7211 11122 7225
rect -753 7206 11122 7211
rect 11358 7211 14331 7442
rect 14567 7211 17462 7447
rect 17698 7211 20593 7447
rect 20829 7220 23747 7447
rect 23983 7376 38423 7456
rect 38933 7464 44972 7680
rect 45482 7700 58251 7768
rect 45482 7464 51626 7700
rect 38933 7396 51626 7464
rect 52136 7464 58251 7700
rect 58761 7464 73229 7768
rect 52136 7396 73229 7464
rect 38933 7376 73229 7396
rect 23983 7220 73229 7376
rect 20829 7211 73229 7220
rect 11358 7206 73229 7211
rect -753 6763 73229 7206
rect -753 6455 35242 6763
rect 35750 6614 73229 6763
rect 35750 6455 67514 6614
rect -753 6371 67514 6455
rect -753 5969 31891 6371
rect 32314 6163 67514 6371
rect 32314 6075 44971 6163
rect 32314 5969 38422 6075
rect -753 5962 38422 5969
rect -753 5960 4747 5962
rect -753 5958 4001 5960
rect -753 5722 3274 5958
rect 3510 5724 4001 5958
rect 4237 5726 4747 5960
rect 4983 5726 5486 5962
rect 5722 5960 38422 5962
rect 5722 5958 8440 5960
rect 5722 5956 7706 5958
rect 5722 5951 6958 5956
rect 5722 5726 6217 5951
rect 4237 5724 6217 5726
rect 3510 5722 6217 5724
rect -753 5715 6217 5722
rect 6453 5720 6958 5951
rect 7194 5722 7706 5956
rect 7942 5724 8440 5958
rect 8676 5771 38422 5960
rect 38932 5890 44971 6075
rect 38932 5771 39871 5890
rect 8676 5724 39871 5771
rect 7942 5722 39871 5724
rect 7194 5720 39871 5722
rect 6453 5715 39871 5720
rect -753 5586 39871 5715
rect 40381 5586 41717 5890
rect 42227 5859 44971 5890
rect 45481 6095 58250 6163
rect 45481 5978 51625 6095
rect 45481 5859 46420 5978
rect 42227 5674 46420 5859
rect 46930 5674 48266 5978
rect 48776 5791 51625 5978
rect 52135 5910 58250 6095
rect 52135 5791 53074 5910
rect 48776 5674 53074 5791
rect 42227 5606 53074 5674
rect 53584 5606 54920 5910
rect 55430 5859 58250 5910
rect 58760 6157 67514 6163
rect 67751 6157 73229 6614
rect 58760 5978 73229 6157
rect 58760 5859 59699 5978
rect 55430 5674 59699 5859
rect 60209 5674 61545 5978
rect 62055 5765 73229 5978
rect 62055 5674 65851 5765
rect 55430 5606 65851 5674
rect 42227 5586 65851 5606
rect -753 5468 65851 5586
rect -753 5195 63847 5468
rect 64207 5426 65851 5468
rect 66224 5426 73229 5765
rect 64207 5195 73229 5426
rect -753 5150 73229 5195
rect -753 4819 72465 5150
rect 72709 4819 73229 5150
rect -753 4531 73229 4819
rect -753 4295 10020 4531
rect 10256 4529 73229 4531
rect 10256 4522 20361 4529
rect 10256 4519 18293 4522
rect 10256 4295 12093 4519
rect -753 4283 12093 4295
rect 12329 4283 14156 4519
rect 14392 4515 18293 4519
rect 14392 4283 16220 4515
rect -753 4279 16220 4283
rect 16456 4286 18293 4515
rect 18529 4293 20361 4522
rect 20597 4524 73229 4529
rect 20597 4293 22434 4524
rect 18529 4288 22434 4293
rect 22670 4515 73229 4524
rect 22670 4288 24501 4515
rect 18529 4286 24501 4288
rect 16456 4279 24501 4286
rect 24737 4279 73229 4515
rect -753 4272 73229 4279
rect -753 3870 31875 4272
rect 32298 3870 73229 4272
rect -753 3560 73229 3870
rect -753 3458 38421 3560
rect -753 3150 35218 3458
rect 35726 3256 38421 3458
rect 38931 3559 58249 3560
rect 38931 3558 51627 3559
rect 38931 3332 44972 3558
rect 38931 3322 41123 3332
rect 38931 3256 39989 3322
rect 35726 3150 39989 3256
rect -753 2812 39989 3150
rect 40293 2822 41123 3322
rect 41427 3254 44972 3332
rect 45482 3330 51627 3558
rect 45482 3320 47674 3330
rect 45482 3254 46540 3320
rect 41427 2822 46540 3254
rect 40293 2812 46540 2822
rect -753 2810 46540 2812
rect 46844 2820 47674 3320
rect 47978 3255 51627 3330
rect 52137 3331 58249 3559
rect 52137 3321 54329 3331
rect 52137 3255 53195 3321
rect 47978 2820 53195 3255
rect 46844 2811 53195 2820
rect 53499 2821 54329 3321
rect 54633 3256 58249 3331
rect 58759 3547 73229 3560
rect 58759 3332 63907 3547
rect 58759 3322 60951 3332
rect 58759 3256 59817 3322
rect 54633 2821 59817 3256
rect 53499 2812 59817 2821
rect 60121 2822 60951 3322
rect 61255 3274 63907 3332
rect 64267 3274 73229 3547
rect 61255 3119 73229 3274
rect 61255 2822 67514 3119
rect 60121 2812 67514 2822
rect 53499 2811 67514 2812
rect 46844 2810 67514 2811
rect -753 2662 67514 2810
rect 67751 2662 73229 3119
rect -753 2270 73229 2662
rect -753 2209 65851 2270
rect -753 1807 31880 2209
rect 32303 2001 65851 2209
rect 66224 2007 73229 2270
rect 66224 2001 72463 2007
rect 32303 1900 72463 2001
rect 32303 1807 38415 1900
rect -753 1596 38415 1807
rect 38925 1899 58243 1900
rect 38925 1898 51621 1899
rect 38925 1596 44966 1898
rect -753 1594 44966 1596
rect 45476 1595 51621 1898
rect 52131 1596 58243 1899
rect 58753 1676 72463 1900
rect 72707 1676 73229 2007
rect 58753 1596 73229 1676
rect 52131 1595 73229 1596
rect 45476 1594 73229 1595
rect -753 694 73229 1594
rect -753 386 35193 694
rect 35701 479 73229 694
rect 35701 386 63903 479
rect -753 295 63903 386
rect -753 231 38414 295
rect -753 226 7565 231
rect -753 -197 1239 226
rect 1875 -197 4439 226
rect 5075 -192 7565 226
rect 8201 -192 10640 231
rect 11276 -192 13830 231
rect 14466 226 38414 231
rect 14466 -192 17055 226
rect 5075 -197 17055 -192
rect 17691 -197 20176 226
rect 20812 224 38414 226
rect 20812 -197 23263 224
rect -753 -199 23263 -197
rect 23899 167 38414 224
rect 23899 -199 31885 167
rect -753 -235 31885 -199
rect 32308 -9 38414 167
rect 38924 294 58242 295
rect 38924 293 51620 294
rect 38924 110 44965 293
rect 38924 -9 39863 110
rect 32308 -194 39863 -9
rect 40373 -194 41709 110
rect 42219 -11 44965 110
rect 45475 108 51620 293
rect 45475 -11 46414 108
rect 42219 -194 46414 -11
rect 32308 -196 46414 -194
rect 46924 -196 48260 108
rect 48770 -10 51620 108
rect 52130 109 58242 294
rect 52130 -10 53069 109
rect 48770 -195 53069 -10
rect 53579 -195 54915 109
rect 55425 -9 58242 109
rect 58752 206 63903 295
rect 64263 206 73229 479
rect 58752 110 73229 206
rect 58752 -9 59691 110
rect 55425 -194 59691 -9
rect 60201 -194 61537 110
rect 62047 -194 73229 110
rect 55425 -195 73229 -194
rect 48770 -196 73229 -195
rect 32308 -235 73229 -196
rect -753 -523 73229 -235
rect -753 -831 41892 -523
rect 42400 -542 73229 -523
rect 42400 -831 48431 -542
rect -753 -850 48431 -831
rect 48939 -567 73229 -542
rect 48939 -850 55137 -567
rect -753 -875 55137 -850
rect 55645 -875 73229 -567
rect -753 -1111 73229 -875
rect -753 -1229 72465 -1111
rect -753 -1686 67514 -1229
rect 67751 -1442 72465 -1229
rect 72709 -1442 73229 -1111
rect 67751 -1686 73229 -1442
rect -753 -1922 73229 -1686
rect -753 -2324 31885 -1922
rect 32308 -2078 73229 -1922
rect 32308 -2324 65851 -2078
rect -753 -2374 65851 -2324
rect -753 -2647 63913 -2374
rect 64273 -2417 65851 -2374
rect 66224 -2417 73229 -2078
rect 64273 -2647 73229 -2417
rect -753 -3642 73229 -2647
rect -753 -3653 7568 -3642
rect -753 -4061 1240 -3653
rect 1879 -4061 4448 -3653
rect 5087 -4050 7568 -3653
rect 8207 -3663 73229 -3642
rect 8207 -3673 13834 -3663
rect 8207 -4050 10632 -3673
rect 5087 -4061 10632 -4050
rect -753 -4081 10632 -4061
rect 11271 -4071 13834 -3673
rect 14473 -3673 73229 -3663
rect 14473 -4071 17011 -3673
rect 11271 -4081 17011 -4071
rect 17650 -4081 20163 -3673
rect 20802 -4081 23319 -3673
rect 23958 -4081 73229 -3673
rect -753 -4363 73229 -4081
rect 28185 -6579 37415 -4363
<< labels >>
flabel locali -2413 2644 -1904 2784 1 FreeSans 800 0 0 0 opcode[2]
port 19 n
flabel locali -2401 -1160 -1892 -1020 1 FreeSans 800 0 0 0 opcode[3]
port 20 n
flabel metal1 -1683 18685 -1609 18752 1 FreeSans 400 0 0 0 B[0]
port 1 n
flabel metal1 -1683 18799 -1609 18866 1 FreeSans 400 0 0 0 B[1]
port 2 n
flabel metal1 -1684 18914 -1610 18981 1 FreeSans 400 0 0 0 B[2]
port 3 n
flabel metal1 -1684 19028 -1610 19095 1 FreeSans 400 0 0 0 B[3]
port 4 n
flabel metal1 -1684 19142 -1610 19209 1 FreeSans 400 0 0 0 B[4]
port 5 n
flabel metal1 -1684 19261 -1610 19328 1 FreeSans 400 0 0 0 B[5]
port 6 n
flabel metal1 -1684 19382 -1610 19449 1 FreeSans 400 0 0 0 B[6]
port 7 n
flabel metal1 -1684 19497 -1610 19564 1 FreeSans 400 0 0 0 B[7]
port 8 n
flabel metal1 -1686 24097 -1612 24164 1 FreeSans 400 0 0 0 A[0]
port 9 n
flabel metal1 -1686 23976 -1612 24043 1 FreeSans 400 0 0 0 A[1]
port 10 n
flabel metal1 -1686 23857 -1612 23924 1 FreeSans 400 0 0 0 A[2]
port 11 n
flabel metal1 -1686 23736 -1612 23803 1 FreeSans 400 0 0 0 A[3]
port 12 n
flabel metal1 -1686 23616 -1612 23683 1 FreeSans 400 0 0 0 A[4]
port 13 n
flabel metal1 -1686 23494 -1612 23561 1 FreeSans 400 0 0 0 A[5]
port 14 n
flabel metal1 -1686 23378 -1612 23445 1 FreeSans 400 0 0 0 A[6]
port 15 n
flabel metal1 -1686 23253 -1612 23320 1 FreeSans 400 0 0 0 A[7]
port 16 n
flabel metal1 -1682 22842 -1176 22979 1 FreeSans 400 0 0 0 opcode[1]
port 17 n
flabel metal1 -1680 22622 -1174 22759 1 FreeSans 400 0 0 0 opcode[0]
port 18 n
flabel metal1 2900 -4479 3022 -4296 1 FreeSans 400 0 0 0 Y[7]
port 21 n
flabel metal1 6047 -4472 6157 -4302 1 FreeSans 400 0 0 0 Y[6]
port 22 n
flabel metal1 9188 -4469 9298 -4299 1 FreeSans 400 0 0 0 Y[5]
port 23 n
flabel metal1 12324 -4464 12434 -4294 1 FreeSans 400 0 0 0 Y[4]
port 24 n
flabel metal1 15532 -4474 15642 -4304 1 FreeSans 400 0 0 0 Y[3]
port 25 n
flabel metal1 18675 -4459 18785 -4289 1 FreeSans 400 0 0 0 Y[2]
port 26 n
flabel metal1 21798 -4461 21908 -4291 1 FreeSans 400 0 0 0 Y[1]
port 27 n
flabel metal1 24945 -4456 25055 -4286 1 FreeSans 400 0 0 0 Y[0]
port 28 n
flabel metal1 38145 25345 38284 25474 1 FreeSans 400 0 0 0 Cout
port 29 n
flabel metal4 28947 24950 35877 26143 1 FreeSans 6400 0 0 0 VDD
port 30 n
flabel metal5 29061 -6255 36677 -4640 1 FreeSans 6400 0 0 0 VSS
port 31 n
<< end >>
