* NGSPICE file created from logic_unit.ext - technology: sky130B

.subckt logic_unit Y[1] Y[2] Y[3] Y[4] Y[5] A[4] A[5] A[6] A[0] A[1] A[2] A[3] A[7]
+ B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] opcode[1] opcode[0] Y[7] Y[6] Y[0] VSS VDD
X0 VDD B[7] a_20252_3694# VDD sky130_fd_pr__pfet_01v8 ad=1.45e+14p pd=1.13448e+09u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X1 VDD a_3891_1714# a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X2 a_3881_n3752# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X3 VSS A[0] a_n25_n6671# VSS sky130_fd_pr__nfet_01v8 ad=6.928e+13p pd=4.5344e+08u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X4 VDD A[7] a_10615_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X5 VDD opcode[0] a_3392_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X6 a_12813_n7362# a_12386_n6669# a_12931_n7362# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X7 a_3891_n1020# a_4290_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X8 VDD B[7] a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X9 a_10852_3062# A[7] a_10615_3699# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X10 VDD a_3891_n1020# a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X11 a_20054_n990# opcode[1] a_20290_n2323# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X12 a_4290_n3726# a_2588_n7362# a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X13 VDD a_747_1714# a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X14 a_10217_n3722# a_6725_n7362# a_10566_n3722# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X15 VDD opcode[1] a_3392_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X16 a_21997_n6357# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X17 a_17916_3694# A[5] a_17798_3694# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X18 a_7083_n990# a_7023_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X19 a_10576_n990# opcode[1] a_10812_n2323# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X20 VDD A[5] a_7669_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X21 a_2588_n7362# a_2043_n6669# a_2588_n8094# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X22 VSS a_6725_n7362# a_11038_n5055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X23 a_7906_3060# A[5] a_7669_3697# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X24 a_7083_1744# a_7023_1718# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X25 VDD A[1] a_3881_n3752# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VDD a_747_n1020# a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X27 Y[6] a_20054_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X28 VDD a_10566_n3722# a_10167_n1016# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X29 VDD a_4290_n3726# a_3891_n1020# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 a_747_1714# a_11952_3694# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X31 a_3951_1740# a_3392_1740# a_4300_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X32 a_20579_n1475# a_20054_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X33 a_15293_n7386# B[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X34 a_1382_n5059# a_737_n3752# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X35 a_1156_1740# a_897_3260# a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X36 a_20526_n2323# a_19146_n990# a_20054_n990# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X37 VSS B[7] a_20134_3694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X38 a_10566_n3722# a_6725_n7362# a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_9668_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X40 VSS opcode[1] a_3392_n994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X41 a_4951_n7390# B[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X42 a_3951_n994# a_3392_n994# a_4300_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X43 a_22839_n3722# a_21997_n6357# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X44 a_9668_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X45 a_1156_n994# a_1681_n1479# a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X46 a_2824_n8094# A[1] a_2588_n7362# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X47 VDD B[4] a_16748_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X48 VSS a_14303_n1479# a_14250_n2327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X49 a_10167_n1016# a_10566_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 a_3891_n1020# a_4290_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 a_13369_1714# a_16630_3696# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X52 a_1146_n3726# opcode[0] a_1382_n5059# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X53 a_10227_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X54 VSS a_20579_n1475# a_20526_n2323# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 a_10227_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X56 Y[1] a_4300_n994# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X57 a_15574_3694# B[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X58 VDD a_7432_n990# Y[2] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X59 a_13238_3694# A[1] a_13120_3694# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X60 VDD a_7432_1744# a_7957_n1475# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X61 VSS B[1] a_2824_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X62 VDD B[1] a_1755_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X63 a_17158_n2327# a_16513_n1020# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X64 VSS a_23723_n1475# a_23670_n2323# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X65 Y[2] a_7432_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 a_7957_n1475# a_7432_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 a_737_n3752# A[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X68 VSS A[4] a_8249_n6669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X69 a_6221_3697# B[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X70 a_5291_3262# a_4701_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X71 a_15293_n7386# B[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X72 a_2470_n7362# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X73 a_9757_3262# a_9167_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X74 VSS B[3] a_15456_3694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X75 VDD opcode[1] a_22290_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X76 VDD a_13120_3694# a_3891_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X77 VDD a_15456_3694# a_10167_1718# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X78 a_16014_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X79 a_21997_n6357# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_4762_n5059# a_3382_n3726# a_4290_n3726# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X81 VDD opcode[0] a_22290_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X82 a_10227_n990# a_10167_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X83 a_10227_1744# a_10167_1718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X84 a_16014_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X85 a_7013_n3748# A[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X86 VDD opcode[0] a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X87 a_7083_n990# a_7023_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 a_13167_n8094# A[6] a_12931_n7362# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X89 a_7083_1744# a_7023_1718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 VSS opcode[0] a_16004_n3726# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X91 VDD opcode[0] a_16004_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X92 Y[6] a_20054_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X93 a_807_1740# a_248_1740# a_1156_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X94 VDD a_13778_1740# a_14303_n1479# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X95 VSS a_8259_3260# a_17394_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X96 VDD opcode[1] a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X97 VSS a_2588_n7362# a_4762_n5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X98 VDD opcode[0] a_248_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X99 a_22849_n990# a_22290_n990# a_23198_n990# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X100 a_14881_n7360# a_14454_n6667# a_14999_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X101 a_11038_n5055# a_9658_n3722# a_10566_n3722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X102 a_20579_n1475# a_20054_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X103 a_4825_n1479# a_4300_1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X104 VSS a_5291_3262# a_11048_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X105 a_13369_n1020# a_13768_n3726# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X106 a_1156_1740# a_897_3260# a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X107 a_22849_1744# a_22290_1744# a_23198_1744# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X108 VDD B[5] a_17916_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 a_807_n994# a_248_n994# a_1156_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X110 VDD a_13778_n994# Y[4] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X111 VDD A[6] a_19635_n3748# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X112 VDD A[2] a_4112_n6671# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X113 VDD opcode[1] a_248_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X114 VSS B[6] a_13167_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 a_10167_n1016# a_10566_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X116 a_1156_n994# a_1681_n1479# a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X117 a_402_n7364# a_814_n7390# a_520_n7364# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=1.74e+12p ps=1.374e+07u w=2e+06u l=300000u
X118 a_16513_n1020# a_16912_n3726# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X119 a_14406_3692# A[2] a_14288_3692# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X120 a_6961_n8094# A[3] a_6725_n7362# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X121 VDD B[5] a_11156_n7386# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X122 a_7422_n3722# a_4657_n7364# a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X123 a_20290_411# a_19230_3112# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X124 a_3843_3262# a_3253_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X125 a_14999_n7360# a_14454_n6667# a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X126 VSS opcode[0] a_238_n3726# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X127 VDD a_13369_1714# a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X128 a_19635_n3748# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X129 a_12931_n8094# a_13225_n7388# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X130 a_7083_n990# a_7957_n1475# a_7432_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X131 a_737_n3752# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X132 VSS opcode[1] a_19146_n990# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X133 a_520_n7364# a_814_n7390# a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X134 a_12070_3694# A[0] a_11952_3694# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X135 a_11156_n7386# B[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X136 a_7073_n3722# a_4657_n7364# a_7422_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X137 a_7083_1744# a_3843_3262# a_7432_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X138 VDD a_13369_n1020# a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X139 a_13419_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X140 a_897_3260# a_307_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X141 a_4701_3699# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X142 VSS opcode[1] a_9668_n990# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X143 a_14881_n7360# a_15293_n7386# a_14999_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X144 a_19645_n1016# a_20044_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X145 VSS opcode[0] a_22290_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X146 Y[0] a_1156_n994# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X147 a_2588_n7362# a_2043_n6669# a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X148 a_19695_n3722# a_19136_n3722# a_20044_n3722# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X149 a_6811_3260# a_6221_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X150 a_20252_3694# A[7] a_20134_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X151 a_23188_n3722# a_14999_n7360# a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X152 VDD A[6] a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X153 VDD A[0] a_737_n3752# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 a_6607_n7362# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X155 VSS B[1] a_13120_3694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X156 a_19705_n990# a_19645_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X157 a_7422_n3722# a_4657_n7364# a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X158 Y[3] a_10576_n990# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X159 a_19705_1744# a_19230_3112# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X160 a_2470_n7362# a_2043_n6669# a_2588_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X161 a_20044_n3722# a_19136_n3722# a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X162 a_22839_n3722# a_14999_n7360# a_23188_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X163 a_11101_n1475# a_10576_1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X164 a_10227_n990# a_10167_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 VSS A[3] a_6180_n6669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X166 a_12813_n7362# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X167 a_13778_1740# a_6811_3260# a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X168 VDD opcode[1] a_6524_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X169 VDD a_7422_n3722# a_7023_n1016# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X170 a_10227_1744# a_10167_1718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X171 a_11205_3262# a_10615_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X172 a_807_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X173 VDD opcode[0] a_6524_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X174 VDD A[3] a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X175 a_16922_1740# a_16014_1740# a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X176 a_13778_n994# a_14303_n1479# a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X177 a_20054_n990# a_20579_n1475# a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X178 a_16922_1740# a_8259_3260# a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X179 a_20054_1744# a_9757_3262# a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X180 a_16912_n3726# a_10862_n7360# a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X181 VDD B[5] a_17916_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 a_807_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X183 a_8259_3260# a_7669_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X184 a_8794_n8094# a_9088_n7388# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X185 a_14999_n7360# a_14454_n6667# a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 a_2588_n7362# a_2043_n6669# a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X187 VSS opcode[0] a_248_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X188 a_16922_n994# a_16014_n994# a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X189 a_23198_n990# a_23723_n1475# a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X190 a_10862_n7360# a_10317_n6667# a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X191 VDD B[6] a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X192 a_16922_n994# a_17447_n1479# a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X193 a_19084_3696# A[6] a_18966_3696# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X194 a_7073_n3722# a_6514_n3722# a_7422_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X195 a_23198_1744# a_11205_3262# a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X196 a_1392_n2327# a_747_n1020# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X197 a_4825_n1479# a_4300_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X198 VDD a_16912_n3726# a_16513_n1020# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X199 a_10576_n990# a_9668_n990# a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X200 Y[2] a_7432_n990# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X201 a_10576_1744# a_9668_1744# a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X202 a_17447_n1479# a_16922_1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X203 VDD a_18966_3696# a_19230_3112# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X204 VDD opcode[1] a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X205 a_10227_n990# a_11101_n1475# a_10576_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 Y[1] a_4300_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X207 a_2470_n7362# a_2882_n7388# a_2588_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X208 a_7422_n3722# opcode[0] a_7658_n5055# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X209 a_16513_1714# a_17798_3694# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X210 VDD opcode[0] a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X211 a_10227_1744# a_5291_3262# a_10576_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X212 VDD A[7] a_14454_n6667# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X213 a_1755_3697# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X214 a_10744_n7360# a_10317_n6667# a_10862_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X215 VDD A[5] a_10317_n6667# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X216 a_12070_3694# A[0] a_11952_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X217 a_797_n3726# a_520_n7364# a_1146_n3726# VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=300000u
X218 a_10157_n3748# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X219 a_814_n7390# B[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X220 VSS opcode[0] a_16014_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X221 a_1156_n994# opcode[1] a_1392_n2327# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X222 a_4701_3699# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X223 VDD opcode[0] a_12870_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X224 a_23424_n5055# a_21997_n6357# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X225 VDD opcode[0] a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X226 VSS B[3] a_4938_3062# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X227 a_7013_n3748# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X228 a_13768_n3726# opcode[0] a_14004_n5059# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X229 VDD a_16630_3696# a_13369_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X230 a_8676_n7362# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.206e+07u as=0p ps=0u w=2e+06u l=300000u
X231 VDD A[6] a_9167_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X232 VDD opcode[1] a_12870_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X233 a_7894_n5055# a_6514_n3722# a_7422_n3722# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X234 a_10217_n3722# a_10157_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X235 a_9404_3062# A[6] a_9167_3699# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X236 VDD opcode[0] a_16014_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X237 a_21997_n6357# A[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X238 a_16912_n3726# opcode[0] a_17148_n5059# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X239 a_1146_n3726# a_520_n7364# a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X240 a_14999_n7360# a_14454_n6667# a_14999_n8092# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X241 a_12813_n7362# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X242 VSS B[2] a_14288_3692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X243 VSS a_2345_3260# a_4772_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X244 a_13768_n3726# a_8794_n7362# a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=300000u
X245 a_12931_n7362# a_12386_n6669# a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X246 a_23188_n3722# opcode[0] a_23424_n5055# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X247 VDD opcode[1] a_16014_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X248 a_13359_n3752# A[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X249 VDD a_14288_3692# a_7023_1718# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X250 a_14240_n5059# a_12860_n3726# a_13768_n3726# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X251 a_3843_3262# a_3253_3699# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X252 VDD B[4] a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X253 a_13778_1740# a_6811_3260# a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X254 a_19146_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X255 a_4772_n2327# a_3392_n994# a_4300_n994# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X256 VDD a_3881_n3752# a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X257 VDD B[5] a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X258 VSS a_4657_n7364# a_7894_n5055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X259 VDD a_10157_n3748# a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X260 VSS A[6] a_12386_n6669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X261 a_11205_3262# a_10615_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X262 VDD opcode[0] a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X263 a_19146_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X264 a_19705_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X265 a_17384_n5059# a_16004_n3726# a_16912_n3726# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X266 a_19705_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X267 a_11048_411# a_9668_1744# a_10576_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X268 a_15235_n8092# A[7] a_14999_n7360# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X269 a_13778_n994# a_14303_n1479# a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X270 a_13419_n3726# a_8794_n7362# a_13768_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X271 a_17394_407# a_16014_1740# a_16922_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X272 a_12813_n7362# a_13225_n7388# a_12931_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X273 VDD a_20134_3694# a_20398_3112# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X274 VDD opcode[1] a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X275 a_3253_3699# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=300000u
X276 a_22849_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X277 VDD opcode[0] a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X278 VSS B[2] a_3490_3062# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X279 a_16630_3696# A[4] a_16748_3696# VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X280 a_22849_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X281 a_6725_n7362# a_6180_n6669# a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X282 a_8676_n7362# B[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X283 a_402_n7364# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X284 VSS a_4825_n1479# a_4772_n2327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X285 VSS B[3] a_6961_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X286 a_16563_n3726# a_10862_n7360# a_16912_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X287 a_10217_n3722# a_10157_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X288 a_1681_n1479# a_1156_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X289 VDD B[2] a_3253_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X290 a_19084_3696# B[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X291 Y[7] a_23198_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X292 a_11048_n2323# a_9668_n990# a_10576_n990# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X293 VDD opcode[1] a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X294 a_814_n7390# B[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X295 VSS a_10862_n7360# a_17384_n5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X296 a_23723_n1475# a_23198_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X297 VDD opcode[1] a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X298 VSS B[7] a_15235_n8092# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X299 a_14406_3692# B[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X300 a_4300_1740# a_2345_3260# a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X301 a_3881_n3752# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X302 Y[0] a_1156_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X303 a_12931_n7362# a_13225_n7388# a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X304 VDD a_18966_3696# a_19230_3112# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X305 VDD opcode[0] a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X306 a_238_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X307 a_3941_n3726# a_3382_n3726# a_4290_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X308 a_5291_3262# a_4701_3699# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X309 VSS opcode[0] a_6514_n3722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X310 a_18966_3696# A[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X311 a_4300_n994# a_4825_n1479# a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X312 VDD B[4] a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X313 VDD A[0] a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X314 a_15456_3694# A[3] a_15574_3694# VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X315 a_6725_n8094# a_7019_n7388# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=300000u
X316 VDD A[0] a_307_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=300000u
X317 VSS opcode[0] a_12870_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X318 a_2588_n8094# a_2882_n7388# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X319 a_544_3060# A[0] a_307_3697# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X320 a_3881_n3752# A[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X321 VDD B[0] a_814_n7390# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X322 a_1755_3697# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X323 VSS B[6] a_18966_3696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X324 VDD A[4] a_6221_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X325 a_12813_n7362# a_13225_n7388# a_12931_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X326 a_6458_3060# A[4] a_6221_3697# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X327 a_22849_n990# a_22789_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X328 VDD opcode[0] a_238_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X329 a_4290_n3726# a_3382_n3726# a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X330 a_22849_1744# a_20398_3112# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X331 a_13359_n3752# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X332 a_1618_n5059# a_238_n3726# a_1146_n3726# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X333 a_402_n7364# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X334 a_14004_n5059# a_13359_n3752# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X335 a_19136_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X336 a_4300_1740# opcode[0] a_4536_407# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X337 a_7957_n1475# a_7432_1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X338 VDD B[3] a_4701_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X339 a_20252_3694# B[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X340 a_747_n1020# a_1146_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X341 VDD A[4] a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X342 a_814_n7390# B[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X343 a_10615_3699# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X344 a_3392_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X345 a_13225_n7388# B[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X346 VSS opcode[0] a_22280_n3722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X347 VSS opcode[0] a_6524_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X348 a_807_1740# a_747_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X349 a_3941_n3726# a_3382_n3726# a_4290_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X350 a_3392_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X351 VDD A[4] a_13359_n3752# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 VSS a_520_n7364# a_1618_n5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X353 a_16563_n3726# a_16004_n3726# a_16912_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X354 a_7669_3697# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X355 VDD B[0] a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X356 VDD opcode[0] a_19136_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X357 a_17158_407# a_16513_1714# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X358 a_14250_407# a_12870_1740# a_13778_1740# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X359 a_807_n994# a_747_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X360 VDD opcode[1] a_6524_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X361 Y[5] a_16922_n994# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X362 VDD a_1146_n3726# a_747_n1020# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X363 a_8794_n7362# a_9088_n7388# a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=300000u
X364 VDD opcode[0] a_6524_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X365 VDD B[6] a_13225_n7388# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X366 VDD B[5] a_7669_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X367 VSS B[0] a_11952_3694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X368 VDD a_20134_3694# a_20398_3112# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 a_20134_3694# A[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X370 VSS opcode[1] a_248_n994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X371 a_10862_n7360# a_10317_n6667# a_10862_n8092# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X372 VDD opcode[1] a_9668_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X373 a_7669_3697# B[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X374 VSS a_897_3260# a_1628_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X375 VDD B[3] a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X376 a_3951_1740# a_3392_1740# a_4300_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X377 VDD opcode[0] a_9668_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X378 VDD a_16922_1740# a_17447_n1479# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X379 a_19635_n3748# A[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X380 a_23198_n990# a_23723_n1475# a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X381 a_7073_n3722# a_7013_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X382 a_747_n1020# a_1146_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X383 a_2345_3260# a_1755_3697# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X384 a_7668_n2323# a_7023_n1016# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X385 a_9088_n7388# B[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X386 a_8676_n7362# a_9088_n7388# a_8794_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X387 a_23198_1744# a_11205_3262# a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X388 VSS B[4] a_16630_3696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X389 a_3951_n994# a_3392_n994# a_4300_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X390 VDD a_16922_n994# Y[5] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X391 a_4300_1740# a_2345_3260# a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X392 a_10862_n7360# a_10317_n6667# a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 VDD a_17798_3694# a_16513_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X394 VDD B[3] a_15574_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X395 a_4657_n7364# a_4112_n6671# a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=1.74e+12p pd=1.374e+07u as=4.06e+12p ps=3.206e+07u w=2e+06u l=300000u
X396 a_6607_n7362# B[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X397 a_4112_n6671# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X398 a_4300_n994# a_4825_n1479# a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X399 a_9088_n7388# B[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X400 VDD a_7013_n3748# a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X401 VDD B[0] a_307_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X402 a_10576_1744# opcode[0] a_10812_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X403 a_7432_n990# opcode[1] a_7668_n2323# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X404 a_13238_3694# B[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X405 Y[3] a_10576_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X406 VDD B[1] a_1755_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X407 VDD B[4] a_6221_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X408 VDD a_15456_3694# a_10167_1718# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X409 a_11101_n1475# a_10576_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X410 a_10744_n7360# a_11156_n7386# a_10862_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X411 VDD opcode[0] a_22280_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X412 VDD a_16513_1714# a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X413 a_12860_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X414 VDD a_4701_3699# a_5291_3262# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X415 a_23434_n2323# a_22789_n1016# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X416 a_737_n3752# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X417 a_15456_3694# A[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X418 a_22290_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X419 a_10217_n3722# a_9658_n3722# a_10566_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X420 VDD opcode[0] a_6514_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X421 a_3891_1714# a_13120_3694# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X422 a_10167_1718# a_15456_3694# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X423 VDD opcode[0] a_16014_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X424 a_13778_n994# opcode[1] a_14014_n2327# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X425 VDD A[6] a_12386_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X426 VDD B[4] a_9088_n7388# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X427 a_22290_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X428 a_4772_407# a_3392_1740# a_4300_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X429 VDD a_16513_n1020# a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X430 a_7904_n2323# a_6524_n990# a_7432_n990# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X431 a_14881_n7360# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X432 VDD opcode[1] a_16014_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X433 a_13429_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X434 a_16922_n994# opcode[1] a_17158_n2327# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X435 a_10862_n7360# a_11156_n7386# a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X436 a_22280_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X437 VSS B[7] a_10852_3062# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X438 VDD opcode[0] a_12860_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X439 VSS opcode[0] a_12860_n3726# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X440 a_7023_n1016# a_7422_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_23198_n990# opcode[1] a_23434_n2323# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X442 a_14250_n2327# a_12870_n994# a_13778_n994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X443 a_10566_n3722# a_9658_n3722# a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X444 a_248_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X445 a_1156_1740# a_248_1740# a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X446 a_14303_n1479# a_13778_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X447 a_13429_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 a_12386_n6669# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X449 VSS A[1] a_2043_n6669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X450 a_9088_n7388# B[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X451 a_807_1740# a_897_3260# a_1156_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X452 a_16573_1740# a_16014_1740# a_16922_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X453 a_1681_n1479# a_1156_1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X454 a_16922_1740# opcode[0] a_17158_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X455 VSS a_7957_n1475# a_7904_n2323# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X456 a_6607_n7362# a_7019_n7388# a_6725_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X457 VDD A[1] a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X458 a_20398_3112# a_20134_3694# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X459 a_1156_n994# a_248_n994# a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X460 a_248_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X461 Y[4] a_13778_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X462 a_3253_3699# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X463 a_22849_n990# a_22290_n990# a_23198_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X464 a_17394_n2327# a_16014_n994# a_16922_n994# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X465 a_10744_n7360# a_11156_n7386# a_10862_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X466 VDD opcode[0] a_22280_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X467 a_897_3260# a_307_3697# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X468 a_807_n994# a_1681_n1479# a_1156_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X469 a_16573_n994# a_16014_n994# a_16922_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X470 a_19695_n3722# a_19136_n3722# a_20044_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X471 a_22849_1744# a_22290_1744# a_23198_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X472 a_19645_n1016# a_20044_n3722# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X473 a_10217_n3722# a_9658_n3722# a_10566_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X474 VDD a_3253_3699# a_3843_3262# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X475 VDD A[6] a_12386_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X476 a_3951_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X477 a_6607_n7362# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X478 a_897_3260# a_307_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X479 a_14406_3692# A[2] a_14288_3692# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X480 VSS B[5] a_17798_3694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X481 a_6725_n7362# a_7019_n7388# a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X482 a_2470_n7362# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X483 a_13429_1740# a_13369_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X484 VSS a_3843_3262# a_7904_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X485 a_2588_n7362# a_2882_n7388# a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X486 a_520_n7364# a_n25_n6671# a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 a_22789_n1016# a_23188_n3722# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X488 a_3951_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X489 VSS a_17447_n1479# a_17394_n2327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X490 a_n25_n6671# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X491 a_7432_n990# a_7957_n1475# a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X492 VDD opcode[0] a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X493 VDD a_17798_3694# a_16513_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X494 VDD A[4] a_8249_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X495 a_7432_1744# a_3843_3262# a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X496 a_13429_n994# a_13369_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X497 a_7422_n3722# a_6514_n3722# a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X498 VDD B[0] a_307_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X499 VSS a_6811_3260# a_14250_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X500 a_7019_n7388# B[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X501 a_6607_n7362# a_7019_n7388# a_6725_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X502 a_11205_3262# a_10615_3699# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X503 VDD B[2] a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X504 VDD a_1755_3697# a_2345_3260# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X505 a_4536_407# a_3891_1714# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X506 a_19695_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X507 a_8249_n6669# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X508 a_7023_1718# a_14288_3692# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X509 a_3951_1740# a_3891_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X510 VDD opcode[0] a_12860_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X511 a_7019_n7388# B[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X512 a_1628_n2327# a_248_n994# a_1156_n994# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X513 a_14014_n2327# a_13369_n1020# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X514 a_2882_n7388# B[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X515 a_22839_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X516 a_16912_n3726# a_16004_n3726# a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X517 VDD A[2] a_7013_n3748# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X518 a_3951_n994# a_3891_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X519 a_19705_n990# a_19645_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X520 VDD opcode[0] a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X521 a_20054_n990# a_20579_n1475# a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X522 a_3941_n3726# a_3881_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X523 a_14999_n7360# a_15293_n7386# a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X524 a_19705_1744# a_19230_3112# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X525 a_4539_n7364# B[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X526 a_16563_n3726# a_16503_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X527 VDD B[7] a_10615_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X528 a_20054_1744# a_9757_3262# a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X529 a_20054_n990# a_19146_n990# a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X530 VDD opcode[0] a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X531 a_13369_n1020# a_13768_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X532 VDD opcode[0] a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X533 VDD A[4] a_8249_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X534 a_20054_1744# a_19146_1744# a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X535 a_13778_1740# opcode[0] a_14014_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X536 a_19705_n990# a_20579_n1475# a_20054_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X537 VDD B[3] a_7019_n7388# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X538 a_19705_1744# a_9757_3262# a_20054_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X539 VSS a_1681_n1479# a_1628_n2327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X540 a_11098_n8092# A[5] a_10862_n7360# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X541 a_17916_3694# B[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X542 VDD opcode[1] a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X543 VDD B[1] a_2882_n7388# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X544 VDD opcode[0] a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 a_7013_n3748# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X546 VSS a_8794_n7362# a_14240_n5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X547 VSS opcode[1] a_6524_n990# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X548 VSS opcode[0] a_19146_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X549 VDD B[2] a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 a_22789_n1016# a_23188_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X551 VDD a_16503_n3752# a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 a_18966_3696# A[6] a_19084_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X553 a_1628_407# a_248_1740# a_1156_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X554 VSS a_11101_n1475# a_11048_n2323# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X555 VDD a_13768_n3726# a_13369_n1020# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X556 a_8259_3260# a_7669_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X557 a_10227_n990# a_9668_n990# a_10576_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X558 a_7019_n7388# B[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X559 a_10227_1744# a_9668_1744# a_10576_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X560 VSS B[5] a_11098_n8092# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X561 a_13768_n3726# a_8794_n7362# a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X562 a_7083_n990# a_6524_n990# a_7432_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X563 a_4825_n1479# a_4300_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X564 a_7083_1744# a_6524_1744# a_7432_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X565 VDD opcode[0] a_12870_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X566 a_14303_n1479# a_13778_1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X567 a_13429_1740# a_13369_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X568 VDD a_23188_n3722# a_22789_n1016# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X569 a_11952_3694# A[0] a_12070_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X570 a_20280_n5055# a_19635_n3748# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X571 a_13369_n1020# a_13768_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X572 VDD A[3] a_4701_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X573 Y[1] a_4300_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X574 a_12870_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X575 VDD opcode[1] a_12870_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X576 a_12813_n7362# B[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 a_4938_3062# A[3] a_4701_3699# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X578 a_10812_411# a_10167_1718# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X579 a_13429_n994# a_13369_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X580 VSS opcode[1] a_22290_n990# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X581 a_13369_1714# a_16630_3696# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X582 a_10862_n8092# a_11156_n7386# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X583 a_12070_3694# B[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X584 a_13225_n7388# B[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X585 a_16513_n1020# a_16912_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X586 a_9167_3699# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X587 a_12870_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X588 a_9757_3262# a_9167_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X589 a_20134_3694# A[7] a_20252_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X590 a_22789_n1016# a_23188_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X591 a_14288_3692# A[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X592 VDD a_11952_3694# a_747_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X593 VDD A[3] a_6180_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X594 VDD B[6] a_9167_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X595 VSS a_11205_3262# a_23670_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X596 a_520_n7364# a_n25_n6671# a_520_n8096# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X597 a_6811_3260# a_6221_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X598 a_13778_1740# a_12870_1740# a_13429_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X599 VDD A[1] a_2043_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X600 a_4657_n7364# a_4112_n6671# a_4657_n8096# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2e+06u l=300000u
X601 VDD opcode[1] a_19146_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X602 VDD opcode[1] a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X603 a_13429_1740# a_12870_1740# a_13778_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X604 VDD opcode[0] a_19146_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X605 a_13778_n994# a_12870_n994# a_13429_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X606 VDD opcode[0] a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X607 a_10167_n1016# a_10566_n3722# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X608 a_6180_n6669# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X609 a_13225_n7388# B[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X610 a_756_n8096# A[0] a_520_n7364# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X611 VDD opcode[0] a_807_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X612 a_13429_n994# a_12870_n994# a_13778_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X613 a_11952_3694# A[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X614 a_16573_1740# a_16014_1740# a_16922_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X615 a_10744_n7360# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X616 a_4893_n8096# A[2] a_4657_n7364# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X617 a_23660_n5055# a_22280_n3722# a_23188_n3722# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X618 VDD a_1156_1740# a_1681_n1479# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X619 VDD opcode[1] a_807_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X620 a_3253_3699# B[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X621 VDD B[6] a_19084_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X622 a_16573_n994# a_16014_n994# a_16922_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X623 a_13359_n3752# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X624 a_402_n7364# B[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X625 VDD opcode[0] a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 a_23198_1744# opcode[0] a_23434_411# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X627 VDD opcode[0] a_3382_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X628 VDD A[3] a_6180_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X629 VDD a_1156_n994# Y[0] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X630 a_797_n3726# a_238_n3726# a_1146_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X631 Y[7] a_23198_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X632 a_4290_n3726# a_2588_n7362# a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X633 a_16503_n3752# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=300000u
X634 VDD opcode[1] a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X635 a_16748_3696# B[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X636 a_23723_n1475# a_23198_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X637 a_7904_411# a_6524_1744# a_7432_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X638 VSS B[2] a_4893_n8096# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X639 a_9757_3262# a_9167_3699# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X640 a_15574_3694# A[3] a_15456_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X641 a_307_3697# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 a_10217_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X643 a_13120_3694# A[1] a_13238_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X644 VDD A[1] a_1755_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X645 a_797_n3726# a_737_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X646 a_2470_n7362# B[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X647 a_1992_3060# A[1] a_1755_3697# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X648 a_1146_n3726# a_238_n3726# a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X649 VDD B[2] a_4951_n7390# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X650 a_3941_n3726# a_2588_n7362# a_4290_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X651 a_14999_n8092# a_15293_n7386# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X652 a_23723_n1475# a_23198_1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X653 VSS B[1] a_1992_3060# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X654 a_8794_n7362# a_8249_n6669# a_8794_n8094# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X655 a_4701_3699# B[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X656 VDD B[7] a_20252_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X657 VSS opcode[1] a_12870_n994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X658 VSS a_9757_3262# a_20526_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X659 VDD B[6] a_9167_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X660 VDD a_11952_3694# a_747_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X661 a_1156_1740# opcode[0] a_1392_407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X662 VDD a_737_n3752# a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X663 VDD B[1] a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X664 a_7073_n3722# a_7013_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X665 a_3951_1740# a_3891_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X666 a_797_n3726# a_238_n3726# a_1146_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X667 VSS A[2] a_4112_n6671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X668 a_4951_n7390# B[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X669 a_19695_n3722# a_19635_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X670 VSS opcode[1] a_16014_n994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X671 VDD A[7] a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 a_10615_3699# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X673 a_3951_n994# a_3891_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X674 Y[4] a_13778_n994# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X675 a_9030_n8094# A[4] a_8794_n7362# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X676 a_10744_n7360# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X677 a_807_1740# a_747_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X678 VDD opcode[1] a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X679 Y[6] a_20054_n990# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X680 a_17798_3694# A[5] a_17916_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X681 a_20398_3112# a_20134_3694# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X682 VDD a_7023_n1016# a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X683 a_797_n3726# a_737_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X684 a_7669_3697# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 VDD opcode[0] a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X686 VDD a_7023_1718# a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X687 VDD a_19635_n3748# a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X688 VSS B[5] a_7906_3060# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X689 a_807_n994# a_747_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X690 a_14881_n7360# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X691 VDD a_20054_n990# Y[6] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X692 a_17916_3694# A[5] a_17798_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X693 Y[7] a_23198_n990# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X694 VDD a_20054_1744# a_20579_n1475# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X695 a_4300_1740# a_3392_1740# a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X696 VDD A[5] a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X697 a_4526_n5059# a_3881_n3752# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X698 VDD opcode[0] a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X699 VDD opcode[1] a_9668_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X700 a_10157_n3748# A[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X701 a_3843_3262# a_3253_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X702 VDD B[6] a_19084_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X703 VDD opcode[0] a_9668_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X704 a_4300_n994# a_3392_n994# a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X705 a_23670_411# a_22290_1744# a_23198_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X706 a_19695_n3722# a_19635_n3748# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X707 a_3951_1740# a_2345_3260# a_4300_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X708 VDD B[7] a_14881_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X709 a_6811_3260# a_6221_3697# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X710 a_7083_n990# a_6524_n990# a_7432_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X711 a_8676_n7362# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X712 a_7083_1744# a_6524_1744# a_7432_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X713 VDD opcode[1] a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X714 Y[3] a_10576_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X715 a_3951_n994# a_4825_n1479# a_4300_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X716 a_4290_n3726# opcode[0] a_4526_n5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X717 VDD opcode[0] a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X718 a_11101_n1475# a_10576_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 a_3941_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X720 VDD opcode[0] a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X721 VDD B[1] a_13238_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X722 VDD a_10576_n990# Y[3] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X723 VSS B[0] a_544_3060# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X724 a_1755_3697# B[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X725 a_20579_n1475# a_20054_1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X726 a_12931_n7362# a_12386_n6669# a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X727 VDD a_10576_1744# a_11101_n1475# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X728 VDD B[1] a_2470_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X729 VDD a_22789_n1016# a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X730 a_20290_n2323# a_19645_n1016# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X731 VSS B[4] a_6458_3060# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X732 a_16573_1740# a_16513_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X733 a_2882_n7388# B[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X734 a_2470_n7362# a_2882_n7388# a_2588_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X735 a_5291_3262# a_4701_3699# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X736 VDD a_20398_3112# a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X737 a_402_n7364# a_n25_n6671# a_520_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 VDD A[0] a_n25_n6671# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X739 a_10566_n3722# a_6725_n7362# a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X740 VDD opcode[1] a_22290_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X741 VDD a_13120_3694# a_3891_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X742 VDD B[4] a_6221_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X743 a_13120_3694# A[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X744 VDD opcode[0] a_22290_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X745 a_22849_n990# a_22789_n1016# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X746 a_4539_n7364# a_4112_n6671# a_4657_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X747 a_16573_n994# a_16513_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X748 VDD B[3] a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X749 VDD A[2] a_4112_n6671# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X750 a_8259_3260# a_7669_3697# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X751 a_22849_1744# a_20398_3112# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X752 a_13419_n3726# a_13359_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X753 VDD a_9167_3699# a_9757_3262# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 a_10167_1718# a_15456_3694# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X755 a_19635_n3748# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X756 a_19695_n3722# a_12931_n7362# a_20044_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 VDD a_10167_n1016# a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X758 a_11156_n7386# B[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X759 a_520_n7364# a_n25_n6671# a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X760 a_807_1740# a_248_1740# a_1156_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X761 VDD a_10167_1718# a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X762 a_6725_n7362# a_6180_n6669# a_6725_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X763 VDD opcode[0] a_248_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X764 a_4657_n7364# a_4112_n6671# a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X765 a_22839_n3722# a_21997_n6357# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X766 a_6524_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X767 VDD a_13359_n3752# a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X768 a_807_n994# a_248_n994# a_1156_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X769 a_6524_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X770 a_14303_n1479# a_13778_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X771 VDD opcode[1] a_248_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X772 VDD B[5] a_7669_3697# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X773 a_23198_n990# a_22290_n990# a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X774 VSS A[7] a_14454_n6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X775 a_20044_n3722# a_12931_n7362# a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X776 VDD opcode[0] a_6514_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X777 a_23198_1744# a_22290_1744# a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X778 VSS A[5] a_10317_n6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X779 a_14881_n7360# a_15293_n7386# a_14999_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X780 a_23434_411# a_20398_3112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X781 Y[4] a_13778_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X782 VDD opcode[0] a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X783 a_17447_n1479# a_16922_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X784 a_4539_n7364# a_4951_n7390# a_4657_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X785 VDD B[0] a_402_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X786 a_23188_n3722# a_14999_n7360# a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X787 VDD opcode[0] a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X788 VDD a_307_3697# a_897_3260# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X789 a_22849_n990# a_23723_n1475# a_23198_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X790 a_23670_n2323# a_22290_n990# a_23198_n990# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X791 a_8794_n7362# a_8249_n6669# a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X792 VDD a_21997_n6357# a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X793 a_14288_3692# A[2] a_14406_3692# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X794 a_17798_3694# A[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X795 a_4657_n8096# a_4951_n7390# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X796 a_13419_n3726# a_13359_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X797 VDD opcode[0] a_9658_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=300000u
X798 a_22849_1744# a_11205_3262# a_23198_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X799 VDD opcode[1] a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X800 Y[5] a_16922_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X801 a_2882_n7388# B[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X802 a_7432_1744# opcode[0] a_7668_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X803 a_6514_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X804 a_16513_1714# a_17798_3694# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X805 a_10576_n990# a_11101_n1475# a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X806 a_16563_n3726# a_16503_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X807 a_307_3697# B[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X808 VSS opcode[0] a_3382_n3726# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X809 a_10576_1744# a_5291_3262# a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X810 a_16503_n3752# A[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X811 VDD opcode[0] a_16004_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X812 VDD B[1] a_13238_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X813 a_7432_n990# a_7957_n1475# a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X814 a_8676_n7362# a_8249_n6669# a_8794_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X815 VDD A[0] a_n25_n6671# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X816 VDD B[3] a_15574_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X817 a_10802_n5055# a_10157_n3748# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X818 a_9658_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_7432_1744# a_3843_3262# a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X820 a_16573_1740# a_16513_1714# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X821 a_2345_3260# a_1755_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X822 a_3891_n1020# a_4290_n3726# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X823 VDD a_6221_3697# a_6811_3260# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X824 VDD a_14288_3692# a_7023_1718# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X825 a_20526_411# a_19146_1744# a_20054_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X826 a_16573_n994# a_16513_n1020# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X827 a_22839_n3722# a_22280_n3722# a_23188_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X828 a_1392_407# a_747_1714# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X829 a_20044_n3722# opcode[0] a_20280_n5055# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X830 a_16004_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X831 VDD B[7] a_10615_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X832 VDD B[6] a_12813_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X833 a_8794_n7362# a_8249_n6669# a_8676_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X834 a_3891_1714# a_13120_3694# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X835 VDD a_19645_n1016# a_19705_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X836 VSS B[4] a_9030_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X837 a_10566_n3722# opcode[0] a_10802_n5055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X838 VDD opcode[0] a_9658_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X839 a_7073_n3722# a_6514_n3722# a_7422_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X840 VDD a_19230_3112# a_19705_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X841 a_19705_n990# a_19146_n990# a_20054_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X842 a_10615_3699# B[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X843 VDD A[5] a_10317_n6667# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X844 a_15293_n7386# B[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X845 a_20044_n3722# a_12931_n7362# a_19695_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X846 a_19705_1744# a_19146_1744# a_20054_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X847 a_12931_n7362# a_12386_n6669# a_12931_n8094# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X848 a_23188_n3722# a_22280_n3722# a_22839_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X849 a_13429_1740# a_6811_3260# a_13778_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X850 a_20516_n5055# a_19136_n3722# a_20044_n3722# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X851 a_13419_n3726# a_12860_n3726# a_13768_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X852 VDD a_10615_3699# a_11205_3262# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X853 a_2043_n6669# A[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X854 a_7658_n5055# a_7013_n3748# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X855 a_19645_n1016# a_20044_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X856 VDD opcode[0] a_7073_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X857 a_16748_3696# A[4] a_16630_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X858 VSS opcode[0] a_3392_1740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X859 a_13429_n994# a_14303_n1479# a_13778_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X860 a_10157_n3748# A[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X861 a_16573_1740# a_8259_3260# a_16922_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X862 VDD A[2] a_3253_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X863 a_19084_3696# A[6] a_18966_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X864 a_10317_n6667# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X865 a_16563_n3726# a_16004_n3726# a_16912_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X866 VDD a_7669_3697# a_8259_3260# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X867 VDD opcode[1] a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X868 VDD B[7] a_15293_n7386# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X869 a_3490_3062# A[2] a_3253_3699# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X870 VDD opcode[0] a_3951_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X871 VDD opcode[0] a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X872 a_22839_n3722# a_22280_n3722# a_23188_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X873 a_16922_1740# a_8259_3260# a_16573_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X874 a_16573_n994# a_17447_n1479# a_16922_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X875 VSS a_12931_n7362# a_20516_n5055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X876 VDD opcode[0] a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X877 a_7432_n990# a_6524_n990# a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X878 VDD a_4300_1740# a_4825_n1479# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X879 VDD opcode[1] a_3951_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X880 VDD A[1] a_2043_n6669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X881 a_7432_1744# a_6524_1744# a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X882 a_10227_n990# a_9668_n990# a_10576_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X883 a_4536_n2327# a_3891_n1020# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X884 VDD a_20044_n3722# a_19645_n1016# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X885 a_7073_n3722# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X886 VDD B[2] a_14406_3692# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X887 a_16922_n994# a_17447_n1479# a_16573_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X888 a_10227_1744# a_9668_1744# a_10576_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X889 VSS a_14999_n7360# a_23660_n5055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X890 a_17148_n5059# a_16503_n3752# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X891 a_19230_3112# a_18966_3696# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X892 a_7083_n990# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X893 a_10576_n990# a_11101_n1475# a_10227_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X894 VDD opcode[0] a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X895 VDD a_4300_n994# Y[1] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X896 a_7083_1744# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X897 a_10576_1744# a_5291_3262# a_10227_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X898 VDD B[0] a_12070_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X899 VDD a_16630_3696# a_13369_1714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X900 VDD opcode[1] a_7083_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X901 Y[2] a_7432_n990# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X902 a_3382_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X903 a_6725_n7362# a_6180_n6669# a_6607_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X904 VDD B[3] a_4701_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X905 VDD opcode[0] a_7083_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X906 a_7957_n1475# a_7432_1744# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X907 VDD A[5] a_16503_n3752# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X908 a_4300_n994# opcode[1] a_4536_n2327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X909 a_2345_3260# a_1755_3697# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X910 a_6221_3697# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X911 a_16563_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X912 a_7023_n1016# a_7422_n3722# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X913 a_9167_3699# A[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X914 VSS opcode[0] a_19136_n3722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X915 VSS B[6] a_9404_3062# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X916 a_13429_1740# a_12870_1740# a_13778_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X917 VDD opcode[0] a_3382_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X918 VSS opcode[0] a_9658_n3722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X919 a_7023_1718# a_14288_3692# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X920 a_6607_n7362# a_6180_n6669# a_6725_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X921 a_16503_n3752# A[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X922 a_13419_n3726# a_12860_n3726# a_13768_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X923 VDD opcode[0] a_3392_1740# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X924 a_19705_n990# a_19146_n990# a_20054_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X925 a_16912_n3726# a_10862_n7360# a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X926 a_13429_n994# a_12870_n994# a_13778_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X927 a_747_n1020# a_1146_n3726# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X928 a_19705_1744# a_19146_1744# a_20054_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X929 VDD A[7] a_14454_n6667# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X930 VDD opcode[0] a_16563_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X931 VDD opcode[1] a_19146_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X932 VSS opcode[0] a_9668_1744# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=300000u
X933 VDD opcode[1] a_3392_n994# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X934 VDD opcode[0] a_19146_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X935 a_16513_n1020# a_16912_n3726# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X936 a_14014_407# a_13369_1714# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X937 VDD opcode[0] a_238_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X938 VDD opcode[0] a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X939 a_13768_n3726# a_12860_n3726# a_13419_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X940 a_1681_n1479# a_1156_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X941 VDD B[2] a_3253_3699# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X942 VDD opcode[1] a_22849_n990# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X943 a_14454_n6667# A[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X944 a_16573_1740# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X945 a_4657_n7364# a_4951_n7390# a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X946 a_4539_n7364# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X947 a_16748_3696# A[4] a_16630_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X948 VDD opcode[0] a_22849_1744# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X949 Y[0] a_1156_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X950 a_1146_n3726# a_520_n7364# a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X951 VDD A[3] a_10157_n3748# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X952 a_17447_n1479# a_16922_1740# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X953 VDD a_23198_n990# Y[7] VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X954 a_16630_3696# A[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X955 a_16573_n994# opcode[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X956 VDD B[4] a_16748_3696# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X957 VDD a_23198_1744# a_23723_n1475# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X958 a_797_n3726# opcode[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X959 VDD B[2] a_14406_3692# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X960 VSS B[0] a_756_n8096# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X961 VDD opcode[0] a_19136_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X962 Y[5] a_16922_n994# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X963 VDD B[5] a_10744_n7360# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X964 a_13238_3694# A[1] a_13120_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X965 a_7668_411# a_7023_1718# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X966 a_4951_n7390# B[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X967 a_4539_n7364# a_4951_n7390# a_4657_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X968 VDD A[2] a_4539_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X969 a_15574_3694# A[3] a_15456_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X970 a_402_n7364# a_814_n7390# a_520_n7364# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X971 a_307_3697# A[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X972 a_7023_n1016# a_7422_n3722# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X973 a_19230_3112# a_18966_3696# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X974 VDD opcode[0] a_797_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X975 a_14881_n7360# B[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X976 a_520_n8096# a_814_n7390# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X977 a_6221_3697# A[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X978 VDD B[0] a_12070_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X979 a_20252_3694# A[7] a_20134_3694# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X980 a_3941_n3726# a_3881_n3752# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X981 a_10744_n7360# B[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X982 a_9167_3699# B[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X983 a_747_1714# a_11952_3694# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X984 VDD A[7] a_21997_n6357# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X985 a_4539_n7364# A[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X986 a_10812_n2323# a_10167_n1016# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X987 a_8676_n7362# a_9088_n7388# a_8794_n7362# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X988 a_20054_1744# opcode[0] a_20290_411# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X989 VDD opcode[0] a_3941_n3726# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X990 a_11156_n7386# B[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X991 VDD opcode[0] a_10217_n3722# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

