magic
tech sky130B
magscale 1 2
timestamp 1736446844
<< nwell >>
rect 0 318 1192 576
rect 1448 318 2640 576
rect 2946 320 4138 578
rect 4394 320 5586 578
rect 803 288 1099 318
rect 2251 288 2547 318
rect 3749 290 4045 320
rect 5197 290 5493 320
rect 5914 318 7106 576
rect 7362 318 8554 576
rect 8860 320 10052 578
rect 10308 320 11500 578
rect 6717 288 7013 318
rect 8165 288 8461 318
rect 9663 290 9959 320
rect 11111 290 11407 320
<< psubdiff >>
rect 538 -712 750 -682
rect 538 -768 578 -712
rect 712 -768 750 -712
rect 538 -790 750 -768
rect 1986 -712 2198 -682
rect 1986 -768 2026 -712
rect 2160 -768 2198 -712
rect 1986 -790 2198 -768
rect 3484 -710 3696 -680
rect 3484 -766 3524 -710
rect 3658 -766 3696 -710
rect 3484 -788 3696 -766
rect 4932 -710 5144 -680
rect 4932 -766 4972 -710
rect 5106 -766 5144 -710
rect 4932 -788 5144 -766
rect 6452 -712 6664 -682
rect 6452 -768 6492 -712
rect 6626 -768 6664 -712
rect 6452 -790 6664 -768
rect 7900 -712 8112 -682
rect 7900 -768 7940 -712
rect 8074 -768 8112 -712
rect 7900 -790 8112 -768
rect 9398 -710 9610 -680
rect 9398 -766 9438 -710
rect 9572 -766 9610 -710
rect 9398 -788 9610 -766
rect 10846 -710 11058 -680
rect 10846 -766 10886 -710
rect 11020 -766 11058 -710
rect 10846 -788 11058 -766
<< nsubdiff >>
rect 298 496 542 534
rect 298 426 354 496
rect 490 426 542 496
rect 298 404 542 426
rect 1746 496 1990 534
rect 1746 426 1802 496
rect 1938 426 1990 496
rect 1746 404 1990 426
rect 3244 498 3488 536
rect 3244 428 3300 498
rect 3436 428 3488 498
rect 3244 406 3488 428
rect 4692 498 4936 536
rect 4692 428 4748 498
rect 4884 428 4936 498
rect 4692 406 4936 428
rect 6212 496 6456 534
rect 6212 426 6268 496
rect 6404 426 6456 496
rect 6212 404 6456 426
rect 7660 496 7904 534
rect 7660 426 7716 496
rect 7852 426 7904 496
rect 7660 404 7904 426
rect 9158 498 9402 536
rect 9158 428 9214 498
rect 9350 428 9402 498
rect 9158 406 9402 428
rect 10606 498 10850 536
rect 10606 428 10662 498
rect 10798 428 10850 498
rect 10606 406 10850 428
<< psubdiffcont >>
rect 578 -768 712 -712
rect 2026 -768 2160 -712
rect 3524 -766 3658 -710
rect 4972 -766 5106 -710
rect 6492 -768 6626 -712
rect 7940 -768 8074 -712
rect 9438 -766 9572 -710
rect 10886 -766 11020 -710
<< nsubdiffcont >>
rect 354 426 490 496
rect 1802 426 1938 496
rect 3300 428 3436 498
rect 4748 428 4884 498
rect 6268 426 6404 496
rect 7716 426 7852 496
rect 9214 428 9350 498
rect 10662 428 10798 498
<< poly >>
rect 95 289 391 325
rect 449 288 745 324
rect 803 288 1099 324
rect 1543 289 1839 325
rect 1897 288 2193 324
rect 2251 288 2547 324
rect 3041 291 3337 327
rect 3395 290 3691 326
rect 3749 290 4045 326
rect 4489 291 4785 327
rect 4843 290 5139 326
rect 5197 290 5493 326
rect 6009 289 6305 325
rect 6363 288 6659 324
rect 6717 288 7013 324
rect 7457 289 7753 325
rect 7811 288 8107 324
rect 8165 288 8461 324
rect 8955 291 9251 327
rect 9309 290 9605 326
rect 9663 290 9959 326
rect 10403 291 10699 327
rect 10757 290 11053 326
rect 11111 290 11407 326
rect 332 -168 390 48
rect 450 -168 510 48
rect 803 36 863 58
rect 800 20 866 36
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -30 866 -14
rect 1780 -168 1838 48
rect 1898 -168 1958 48
rect 2251 36 2311 58
rect 2248 20 2314 36
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 2248 -30 2314 -14
rect 3278 -166 3336 50
rect 3396 -166 3456 50
rect 3749 38 3809 60
rect 3746 22 3812 38
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 3746 -28 3812 -12
rect 4726 -166 4784 50
rect 4844 -166 4904 50
rect 5197 38 5257 60
rect 5194 22 5260 38
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 5194 -28 5260 -12
rect 6246 -168 6304 48
rect 6364 -168 6424 48
rect 6717 36 6777 58
rect 6714 20 6780 36
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 6714 -30 6780 -14
rect 7694 -168 7752 48
rect 7812 -168 7872 48
rect 8165 36 8225 58
rect 8162 20 8228 36
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 8162 -30 8228 -14
rect 9192 -166 9250 50
rect 9310 -166 9370 50
rect 9663 38 9723 60
rect 9660 22 9726 38
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 9660 -28 9726 -12
rect 10640 -166 10698 50
rect 10758 -166 10818 50
rect 11111 38 11171 60
rect 11108 22 11174 38
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 11108 -28 11174 -12
<< polycont >>
rect 816 -14 850 20
rect 2264 -14 2298 20
rect 3762 -12 3796 22
rect 5210 -12 5244 22
rect 6730 -14 6764 20
rect 8178 -14 8212 20
rect 9676 -12 9710 22
rect 11124 -12 11158 22
<< locali >>
rect 338 496 506 512
rect 338 426 354 496
rect 490 426 506 496
rect 338 410 506 426
rect 1786 496 1954 512
rect 1786 426 1802 496
rect 1938 426 1954 496
rect 1786 410 1954 426
rect 3284 498 3452 514
rect 3284 428 3300 498
rect 3436 428 3452 498
rect 3284 412 3452 428
rect 4732 498 4900 514
rect 4732 428 4748 498
rect 4884 428 4900 498
rect 4732 412 4900 428
rect 6252 496 6420 512
rect 6252 426 6268 496
rect 6404 426 6420 496
rect 6252 410 6420 426
rect 7700 496 7868 512
rect 7700 426 7716 496
rect 7852 426 7868 496
rect 7700 410 7868 426
rect 9198 498 9366 514
rect 9198 428 9214 498
rect 9350 428 9366 498
rect 9198 412 9366 428
rect 10646 498 10814 514
rect 10646 428 10662 498
rect 10798 428 10814 498
rect 10646 412 10814 428
rect 875 306 1145 340
rect 875 240 909 306
rect 1111 240 1145 306
rect 2323 306 2593 340
rect 2323 240 2357 306
rect 2559 240 2593 306
rect 3821 308 4091 342
rect 3821 242 3855 308
rect 4057 242 4091 308
rect 5269 308 5539 342
rect 5269 242 5303 308
rect 5505 242 5539 308
rect 6789 306 7059 340
rect 6789 240 6823 306
rect 7025 240 7059 306
rect 8237 306 8507 340
rect 8237 240 8271 306
rect 8473 240 8507 306
rect 9735 308 10005 342
rect 9735 242 9769 308
rect 9971 242 10005 308
rect 11183 308 11453 342
rect 11183 242 11217 308
rect 11419 242 11453 308
rect 800 -14 816 20
rect 850 -14 866 20
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 562 -712 730 -694
rect 562 -768 578 -712
rect 712 -768 730 -712
rect 562 -784 730 -768
rect 2010 -712 2178 -694
rect 2010 -768 2026 -712
rect 2160 -768 2178 -712
rect 2010 -784 2178 -768
rect 3508 -710 3676 -692
rect 3508 -766 3524 -710
rect 3658 -766 3676 -710
rect 3508 -782 3676 -766
rect 4956 -710 5124 -692
rect 4956 -766 4972 -710
rect 5106 -766 5124 -710
rect 4956 -782 5124 -766
rect 6476 -712 6644 -694
rect 6476 -768 6492 -712
rect 6626 -768 6644 -712
rect 6476 -784 6644 -768
rect 7924 -712 8092 -694
rect 7924 -768 7940 -712
rect 8074 -768 8092 -712
rect 7924 -784 8092 -768
rect 9422 -710 9590 -692
rect 9422 -766 9438 -710
rect 9572 -766 9590 -710
rect 9422 -782 9590 -766
rect 10870 -710 11038 -692
rect 10870 -766 10886 -710
rect 11020 -766 11038 -710
rect 10870 -782 11038 -766
<< viali >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 816 -14 850 20
rect 2264 -14 2298 20
rect 3762 -12 3796 22
rect 5210 -12 5244 22
rect 6730 -14 6764 20
rect 8178 -14 8212 20
rect 9676 -12 9710 22
rect 11124 -12 11158 22
rect 618 -764 670 -718
rect 2066 -764 2118 -718
rect 3564 -762 3616 -716
rect 5012 -762 5064 -716
rect 6532 -764 6584 -718
rect 7980 -764 8032 -718
rect 9478 -762 9530 -716
rect 10926 -762 10978 -716
<< metal1 >>
rect 354 494 490 514
rect 354 432 390 494
rect 450 432 490 494
rect 354 404 490 432
rect 1802 494 1938 514
rect 1802 432 1838 494
rect 1898 432 1938 494
rect 1802 404 1938 432
rect 3300 496 3436 516
rect 3300 434 3336 496
rect 3396 434 3436 496
rect 3300 406 3436 434
rect 4748 496 4884 516
rect 4748 434 4784 496
rect 4844 434 4884 496
rect 4748 406 4884 434
rect 6268 494 6404 514
rect 6268 432 6304 494
rect 6364 432 6404 494
rect 50 374 1027 404
rect 50 250 82 374
rect 286 250 318 374
rect 522 250 554 374
rect 758 250 790 374
rect 993 241 1027 374
rect 1498 374 2475 404
rect 1498 250 1530 374
rect 1734 250 1766 374
rect 1970 250 2002 374
rect 2206 250 2238 374
rect 2441 241 2475 374
rect 2996 376 3973 406
rect 2996 252 3028 376
rect 3232 252 3264 376
rect 3468 252 3500 376
rect 3704 252 3736 376
rect 3939 243 3973 376
rect 4444 376 5421 406
rect 6268 404 6404 432
rect 7716 494 7852 514
rect 7716 432 7752 494
rect 7812 432 7852 494
rect 7716 404 7852 432
rect 9214 496 9350 516
rect 9214 434 9250 496
rect 9310 434 9350 496
rect 9214 406 9350 434
rect 10662 496 10798 516
rect 10662 434 10698 496
rect 10758 434 10798 496
rect 10662 406 10798 434
rect 4444 252 4476 376
rect 4680 252 4712 376
rect 4916 252 4948 376
rect 5152 252 5184 376
rect 5387 243 5421 376
rect 5964 374 6941 404
rect 5964 250 5996 374
rect 6200 250 6232 374
rect 6436 250 6468 374
rect 6672 250 6704 374
rect 6907 241 6941 374
rect 7412 374 8389 404
rect 7412 250 7444 374
rect 7648 250 7680 374
rect 7884 250 7916 374
rect 8120 250 8152 374
rect 8355 241 8389 374
rect 8910 376 9887 406
rect 8910 252 8942 376
rect 9146 252 9178 376
rect 9382 252 9414 376
rect 9618 252 9650 376
rect 9853 243 9887 376
rect 10358 376 11335 406
rect 10358 252 10390 376
rect 10594 252 10626 376
rect 10830 252 10862 376
rect 11066 252 11098 376
rect 11301 243 11335 376
rect 166 -26 202 84
rect 402 -26 438 84
rect 638 -25 674 86
rect 800 20 866 27
rect 800 -14 816 20
rect 850 -14 866 20
rect 800 -25 866 -14
rect 638 -26 866 -25
rect 166 -55 866 -26
rect 166 -56 748 -55
rect 286 -194 320 -56
rect 682 -138 748 -56
rect 1110 -165 1145 96
rect 1614 -26 1650 84
rect 1850 -26 1886 84
rect 2086 -25 2122 86
rect 2248 20 2314 27
rect 2248 -14 2264 20
rect 2298 -14 2314 20
rect 2248 -25 2314 -14
rect 2086 -26 2314 -25
rect 1614 -55 2314 -26
rect 1614 -56 2196 -55
rect 756 -194 1145 -165
rect 1734 -194 1768 -56
rect 2130 -138 2196 -56
rect 2558 -165 2593 96
rect 3112 -24 3148 86
rect 3348 -24 3384 86
rect 3584 -23 3620 88
rect 3746 22 3812 29
rect 3746 -12 3762 22
rect 3796 -12 3812 22
rect 3746 -23 3812 -12
rect 3584 -24 3812 -23
rect 3112 -53 3812 -24
rect 3112 -54 3694 -53
rect 2204 -194 2593 -165
rect 3232 -192 3266 -54
rect 3628 -136 3694 -54
rect 4056 -163 4091 98
rect 4560 -24 4596 86
rect 4796 -24 4832 86
rect 5032 -23 5068 88
rect 5194 22 5260 29
rect 5194 -12 5210 22
rect 5244 -12 5260 22
rect 5194 -23 5260 -12
rect 5032 -24 5260 -23
rect 4560 -53 5260 -24
rect 4560 -54 5142 -53
rect 3702 -192 4091 -163
rect 4680 -192 4714 -54
rect 5076 -136 5142 -54
rect 5504 -163 5539 98
rect 6080 -26 6116 84
rect 6316 -26 6352 84
rect 6552 -25 6588 86
rect 6714 20 6780 27
rect 6714 -14 6730 20
rect 6764 -14 6780 20
rect 6714 -25 6780 -14
rect 6552 -26 6780 -25
rect 6080 -55 6780 -26
rect 6080 -56 6662 -55
rect 5150 -192 5539 -163
rect 1041 -274 1145 -194
rect 2489 -274 2593 -194
rect 3987 -272 4091 -192
rect 5435 -272 5539 -192
rect 6200 -194 6234 -56
rect 6596 -138 6662 -56
rect 7024 -165 7059 96
rect 7528 -26 7564 84
rect 7764 -26 7800 84
rect 8000 -25 8036 86
rect 8162 20 8228 27
rect 8162 -14 8178 20
rect 8212 -14 8228 20
rect 8162 -25 8228 -14
rect 8000 -26 8228 -25
rect 7528 -55 8228 -26
rect 7528 -56 8110 -55
rect 6670 -194 7059 -165
rect 7648 -194 7682 -56
rect 8044 -138 8110 -56
rect 8472 -165 8507 96
rect 9026 -24 9062 86
rect 9262 -24 9298 86
rect 9498 -23 9534 88
rect 9660 22 9726 29
rect 9660 -12 9676 22
rect 9710 -12 9726 22
rect 9660 -23 9726 -12
rect 9498 -24 9726 -23
rect 9026 -53 9726 -24
rect 9026 -54 9608 -53
rect 8118 -194 8507 -165
rect 9146 -192 9180 -54
rect 9542 -136 9608 -54
rect 9970 -163 10005 98
rect 10474 -24 10510 86
rect 10710 -24 10746 86
rect 10946 -23 10982 88
rect 11108 22 11174 29
rect 11108 -12 11124 22
rect 11158 -12 11174 22
rect 11108 -23 11174 -12
rect 10946 -24 11174 -23
rect 10474 -53 11174 -24
rect 10474 -54 11056 -53
rect 9616 -192 10005 -163
rect 10594 -192 10628 -54
rect 10990 -136 11056 -54
rect 11418 -163 11453 98
rect 11064 -192 11453 -163
rect 6955 -274 7059 -194
rect 8403 -274 8507 -194
rect 9901 -272 10005 -192
rect 11349 -272 11453 -192
rect 140 -409 240 -309
rect 639 -364 674 -317
rect 28 -537 128 -437
rect 50 -686 104 -537
rect 164 -601 218 -409
rect 639 -530 682 -364
rect 1588 -409 1688 -309
rect 2087 -364 2122 -317
rect 560 -533 682 -530
rect 522 -573 682 -533
rect 1476 -537 1576 -437
rect 164 -657 395 -601
rect 447 -686 513 -601
rect 50 -694 513 -686
rect 50 -726 514 -694
rect 606 -710 682 -573
rect 1498 -686 1552 -537
rect 1612 -601 1666 -409
rect 2087 -530 2130 -364
rect 3086 -407 3186 -307
rect 3585 -362 3620 -315
rect 2008 -533 2130 -530
rect 1970 -573 2130 -533
rect 2974 -535 3074 -435
rect 1612 -657 1843 -601
rect 1895 -686 1961 -601
rect 1498 -694 1961 -686
rect 602 -770 612 -710
rect 674 -770 684 -710
rect 1498 -726 1962 -694
rect 2054 -710 2130 -573
rect 2996 -684 3050 -535
rect 3110 -599 3164 -407
rect 3585 -528 3628 -362
rect 4534 -407 4634 -307
rect 5033 -362 5068 -315
rect 3506 -531 3628 -528
rect 3468 -571 3628 -531
rect 4422 -535 4522 -435
rect 3110 -655 3341 -599
rect 3393 -684 3459 -599
rect 2996 -692 3459 -684
rect 2050 -770 2060 -710
rect 2122 -770 2132 -710
rect 2996 -724 3460 -692
rect 3552 -708 3628 -571
rect 4444 -684 4498 -535
rect 4558 -599 4612 -407
rect 5033 -528 5076 -362
rect 6054 -409 6154 -309
rect 6553 -364 6588 -317
rect 4954 -531 5076 -528
rect 4916 -571 5076 -531
rect 5942 -537 6042 -437
rect 4558 -655 4789 -599
rect 4841 -684 4907 -599
rect 4444 -692 4907 -684
rect 3548 -768 3558 -708
rect 3620 -768 3630 -708
rect 4444 -724 4908 -692
rect 5000 -708 5076 -571
rect 5964 -686 6018 -537
rect 6078 -601 6132 -409
rect 6553 -530 6596 -364
rect 7502 -409 7602 -309
rect 8001 -364 8036 -317
rect 6474 -533 6596 -530
rect 6436 -573 6596 -533
rect 7390 -537 7490 -437
rect 6078 -657 6309 -601
rect 6361 -686 6427 -601
rect 5964 -694 6427 -686
rect 4996 -768 5006 -708
rect 5068 -768 5078 -708
rect 5964 -726 6428 -694
rect 6520 -710 6596 -573
rect 7412 -686 7466 -537
rect 7526 -601 7580 -409
rect 8001 -530 8044 -364
rect 9000 -407 9100 -307
rect 9499 -362 9534 -315
rect 7922 -533 8044 -530
rect 7884 -573 8044 -533
rect 8888 -535 8988 -435
rect 7526 -657 7757 -601
rect 7809 -686 7875 -601
rect 7412 -694 7875 -686
rect 6516 -770 6526 -710
rect 6588 -770 6598 -710
rect 7412 -726 7876 -694
rect 7968 -710 8044 -573
rect 8910 -684 8964 -535
rect 9024 -599 9078 -407
rect 9499 -528 9542 -362
rect 10448 -407 10548 -307
rect 10947 -362 10982 -315
rect 9420 -531 9542 -528
rect 9382 -571 9542 -531
rect 10336 -535 10436 -435
rect 9024 -655 9255 -599
rect 9307 -684 9373 -599
rect 8910 -692 9373 -684
rect 7964 -770 7974 -710
rect 8036 -770 8046 -710
rect 8910 -724 9374 -692
rect 9466 -708 9542 -571
rect 10358 -684 10412 -535
rect 10472 -599 10526 -407
rect 10947 -528 10990 -362
rect 10868 -531 10990 -528
rect 10830 -571 10990 -531
rect 10472 -655 10703 -599
rect 10755 -684 10821 -599
rect 10358 -692 10821 -684
rect 9462 -768 9472 -708
rect 9534 -768 9544 -708
rect 10358 -724 10822 -692
rect 10914 -708 10990 -571
rect 10910 -768 10920 -708
rect 10982 -768 10992 -708
<< via1 >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 612 -718 674 -710
rect 612 -764 618 -718
rect 618 -764 670 -718
rect 670 -764 674 -718
rect 612 -770 674 -764
rect 2060 -718 2122 -710
rect 2060 -764 2066 -718
rect 2066 -764 2118 -718
rect 2118 -764 2122 -718
rect 2060 -770 2122 -764
rect 3558 -716 3620 -708
rect 3558 -762 3564 -716
rect 3564 -762 3616 -716
rect 3616 -762 3620 -716
rect 3558 -768 3620 -762
rect 5006 -716 5068 -708
rect 5006 -762 5012 -716
rect 5012 -762 5064 -716
rect 5064 -762 5068 -716
rect 5006 -768 5068 -762
rect 6526 -718 6588 -710
rect 6526 -764 6532 -718
rect 6532 -764 6584 -718
rect 6584 -764 6588 -718
rect 6526 -770 6588 -764
rect 7974 -718 8036 -710
rect 7974 -764 7980 -718
rect 7980 -764 8032 -718
rect 8032 -764 8036 -718
rect 7974 -770 8036 -764
rect 9472 -716 9534 -708
rect 9472 -762 9478 -716
rect 9478 -762 9530 -716
rect 9530 -762 9534 -716
rect 9472 -768 9534 -762
rect 10920 -716 10982 -708
rect 10920 -762 10926 -716
rect 10926 -762 10978 -716
rect 10978 -762 10982 -716
rect 10920 -768 10982 -762
<< metal2 >>
rect 390 494 450 504
rect 390 422 450 432
rect 1838 494 1898 504
rect 1838 422 1898 432
rect 3336 496 3396 506
rect 3336 424 3396 434
rect 4784 496 4844 506
rect 4784 424 4844 434
rect 6304 494 6364 504
rect 6304 422 6364 432
rect 7752 494 7812 504
rect 7752 422 7812 432
rect 9250 496 9310 506
rect 9250 424 9310 434
rect 10698 496 10758 506
rect 10698 424 10758 434
rect 3558 -700 3620 -698
rect 5006 -700 5068 -698
rect 9472 -700 9534 -698
rect 10920 -700 10982 -698
rect 612 -702 674 -700
rect 2060 -702 2122 -700
rect 612 -710 676 -702
rect 674 -712 676 -710
rect 612 -784 676 -774
rect 2060 -710 2124 -702
rect 2122 -712 2124 -710
rect 2060 -784 2124 -774
rect 3558 -708 3622 -700
rect 3620 -710 3622 -708
rect 3558 -782 3622 -772
rect 5006 -708 5070 -700
rect 5068 -710 5070 -708
rect 5006 -782 5070 -772
rect 6526 -702 6588 -700
rect 7974 -702 8036 -700
rect 6526 -710 6590 -702
rect 6588 -712 6590 -710
rect 6526 -784 6590 -774
rect 7974 -710 8038 -702
rect 8036 -712 8038 -710
rect 7974 -784 8038 -774
rect 9472 -708 9536 -700
rect 9534 -710 9536 -708
rect 9472 -782 9536 -772
rect 10920 -708 10984 -700
rect 10982 -710 10984 -708
rect 10920 -782 10984 -772
<< via2 >>
rect 390 432 450 494
rect 1838 432 1898 494
rect 3336 434 3396 496
rect 4784 434 4844 496
rect 6304 432 6364 494
rect 7752 432 7812 494
rect 9250 434 9310 496
rect 10698 434 10758 496
rect 612 -770 674 -712
rect 674 -770 676 -712
rect 612 -774 676 -770
rect 2060 -770 2122 -712
rect 2122 -770 2124 -712
rect 2060 -774 2124 -770
rect 3558 -768 3620 -710
rect 3620 -768 3622 -710
rect 3558 -772 3622 -768
rect 5006 -768 5068 -710
rect 5068 -768 5070 -710
rect 5006 -772 5070 -768
rect 6526 -770 6588 -712
rect 6588 -770 6590 -712
rect 6526 -774 6590 -770
rect 7974 -770 8036 -712
rect 8036 -770 8038 -712
rect 7974 -774 8038 -770
rect 9472 -768 9534 -710
rect 9534 -768 9536 -710
rect 9472 -772 9536 -768
rect 10920 -768 10982 -710
rect 10982 -768 10984 -710
rect 10920 -772 10984 -768
<< metal3 >>
rect 374 498 472 516
rect 374 426 384 498
rect 454 426 472 498
rect 374 418 472 426
rect 1822 498 1920 516
rect 1822 426 1832 498
rect 1902 426 1920 498
rect 1822 418 1920 426
rect 3320 500 3418 518
rect 3320 428 3330 500
rect 3400 428 3418 500
rect 3320 420 3418 428
rect 4768 500 4866 518
rect 4768 428 4778 500
rect 4848 428 4866 500
rect 4768 420 4866 428
rect 6288 498 6386 516
rect 6288 426 6298 498
rect 6368 426 6386 498
rect 6288 418 6386 426
rect 7736 498 7834 516
rect 7736 426 7746 498
rect 7816 426 7834 498
rect 7736 418 7834 426
rect 9234 500 9332 518
rect 9234 428 9244 500
rect 9314 428 9332 500
rect 9234 420 9332 428
rect 10682 500 10780 518
rect 10682 428 10692 500
rect 10762 428 10780 500
rect 10682 420 10780 428
rect 592 -706 694 -690
rect 592 -774 606 -706
rect 680 -774 694 -706
rect 592 -788 694 -774
rect 2040 -706 2142 -690
rect 2040 -774 2054 -706
rect 2128 -774 2142 -706
rect 2040 -788 2142 -774
rect 3538 -704 3640 -688
rect 3538 -772 3552 -704
rect 3626 -772 3640 -704
rect 3538 -786 3640 -772
rect 4986 -704 5088 -688
rect 4986 -772 5000 -704
rect 5074 -772 5088 -704
rect 4986 -786 5088 -772
rect 6506 -706 6608 -690
rect 6506 -774 6520 -706
rect 6594 -774 6608 -706
rect 6506 -788 6608 -774
rect 7954 -706 8056 -690
rect 7954 -774 7968 -706
rect 8042 -774 8056 -706
rect 7954 -788 8056 -774
rect 9452 -704 9554 -688
rect 9452 -772 9466 -704
rect 9540 -772 9554 -704
rect 9452 -786 9554 -772
rect 10900 -704 11002 -688
rect 10900 -772 10914 -704
rect 10988 -772 11002 -704
rect 10900 -786 11002 -772
<< via3 >>
rect 384 494 454 498
rect 384 432 390 494
rect 390 432 450 494
rect 450 432 454 494
rect 384 426 454 432
rect 1832 494 1902 498
rect 1832 432 1838 494
rect 1838 432 1898 494
rect 1898 432 1902 494
rect 1832 426 1902 432
rect 3330 496 3400 500
rect 3330 434 3336 496
rect 3336 434 3396 496
rect 3396 434 3400 496
rect 3330 428 3400 434
rect 4778 496 4848 500
rect 4778 434 4784 496
rect 4784 434 4844 496
rect 4844 434 4848 496
rect 4778 428 4848 434
rect 6298 494 6368 498
rect 6298 432 6304 494
rect 6304 432 6364 494
rect 6364 432 6368 494
rect 6298 426 6368 432
rect 7746 494 7816 498
rect 7746 432 7752 494
rect 7752 432 7812 494
rect 7812 432 7816 494
rect 7746 426 7816 432
rect 9244 496 9314 500
rect 9244 434 9250 496
rect 9250 434 9310 496
rect 9310 434 9314 496
rect 9244 428 9314 434
rect 10692 496 10762 500
rect 10692 434 10698 496
rect 10698 434 10758 496
rect 10758 434 10762 496
rect 10692 428 10762 434
rect 606 -712 680 -706
rect 606 -774 612 -712
rect 612 -774 676 -712
rect 676 -774 680 -712
rect 2054 -712 2128 -706
rect 2054 -774 2060 -712
rect 2060 -774 2124 -712
rect 2124 -774 2128 -712
rect 3552 -710 3626 -704
rect 3552 -772 3558 -710
rect 3558 -772 3622 -710
rect 3622 -772 3626 -710
rect 5000 -710 5074 -704
rect 5000 -772 5006 -710
rect 5006 -772 5070 -710
rect 5070 -772 5074 -710
rect 6520 -712 6594 -706
rect 6520 -774 6526 -712
rect 6526 -774 6590 -712
rect 6590 -774 6594 -712
rect 7968 -712 8042 -706
rect 7968 -774 7974 -712
rect 7974 -774 8038 -712
rect 8038 -774 8042 -712
rect 9466 -710 9540 -704
rect 9466 -772 9472 -710
rect 9472 -772 9536 -710
rect 9536 -772 9540 -710
rect 10914 -710 10988 -704
rect 10914 -772 10920 -710
rect 10920 -772 10984 -710
rect 10984 -772 10988 -710
<< metal4 >>
rect 28 500 11162 556
rect 28 498 3330 500
rect 28 426 384 498
rect 454 426 1832 498
rect 1902 428 3330 498
rect 3400 428 4778 500
rect 4848 498 9244 500
rect 4848 428 6298 498
rect 1902 426 6298 428
rect 6368 426 7746 498
rect 7816 428 9244 498
rect 9314 428 10692 500
rect 10762 428 11162 500
rect 7816 426 11162 428
rect 28 398 11162 426
rect 3424 -678 3756 -676
rect 4872 -678 5204 -676
rect 9338 -678 9670 -676
rect 10786 -678 11118 -676
rect 32 -704 11156 -678
rect 32 -706 3552 -704
rect 32 -774 606 -706
rect 680 -774 2054 -706
rect 2128 -772 3552 -706
rect 3626 -772 5000 -704
rect 5074 -706 9466 -704
rect 5074 -772 6520 -706
rect 2128 -774 6520 -772
rect 6594 -774 7968 -706
rect 8042 -772 9466 -706
rect 9540 -772 10914 -704
rect 10988 -772 11156 -704
rect 8042 -774 11156 -772
rect 32 -812 11156 -774
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_0
timestamp 1735468497
transform 1 0 3426 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_1
timestamp 1735468497
transform 1 0 1928 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_2
timestamp 1735468497
transform 1 0 1810 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_3
timestamp 1735468497
transform 1 0 3308 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_4
timestamp 1735468497
transform 1 0 4756 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_5
timestamp 1735468497
transform 1 0 4874 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_6
timestamp 1735468497
transform 1 0 362 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_7
timestamp 1735468497
transform 1 0 480 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_8
timestamp 1735468497
transform 1 0 10788 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_9
timestamp 1735468497
transform 1 0 10670 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_10
timestamp 1735468497
transform 1 0 9222 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_11
timestamp 1735468497
transform 1 0 9340 0 1 -398
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_12
timestamp 1735468497
transform 1 0 7724 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_13
timestamp 1735468497
transform 1 0 7842 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_14
timestamp 1735468497
transform 1 0 6394 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_M82KHF  sky130_fd_pr__nfet_01v8_M82KHF_15
timestamp 1735468497
transform 1 0 6276 0 1 -400
box -88 -257 88 257
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_0
timestamp 1735468497
transform 1 0 2163 0 1 -238
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_1
timestamp 1735468497
transform 1 0 3661 0 1 -236
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_2
timestamp 1735468497
transform 1 0 5109 0 1 -236
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_3
timestamp 1735468497
transform 1 0 715 0 1 -238
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_4
timestamp 1735468497
transform 1 0 11023 0 1 -236
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_5
timestamp 1735468497
transform 1 0 9575 0 1 -236
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_6
timestamp 1735468497
transform 1 0 8077 0 1 -238
box -88 -157 88 157
use sky130_fd_pr__nfet_01v8_UMD3L6  sky130_fd_pr__nfet_01v8_UMD3L6_7
timestamp 1735468497
transform 1 0 6629 0 1 -238
box -88 -157 88 157
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_0
timestamp 1735468497
transform 1 0 2045 0 1 168
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_1
timestamp 1735468497
transform 1 0 3543 0 1 170
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_2
timestamp 1735468497
transform 1 0 4991 0 1 170
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_3
timestamp 1735468497
transform 1 0 597 0 1 168
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_4
timestamp 1735468497
transform 1 0 10905 0 1 170
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_5
timestamp 1735468497
transform 1 0 9457 0 1 170
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_6
timestamp 1735468497
transform 1 0 7959 0 1 168
box -596 -162 596 162
use sky130_fd_pr__pfet_01v8_A6G7W3  sky130_fd_pr__pfet_01v8_A6G7W3_7
timestamp 1735468497
transform 1 0 6511 0 1 168
box -596 -162 596 162
<< labels >>
flabel metal4 5504 -790 5734 -706 1 FreeSerif 640 0 0 0 VSS
port 1 n
flabel metal4 5566 432 5778 540 1 FreeSerif 640 0 0 0 VDD
port 2 n
flabel metal1 152 -390 228 -320 1 FreeSerif 400 0 0 0 A[0]
port 3 n
flabel metal1 1600 -396 1676 -326 1 FreeSerif 400 0 0 0 A[1]
port 4 n
flabel metal1 3102 -390 3178 -320 1 FreeSerif 400 0 0 0 A[2]
port 5 n
flabel metal1 4548 -392 4624 -322 1 FreeSerif 400 0 0 0 A[3]
port 6 n
flabel metal1 6070 -390 6146 -320 1 FreeSerif 400 0 0 0 A[4]
port 7 n
flabel metal1 7520 -386 7596 -316 1 FreeSerif 400 0 0 0 A[5]
port 8 n
flabel metal1 9014 -392 9090 -322 1 FreeSerif 400 0 0 0 A[6]
port 9 n
flabel metal1 10460 -392 10536 -322 1 FreeSerif 400 0 0 0 A[7]
port 10 n
flabel metal1 10348 -516 10424 -446 1 FreeSerif 400 0 0 0 B[7]
port 11 n
flabel metal1 8900 -516 8976 -446 1 FreeSerif 400 0 0 0 B[6]
port 12 n
flabel metal1 7400 -520 7476 -450 1 FreeSerif 400 0 0 0 B[5]
port 13 n
flabel metal1 4434 -518 4510 -448 1 FreeSerif 400 0 0 0 B[3]
port 14 n
flabel metal1 5952 -518 6028 -448 1 FreeSerif 400 0 0 0 B[4]
port 15 n
flabel metal1 2988 -520 3064 -450 1 FreeSerif 400 0 0 0 B[2]
port 16 n
flabel metal1 1492 -518 1568 -448 1 FreeSerif 400 0 0 0 B[1]
port 17 n
flabel metal1 44 -518 120 -448 1 FreeSerif 400 0 0 0 B[0]
port 18 n
flabel metal1 1058 -258 1134 -188 1 FreeSerif 400 0 0 0 Y[0]
port 19 n
flabel metal1 2500 -254 2576 -184 1 FreeSerif 400 0 0 0 Y[1]
port 20 n
flabel metal1 4004 -252 4080 -182 1 FreeSerif 400 0 0 0 Y[2]
port 21 n
flabel metal1 5454 -254 5530 -184 1 FreeSerif 400 0 0 0 Y[3]
port 22 n
flabel metal1 6970 -252 7046 -182 1 FreeSerif 400 0 0 0 Y[4]
port 23 n
flabel metal1 8422 -254 8498 -184 1 FreeSerif 400 0 0 0 Y[5]
port 24 n
flabel metal1 9912 -262 9988 -192 1 FreeSerif 400 0 0 0 Y[6]
port 25 n
flabel metal1 11362 -256 11438 -186 1 FreeSerif 400 0 0 0 Y[7]
port 26 n
<< end >>
