* NGSPICE file created from logic_or_pex.ext - technology: sky130B

.subckt logic_or A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3]
+ Y[4] Y[5] Y[6] Y[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
X0 a_1780_788.t2 A[1].t0 a_1662_788.t1 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 VDD.t67 B[4].t0 a_5290_790.t3 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2 a_6340_788.t2 A[5].t0 a_6458_788.t2 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3 VDD.t65 a_494_788.t5 Y[0].t2 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4 VSS.t13 B[1].t0 a_1662_788.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 a_6340_788.t3 A[5].t1 VSS.t8 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 a_8794_788.t3 A[7].t0 a_8676_788.t1 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 a_7508_790.t3 A[6].t0 VSS.t12 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 VDD.t91 B[4].t1 a_5290_790.t2 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 Y[6].t3 a_7508_790.t5 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 a_612_788.t4 A[0].t0 a_494_788.t2 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_612_788.t5 B[0].t0 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 a_3998_788.t1 A[3].t0 VSS.t9 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 Y[0].t1 a_494_788.t6 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 VDD.t51 a_2830_786.t5 Y[2].t3 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 Y[4].t0 a_5172_790.t5 VSS.t16 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 a_1662_788.t0 A[1].t1 a_1780_788.t1 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 VDD.t7 B[2].t0 a_2948_786.t5 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_5290_790.t1 B[4].t2 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_1662_788.t3 A[1].t2 VSS.t19 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X20 VDD.t24 B[0].t1 a_612_788.t0 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X21 Y[2].t0 a_2830_786.t6 VSS.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X22 a_494_788.t4 A[0].t1 a_612_788.t3 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 VDD.t79 B[6].t0 a_7626_790.t5 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 VDD.t61 a_5172_790.t6 Y[4].t3 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 VDD.t13 a_7508_790.t6 Y[6].t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 a_5290_790.t5 A[4].t0 a_5172_790.t4 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X27 VDD.t76 a_1662_788.t5 Y[1].t3 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 VDD.t83 B[7].t0 a_8794_788.t4 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X29 Y[7].t0 a_8676_788.t5 VSS.t17 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 a_1780_788.t0 A[1].t3 a_1662_788.t2 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X31 Y[0].t3 a_494_788.t7 VSS.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 a_2948_786.t4 B[2].t1 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X33 a_7508_790.t1 A[6].t1 a_7626_790.t2 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X34 VSS.t11 B[4].t3 a_5172_790.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X35 VDD.t115 B[7].t1 a_8794_788.t5 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X36 VDD.t28 a_6340_788.t5 Y[5].t3 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X37 a_612_788.t2 A[0].t2 a_494_788.t1 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 VDD.t117 B[5].t0 a_6458_788.t5 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_7626_790.t1 A[6].t2 a_7508_790.t4 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X40 Y[4].t2 a_5172_790.t7 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 a_1780_788.t3 B[1].t1 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X42 VSS.t10 B[0].t2 a_494_788.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 VDD.t104 B[3].t0 a_4116_788.t2 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X44 a_5172_790.t3 A[4].t1 a_5290_790.t4 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X45 Y[1].t2 a_1662_788.t6 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 a_8794_788.t0 B[7].t2 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X47 a_7626_790.t0 A[6].t3 a_7508_790.t2 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 a_5172_790.t0 A[4].t2 VSS.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X49 VSS.t22 B[7].t3 a_8676_788.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 VDD.t41 B[2].t2 a_2948_786.t3 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X51 VDD.t119 B[1].t2 a_1780_788.t5 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 a_6458_788.t1 B[5].t1 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 a_2830_786.t4 A[2].t0 VSS.t23 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X54 a_5290_790.t0 A[4].t3 a_5172_790.t1 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 VDD.t101 B[1].t3 a_1780_788.t4 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X56 a_494_788.t0 A[0].t3 VSS.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 VDD.t72 a_1662_788.t7 Y[1].t1 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X58 VDD.t49 a_3998_788.t5 Y[3].t3 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X59 VDD.t108 a_5172_790.t8 Y[4].t1 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X60 a_4116_788.t1 B[3].t1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X61 VSS.t18 B[2].t3 a_2830_786.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 a_8676_788.t2 A[7].t1 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_2948_786.t2 A[2].t1 a_2830_786.t2 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X64 a_4116_788.t5 A[3].t1 a_3998_788.t4 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X65 VDD.t39 a_3998_788.t6 Y[3].t2 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 VDD.t88 a_8676_788.t6 Y[7].t3 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 VDD.t5 B[5].t2 a_6458_788.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X68 VDD.t10 B[6].t1 a_7626_790.t4 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X69 VSS.t0 B[3].t2 a_3998_788.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X70 VDD.t94 B[3].t3 a_4116_788.t0 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X71 Y[3].t1 a_3998_788.t7 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X72 Y[5].t0 a_6340_788.t6 VSS.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 a_8794_788.t2 A[7].t2 a_8676_788.t0 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 Y[3].t0 a_3998_788.t8 VSS.t21 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 Y[5].t2 a_6340_788.t7 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 Y[7].t2 a_8676_788.t7 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 a_3998_788.t2 A[3].t2 a_4116_788.t4 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X78 a_2830_786.t1 A[2].t2 a_2948_786.t1 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X79 a_6458_788.t4 A[5].t2 a_6340_788.t1 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X80 a_7626_790.t3 B[6].t2 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X81 VDD.t63 a_2830_786.t7 Y[2].t2 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X82 Y[1].t0 a_1662_788.t8 VSS.t14 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X83 VSS.t15 B[5].t3 a_6340_788.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 a_8676_788.t3 A[7].t3 a_8794_788.t1 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X85 VSS.t4 B[6].t3 a_7508_790.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X86 VDD.t15 a_7508_790.t7 Y[6].t1 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X87 a_6458_788.t3 A[5].t3 a_6340_788.t0 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 VDD.t26 a_6340_788.t8 Y[5].t1 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 VDD.t47 B[0].t3 a_612_788.t1 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 Y[6].t0 a_7508_790.t8 VSS.t20 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X91 VDD.t56 a_8676_788.t8 Y[7].t1 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X92 a_2948_786.t0 A[2].t3 a_2830_786.t0 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 a_4116_788.t3 A[3].t3 a_3998_788.t3 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X94 VDD.t86 a_494_788.t8 Y[0].t0 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X95 Y[2].t1 a_2830_786.t8 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 A[1].t3 A[1].t2 575.234
R1 A[1].n0 A[1].t0 284.688
R2 A[1].n0 A[1].t1 160.666
R3 A[1].n1 A[1].t3 160.666
R4 A[1] A[1].n1 159.954
R5 A[1].n1 A[1].n0 115.593
R6 a_1662_788.t8 a_1662_788.n2 404.877
R7 a_1662_788.n1 a_1662_788.t5 210.902
R8 a_1662_788.n3 a_1662_788.t8 136.943
R9 a_1662_788.n2 a_1662_788.n1 107.801
R10 a_1662_788.n1 a_1662_788.t6 80.333
R11 a_1662_788.n2 a_1662_788.t7 80.333
R12 a_1662_788.n0 a_1662_788.t4 17.4
R13 a_1662_788.n0 a_1662_788.t3 17.4
R14 a_1662_788.n4 a_1662_788.t2 15.036
R15 a_1662_788.n5 a_1662_788.t1 14.282
R16 a_1662_788.t0 a_1662_788.n5 14.282
R17 a_1662_788.n5 a_1662_788.n4 1.654
R18 a_1662_788.n3 a_1662_788.n0 0.672
R19 a_1662_788.n4 a_1662_788.n3 0.665
R20 a_1780_788.n1 a_1780_788.t4 14.282
R21 a_1780_788.n1 a_1780_788.t2 14.282
R22 a_1780_788.n0 a_1780_788.t1 14.282
R23 a_1780_788.n0 a_1780_788.t0 14.282
R24 a_1780_788.n3 a_1780_788.t5 14.282
R25 a_1780_788.t3 a_1780_788.n3 14.282
R26 a_1780_788.n2 a_1780_788.n0 2.538
R27 a_1780_788.n3 a_1780_788.n2 2.375
R28 a_1780_788.n2 a_1780_788.n1 0.001
R29 VDD.n33 VDD.n32 604.435
R30 VDD.n91 VDD.n90 604.408
R31 VDD.n19 VDD.n18 600.509
R32 VDD.n47 VDD.n46 600.503
R33 VDD.n77 VDD.n76 600.482
R34 VDD.n5 VDD.n4 563.326
R35 VDD.t73 VDD.t75 406.159
R36 VDD.t69 VDD.t62 406.159
R37 VDD.n90 VDD.t71 404.97
R38 VDD.n76 VDD.t50 404.97
R39 VDD.t53 VDD.t107 397.517
R40 VDD.t57 VDD.t87 397.517
R41 VDD.n46 VDD.t55 396.391
R42 VDD.t44 VDD.t14 396.113
R43 VDD.t109 VDD.t27 396.113
R44 VDD.n32 VDD.t12 394.999
R45 VDD.n18 VDD.t25 394.999
R46 VDD.n3 VDD.t60 394.148
R47 VDD.n87 VDD.n86 222.796
R48 VDD.n73 VDD.n72 222.796
R49 VDD.n61 VDD.n60 222.796
R50 VDD.n105 VDD.n104 222.796
R51 VDD.t105 VDD.t48 191.952
R52 VDD.t105 VDD.t38 191.952
R53 VDD.t21 VDD.t64 190
R54 VDD.t21 VDD.t85 190
R55 VDD.t100 VDD.t97 144.087
R56 VDD.t97 VDD.t96 144.087
R57 VDD.t96 VDD.t95 144.087
R58 VDD.t93 VDD.t32 144.087
R59 VDD.t32 VDD.t52 144.087
R60 VDD.t52 VDD.t20 144.087
R61 VDD.t90 VDD.t92 144.087
R62 VDD.t92 VDD.t77 144.087
R63 VDD.t77 VDD.t35 144.087
R64 VDD.t78 VDD.t59 144.087
R65 VDD.t59 VDD.t89 144.087
R66 VDD.t89 VDD.t111 144.087
R67 VDD.t23 VDD.t37 144.087
R68 VDD.t37 VDD.t102 144.087
R69 VDD.t102 VDD.t31 144.087
R70 VDD.t40 VDD.t36 143.717
R71 VDD.t36 VDD.t11 143.717
R72 VDD.t11 VDD.t8 143.717
R73 VDD.t114 VDD.t30 143.717
R74 VDD.t30 VDD.t19 143.717
R75 VDD.t19 VDD.t18 143.717
R76 VDD.t4 VDD.t68 143.717
R77 VDD.t68 VDD.t84 143.717
R78 VDD.t84 VDD.t29 143.717
R79 VDD.n87 VDD.t100 137.982
R80 VDD.n61 VDD.t93 137.982
R81 VDD.n0 VDD.t90 137.982
R82 VDD.n29 VDD.t78 137.982
R83 VDD.n104 VDD.t23 137.982
R84 VDD.n73 VDD.t40 137.628
R85 VDD.n43 VDD.t114 137.628
R86 VDD.n15 VDD.t4 137.628
R87 VDD.n88 VDD.t98 61.054
R88 VDD.n62 VDD.t2 61.054
R89 VDD.n1 VDD.t42 61.054
R90 VDD.n30 VDD.t0 61.054
R91 VDD.t112 VDD.n103 61.054
R92 VDD.n74 VDD.t80 60.898
R93 VDD.n44 VDD.t16 60.898
R94 VDD.n16 VDD.t33 60.898
R95 VDD.n4 VDD.n3 41.219
R96 VDD.n92 VDD.n91 37.853
R97 VDD.n64 VDD.t105 37.853
R98 VDD.t21 VDD.n101 37.853
R99 VDD.n78 VDD.n77 37.756
R100 VDD.n91 VDD.n89 29.305
R101 VDD.t105 VDD.n63 29.305
R102 VDD.n6 VDD.n5 29.305
R103 VDD.n34 VDD.n33 29.305
R104 VDD.n102 VDD.t21 29.305
R105 VDD.n77 VDD.n75 29.23
R106 VDD.n48 VDD.n47 29.23
R107 VDD.n20 VDD.n19 29.23
R108 VDD.n95 VDD.t76 28.57
R109 VDD.n81 VDD.t63 28.57
R110 VDD.n67 VDD.t49 28.57
R111 VDD.n10 VDD.t61 28.57
R112 VDD.n38 VDD.t15 28.57
R113 VDD.n52 VDD.t88 28.57
R114 VDD.n24 VDD.t28 28.57
R115 VDD.n107 VDD.t65 28.57
R116 VDD.n94 VDD.t74 28.565
R117 VDD.n94 VDD.t72 28.565
R118 VDD.n80 VDD.t70 28.565
R119 VDD.n80 VDD.t51 28.565
R120 VDD.n66 VDD.t106 28.565
R121 VDD.n66 VDD.t39 28.565
R122 VDD.n9 VDD.t54 28.565
R123 VDD.n9 VDD.t108 28.565
R124 VDD.n37 VDD.t45 28.565
R125 VDD.n37 VDD.t13 28.565
R126 VDD.n51 VDD.t58 28.565
R127 VDD.n51 VDD.t56 28.565
R128 VDD.n23 VDD.t110 28.565
R129 VDD.n23 VDD.t26 28.565
R130 VDD.n106 VDD.t22 28.565
R131 VDD.n106 VDD.t86 28.565
R132 VDD.n96 VDD.t119 14.284
R133 VDD.n82 VDD.t7 14.284
R134 VDD.n68 VDD.t104 14.284
R135 VDD.n11 VDD.t67 14.284
R136 VDD.n39 VDD.t10 14.284
R137 VDD.n53 VDD.t83 14.284
R138 VDD.n25 VDD.t117 14.284
R139 VDD.n108 VDD.t47 14.284
R140 VDD.n97 VDD.t99 14.282
R141 VDD.n97 VDD.t101 14.282
R142 VDD.n83 VDD.t81 14.282
R143 VDD.n83 VDD.t41 14.282
R144 VDD.n69 VDD.t3 14.282
R145 VDD.n69 VDD.t94 14.282
R146 VDD.n12 VDD.t43 14.282
R147 VDD.n12 VDD.t91 14.282
R148 VDD.n40 VDD.t1 14.282
R149 VDD.n40 VDD.t79 14.282
R150 VDD.n54 VDD.t17 14.282
R151 VDD.n54 VDD.t115 14.282
R152 VDD.n26 VDD.t34 14.282
R153 VDD.n26 VDD.t5 14.282
R154 VDD.n109 VDD.t113 14.282
R155 VDD.n109 VDD.t24 14.282
R156 VDD.n92 VDD.t118 13.431
R157 VDD.n64 VDD.t103 13.431
R158 VDD.n7 VDD.t66 13.431
R159 VDD.n35 VDD.t9 13.431
R160 VDD.n101 VDD.t46 13.431
R161 VDD.n78 VDD.t6 13.397
R162 VDD.n49 VDD.t82 13.397
R163 VDD.n21 VDD.t116 13.397
R164 VDD.t98 VDD.n87 6.105
R165 VDD.t2 VDD.n61 6.105
R166 VDD.t42 VDD.n0 6.105
R167 VDD.t0 VDD.n29 6.105
R168 VDD.n104 VDD.t112 6.105
R169 VDD.t80 VDD.n73 6.089
R170 VDD.t16 VDD.n43 6.089
R171 VDD.t33 VDD.n15 6.089
R172 VDD.n93 VDD.n92 5.506
R173 VDD.n79 VDD.n78 5.506
R174 VDD.n65 VDD.n64 5.506
R175 VDD.n8 VDD.n7 5.506
R176 VDD.n36 VDD.n35 5.506
R177 VDD.n50 VDD.n49 5.506
R178 VDD.n22 VDD.n21 5.506
R179 VDD.n101 VDD.n100 5.506
R180 VDD.n3 VDD.t53 3.368
R181 VDD.n39 VDD.n38 2.225
R182 VDD.n11 VDD.n10 2.221
R183 VDD.n108 VDD.n107 2.221
R184 VDD.n25 VDD.n24 2.218
R185 VDD.n53 VDD.n52 2.214
R186 VDD.n96 VDD.n95 2.199
R187 VDD.n68 VDD.n67 2.199
R188 VDD.n82 VDD.n81 2.192
R189 VDD.n95 VDD.n94 1.651
R190 VDD.n81 VDD.n80 1.651
R191 VDD.n67 VDD.n66 1.651
R192 VDD.n10 VDD.n9 1.607
R193 VDD.n52 VDD.n51 1.607
R194 VDD.n107 VDD.n106 1.607
R195 VDD.n38 VDD.n37 1.599
R196 VDD.n24 VDD.n23 1.599
R197 VDD.n84 VDD.n82 1.161
R198 VDD.n55 VDD.n53 1.161
R199 VDD.n27 VDD.n25 1.161
R200 VDD.n98 VDD.n96 1.154
R201 VDD.n70 VDD.n68 1.154
R202 VDD.n13 VDD.n11 1.154
R203 VDD.n41 VDD.n39 1.154
R204 VDD.n110 VDD.n108 1.154
R205 VDD.n84 VDD.n83 1.107
R206 VDD.n55 VDD.n54 1.107
R207 VDD.n27 VDD.n26 1.107
R208 VDD.n98 VDD.n97 1.1
R209 VDD.n70 VDD.n69 1.1
R210 VDD.n13 VDD.n12 1.1
R211 VDD.n41 VDD.n40 1.1
R212 VDD.n110 VDD.n109 1.1
R213 VDD.n89 VDD.n88 1.008
R214 VDD.n63 VDD.n62 1.008
R215 VDD.n103 VDD.n102 1.008
R216 VDD.n75 VDD.n74 1.006
R217 VDD.n112 VDD.n111 0.284
R218 VDD.n57 VDD.n56 0.283
R219 VDD.n58 VDD.n57 0.28
R220 VDD.n59 VDD.n58 0.28
R221 VDD.n114 VDD.n113 0.28
R222 VDD.n113 VDD.n112 0.28
R223 VDD.n99 VDD.n98 0.241
R224 VDD.n85 VDD.n84 0.241
R225 VDD.n71 VDD.n70 0.241
R226 VDD.n14 VDD.n13 0.241
R227 VDD.n42 VDD.n41 0.241
R228 VDD.n56 VDD.n55 0.241
R229 VDD.n28 VDD.n27 0.241
R230 VDD.n111 VDD.n110 0.241
R231 VDD VDD.n59 0.223
R232 VDD.n99 VDD.n93 0.182
R233 VDD.n85 VDD.n79 0.182
R234 VDD.n71 VDD.n65 0.182
R235 VDD.n14 VDD.n8 0.182
R236 VDD.n42 VDD.n36 0.182
R237 VDD.n56 VDD.n50 0.182
R238 VDD.n28 VDD.n22 0.182
R239 VDD.n111 VDD.n100 0.182
R240 VDD.n90 VDD.t73 0.124
R241 VDD.n76 VDD.t69 0.124
R242 VDD.n46 VDD.t57 0.106
R243 VDD.n32 VDD.t44 0.101
R244 VDD.n18 VDD.t109 0.101
R245 VDD.n93 VDD.n89 0.065
R246 VDD.n79 VDD.n75 0.065
R247 VDD.n65 VDD.n63 0.065
R248 VDD.n8 VDD.n6 0.065
R249 VDD.n36 VDD.n34 0.065
R250 VDD.n50 VDD.n48 0.065
R251 VDD.n22 VDD.n20 0.065
R252 VDD.n102 VDD.n100 0.065
R253 VDD VDD.n114 0.042
R254 VDD.n114 VDD.n71 0.006
R255 VDD.n112 VDD.n99 0.003
R256 VDD.n113 VDD.n85 0.003
R257 VDD.n59 VDD.n14 0.003
R258 VDD.n57 VDD.n42 0.003
R259 VDD.n58 VDD.n28 0.002
R260 VDD.n88 VDD.n86 0.001
R261 VDD.n74 VDD.n72 0.001
R262 VDD.n62 VDD.n60 0.001
R263 VDD.n2 VDD.n1 0.001
R264 VDD.n31 VDD.n30 0.001
R265 VDD.n45 VDD.n44 0.001
R266 VDD.n17 VDD.n16 0.001
R267 VDD.n105 VDD.n103 0.001
R268 VDD.n99 VDD.n86 0.001
R269 VDD.n85 VDD.n72 0.001
R270 VDD.n71 VDD.n60 0.001
R271 VDD.n14 VDD.n2 0.001
R272 VDD.n42 VDD.n31 0.001
R273 VDD.n56 VDD.n45 0.001
R274 VDD.n28 VDD.n17 0.001
R275 VDD.n111 VDD.n105 0.001
R276 B[4].t1 B[4].t3 802.481
R277 B[4] B[4].n1 627.607
R278 B[4].n0 B[4].t0 284.688
R279 B[4].n1 B[4].t1 192.799
R280 B[4].n0 B[4].t2 160.666
R281 B[4].n1 B[4].n0 91.889
R282 a_5290_790.n0 a_5290_790.t2 14.282
R283 a_5290_790.n0 a_5290_790.t5 14.282
R284 a_5290_790.n1 a_5290_790.t3 14.282
R285 a_5290_790.n1 a_5290_790.t1 14.282
R286 a_5290_790.n3 a_5290_790.t4 14.282
R287 a_5290_790.t0 a_5290_790.n3 14.282
R288 a_5290_790.n3 a_5290_790.n2 2.538
R289 a_5290_790.n2 a_5290_790.n1 2.375
R290 a_5290_790.n2 a_5290_790.n0 0.001
R291 A[5].t3 A[5].t1 575.234
R292 A[5].n0 A[5].t2 285.543
R293 A[5].n0 A[5].t0 160.666
R294 A[5].n1 A[5].t3 160.666
R295 A[5] A[5].n1 159.202
R296 A[5].n1 A[5].n0 114.089
R297 a_6458_788.n0 a_6458_788.t2 14.282
R298 a_6458_788.n0 a_6458_788.t3 14.282
R299 a_6458_788.n1 a_6458_788.t5 14.282
R300 a_6458_788.n1 a_6458_788.t1 14.282
R301 a_6458_788.t0 a_6458_788.n3 14.282
R302 a_6458_788.n3 a_6458_788.t4 14.282
R303 a_6458_788.n2 a_6458_788.n0 2.554
R304 a_6458_788.n2 a_6458_788.n1 2.361
R305 a_6458_788.n3 a_6458_788.n2 0.001
R306 a_6340_788.t6 a_6340_788.n2 405.372
R307 a_6340_788.n1 a_6340_788.t5 207.38
R308 a_6340_788.n3 a_6340_788.t6 138.55
R309 a_6340_788.n2 a_6340_788.n1 112.003
R310 a_6340_788.n1 a_6340_788.t7 80.333
R311 a_6340_788.n2 a_6340_788.t8 80.333
R312 a_6340_788.n0 a_6340_788.t4 17.4
R313 a_6340_788.n0 a_6340_788.t3 17.4
R314 a_6340_788.n4 a_6340_788.t0 15.029
R315 a_6340_788.n5 a_6340_788.t1 14.282
R316 a_6340_788.t2 a_6340_788.n5 14.282
R317 a_6340_788.n5 a_6340_788.n4 1.647
R318 a_6340_788.n3 a_6340_788.n0 0.679
R319 a_6340_788.n4 a_6340_788.n3 0.665
R320 a_494_788.t7 a_494_788.n3 406.221
R321 a_494_788.n2 a_494_788.t5 190.962
R322 a_494_788.n4 a_494_788.t7 138.55
R323 a_494_788.n3 a_494_788.n2 111.349
R324 a_494_788.n2 a_494_788.t6 80.333
R325 a_494_788.n3 a_494_788.t8 80.333
R326 a_494_788.n1 a_494_788.t3 17.4
R327 a_494_788.n1 a_494_788.t0 17.4
R328 a_494_788.t1 a_494_788.n5 15.036
R329 a_494_788.n0 a_494_788.t2 14.282
R330 a_494_788.n0 a_494_788.t4 14.282
R331 a_494_788.n5 a_494_788.n0 1.654
R332 a_494_788.n4 a_494_788.n1 0.679
R333 a_494_788.n5 a_494_788.n4 0.665
R334 Y[0].n0 Y[0].t0 28.57
R335 Y[0].n1 Y[0].t2 28.565
R336 Y[0].n1 Y[0].t1 28.565
R337 Y[0].n0 Y[0].t3 17.639
R338 Y[0].n2 Y[0].n1 0.712
R339 Y[0].n2 Y[0].n0 0.605
R340 Y[0] Y[0].n2 0.188
R341 Y[0] Y[0].n3 0.057
R342 Y[0].n3 Y[0] 0.052
R343 Y[0].n3 Y[0] 0.022
R344 B[1].t3 B[1].t0 800.875
R345 B[1] B[1].n1 627.607
R346 B[1].n0 B[1].t2 284.688
R347 B[1].n1 B[1].t3 192.799
R348 B[1].n0 B[1].t1 160.666
R349 B[1].n1 B[1].n0 91.889
R350 VSS.n20 VSS.t19 18.459
R351 VSS.n23 VSS.t23 18.459
R352 VSS.n26 VSS.t9 18.459
R353 VSS.n5 VSS.t12 18.459
R354 VSS.n7 VSS.t3 18.459
R355 VSS.n1 VSS.t2 18.452
R356 VSS.n3 VSS.t8 18.452
R357 VSS.n14 VSS.t1 18.452
R358 VSS.n19 VSS.t14 17.4
R359 VSS.n19 VSS.t13 17.4
R360 VSS.n22 VSS.t7 17.4
R361 VSS.n22 VSS.t18 17.4
R362 VSS.n25 VSS.t21 17.4
R363 VSS.n25 VSS.t0 17.4
R364 VSS.n0 VSS.t16 17.4
R365 VSS.n0 VSS.t11 17.4
R366 VSS.n2 VSS.t5 17.4
R367 VSS.n2 VSS.t15 17.4
R368 VSS.n4 VSS.t20 17.4
R369 VSS.n4 VSS.t4 17.4
R370 VSS.n6 VSS.t17 17.4
R371 VSS.n6 VSS.t22 17.4
R372 VSS.n13 VSS.t6 17.4
R373 VSS.n13 VSS.t10 17.4
R374 VSS.n12 VSS.n11 3.425
R375 VSS.n18 VSS.n17 3.41
R376 VSS.n15 VSS.n12 0.854
R377 VSS.n20 VSS.n19 0.533
R378 VSS.n23 VSS.n22 0.533
R379 VSS.n26 VSS.n25 0.533
R380 VSS.n5 VSS.n4 0.533
R381 VSS.n7 VSS.n6 0.533
R382 VSS.n1 VSS.n0 0.526
R383 VSS.n3 VSS.n2 0.526
R384 VSS.n14 VSS.n13 0.526
R385 VSS.n8 VSS.n7 0.449
R386 VSS.n9 VSS.n8 0.278
R387 VSS.n10 VSS.n9 0.278
R388 VSS.n27 VSS.n24 0.278
R389 VSS.n24 VSS.n21 0.278
R390 VSS.n21 VSS.n18 0.267
R391 VSS.n21 VSS.n20 0.172
R392 VSS.n24 VSS.n23 0.172
R393 VSS.n27 VSS.n26 0.172
R394 VSS.n10 VSS.n1 0.172
R395 VSS.n9 VSS.n3 0.172
R396 VSS.n8 VSS.n5 0.172
R397 VSS.n15 VSS.n14 0.17
R398 VSS VSS.n27 0.148
R399 VSS VSS.n10 0.097
R400 VSS.n18 VSS.n11 0.011
R401 VSS.n17 VSS.n12 0.003
R402 VSS.n16 VSS.n15 0.003
R403 VSS.n16 VSS.n11 0.001
R404 VSS.n17 VSS.n16 0.001
R405 A[7].t0 A[7].t1 573.627
R406 A[7].n0 A[7].t2 285.543
R407 A[7].n0 A[7].t3 160.666
R408 A[7].n1 A[7].t0 160.666
R409 A[7] A[7].n1 159.202
R410 A[7].n1 A[7].n0 114.089
R411 a_8676_788.t5 a_8676_788.n2 406.651
R412 a_8676_788.n1 a_8676_788.t6 207.856
R413 a_8676_788.n3 a_8676_788.t5 136.943
R414 a_8676_788.n2 a_8676_788.n1 111.349
R415 a_8676_788.n1 a_8676_788.t7 80.333
R416 a_8676_788.n2 a_8676_788.t8 80.333
R417 a_8676_788.n0 a_8676_788.t4 17.4
R418 a_8676_788.n0 a_8676_788.t2 17.4
R419 a_8676_788.n4 a_8676_788.t1 15.029
R420 a_8676_788.t0 a_8676_788.n5 14.282
R421 a_8676_788.n5 a_8676_788.t3 14.282
R422 a_8676_788.n5 a_8676_788.n4 1.647
R423 a_8676_788.n3 a_8676_788.n0 0.672
R424 a_8676_788.n4 a_8676_788.n3 0.665
R425 a_8794_788.n1 a_8794_788.t5 14.282
R426 a_8794_788.n1 a_8794_788.t2 14.282
R427 a_8794_788.n0 a_8794_788.t1 14.282
R428 a_8794_788.n0 a_8794_788.t3 14.282
R429 a_8794_788.n3 a_8794_788.t4 14.282
R430 a_8794_788.t0 a_8794_788.n3 14.282
R431 a_8794_788.n2 a_8794_788.n0 2.554
R432 a_8794_788.n3 a_8794_788.n2 2.361
R433 a_8794_788.n2 a_8794_788.n1 0.001
R434 A[6].t3 A[6].t0 575.234
R435 A[6].n0 A[6].t2 284.688
R436 A[6].n0 A[6].t1 160.666
R437 A[6].n1 A[6].t3 160.666
R438 A[6] A[6].n1 159.954
R439 A[6].n1 A[6].n0 115.593
R440 a_7508_790.t8 a_7508_790.n2 406.978
R441 a_7508_790.n1 a_7508_790.t7 207.38
R442 a_7508_790.n3 a_7508_790.t8 136.943
R443 a_7508_790.n2 a_7508_790.n1 112.003
R444 a_7508_790.n1 a_7508_790.t5 80.333
R445 a_7508_790.n2 a_7508_790.t6 80.333
R446 a_7508_790.n0 a_7508_790.t0 17.4
R447 a_7508_790.n0 a_7508_790.t3 17.4
R448 a_7508_790.n4 a_7508_790.t2 15.036
R449 a_7508_790.n5 a_7508_790.t4 14.282
R450 a_7508_790.t1 a_7508_790.n5 14.282
R451 a_7508_790.n5 a_7508_790.n4 1.654
R452 a_7508_790.n3 a_7508_790.n0 0.672
R453 a_7508_790.n4 a_7508_790.n3 0.665
R454 Y[6].n0 Y[6].t2 28.57
R455 Y[6].n1 Y[6].t1 28.565
R456 Y[6].n1 Y[6].t3 28.565
R457 Y[6].n0 Y[6].t0 17.638
R458 Y[6].n2 Y[6].n1 0.716
R459 Y[6].n2 Y[6].n0 0.607
R460 Y[6] Y[6].n2 0.188
R461 Y[6] Y[6].n3 0.057
R462 Y[6].n3 Y[6] 0.052
R463 Y[6].n3 Y[6] 0.022
R464 A[0].t2 A[0].t3 576.841
R465 A[0].n0 A[0].t0 284.688
R466 A[0].n0 A[0].t1 160.666
R467 A[0].n1 A[0].t2 160.666
R468 A[0] A[0].n1 159.954
R469 A[0].n1 A[0].n0 115.593
R470 a_612_788.n0 a_612_788.t3 14.282
R471 a_612_788.n0 a_612_788.t2 14.282
R472 a_612_788.n1 a_612_788.t1 14.282
R473 a_612_788.n1 a_612_788.t5 14.282
R474 a_612_788.t0 a_612_788.n3 14.282
R475 a_612_788.n3 a_612_788.t4 14.282
R476 a_612_788.n2 a_612_788.n0 2.538
R477 a_612_788.n2 a_612_788.n1 2.375
R478 a_612_788.n3 a_612_788.n2 0.001
R479 B[0].t1 B[0].t2 802.481
R480 B[0] B[0].n1 627.607
R481 B[0].n0 B[0].t3 284.688
R482 B[0].n1 B[0].t1 192.799
R483 B[0].n0 B[0].t0 160.666
R484 B[0].n1 B[0].n0 91.889
R485 A[3].t3 A[3].t0 575.234
R486 A[3].n0 A[3].t1 284.688
R487 A[3].n0 A[3].t2 160.666
R488 A[3].n1 A[3].t3 160.666
R489 A[3] A[3].n1 159.954
R490 A[3].n1 A[3].n0 115.593
R491 a_3998_788.t8 a_3998_788.n2 406.053
R492 a_3998_788.n1 a_3998_788.t5 187.473
R493 a_3998_788.n3 a_3998_788.t8 136.943
R494 a_3998_788.n2 a_3998_788.n1 107.801
R495 a_3998_788.n1 a_3998_788.t7 80.333
R496 a_3998_788.n2 a_3998_788.t6 80.333
R497 a_3998_788.n0 a_3998_788.t0 17.4
R498 a_3998_788.n0 a_3998_788.t1 17.4
R499 a_3998_788.n4 a_3998_788.t3 15.036
R500 a_3998_788.n5 a_3998_788.t4 14.282
R501 a_3998_788.t2 a_3998_788.n5 14.282
R502 a_3998_788.n5 a_3998_788.n4 1.654
R503 a_3998_788.n3 a_3998_788.n0 0.672
R504 a_3998_788.n4 a_3998_788.n3 0.665
R505 a_2830_786.t6 a_2830_786.n3 404.877
R506 a_2830_786.n2 a_2830_786.t7 210.902
R507 a_2830_786.n4 a_2830_786.t6 136.943
R508 a_2830_786.n3 a_2830_786.n2 107.801
R509 a_2830_786.n2 a_2830_786.t8 80.333
R510 a_2830_786.n3 a_2830_786.t5 80.333
R511 a_2830_786.n1 a_2830_786.t3 17.4
R512 a_2830_786.n1 a_2830_786.t4 17.4
R513 a_2830_786.t0 a_2830_786.n5 15.029
R514 a_2830_786.n0 a_2830_786.t2 14.282
R515 a_2830_786.n0 a_2830_786.t1 14.282
R516 a_2830_786.n5 a_2830_786.n0 1.647
R517 a_2830_786.n4 a_2830_786.n1 0.672
R518 a_2830_786.n5 a_2830_786.n4 0.665
R519 Y[2].n0 Y[2].t3 28.57
R520 Y[2].n1 Y[2].t2 28.565
R521 Y[2].n1 Y[2].t1 28.565
R522 Y[2].n0 Y[2].t0 17.638
R523 Y[2].n2 Y[2].n1 0.69
R524 Y[2].n2 Y[2].n0 0.6
R525 Y[2] Y[2].n2 0.188
R526 Y[2] Y[2].n3 0.057
R527 Y[2].n3 Y[2] 0.052
R528 Y[2].n3 Y[2] 0.022
R529 a_5172_790.t5 a_5172_790.n3 403.87
R530 a_5172_790.n2 a_5172_790.t6 191.682
R531 a_5172_790.n4 a_5172_790.t5 138.55
R532 a_5172_790.n3 a_5172_790.n2 111.349
R533 a_5172_790.n2 a_5172_790.t7 80.333
R534 a_5172_790.n3 a_5172_790.t8 80.333
R535 a_5172_790.n1 a_5172_790.t2 17.4
R536 a_5172_790.n1 a_5172_790.t0 17.4
R537 a_5172_790.t1 a_5172_790.n5 15.036
R538 a_5172_790.n0 a_5172_790.t4 14.282
R539 a_5172_790.n0 a_5172_790.t3 14.282
R540 a_5172_790.n5 a_5172_790.n0 1.654
R541 a_5172_790.n4 a_5172_790.n1 0.679
R542 a_5172_790.n5 a_5172_790.n4 0.665
R543 Y[4].n0 Y[4].t1 28.57
R544 Y[4].n1 Y[4].t3 28.565
R545 Y[4].n1 Y[4].t2 28.565
R546 Y[4].n0 Y[4].t0 17.636
R547 Y[4].n2 Y[4].n1 0.712
R548 Y[4].n2 Y[4].n0 0.605
R549 Y[4] Y[4].n2 0.188
R550 Y[4] Y[4].n3 0.057
R551 Y[4].n3 Y[4] 0.052
R552 Y[4].n3 Y[4] 0.022
R553 B[2].t2 B[2].t3 799.268
R554 B[2] B[2].n1 627.607
R555 B[2].n0 B[2].t0 285.543
R556 B[2].n1 B[2].t2 194.406
R557 B[2].n0 B[2].t1 160.666
R558 B[2].n1 B[2].n0 91.137
R559 a_2948_786.n0 a_2948_786.t3 14.282
R560 a_2948_786.n0 a_2948_786.t2 14.282
R561 a_2948_786.n1 a_2948_786.t5 14.282
R562 a_2948_786.n1 a_2948_786.t4 14.282
R563 a_2948_786.n3 a_2948_786.t1 14.282
R564 a_2948_786.t0 a_2948_786.n3 14.282
R565 a_2948_786.n3 a_2948_786.n2 2.554
R566 a_2948_786.n2 a_2948_786.n1 2.361
R567 a_2948_786.n2 a_2948_786.n0 0.001
R568 B[6].t0 B[6].t3 800.875
R569 B[6] B[6].n1 627.607
R570 B[6].n0 B[6].t1 284.688
R571 B[6].n1 B[6].t0 192.799
R572 B[6].n0 B[6].t2 160.666
R573 B[6].n1 B[6].n0 91.889
R574 a_7626_790.n0 a_7626_790.t5 14.282
R575 a_7626_790.n0 a_7626_790.t1 14.282
R576 a_7626_790.n1 a_7626_790.t4 14.282
R577 a_7626_790.n1 a_7626_790.t3 14.282
R578 a_7626_790.t2 a_7626_790.n3 14.282
R579 a_7626_790.n3 a_7626_790.t0 14.282
R580 a_7626_790.n3 a_7626_790.n2 2.538
R581 a_7626_790.n2 a_7626_790.n1 2.375
R582 a_7626_790.n2 a_7626_790.n0 0.001
R583 A[4].t3 A[4].t2 576.841
R584 A[4].n0 A[4].t0 284.688
R585 A[4].n0 A[4].t1 160.666
R586 A[4].n1 A[4].t3 160.666
R587 A[4] A[4].n1 159.954
R588 A[4].n1 A[4].n0 115.593
R589 Y[1].n0 Y[1].t1 28.57
R590 Y[1].n1 Y[1].t3 28.565
R591 Y[1].n1 Y[1].t2 28.565
R592 Y[1].n0 Y[1].t0 17.638
R593 Y[1].n2 Y[1].n1 0.69
R594 Y[1].n2 Y[1].n0 0.6
R595 Y[1] Y[1].n2 0.188
R596 Y[1] Y[1].n3 0.057
R597 Y[1].n3 Y[1] 0.052
R598 Y[1].n3 Y[1] 0.022
R599 B[7].t1 B[7].t3 799.268
R600 B[7] B[7].n1 627.607
R601 B[7].n0 B[7].t0 285.543
R602 B[7].n1 B[7].t1 194.406
R603 B[7].n0 B[7].t2 160.666
R604 B[7].n1 B[7].n0 91.137
R605 Y[7].n0 Y[7].t1 28.57
R606 Y[7].n1 Y[7].t3 28.565
R607 Y[7].n1 Y[7].t2 28.565
R608 Y[7].n0 Y[7].t0 17.638
R609 Y[7].n2 Y[7].n1 0.712
R610 Y[7].n2 Y[7].n0 0.605
R611 Y[7] Y[7].n2 0.188
R612 Y[7] Y[7].n3 0.057
R613 Y[7].n3 Y[7] 0.052
R614 Y[7].n3 Y[7] 0.022
R615 Y[5].n0 Y[5].t1 28.57
R616 Y[5].n1 Y[5].t3 28.565
R617 Y[5].n1 Y[5].t2 28.565
R618 Y[5].n0 Y[5].t0 17.638
R619 Y[5].n2 Y[5].n1 0.716
R620 Y[5].n2 Y[5].n0 0.607
R621 Y[5] Y[5].n2 0.188
R622 Y[5] Y[5].n3 0.057
R623 Y[5].n3 Y[5] 0.052
R624 Y[5].n3 Y[5] 0.022
R625 B[5].t2 B[5].t3 800.874
R626 B[5] B[5].n1 627.607
R627 B[5].n0 B[5].t0 285.543
R628 B[5].n1 B[5].t2 194.406
R629 B[5].n0 B[5].t1 160.666
R630 B[5].n1 B[5].n0 91.137
R631 B[3].t3 B[3].t2 800.875
R632 B[3] B[3].n1 627.607
R633 B[3].n0 B[3].t0 284.688
R634 B[3].n1 B[3].t3 192.799
R635 B[3].n0 B[3].t1 160.666
R636 B[3].n1 B[3].n0 91.889
R637 a_4116_788.n1 a_4116_788.t0 14.282
R638 a_4116_788.n1 a_4116_788.t5 14.282
R639 a_4116_788.n0 a_4116_788.t4 14.282
R640 a_4116_788.n0 a_4116_788.t3 14.282
R641 a_4116_788.t2 a_4116_788.n3 14.282
R642 a_4116_788.n3 a_4116_788.t1 14.282
R643 a_4116_788.n2 a_4116_788.n0 2.538
R644 a_4116_788.n3 a_4116_788.n2 2.375
R645 a_4116_788.n2 a_4116_788.n1 0.001
R646 A[2].t3 A[2].t0 573.627
R647 A[2].n0 A[2].t1 285.543
R648 A[2].n0 A[2].t2 160.666
R649 A[2].n1 A[2].t3 160.666
R650 A[2] A[2].n1 159.202
R651 A[2].n1 A[2].n0 114.089
R652 Y[3].n0 Y[3].t2 28.57
R653 Y[3].n1 Y[3].t3 28.565
R654 Y[3].n1 Y[3].t1 28.565
R655 Y[3].n0 Y[3].t0 17.639
R656 Y[3].n2 Y[3].n1 0.69
R657 Y[3].n2 Y[3].n0 0.6
R658 Y[3] Y[3].n2 0.188
R659 Y[3] Y[3].n3 0.057
R660 Y[3].n3 Y[3] 0.052
R661 Y[3].n3 Y[3] 0.022
C0 A[7] Y[5] 0.00fF
C1 A[2] B[1] 0.01fF
C2 B[2] A[2] 0.44fF
C3 VDD A[1] 0.24fF
C4 VDD B[3] 0.48fF
C5 VDD B[5] 0.48fF
C6 A[2] Y[0] 0.00fF
C7 A[7] Y[7] 0.01fF
C8 A[7] B[6] 0.01fF
C9 B[3] A[4] 0.01fF
C10 Y[0] A[0] 0.01fF
C11 B[7] VDD 0.47fF
C12 VDD A[4] 0.24fF
C13 A[1] B[1] 0.44fF
C14 Y[4] B[3] 0.00fF
C15 Y[4] B[5] 0.00fF
C16 Y[2] A[3] 0.00fF
C17 VDD B[1] 0.48fF
C18 B[2] B[3] 0.01fF
C19 Y[4] VDD 0.88fF
C20 B[3] A[5] 0.00fF
C21 A[6] B[4] 0.00fF
C22 B[2] VDD 0.48fF
C23 A[5] B[5] 0.44fF
C24 VDD A[5] 0.24fF
C25 Y[0] A[1] 0.00fF
C26 Y[3] B[4] 0.00fF
C27 Y[0] VDD 0.87fF
C28 Y[6] B[5] 0.00fF
C29 A[2] Y[2] 0.01fF
C30 Y[6] VDD 0.88fF
C31 Y[5] B[5] 0.03fF
C32 Y[4] A[4] 0.01fF
C33 A[7] A[6] 0.01fF
C34 Y[5] VDD 0.88fF
C35 Y[1] B[0] 0.00fF
C36 B[2] A[4] 0.00fF
C37 A[5] A[4] 0.01fF
C38 B[2] B[1] 0.01fF
C39 Y[4] A[5] 0.00fF
C40 Y[1] A[3] 0.00fF
C41 Y[3] A[3] 0.01fF
C42 Y[6] B[7] 0.00fF
C43 Y[0] B[1] 0.00fF
C44 Y[5] A[4] 0.00fF
C45 Y[7] VDD 0.88fF
C46 B[6] B[5] 0.01fF
C47 Y[6] A[5] 0.00fF
C48 VDD B[6] 0.48fF
C49 Y[5] Y[4] 0.01fF
C50 Y[2] A[1] 0.00fF
C51 Y[2] B[3] 0.00fF
C52 A[2] Y[1] 0.00fF
C53 A[2] Y[3] 0.00fF
C54 Y[2] VDD 0.88fF
C55 Y[5] A[5] 0.01fF
C56 Y[5] Y[6] 0.01fF
C57 Y[7] B[7] 0.03fF
C58 B[7] B[6] 0.01fF
C59 Y[1] A[0] 0.00fF
C60 Y[2] A[4] 0.00fF
C61 Y[2] B[1] 0.00fF
C62 A[6] B[5] 0.01fF
C63 VDD A[6] 0.24fF
C64 B[2] Y[2] 0.03fF
C65 Y[1] A[1] 0.01fF
C66 Y[3] B[3] 0.03fF
C67 Y[6] Y[7] 0.01fF
C68 Y[1] VDD 0.88fF
C69 Y[3] VDD 0.88fF
C70 Y[6] B[6] 0.03fF
C71 A[2] B[0] 0.00fF
C72 Y[5] B[6] 0.00fF
C73 A[2] A[3] 0.01fF
C74 Y[4] A[6] 0.00fF
C75 Y[3] A[4] 0.00fF
C76 Y[1] B[1] 0.03fF
C77 A[6] A[5] 0.01fF
C78 B[0] A[0] 0.44fF
C79 B[3] B[4] 0.01fF
C80 Y[3] Y[4] 0.01fF
C81 B[4] B[5] 0.01fF
C82 B[2] Y[1] 0.00fF
C83 VDD B[4] 0.49fF
C84 B[2] Y[3] 0.00fF
C85 Y[7] B[6] 0.00fF
C86 Y[3] A[5] 0.00fF
C87 Y[6] A[6] 0.01fF
C88 Y[0] Y[1] 0.01fF
C89 B[0] A[1] 0.01fF
C90 Y[5] A[6] 0.00fF
C91 B[0] VDD 0.40fF
C92 A[7] B[5] 0.00fF
C93 A[7] VDD 0.24fF
C94 B[4] A[4] 0.44fF
C95 A[3] B[3] 0.44fF
C96 VDD A[3] 0.24fF
C97 Y[4] B[4] 0.03fF
C98 A[5] B[4] 0.01fF
C99 Y[7] A[6] 0.00fF
C100 A[2] A[1] 0.01fF
C101 A[7] B[7] 0.44fF
C102 A[6] B[6] 0.44fF
C103 B[0] B[1] 0.01fF
C104 A[2] VDD 0.24fF
C105 A[3] A[4] 0.01fF
C106 Y[5] B[4] 0.00fF
C107 A[3] B[1] 0.00fF
C108 Y[2] Y[1] 0.01fF
C109 Y[3] Y[2] 0.01fF
C110 Y[4] A[3] 0.00fF
C111 Y[0] B[0] 0.03fF
C112 B[2] A[3] 0.01fF
C113 A[0] A[1] 0.01fF
C114 A[7] Y[6] 0.00fF
C115 VDD A[0] 0.15fF
.ends

