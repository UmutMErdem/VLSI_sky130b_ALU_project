magic
tech sky130B
magscale 1 2
timestamp 1733697342
<< nwell >>
rect 1 6 839 330
<< nmos >>
rect 332 -376 392 -176
rect 450 -376 510 -176
<< pmos >>
rect 95 68 155 268
rect 213 68 273 268
rect 331 68 391 268
rect 449 68 509 268
rect 567 68 627 268
rect 685 68 745 268
<< ndiff >>
rect 274 -188 332 -176
rect 274 -364 286 -188
rect 320 -364 332 -188
rect 274 -376 332 -364
rect 392 -188 450 -176
rect 392 -364 404 -188
rect 438 -364 450 -188
rect 392 -376 450 -364
rect 510 -188 568 -176
rect 510 -364 522 -188
rect 556 -364 568 -188
rect 510 -376 568 -364
<< pdiff >>
rect 37 256 95 268
rect 37 80 49 256
rect 83 80 95 256
rect 37 68 95 80
rect 155 256 213 268
rect 155 80 167 256
rect 201 80 213 256
rect 155 68 213 80
rect 273 256 331 268
rect 273 80 285 256
rect 319 80 331 256
rect 273 68 331 80
rect 391 256 449 268
rect 391 80 403 256
rect 437 80 449 256
rect 391 68 449 80
rect 509 256 567 268
rect 509 80 521 256
rect 555 80 567 256
rect 509 68 567 80
rect 627 256 685 268
rect 627 80 639 256
rect 673 80 685 256
rect 627 68 685 80
rect 745 256 803 268
rect 745 80 757 256
rect 791 80 803 256
rect 745 68 803 80
<< ndiffc >>
rect 286 -364 320 -188
rect 404 -364 438 -188
rect 522 -364 556 -188
<< pdiffc >>
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
<< poly >>
rect 95 289 391 325
rect 95 268 155 289
rect 213 268 273 289
rect 331 268 391 289
rect 449 288 745 324
rect 449 268 509 288
rect 567 268 627 288
rect 685 268 745 288
rect 95 42 155 68
rect 213 42 273 68
rect 331 42 391 68
rect 449 42 509 68
rect 567 42 627 68
rect 685 42 745 68
rect 332 -150 390 42
rect 450 -150 508 42
rect 332 -176 392 -150
rect 450 -176 510 -150
rect 332 -398 392 -376
rect 450 -398 510 -376
rect 329 -414 395 -398
rect 329 -448 345 -414
rect 379 -448 395 -414
rect 329 -464 395 -448
rect 447 -414 513 -398
rect 447 -448 463 -414
rect 497 -448 513 -414
rect 447 -464 513 -448
<< polycont >>
rect 345 -448 379 -414
rect 463 -448 497 -414
<< locali >>
rect 49 256 83 272
rect 49 64 83 80
rect 167 256 201 272
rect 167 64 201 80
rect 285 256 319 272
rect 285 64 319 80
rect 403 256 437 272
rect 403 64 437 80
rect 521 256 555 272
rect 521 64 555 80
rect 639 256 673 272
rect 639 64 673 80
rect 757 256 791 272
rect 757 64 791 80
rect 286 -188 320 -172
rect 286 -380 320 -364
rect 404 -188 438 -172
rect 404 -380 438 -364
rect 522 -188 556 -172
rect 522 -380 556 -364
rect 329 -448 345 -414
rect 379 -448 395 -414
rect 447 -448 463 -414
rect 497 -448 513 -414
<< viali >>
rect 49 80 83 256
rect 167 80 201 256
rect 285 80 319 256
rect 403 80 437 256
rect 521 80 555 256
rect 639 80 673 256
rect 757 80 791 256
rect 286 -364 320 -188
rect 404 -364 438 -188
rect 522 -364 556 -188
rect 345 -448 379 -414
rect 463 -448 497 -414
<< metal1 >>
rect 386 522 446 532
rect 386 452 446 462
rect 394 404 434 452
rect 50 374 790 404
rect 50 268 82 374
rect 286 268 318 374
rect 522 268 554 374
rect 758 268 790 374
rect 43 256 89 268
rect 43 80 49 256
rect 83 80 89 256
rect 43 68 89 80
rect 161 256 207 268
rect 161 80 167 256
rect 201 80 207 256
rect 161 68 207 80
rect 279 256 325 268
rect 279 80 285 256
rect 319 80 325 256
rect 279 68 325 80
rect 397 256 443 268
rect 397 80 403 256
rect 437 80 443 256
rect 397 68 443 80
rect 515 256 561 268
rect 515 80 521 256
rect 555 80 561 256
rect 515 68 561 80
rect 633 256 679 268
rect 633 80 639 256
rect 673 80 679 256
rect 633 68 679 80
rect 751 256 797 268
rect 751 80 757 256
rect 791 80 797 256
rect 751 68 797 80
rect 166 -26 202 68
rect 402 -26 438 68
rect 638 -24 674 68
rect 638 -26 836 -24
rect 166 -56 836 -26
rect 286 -176 320 -56
rect 642 -58 836 -56
rect 736 -124 836 -58
rect 280 -188 326 -176
rect 280 -364 286 -188
rect 320 -364 326 -188
rect 280 -376 326 -364
rect 398 -188 444 -176
rect 398 -364 404 -188
rect 438 -364 444 -188
rect 398 -376 444 -364
rect 516 -188 562 -176
rect 516 -364 522 -188
rect 556 -340 562 -188
rect 694 -340 704 -332
rect 556 -364 704 -340
rect 516 -376 704 -364
rect 522 -380 704 -376
rect 58 -408 158 -380
rect 694 -392 704 -380
rect 764 -392 774 -332
rect 58 -414 392 -408
rect 58 -448 345 -414
rect 379 -448 392 -414
rect 58 -456 392 -448
rect 450 -414 512 -408
rect 450 -448 463 -414
rect 497 -448 512 -414
rect 58 -480 158 -456
rect 58 -544 158 -522
rect 450 -544 512 -448
rect 58 -592 512 -544
rect 58 -622 158 -592
<< via1 >>
rect 386 462 446 522
rect 704 -392 764 -332
<< metal2 >>
rect 366 452 376 532
rect 456 452 466 532
rect 694 -322 774 -312
rect 694 -412 774 -402
<< via2 >>
rect 376 522 456 532
rect 376 462 386 522
rect 386 462 446 522
rect 446 462 456 522
rect 376 452 456 462
rect 694 -332 774 -322
rect 694 -392 704 -332
rect 704 -392 764 -332
rect 764 -392 774 -332
rect 694 -402 774 -392
<< metal3 >>
rect 360 610 472 620
rect 360 530 366 610
rect 466 530 472 610
rect 366 432 466 442
rect 674 -412 684 -312
rect 784 -412 794 -312
<< via3 >>
rect 366 532 466 610
rect 366 452 376 532
rect 376 452 456 532
rect 456 452 466 532
rect 366 442 466 452
rect 684 -322 784 -312
rect 684 -402 694 -322
rect 694 -402 774 -322
rect 774 -402 784 -322
rect 684 -412 784 -402
<< metal4 >>
rect 316 610 540 642
rect 316 494 366 610
rect 365 442 366 494
rect 466 494 540 610
rect 466 442 467 494
rect 365 441 467 442
rect 742 -311 910 -302
rect 683 -312 910 -311
rect 683 -412 684 -312
rect 784 -412 910 -312
rect 683 -413 910 -412
rect 742 -492 910 -413
<< labels >>
flabel metal4 760 -452 880 -348 1 FreeSans 480 0 0 0 VSS
port 1 n
flabel metal1 58 -622 158 -522 1 FreeSans 480 0 0 0 B
port 3 n
flabel metal1 58 -480 158 -380 1 FreeSans 480 0 0 0 A
port 2 n
flabel metal1 736 -124 836 -24 1 FreeSans 480 0 0 0 Y
port 5 n
flabel metal4 322 498 522 640 1 FreeSans 480 0 0 0 VDD
port 4 n
<< end >>
