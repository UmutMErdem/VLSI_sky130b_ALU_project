magic
tech sky130B
magscale 1 2
timestamp 1736542081
<< nwell >>
rect 546 772 1022 964
rect 2614 774 3090 964
rect 356 476 1200 772
rect 2424 478 3268 774
rect 4683 772 5159 964
rect 6751 774 7227 964
rect 8820 774 9296 966
rect 10888 776 11364 966
rect 4493 476 5337 772
rect 6561 478 7405 774
rect 8630 478 9474 774
rect 10698 480 11542 776
rect 12957 774 13433 966
rect 15025 776 15501 966
rect 12767 478 13611 774
rect 14835 480 15679 776
rect -31 181 265 198
rect -77 153 265 181
rect 807 173 1096 196
rect 2037 183 2333 200
rect 302 -60 1140 173
rect 1991 155 2333 183
rect 2875 175 3164 198
rect 4106 181 4402 198
rect 2370 -58 3208 175
rect 4060 153 4402 181
rect 4944 173 5233 196
rect 6174 183 6470 200
rect 4439 -60 5277 173
rect 6128 155 6470 183
rect 7012 175 7301 198
rect 8243 183 8539 200
rect 6507 -58 7345 175
rect 8197 155 8539 183
rect 9081 175 9370 198
rect 10311 185 10607 202
rect 8576 -58 9414 175
rect 10265 157 10607 185
rect 11149 177 11438 200
rect 12380 183 12676 200
rect 10644 -56 11482 177
rect 12334 155 12676 183
rect 13218 175 13507 198
rect 14448 185 14744 202
rect 12713 -58 13551 175
rect 14402 157 14744 185
rect 15286 177 15575 200
rect 14781 -56 15619 177
<< psubdiff >>
rect 600 -1386 852 -1366
rect 600 -1442 658 -1386
rect 790 -1442 852 -1386
rect 600 -1464 852 -1442
rect 2668 -1384 2920 -1364
rect 2668 -1440 2726 -1384
rect 2858 -1440 2920 -1384
rect 2668 -1462 2920 -1440
rect 4737 -1386 4989 -1366
rect 4737 -1442 4795 -1386
rect 4927 -1442 4989 -1386
rect 4737 -1464 4989 -1442
rect 6805 -1384 7057 -1364
rect 6805 -1440 6863 -1384
rect 6995 -1440 7057 -1384
rect 6805 -1462 7057 -1440
rect 8874 -1384 9126 -1364
rect 8874 -1440 8932 -1384
rect 9064 -1440 9126 -1384
rect 8874 -1462 9126 -1440
rect 10942 -1382 11194 -1362
rect 10942 -1438 11000 -1382
rect 11132 -1438 11194 -1382
rect 10942 -1460 11194 -1438
rect 13011 -1384 13263 -1364
rect 13011 -1440 13069 -1384
rect 13201 -1440 13263 -1384
rect 13011 -1462 13263 -1440
rect 15079 -1382 15331 -1362
rect 15079 -1438 15137 -1382
rect 15269 -1438 15331 -1382
rect 15079 -1460 15331 -1438
<< nsubdiff >>
rect 584 874 984 926
rect 584 830 708 874
rect 830 830 984 874
rect 584 782 984 830
rect 2652 876 3052 928
rect 2652 832 2776 876
rect 2898 832 3052 876
rect 2652 784 3052 832
rect 4721 874 5121 926
rect 4721 830 4845 874
rect 4967 830 5121 874
rect 4721 782 5121 830
rect 6789 876 7189 928
rect 6789 832 6913 876
rect 7035 832 7189 876
rect 6789 784 7189 832
rect 8858 876 9258 928
rect 8858 832 8982 876
rect 9104 832 9258 876
rect 8858 784 9258 832
rect 10926 878 11326 930
rect 10926 834 11050 878
rect 11172 834 11326 878
rect 10926 786 11326 834
rect 12995 876 13395 928
rect 12995 832 13119 876
rect 13241 832 13395 876
rect 12995 784 13395 832
rect 15063 878 15463 930
rect 15063 834 15187 878
rect 15309 834 15463 878
rect 15063 786 15463 834
<< psubdiffcont >>
rect 658 -1442 790 -1386
rect 2726 -1440 2858 -1384
rect 4795 -1442 4927 -1386
rect 6863 -1440 6995 -1384
rect 8932 -1440 9064 -1384
rect 11000 -1438 11132 -1382
rect 13069 -1440 13201 -1384
rect 15137 -1438 15269 -1382
<< nsubdiffcont >>
rect 708 830 830 874
rect 2776 832 2898 876
rect 4845 830 4967 874
rect 6913 832 7035 876
rect 8982 832 9104 876
rect 11050 834 11172 878
rect 13119 832 13241 876
rect 15187 834 15309 878
<< poly >>
rect 453 630 749 681
rect 2521 632 2817 683
rect 4590 630 4886 681
rect 6658 632 6954 683
rect 8727 632 9023 683
rect 10795 634 11091 685
rect 12864 632 13160 683
rect 14932 634 15228 685
rect 1290 432 1586 483
rect 3358 434 3654 485
rect 5427 432 5723 483
rect 7495 434 7791 485
rect 9564 434 9860 485
rect 11632 436 11928 487
rect 13701 434 13997 485
rect 15769 436 16065 487
rect -31 147 513 198
rect 1408 196 1467 214
rect 94 -132 154 147
rect 807 145 1350 196
rect 1392 145 1467 196
rect 2037 149 2581 200
rect 3476 198 3535 216
rect 1392 58 1452 145
rect 1324 48 1452 58
rect 1324 14 1340 48
rect 1374 14 1452 48
rect 396 -55 692 5
rect 750 -54 1046 6
rect 1324 4 1452 14
rect 750 -55 810 -54
rect 868 -55 928 -54
rect 986 -55 1046 -54
rect -70 -146 154 -132
rect -70 -180 -54 -146
rect -20 -180 154 -146
rect -70 -192 154 -180
rect 94 -705 154 -192
rect 364 -645 431 -638
rect 514 -645 574 -497
rect 364 -654 574 -645
rect 364 -688 380 -654
rect 414 -688 574 -654
rect 364 -704 574 -688
rect 94 -721 245 -705
rect 94 -755 195 -721
rect 229 -755 245 -721
rect 94 -771 245 -755
rect 94 -800 154 -771
rect 514 -801 574 -704
rect 868 -645 928 -497
rect 1011 -645 1078 -638
rect 868 -654 1078 -645
rect 868 -688 1028 -654
rect 1062 -688 1078 -654
rect 868 -704 1078 -688
rect 630 -738 696 -722
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 630 -788 696 -772
rect 748 -737 814 -722
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 748 -787 814 -771
rect 632 -800 692 -788
rect 750 -799 810 -787
rect 868 -801 928 -704
rect 1392 -706 1452 4
rect 2162 -130 2222 149
rect 2875 147 3418 198
rect 3460 147 3535 198
rect 4106 147 4650 198
rect 5545 196 5604 214
rect 3460 60 3520 147
rect 3392 50 3520 60
rect 3392 16 3408 50
rect 3442 16 3520 50
rect 2464 -53 2760 7
rect 2818 -52 3114 8
rect 3392 6 3520 16
rect 2818 -53 2878 -52
rect 2936 -53 2996 -52
rect 3054 -53 3114 -52
rect 1998 -144 2222 -130
rect 1998 -178 2014 -144
rect 2048 -178 2222 -144
rect 1998 -190 2222 -178
rect 1302 -722 1452 -706
rect 1302 -756 1318 -722
rect 1352 -756 1452 -722
rect 1302 -772 1452 -756
rect 1392 -800 1452 -772
rect 2162 -703 2222 -190
rect 2432 -643 2499 -636
rect 2582 -643 2642 -495
rect 2432 -652 2642 -643
rect 2432 -686 2448 -652
rect 2482 -686 2642 -652
rect 2432 -702 2642 -686
rect 2162 -719 2313 -703
rect 2162 -753 2263 -719
rect 2297 -753 2313 -719
rect 2162 -769 2313 -753
rect 2162 -798 2222 -769
rect 2582 -799 2642 -702
rect 2936 -643 2996 -495
rect 3079 -643 3146 -636
rect 2936 -652 3146 -643
rect 2936 -686 3096 -652
rect 3130 -686 3146 -652
rect 2936 -702 3146 -686
rect 2698 -736 2764 -720
rect 2698 -770 2714 -736
rect 2748 -770 2764 -736
rect 2698 -786 2764 -770
rect 2816 -735 2882 -720
rect 2816 -769 2832 -735
rect 2866 -769 2882 -735
rect 2816 -785 2882 -769
rect 2700 -798 2760 -786
rect 2818 -797 2878 -785
rect 2936 -799 2996 -702
rect 3460 -704 3520 6
rect 4231 -132 4291 147
rect 4944 145 5487 196
rect 5529 145 5604 196
rect 6174 149 6718 200
rect 7613 198 7672 216
rect 5529 58 5589 145
rect 5461 48 5589 58
rect 5461 14 5477 48
rect 5511 14 5589 48
rect 4533 -55 4829 5
rect 4887 -54 5183 6
rect 5461 4 5589 14
rect 4887 -55 4947 -54
rect 5005 -55 5065 -54
rect 5123 -55 5183 -54
rect 4067 -146 4291 -132
rect 4067 -180 4083 -146
rect 4117 -180 4291 -146
rect 4067 -192 4291 -180
rect 3370 -720 3520 -704
rect 3370 -754 3386 -720
rect 3420 -754 3520 -720
rect 3370 -770 3520 -754
rect 3460 -798 3520 -770
rect 4231 -705 4291 -192
rect 4501 -645 4568 -638
rect 4651 -645 4711 -497
rect 4501 -654 4711 -645
rect 4501 -688 4517 -654
rect 4551 -688 4711 -654
rect 4501 -704 4711 -688
rect 4231 -721 4382 -705
rect 4231 -755 4332 -721
rect 4366 -755 4382 -721
rect 4231 -771 4382 -755
rect 4231 -800 4291 -771
rect 4651 -801 4711 -704
rect 5005 -645 5065 -497
rect 5148 -645 5215 -638
rect 5005 -654 5215 -645
rect 5005 -688 5165 -654
rect 5199 -688 5215 -654
rect 5005 -704 5215 -688
rect 4767 -738 4833 -722
rect 4767 -772 4783 -738
rect 4817 -772 4833 -738
rect 4767 -788 4833 -772
rect 4885 -737 4951 -722
rect 4885 -771 4901 -737
rect 4935 -771 4951 -737
rect 4885 -787 4951 -771
rect 4769 -800 4829 -788
rect 4887 -799 4947 -787
rect 5005 -801 5065 -704
rect 5529 -706 5589 4
rect 6299 -130 6359 149
rect 7012 147 7555 198
rect 7597 147 7672 198
rect 8243 149 8787 200
rect 9682 198 9741 216
rect 7597 60 7657 147
rect 7529 50 7657 60
rect 7529 16 7545 50
rect 7579 16 7657 50
rect 6601 -53 6897 7
rect 6955 -52 7251 8
rect 7529 6 7657 16
rect 6955 -53 7015 -52
rect 7073 -53 7133 -52
rect 7191 -53 7251 -52
rect 6135 -144 6359 -130
rect 6135 -178 6151 -144
rect 6185 -178 6359 -144
rect 6135 -190 6359 -178
rect 5439 -722 5589 -706
rect 5439 -756 5455 -722
rect 5489 -756 5589 -722
rect 5439 -772 5589 -756
rect 5529 -800 5589 -772
rect 6299 -703 6359 -190
rect 6569 -643 6636 -636
rect 6719 -643 6779 -495
rect 6569 -652 6779 -643
rect 6569 -686 6585 -652
rect 6619 -686 6779 -652
rect 6569 -702 6779 -686
rect 6299 -719 6450 -703
rect 6299 -753 6400 -719
rect 6434 -753 6450 -719
rect 6299 -769 6450 -753
rect 6299 -798 6359 -769
rect 6719 -799 6779 -702
rect 7073 -643 7133 -495
rect 7216 -643 7283 -636
rect 7073 -652 7283 -643
rect 7073 -686 7233 -652
rect 7267 -686 7283 -652
rect 7073 -702 7283 -686
rect 6835 -736 6901 -720
rect 6835 -770 6851 -736
rect 6885 -770 6901 -736
rect 6835 -786 6901 -770
rect 6953 -735 7019 -720
rect 6953 -769 6969 -735
rect 7003 -769 7019 -735
rect 6953 -785 7019 -769
rect 6837 -798 6897 -786
rect 6955 -797 7015 -785
rect 7073 -799 7133 -702
rect 7597 -704 7657 6
rect 8368 -130 8428 149
rect 9081 147 9624 198
rect 9666 147 9741 198
rect 10311 151 10855 202
rect 11750 200 11809 218
rect 9666 60 9726 147
rect 9598 50 9726 60
rect 9598 16 9614 50
rect 9648 16 9726 50
rect 8670 -53 8966 7
rect 9024 -52 9320 8
rect 9598 6 9726 16
rect 9024 -53 9084 -52
rect 9142 -53 9202 -52
rect 9260 -53 9320 -52
rect 8204 -144 8428 -130
rect 8204 -178 8220 -144
rect 8254 -178 8428 -144
rect 8204 -190 8428 -178
rect 7507 -720 7657 -704
rect 7507 -754 7523 -720
rect 7557 -754 7657 -720
rect 7507 -770 7657 -754
rect 7597 -798 7657 -770
rect 8368 -703 8428 -190
rect 8638 -643 8705 -636
rect 8788 -643 8848 -495
rect 8638 -652 8848 -643
rect 8638 -686 8654 -652
rect 8688 -686 8848 -652
rect 8638 -702 8848 -686
rect 8368 -719 8519 -703
rect 8368 -753 8469 -719
rect 8503 -753 8519 -719
rect 8368 -769 8519 -753
rect 8368 -798 8428 -769
rect 8788 -799 8848 -702
rect 9142 -643 9202 -495
rect 9285 -643 9352 -636
rect 9142 -652 9352 -643
rect 9142 -686 9302 -652
rect 9336 -686 9352 -652
rect 9142 -702 9352 -686
rect 8904 -736 8970 -720
rect 8904 -770 8920 -736
rect 8954 -770 8970 -736
rect 8904 -786 8970 -770
rect 9022 -735 9088 -720
rect 9022 -769 9038 -735
rect 9072 -769 9088 -735
rect 9022 -785 9088 -769
rect 8906 -798 8966 -786
rect 9024 -797 9084 -785
rect 9142 -799 9202 -702
rect 9666 -704 9726 6
rect 10436 -128 10496 151
rect 11149 149 11692 200
rect 11734 149 11809 200
rect 12380 149 12924 200
rect 13819 198 13878 216
rect 11734 62 11794 149
rect 11666 52 11794 62
rect 11666 18 11682 52
rect 11716 18 11794 52
rect 10738 -51 11034 9
rect 11092 -50 11388 10
rect 11666 8 11794 18
rect 11092 -51 11152 -50
rect 11210 -51 11270 -50
rect 11328 -51 11388 -50
rect 10272 -142 10496 -128
rect 10272 -176 10288 -142
rect 10322 -176 10496 -142
rect 10272 -188 10496 -176
rect 9576 -720 9726 -704
rect 9576 -754 9592 -720
rect 9626 -754 9726 -720
rect 9576 -770 9726 -754
rect 9666 -798 9726 -770
rect 10436 -701 10496 -188
rect 10706 -641 10773 -634
rect 10856 -641 10916 -493
rect 10706 -650 10916 -641
rect 10706 -684 10722 -650
rect 10756 -684 10916 -650
rect 10706 -700 10916 -684
rect 10436 -717 10587 -701
rect 10436 -751 10537 -717
rect 10571 -751 10587 -717
rect 10436 -767 10587 -751
rect 10436 -796 10496 -767
rect 10856 -797 10916 -700
rect 11210 -641 11270 -493
rect 11353 -641 11420 -634
rect 11210 -650 11420 -641
rect 11210 -684 11370 -650
rect 11404 -684 11420 -650
rect 11210 -700 11420 -684
rect 10972 -734 11038 -718
rect 10972 -768 10988 -734
rect 11022 -768 11038 -734
rect 10972 -784 11038 -768
rect 11090 -733 11156 -718
rect 11090 -767 11106 -733
rect 11140 -767 11156 -733
rect 11090 -783 11156 -767
rect 10974 -796 11034 -784
rect 11092 -795 11152 -783
rect 11210 -797 11270 -700
rect 11734 -702 11794 8
rect 12505 -130 12565 149
rect 13218 147 13761 198
rect 13803 147 13878 198
rect 14448 151 14992 202
rect 15887 200 15946 218
rect 13803 60 13863 147
rect 13735 50 13863 60
rect 13735 16 13751 50
rect 13785 16 13863 50
rect 12807 -53 13103 7
rect 13161 -52 13457 8
rect 13735 6 13863 16
rect 13161 -53 13221 -52
rect 13279 -53 13339 -52
rect 13397 -53 13457 -52
rect 12341 -144 12565 -130
rect 12341 -178 12357 -144
rect 12391 -178 12565 -144
rect 12341 -190 12565 -178
rect 11644 -718 11794 -702
rect 11644 -752 11660 -718
rect 11694 -752 11794 -718
rect 11644 -768 11794 -752
rect 11734 -796 11794 -768
rect 12505 -703 12565 -190
rect 12775 -643 12842 -636
rect 12925 -643 12985 -495
rect 12775 -652 12985 -643
rect 12775 -686 12791 -652
rect 12825 -686 12985 -652
rect 12775 -702 12985 -686
rect 12505 -719 12656 -703
rect 12505 -753 12606 -719
rect 12640 -753 12656 -719
rect 12505 -769 12656 -753
rect 12505 -798 12565 -769
rect 12925 -799 12985 -702
rect 13279 -643 13339 -495
rect 13422 -643 13489 -636
rect 13279 -652 13489 -643
rect 13279 -686 13439 -652
rect 13473 -686 13489 -652
rect 13279 -702 13489 -686
rect 13041 -736 13107 -720
rect 13041 -770 13057 -736
rect 13091 -770 13107 -736
rect 13041 -786 13107 -770
rect 13159 -735 13225 -720
rect 13159 -769 13175 -735
rect 13209 -769 13225 -735
rect 13159 -785 13225 -769
rect 13043 -798 13103 -786
rect 13161 -797 13221 -785
rect 13279 -799 13339 -702
rect 13803 -704 13863 6
rect 14573 -128 14633 151
rect 15286 149 15829 200
rect 15871 149 15946 200
rect 15871 62 15931 149
rect 15803 52 15931 62
rect 15803 18 15819 52
rect 15853 18 15931 52
rect 14875 -51 15171 9
rect 15229 -50 15525 10
rect 15803 8 15931 18
rect 15229 -51 15289 -50
rect 15347 -51 15407 -50
rect 15465 -51 15525 -50
rect 14409 -142 14633 -128
rect 14409 -176 14425 -142
rect 14459 -176 14633 -142
rect 14409 -188 14633 -176
rect 13713 -720 13863 -704
rect 13713 -754 13729 -720
rect 13763 -754 13863 -720
rect 13713 -770 13863 -754
rect 13803 -798 13863 -770
rect 14573 -701 14633 -188
rect 14843 -641 14910 -634
rect 14993 -641 15053 -493
rect 14843 -650 15053 -641
rect 14843 -684 14859 -650
rect 14893 -684 15053 -650
rect 14843 -700 15053 -684
rect 14573 -717 14724 -701
rect 14573 -751 14674 -717
rect 14708 -751 14724 -717
rect 14573 -767 14724 -751
rect 14573 -796 14633 -767
rect 14993 -797 15053 -700
rect 15347 -641 15407 -493
rect 15490 -641 15557 -634
rect 15347 -650 15557 -641
rect 15347 -684 15507 -650
rect 15541 -684 15557 -650
rect 15347 -700 15557 -684
rect 15109 -734 15175 -718
rect 15109 -768 15125 -734
rect 15159 -768 15175 -734
rect 15109 -784 15175 -768
rect 15227 -733 15293 -718
rect 15227 -767 15243 -733
rect 15277 -767 15293 -733
rect 15227 -783 15293 -767
rect 15111 -796 15171 -784
rect 15229 -795 15289 -783
rect 15347 -797 15407 -700
rect 15871 -702 15931 8
rect 15781 -718 15931 -702
rect 15781 -752 15797 -718
rect 15831 -752 15931 -718
rect 15781 -768 15931 -752
rect 15871 -796 15931 -768
<< polycont >>
rect 1340 14 1374 48
rect -54 -180 -20 -146
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1028 -688 1062 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 3408 16 3442 50
rect 2014 -178 2048 -144
rect 1318 -756 1352 -722
rect 2448 -686 2482 -652
rect 2263 -753 2297 -719
rect 3096 -686 3130 -652
rect 2714 -770 2748 -736
rect 2832 -769 2866 -735
rect 5477 14 5511 48
rect 4083 -180 4117 -146
rect 3386 -754 3420 -720
rect 4517 -688 4551 -654
rect 4332 -755 4366 -721
rect 5165 -688 5199 -654
rect 4783 -772 4817 -738
rect 4901 -771 4935 -737
rect 7545 16 7579 50
rect 6151 -178 6185 -144
rect 5455 -756 5489 -722
rect 6585 -686 6619 -652
rect 6400 -753 6434 -719
rect 7233 -686 7267 -652
rect 6851 -770 6885 -736
rect 6969 -769 7003 -735
rect 9614 16 9648 50
rect 8220 -178 8254 -144
rect 7523 -754 7557 -720
rect 8654 -686 8688 -652
rect 8469 -753 8503 -719
rect 9302 -686 9336 -652
rect 8920 -770 8954 -736
rect 9038 -769 9072 -735
rect 11682 18 11716 52
rect 10288 -176 10322 -142
rect 9592 -754 9626 -720
rect 10722 -684 10756 -650
rect 10537 -751 10571 -717
rect 11370 -684 11404 -650
rect 10988 -768 11022 -734
rect 11106 -767 11140 -733
rect 13751 16 13785 50
rect 12357 -178 12391 -144
rect 11660 -752 11694 -718
rect 12791 -686 12825 -652
rect 12606 -753 12640 -719
rect 13439 -686 13473 -652
rect 13057 -770 13091 -736
rect 13175 -769 13209 -735
rect 15819 18 15853 52
rect 14425 -176 14459 -142
rect 13729 -754 13763 -720
rect 14859 -684 14893 -650
rect 14674 -751 14708 -717
rect 15507 -684 15541 -650
rect 15125 -768 15159 -734
rect 15243 -767 15277 -733
rect 15797 -752 15831 -718
<< locali >>
rect 674 874 876 894
rect 674 830 708 874
rect 830 830 876 874
rect 674 820 760 830
rect 798 820 876 830
rect 674 802 876 820
rect 2742 876 2944 896
rect 2742 832 2776 876
rect 2898 832 2944 876
rect 2742 822 2828 832
rect 2866 822 2944 832
rect 2742 804 2944 822
rect 4811 874 5013 894
rect 4811 830 4845 874
rect 4967 830 5013 874
rect 4811 820 4897 830
rect 4935 820 5013 830
rect 4811 802 5013 820
rect 6879 876 7081 896
rect 6879 832 6913 876
rect 7035 832 7081 876
rect 6879 822 6965 832
rect 7003 822 7081 832
rect 6879 804 7081 822
rect 8948 876 9150 896
rect 8948 832 8982 876
rect 9104 832 9150 876
rect 8948 822 9034 832
rect 9072 822 9150 832
rect 8948 804 9150 822
rect 11016 878 11218 898
rect 11016 834 11050 878
rect 11172 834 11218 878
rect 11016 824 11102 834
rect 11140 824 11218 834
rect 11016 806 11218 824
rect 13085 876 13287 896
rect 13085 832 13119 876
rect 13241 832 13287 876
rect 13085 822 13171 832
rect 13209 822 13287 832
rect 13085 804 13287 822
rect 15153 878 15355 898
rect 15153 834 15187 878
rect 15309 834 15355 878
rect 15153 824 15239 834
rect 15277 824 15355 834
rect 15153 806 15355 824
rect 761 656 1031 691
rect 761 613 795 656
rect 997 613 1031 656
rect 2829 658 3099 693
rect 2829 615 2863 658
rect 3065 615 3099 658
rect 4898 656 5168 691
rect 4898 613 4932 656
rect 5134 613 5168 656
rect 6966 658 7236 693
rect 6966 615 7000 658
rect 7202 615 7236 658
rect 9035 658 9305 693
rect 9035 615 9069 658
rect 9271 615 9305 658
rect 11103 660 11373 695
rect 11103 617 11137 660
rect 11339 617 11373 660
rect 13172 658 13442 693
rect 13172 615 13206 658
rect 13408 615 13442 658
rect 15240 660 15510 695
rect 15240 617 15274 660
rect 15476 617 15510 660
rect -77 457 193 492
rect -77 415 -43 457
rect 159 415 193 457
rect 1991 459 2261 494
rect 1991 417 2025 459
rect 2227 417 2261 459
rect 4060 457 4330 492
rect 4060 415 4094 457
rect 4296 415 4330 457
rect 6128 459 6398 494
rect 6128 417 6162 459
rect 6364 417 6398 459
rect 8197 459 8467 494
rect 8197 417 8231 459
rect 8433 417 8467 459
rect 10265 461 10535 496
rect 10265 419 10299 461
rect 10501 419 10535 461
rect 12334 459 12604 494
rect 12334 417 12368 459
rect 12570 417 12604 459
rect 14402 461 14672 496
rect 14402 419 14436 461
rect 14638 419 14672 461
rect 1324 14 1330 48
rect 1384 14 1390 48
rect 3392 16 3398 50
rect 3452 16 3458 50
rect 5461 14 5467 48
rect 5521 14 5527 48
rect 7529 16 7535 50
rect 7589 16 7595 50
rect 9598 16 9604 50
rect 9658 16 9664 50
rect 11666 18 11672 52
rect 11726 18 11732 52
rect 13735 16 13741 50
rect 13795 16 13801 50
rect 15803 18 15809 52
rect 15863 18 15869 52
rect 467 -524 503 -419
rect 702 -524 738 -419
rect 940 -524 976 -420
rect 467 -564 1562 -524
rect 486 -565 1562 -564
rect 364 -654 431 -638
rect 364 -688 380 -654
rect 414 -688 431 -654
rect 364 -704 431 -688
rect 195 -721 229 -705
rect 195 -771 229 -755
rect 541 -806 575 -565
rect 2535 -522 2571 -417
rect 2770 -522 2806 -417
rect 3008 -522 3044 -418
rect 2535 -562 3630 -522
rect 2554 -563 3630 -562
rect 1011 -654 1078 -638
rect 1011 -688 1028 -654
rect 1062 -688 1078 -654
rect 1011 -704 1078 -688
rect 2432 -652 2499 -636
rect 2432 -686 2448 -652
rect 2482 -686 2499 -652
rect 2432 -702 2499 -686
rect 1318 -722 1352 -706
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 1318 -772 1352 -756
rect 2263 -719 2297 -703
rect 2263 -769 2297 -753
rect 2609 -804 2643 -563
rect 4604 -524 4640 -419
rect 4839 -524 4875 -419
rect 5077 -524 5113 -420
rect 4604 -564 5699 -524
rect 4623 -565 5699 -564
rect 3079 -652 3146 -636
rect 3079 -686 3096 -652
rect 3130 -686 3146 -652
rect 3079 -702 3146 -686
rect 4501 -654 4568 -638
rect 4501 -688 4517 -654
rect 4551 -688 4568 -654
rect 4501 -704 4568 -688
rect 3386 -720 3420 -704
rect 2698 -770 2714 -736
rect 2748 -770 2764 -736
rect 2816 -769 2832 -735
rect 2866 -769 2882 -735
rect 3386 -770 3420 -754
rect 4332 -721 4366 -705
rect 4332 -771 4366 -755
rect 541 -809 613 -806
rect 2609 -807 2681 -804
rect 4678 -806 4712 -565
rect 6672 -522 6708 -417
rect 6907 -522 6943 -417
rect 7145 -522 7181 -418
rect 6672 -562 7767 -522
rect 6691 -563 7767 -562
rect 5148 -654 5215 -638
rect 5148 -688 5165 -654
rect 5199 -688 5215 -654
rect 5148 -704 5215 -688
rect 6569 -652 6636 -636
rect 6569 -686 6585 -652
rect 6619 -686 6636 -652
rect 6569 -702 6636 -686
rect 5455 -722 5489 -706
rect 4767 -772 4783 -738
rect 4817 -772 4833 -738
rect 4885 -771 4901 -737
rect 4935 -771 4951 -737
rect 5455 -772 5489 -756
rect 6400 -719 6434 -703
rect 6400 -769 6434 -753
rect 6746 -804 6780 -563
rect 8741 -522 8777 -417
rect 8976 -522 9012 -417
rect 9214 -522 9250 -418
rect 8741 -562 9836 -522
rect 8760 -563 9836 -562
rect 7216 -652 7283 -636
rect 7216 -686 7233 -652
rect 7267 -686 7283 -652
rect 7216 -702 7283 -686
rect 8638 -652 8705 -636
rect 8638 -686 8654 -652
rect 8688 -686 8705 -652
rect 8638 -702 8705 -686
rect 7523 -720 7557 -704
rect 6835 -770 6851 -736
rect 6885 -770 6901 -736
rect 6953 -769 6969 -735
rect 7003 -769 7019 -735
rect 7523 -770 7557 -754
rect 8469 -719 8503 -703
rect 8469 -769 8503 -753
rect 8815 -804 8849 -563
rect 10809 -520 10845 -415
rect 11044 -520 11080 -415
rect 11282 -520 11318 -416
rect 10809 -560 11904 -520
rect 10828 -561 11904 -560
rect 9285 -652 9352 -636
rect 9285 -686 9302 -652
rect 9336 -686 9352 -652
rect 9285 -702 9352 -686
rect 10706 -650 10773 -634
rect 10706 -684 10722 -650
rect 10756 -684 10773 -650
rect 10706 -700 10773 -684
rect 9592 -720 9626 -704
rect 8904 -770 8920 -736
rect 8954 -770 8970 -736
rect 9022 -769 9038 -735
rect 9072 -769 9088 -735
rect 9592 -770 9626 -754
rect 10537 -717 10571 -701
rect 10537 -767 10571 -751
rect 10883 -802 10917 -561
rect 12878 -522 12914 -417
rect 13113 -522 13149 -417
rect 13351 -522 13387 -418
rect 12878 -562 13973 -522
rect 12897 -563 13973 -562
rect 11353 -650 11420 -634
rect 11353 -684 11370 -650
rect 11404 -684 11420 -650
rect 11353 -700 11420 -684
rect 12775 -652 12842 -636
rect 12775 -686 12791 -652
rect 12825 -686 12842 -652
rect 12775 -702 12842 -686
rect 11660 -718 11694 -702
rect 10972 -768 10988 -734
rect 11022 -768 11038 -734
rect 11090 -767 11106 -733
rect 11140 -767 11156 -733
rect 11660 -768 11694 -752
rect 12606 -719 12640 -703
rect 12606 -769 12640 -753
rect 541 -852 620 -809
rect 2609 -850 2688 -807
rect 4678 -809 4750 -806
rect 6746 -807 6818 -804
rect 8815 -807 8887 -804
rect 10883 -805 10955 -802
rect 12952 -804 12986 -563
rect 14946 -520 14982 -415
rect 15181 -520 15217 -415
rect 15419 -520 15455 -416
rect 14946 -560 16041 -520
rect 14965 -561 16041 -560
rect 13422 -652 13489 -636
rect 13422 -686 13439 -652
rect 13473 -686 13489 -652
rect 13422 -702 13489 -686
rect 14843 -650 14910 -634
rect 14843 -684 14859 -650
rect 14893 -684 14910 -650
rect 14843 -700 14910 -684
rect 13729 -720 13763 -704
rect 13041 -770 13057 -736
rect 13091 -770 13107 -736
rect 13159 -769 13175 -735
rect 13209 -769 13225 -735
rect 13729 -770 13763 -754
rect 14674 -717 14708 -701
rect 14674 -767 14708 -751
rect 15020 -802 15054 -561
rect 15490 -650 15557 -634
rect 15490 -684 15507 -650
rect 15541 -684 15557 -650
rect 15490 -700 15557 -684
rect 15797 -718 15831 -702
rect 15109 -768 15125 -734
rect 15159 -768 15175 -734
rect 15227 -767 15243 -733
rect 15277 -767 15293 -733
rect 15797 -768 15831 -752
rect 4678 -852 4757 -809
rect 6746 -850 6825 -807
rect 8815 -850 8894 -807
rect 10883 -848 10962 -805
rect 12952 -807 13024 -804
rect 15020 -805 15092 -802
rect 12952 -850 13031 -807
rect 15020 -848 15099 -805
rect 468 -1265 503 -1198
rect 939 -1265 974 -1198
rect 468 -1300 974 -1265
rect 2536 -1263 2571 -1196
rect 3007 -1263 3042 -1196
rect 2536 -1298 3042 -1263
rect 4605 -1265 4640 -1198
rect 5076 -1265 5111 -1198
rect 4605 -1300 5111 -1265
rect 6673 -1263 6708 -1196
rect 7144 -1263 7179 -1196
rect 6673 -1298 7179 -1263
rect 8742 -1263 8777 -1196
rect 9213 -1263 9248 -1196
rect 8742 -1298 9248 -1263
rect 10810 -1261 10845 -1194
rect 11281 -1261 11316 -1194
rect 10810 -1296 11316 -1261
rect 12879 -1263 12914 -1196
rect 13350 -1263 13385 -1196
rect 12879 -1298 13385 -1263
rect 14947 -1261 14982 -1194
rect 15418 -1261 15453 -1194
rect 14947 -1296 15453 -1261
rect 642 -1386 698 -1370
rect 748 -1386 806 -1370
rect 642 -1442 658 -1386
rect 790 -1442 806 -1386
rect 642 -1458 806 -1442
rect 2710 -1384 2766 -1368
rect 2816 -1384 2874 -1368
rect 2710 -1440 2726 -1384
rect 2858 -1440 2874 -1384
rect 2710 -1456 2874 -1440
rect 4779 -1386 4835 -1370
rect 4885 -1386 4943 -1370
rect 4779 -1442 4795 -1386
rect 4927 -1442 4943 -1386
rect 4779 -1458 4943 -1442
rect 6847 -1384 6903 -1368
rect 6953 -1384 7011 -1368
rect 6847 -1440 6863 -1384
rect 6995 -1440 7011 -1384
rect 6847 -1456 7011 -1440
rect 8916 -1384 8972 -1368
rect 9022 -1384 9080 -1368
rect 8916 -1440 8932 -1384
rect 9064 -1440 9080 -1384
rect 8916 -1456 9080 -1440
rect 10984 -1382 11040 -1366
rect 11090 -1382 11148 -1366
rect 10984 -1438 11000 -1382
rect 11132 -1438 11148 -1382
rect 10984 -1454 11148 -1438
rect 13053 -1384 13109 -1368
rect 13159 -1384 13217 -1368
rect 13053 -1440 13069 -1384
rect 13201 -1440 13217 -1384
rect 13053 -1456 13217 -1440
rect 15121 -1382 15177 -1366
rect 15227 -1382 15285 -1366
rect 15121 -1438 15137 -1382
rect 15269 -1438 15285 -1382
rect 15121 -1454 15285 -1438
<< viali >>
rect 760 830 798 858
rect 760 820 798 830
rect 2828 832 2866 860
rect 2828 822 2866 832
rect 4897 830 4935 858
rect 4897 820 4935 830
rect 6965 832 7003 860
rect 6965 822 7003 832
rect 9034 832 9072 860
rect 9034 822 9072 832
rect 11102 834 11140 862
rect 11102 824 11140 834
rect 13171 832 13209 860
rect 13171 822 13209 832
rect 15239 834 15277 862
rect 15239 824 15277 834
rect 1330 48 1384 58
rect 3398 50 3452 60
rect 1330 14 1340 48
rect 1340 14 1374 48
rect 1374 14 1384 48
rect 3398 16 3408 50
rect 3408 16 3442 50
rect 3442 16 3452 50
rect 5467 48 5521 58
rect 7535 50 7589 60
rect 9604 50 9658 60
rect 11672 52 11726 62
rect 1330 4 1384 14
rect 3398 6 3452 16
rect 5467 14 5477 48
rect 5477 14 5511 48
rect 5511 14 5521 48
rect 7535 16 7545 50
rect 7545 16 7579 50
rect 7579 16 7589 50
rect 9604 16 9614 50
rect 9614 16 9648 50
rect 9648 16 9658 50
rect 11672 18 11682 52
rect 11682 18 11716 52
rect 11716 18 11726 52
rect 13741 50 13795 60
rect 15809 52 15863 62
rect 5467 4 5521 14
rect 7535 6 7589 16
rect 9604 6 9658 16
rect 11672 8 11726 18
rect 13741 16 13751 50
rect 13751 16 13785 50
rect 13785 16 13795 50
rect 15809 18 15819 52
rect 15819 18 15853 52
rect 15853 18 15863 52
rect 13741 6 13795 16
rect 15809 8 15863 18
rect -70 -146 -4 -132
rect -70 -180 -54 -146
rect -54 -180 -20 -146
rect -20 -180 -4 -146
rect -70 -192 -4 -180
rect 1998 -144 2064 -130
rect 1998 -178 2014 -144
rect 2014 -178 2048 -144
rect 2048 -178 2064 -144
rect 1998 -190 2064 -178
rect 4067 -146 4133 -132
rect 4067 -180 4083 -146
rect 4083 -180 4117 -146
rect 4117 -180 4133 -146
rect 4067 -192 4133 -180
rect 6135 -144 6201 -130
rect 6135 -178 6151 -144
rect 6151 -178 6185 -144
rect 6185 -178 6201 -144
rect 6135 -190 6201 -178
rect 8204 -144 8270 -130
rect 8204 -178 8220 -144
rect 8220 -178 8254 -144
rect 8254 -178 8270 -144
rect 8204 -190 8270 -178
rect 10272 -142 10338 -128
rect 10272 -176 10288 -142
rect 10288 -176 10322 -142
rect 10322 -176 10338 -142
rect 10272 -188 10338 -176
rect 12341 -144 12407 -130
rect 12341 -178 12357 -144
rect 12357 -178 12391 -144
rect 12391 -178 12407 -144
rect 12341 -190 12407 -178
rect 14409 -142 14475 -128
rect 14409 -176 14425 -142
rect 14425 -176 14459 -142
rect 14459 -176 14475 -142
rect 14409 -188 14475 -176
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1562 -596 1664 -494
rect 1028 -688 1062 -654
rect 2448 -686 2482 -652
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
rect 2263 -753 2297 -719
rect 3630 -594 3732 -492
rect 3096 -686 3130 -652
rect 4517 -688 4551 -654
rect 2714 -770 2748 -736
rect 2832 -769 2866 -735
rect 3386 -754 3420 -720
rect 4332 -755 4366 -721
rect 5699 -596 5801 -494
rect 5165 -688 5199 -654
rect 6585 -686 6619 -652
rect 4783 -772 4817 -738
rect 4901 -771 4935 -737
rect 5455 -756 5489 -722
rect 6400 -753 6434 -719
rect 7767 -594 7869 -492
rect 7233 -686 7267 -652
rect 8654 -686 8688 -652
rect 6851 -770 6885 -736
rect 6969 -769 7003 -735
rect 7523 -754 7557 -720
rect 8469 -753 8503 -719
rect 9836 -594 9938 -492
rect 9302 -686 9336 -652
rect 10722 -684 10756 -650
rect 8920 -770 8954 -736
rect 9038 -769 9072 -735
rect 9592 -754 9626 -720
rect 10537 -751 10571 -717
rect 11904 -592 12006 -490
rect 11370 -684 11404 -650
rect 12791 -686 12825 -652
rect 10988 -768 11022 -734
rect 11106 -767 11140 -733
rect 11660 -752 11694 -718
rect 12606 -753 12640 -719
rect 13973 -594 14075 -492
rect 13439 -686 13473 -652
rect 14859 -684 14893 -650
rect 13057 -770 13091 -736
rect 13175 -769 13209 -735
rect 13729 -754 13763 -720
rect 14674 -751 14708 -717
rect 16041 -592 16143 -490
rect 15507 -684 15541 -650
rect 15125 -768 15159 -734
rect 15243 -767 15277 -733
rect 15797 -752 15831 -718
rect 698 -1386 748 -1364
rect 698 -1406 748 -1386
rect 2766 -1384 2816 -1362
rect 2766 -1404 2816 -1384
rect 4835 -1386 4885 -1364
rect 4835 -1406 4885 -1386
rect 6903 -1384 6953 -1362
rect 6903 -1404 6953 -1384
rect 8972 -1384 9022 -1362
rect 8972 -1404 9022 -1384
rect 11040 -1382 11090 -1360
rect 11040 -1402 11090 -1382
rect 13109 -1384 13159 -1362
rect 13109 -1404 13159 -1384
rect 15177 -1382 15227 -1360
rect 15177 -1402 15227 -1382
<< metal1 >>
rect 740 844 750 866
rect 712 812 750 844
rect 804 844 814 866
rect 2808 846 2818 868
rect 804 812 846 844
rect 712 761 846 812
rect 2780 814 2818 846
rect 2872 846 2882 868
rect 2872 814 2914 846
rect 4877 844 4887 866
rect 2780 763 2914 814
rect 4849 812 4887 844
rect 4941 844 4951 866
rect 6945 846 6955 868
rect 4941 812 4983 844
rect 41 718 1514 761
rect 41 415 75 718
rect 407 613 441 718
rect 643 613 677 718
rect 879 613 913 718
rect 1115 613 1149 718
rect 1480 415 1514 718
rect 2109 720 3582 763
rect 4849 761 4983 812
rect 6917 814 6955 846
rect 7009 846 7019 868
rect 9014 846 9024 868
rect 7009 814 7051 846
rect 6917 763 7051 814
rect 8986 814 9024 846
rect 9078 846 9088 868
rect 11082 848 11092 870
rect 9078 814 9120 846
rect 8986 763 9120 814
rect 11054 816 11092 848
rect 11146 848 11156 870
rect 11146 816 11188 848
rect 13151 846 13161 868
rect 11054 765 11188 816
rect 13123 814 13161 846
rect 13215 846 13225 868
rect 15219 848 15229 870
rect 13215 814 13257 846
rect 2109 417 2143 720
rect 2475 615 2509 720
rect 2711 615 2745 720
rect 2947 615 2981 720
rect 3183 615 3217 720
rect 3548 417 3582 720
rect 4178 718 5651 761
rect 4178 415 4212 718
rect 4544 613 4578 718
rect 4780 613 4814 718
rect 5016 613 5050 718
rect 5252 613 5286 718
rect 5617 415 5651 718
rect 6246 720 7719 763
rect 6246 417 6280 720
rect 6612 615 6646 720
rect 6848 615 6882 720
rect 7084 615 7118 720
rect 7320 615 7354 720
rect 7685 417 7719 720
rect 8315 720 9788 763
rect 8315 417 8349 720
rect 8681 615 8715 720
rect 8917 615 8951 720
rect 9153 615 9187 720
rect 9389 615 9423 720
rect 9754 417 9788 720
rect 10383 722 11856 765
rect 13123 763 13257 814
rect 15191 816 15229 848
rect 15283 848 15293 870
rect 15283 816 15325 848
rect 15191 765 15325 816
rect 10383 419 10417 722
rect 10749 617 10783 722
rect 10985 617 11019 722
rect 11221 617 11255 722
rect 11457 617 11491 722
rect 11822 419 11856 722
rect 12452 720 13925 763
rect 12452 417 12486 720
rect 12818 615 12852 720
rect 13054 615 13088 720
rect 13290 615 13324 720
rect 13526 615 13560 720
rect 13891 417 13925 720
rect 14520 722 15993 765
rect 14520 419 14554 722
rect 14886 617 14920 722
rect 15122 617 15156 722
rect 15358 617 15392 722
rect 15594 617 15628 722
rect 15959 419 15993 722
rect 186 378 193 403
rect 311 378 410 403
rect -77 181 -43 235
rect 304 227 410 378
rect 761 247 795 337
rect 525 235 565 247
rect 637 235 683 247
rect 755 235 795 247
rect 525 181 559 235
rect 761 181 795 235
rect 1143 227 1247 403
rect 2254 380 2261 405
rect 2379 380 2478 405
rect -77 146 82 181
rect 525 146 795 181
rect 1362 181 1396 249
rect 1598 181 1632 249
rect 1362 146 1632 181
rect 1991 183 2025 237
rect 2372 229 2478 380
rect 2829 249 2863 339
rect 2593 237 2633 249
rect 2705 237 2751 249
rect 2823 237 2863 249
rect 2593 183 2627 237
rect 2829 183 2863 237
rect 3211 229 3315 405
rect 4323 378 4330 403
rect 4448 378 4547 403
rect 1991 148 2150 183
rect 2593 148 2863 183
rect 3430 183 3464 251
rect 3666 183 3700 251
rect 3430 148 3700 183
rect 4060 181 4094 235
rect 4441 227 4547 378
rect 4898 247 4932 337
rect 4662 235 4702 247
rect 4774 235 4820 247
rect 4892 235 4932 247
rect 4662 181 4696 235
rect 4898 181 4932 235
rect 5280 227 5384 403
rect 6391 380 6398 405
rect 6516 380 6615 405
rect -132 -2 -58 64
rect 8 -2 18 64
rect -132 -132 8 -126
rect -132 -192 -70 -132
rect -4 -192 8 -132
rect -132 -198 8 -192
rect 48 -638 82 146
rect 761 84 795 146
rect 350 46 1092 84
rect 350 -92 384 46
rect 586 -96 620 46
rect 822 -98 856 46
rect 1058 -98 1092 46
rect 1318 58 1396 64
rect 1318 4 1330 58
rect 1384 4 1396 58
rect 1318 -2 1396 4
rect 350 -393 385 -359
rect 585 -393 620 -359
rect 822 -393 857 -359
rect 1058 -381 1092 -359
rect 1464 -637 1498 146
rect 1936 0 2010 66
rect 2076 0 2086 66
rect 1936 -130 2076 -124
rect 1936 -190 1998 -130
rect 2064 -190 2076 -130
rect 1936 -196 2076 -190
rect 1550 -494 1676 -488
rect 1550 -596 1562 -494
rect 1664 -596 1676 -494
rect 1550 -602 1676 -596
rect 1191 -638 1498 -637
rect 48 -643 364 -638
rect 1078 -643 1498 -638
rect 48 -654 431 -643
rect 48 -681 380 -654
rect 48 -828 82 -681
rect 364 -688 380 -681
rect 414 -688 431 -654
rect 364 -694 431 -688
rect 1011 -654 1498 -643
rect 1011 -688 1028 -654
rect 1062 -681 1498 -654
rect 1062 -688 1078 -681
rect 1191 -682 1498 -681
rect 1011 -694 1078 -688
rect 189 -721 245 -709
rect 189 -755 195 -721
rect 229 -722 245 -721
rect 1302 -722 1358 -710
rect 229 -738 696 -722
rect 229 -755 646 -738
rect 189 -771 646 -755
rect 630 -772 646 -771
rect 680 -772 696 -738
rect 630 -779 696 -772
rect 748 -737 1318 -722
rect 748 -771 764 -737
rect 798 -756 1318 -737
rect 1352 -756 1358 -722
rect 798 -771 1358 -756
rect 748 -781 815 -771
rect 1302 -772 1358 -771
rect 1464 -828 1498 -682
rect 2116 -636 2150 148
rect 2829 86 2863 148
rect 2418 48 3160 86
rect 2418 -90 2452 48
rect 2654 -94 2688 48
rect 2890 -96 2924 48
rect 3126 -96 3160 48
rect 3386 60 3464 66
rect 3386 6 3398 60
rect 3452 6 3464 60
rect 3386 0 3464 6
rect 2418 -391 2453 -357
rect 2653 -391 2688 -357
rect 2890 -391 2925 -357
rect 3126 -379 3160 -357
rect 3532 -635 3566 148
rect 4060 146 4219 181
rect 4662 146 4932 181
rect 5499 181 5533 249
rect 5735 181 5769 249
rect 5499 146 5769 181
rect 6128 183 6162 237
rect 6509 229 6615 380
rect 6966 249 7000 339
rect 6730 237 6770 249
rect 6842 237 6888 249
rect 6960 237 7000 249
rect 6730 183 6764 237
rect 6966 183 7000 237
rect 7348 229 7452 405
rect 8460 380 8467 405
rect 8585 380 8684 405
rect 6128 148 6287 183
rect 6730 148 7000 183
rect 7567 183 7601 251
rect 7803 183 7837 251
rect 7567 148 7837 183
rect 8197 183 8231 237
rect 8578 229 8684 380
rect 9035 249 9069 339
rect 8799 237 8839 249
rect 8911 237 8957 249
rect 9029 237 9069 249
rect 8799 183 8833 237
rect 9035 183 9069 237
rect 9417 229 9521 405
rect 10528 382 10535 407
rect 10653 382 10752 407
rect 8197 148 8356 183
rect 8799 148 9069 183
rect 9636 183 9670 251
rect 9872 183 9906 251
rect 9636 148 9906 183
rect 10265 185 10299 239
rect 10646 231 10752 382
rect 11103 251 11137 341
rect 10867 239 10907 251
rect 10979 239 11025 251
rect 11097 239 11137 251
rect 10867 185 10901 239
rect 11103 185 11137 239
rect 11485 231 11589 407
rect 12597 380 12604 405
rect 12722 380 12821 405
rect 10265 150 10424 185
rect 10867 150 11137 185
rect 11704 185 11738 253
rect 11940 185 11974 253
rect 11704 150 11974 185
rect 12334 183 12368 237
rect 12715 229 12821 380
rect 13172 249 13206 339
rect 12936 237 12976 249
rect 13048 237 13094 249
rect 13166 237 13206 249
rect 12936 183 12970 237
rect 13172 183 13206 237
rect 13554 229 13658 405
rect 14665 382 14672 407
rect 14790 382 14889 407
rect 4005 -2 4079 64
rect 4145 -2 4155 64
rect 4005 -132 4145 -126
rect 4005 -192 4067 -132
rect 4133 -192 4145 -132
rect 4005 -198 4145 -192
rect 3618 -492 3744 -486
rect 3618 -594 3630 -492
rect 3732 -594 3744 -492
rect 3618 -600 3744 -594
rect 3259 -636 3566 -635
rect 2116 -641 2432 -636
rect 3146 -641 3566 -636
rect 2116 -652 2499 -641
rect 2116 -679 2448 -652
rect 2116 -826 2150 -679
rect 2432 -686 2448 -679
rect 2482 -686 2499 -652
rect 2432 -692 2499 -686
rect 3079 -652 3566 -641
rect 3079 -686 3096 -652
rect 3130 -679 3566 -652
rect 3130 -686 3146 -679
rect 3259 -680 3566 -679
rect 3079 -692 3146 -686
rect 2257 -719 2313 -707
rect 2257 -753 2263 -719
rect 2297 -720 2313 -719
rect 3370 -720 3426 -708
rect 2297 -736 2764 -720
rect 2297 -753 2714 -736
rect 2257 -769 2714 -753
rect 2698 -770 2714 -769
rect 2748 -770 2764 -736
rect 2698 -777 2764 -770
rect 2816 -735 3386 -720
rect 2816 -769 2832 -735
rect 2866 -754 3386 -735
rect 3420 -754 3426 -720
rect 2866 -769 3426 -754
rect 2816 -779 2883 -769
rect 3370 -770 3426 -769
rect 3532 -826 3566 -680
rect 4185 -638 4219 146
rect 4898 84 4932 146
rect 4487 46 5229 84
rect 4487 -92 4521 46
rect 4723 -96 4757 46
rect 4959 -98 4993 46
rect 5195 -98 5229 46
rect 5455 58 5533 64
rect 5455 4 5467 58
rect 5521 4 5533 58
rect 5455 -2 5533 4
rect 4487 -393 4522 -359
rect 4722 -393 4757 -359
rect 4959 -393 4994 -359
rect 5195 -381 5229 -359
rect 5601 -637 5635 146
rect 6073 0 6147 66
rect 6213 0 6223 66
rect 6073 -130 6213 -124
rect 6073 -190 6135 -130
rect 6201 -190 6213 -130
rect 6073 -196 6213 -190
rect 5687 -494 5813 -488
rect 5687 -596 5699 -494
rect 5801 -596 5813 -494
rect 5687 -602 5813 -596
rect 5328 -638 5635 -637
rect 4185 -643 4501 -638
rect 5215 -643 5635 -638
rect 4185 -654 4568 -643
rect 4185 -681 4517 -654
rect 4185 -828 4219 -681
rect 4501 -688 4517 -681
rect 4551 -688 4568 -654
rect 4501 -694 4568 -688
rect 5148 -654 5635 -643
rect 5148 -688 5165 -654
rect 5199 -681 5635 -654
rect 5199 -688 5215 -681
rect 5328 -682 5635 -681
rect 5148 -694 5215 -688
rect 4326 -721 4382 -709
rect 4326 -755 4332 -721
rect 4366 -722 4382 -721
rect 5439 -722 5495 -710
rect 4366 -738 4833 -722
rect 4366 -755 4783 -738
rect 4326 -771 4783 -755
rect 4767 -772 4783 -771
rect 4817 -772 4833 -738
rect 4767 -779 4833 -772
rect 4885 -737 5455 -722
rect 4885 -771 4901 -737
rect 4935 -756 5455 -737
rect 5489 -756 5495 -722
rect 4935 -771 5495 -756
rect 4885 -781 4952 -771
rect 5439 -772 5495 -771
rect 5601 -828 5635 -682
rect 6253 -636 6287 148
rect 6966 86 7000 148
rect 6555 48 7297 86
rect 6555 -90 6589 48
rect 6791 -94 6825 48
rect 7027 -96 7061 48
rect 7263 -96 7297 48
rect 7523 60 7601 66
rect 7523 6 7535 60
rect 7589 6 7601 60
rect 7523 0 7601 6
rect 6555 -391 6590 -357
rect 6790 -391 6825 -357
rect 7027 -391 7062 -357
rect 7263 -379 7297 -357
rect 7669 -635 7703 148
rect 8142 0 8216 66
rect 8282 0 8292 66
rect 8142 -130 8282 -124
rect 8142 -190 8204 -130
rect 8270 -190 8282 -130
rect 8142 -196 8282 -190
rect 7755 -492 7881 -486
rect 7755 -594 7767 -492
rect 7869 -594 7881 -492
rect 7755 -600 7881 -594
rect 7396 -636 7703 -635
rect 6253 -641 6569 -636
rect 7283 -641 7703 -636
rect 6253 -652 6636 -641
rect 6253 -679 6585 -652
rect 6253 -826 6287 -679
rect 6569 -686 6585 -679
rect 6619 -686 6636 -652
rect 6569 -692 6636 -686
rect 7216 -652 7703 -641
rect 7216 -686 7233 -652
rect 7267 -679 7703 -652
rect 7267 -686 7283 -679
rect 7396 -680 7703 -679
rect 7216 -692 7283 -686
rect 6394 -719 6450 -707
rect 6394 -753 6400 -719
rect 6434 -720 6450 -719
rect 7507 -720 7563 -708
rect 6434 -736 6901 -720
rect 6434 -753 6851 -736
rect 6394 -769 6851 -753
rect 6835 -770 6851 -769
rect 6885 -770 6901 -736
rect 6835 -777 6901 -770
rect 6953 -735 7523 -720
rect 6953 -769 6969 -735
rect 7003 -754 7523 -735
rect 7557 -754 7563 -720
rect 7003 -769 7563 -754
rect 6953 -779 7020 -769
rect 7507 -770 7563 -769
rect 7669 -826 7703 -680
rect 8322 -636 8356 148
rect 9035 86 9069 148
rect 8624 48 9366 86
rect 8624 -90 8658 48
rect 8860 -94 8894 48
rect 9096 -96 9130 48
rect 9332 -96 9366 48
rect 9592 60 9670 66
rect 9592 6 9604 60
rect 9658 6 9670 60
rect 9592 0 9670 6
rect 8624 -391 8659 -357
rect 8859 -391 8894 -357
rect 9096 -391 9131 -357
rect 9332 -379 9366 -357
rect 9738 -635 9772 148
rect 10210 2 10284 68
rect 10350 2 10360 68
rect 10210 -128 10350 -122
rect 10210 -188 10272 -128
rect 10338 -188 10350 -128
rect 10210 -194 10350 -188
rect 9824 -492 9950 -486
rect 9824 -594 9836 -492
rect 9938 -594 9950 -492
rect 9824 -600 9950 -594
rect 9465 -636 9772 -635
rect 8322 -641 8638 -636
rect 9352 -641 9772 -636
rect 8322 -652 8705 -641
rect 8322 -679 8654 -652
rect 8322 -826 8356 -679
rect 8638 -686 8654 -679
rect 8688 -686 8705 -652
rect 8638 -692 8705 -686
rect 9285 -652 9772 -641
rect 9285 -686 9302 -652
rect 9336 -679 9772 -652
rect 9336 -686 9352 -679
rect 9465 -680 9772 -679
rect 9285 -692 9352 -686
rect 8463 -719 8519 -707
rect 8463 -753 8469 -719
rect 8503 -720 8519 -719
rect 9576 -720 9632 -708
rect 8503 -736 8970 -720
rect 8503 -753 8920 -736
rect 8463 -769 8920 -753
rect 8904 -770 8920 -769
rect 8954 -770 8970 -736
rect 8904 -777 8970 -770
rect 9022 -735 9592 -720
rect 9022 -769 9038 -735
rect 9072 -754 9592 -735
rect 9626 -754 9632 -720
rect 9072 -769 9632 -754
rect 9022 -779 9089 -769
rect 9576 -770 9632 -769
rect 9738 -826 9772 -680
rect 10390 -634 10424 150
rect 11103 88 11137 150
rect 10692 50 11434 88
rect 10692 -88 10726 50
rect 10928 -92 10962 50
rect 11164 -94 11198 50
rect 11400 -94 11434 50
rect 11660 62 11738 68
rect 11660 8 11672 62
rect 11726 8 11738 62
rect 11660 2 11738 8
rect 10692 -389 10727 -355
rect 10927 -389 10962 -355
rect 11164 -389 11199 -355
rect 11400 -377 11434 -355
rect 11806 -633 11840 150
rect 12334 148 12493 183
rect 12936 148 13206 183
rect 13773 183 13807 251
rect 14009 183 14043 251
rect 13773 148 14043 183
rect 14402 185 14436 239
rect 14783 231 14889 382
rect 15240 251 15274 341
rect 15004 239 15044 251
rect 15116 239 15162 251
rect 15234 239 15274 251
rect 15004 185 15038 239
rect 15240 185 15274 239
rect 15622 231 15726 407
rect 14402 150 14561 185
rect 15004 150 15274 185
rect 15841 185 15875 253
rect 16077 185 16111 253
rect 15841 150 16111 185
rect 12279 0 12353 66
rect 12419 0 12429 66
rect 12279 -130 12419 -124
rect 12279 -190 12341 -130
rect 12407 -190 12419 -130
rect 12279 -196 12419 -190
rect 11892 -490 12018 -484
rect 11892 -592 11904 -490
rect 12006 -592 12018 -490
rect 11892 -598 12018 -592
rect 11533 -634 11840 -633
rect 10390 -639 10706 -634
rect 11420 -639 11840 -634
rect 10390 -650 10773 -639
rect 10390 -677 10722 -650
rect 10390 -824 10424 -677
rect 10706 -684 10722 -677
rect 10756 -684 10773 -650
rect 10706 -690 10773 -684
rect 11353 -650 11840 -639
rect 11353 -684 11370 -650
rect 11404 -677 11840 -650
rect 11404 -684 11420 -677
rect 11533 -678 11840 -677
rect 11353 -690 11420 -684
rect 10531 -717 10587 -705
rect 10531 -751 10537 -717
rect 10571 -718 10587 -717
rect 11644 -718 11700 -706
rect 10571 -734 11038 -718
rect 10571 -751 10988 -734
rect 10531 -767 10988 -751
rect 10972 -768 10988 -767
rect 11022 -768 11038 -734
rect 10972 -775 11038 -768
rect 11090 -733 11660 -718
rect 11090 -767 11106 -733
rect 11140 -752 11660 -733
rect 11694 -752 11700 -718
rect 11140 -767 11700 -752
rect 11090 -777 11157 -767
rect 11644 -768 11700 -767
rect 11806 -824 11840 -678
rect 12459 -636 12493 148
rect 13172 86 13206 148
rect 12761 48 13503 86
rect 12761 -90 12795 48
rect 12997 -94 13031 48
rect 13233 -96 13267 48
rect 13469 -96 13503 48
rect 13729 60 13807 66
rect 13729 6 13741 60
rect 13795 6 13807 60
rect 13729 0 13807 6
rect 12761 -391 12796 -357
rect 12996 -391 13031 -357
rect 13233 -391 13268 -357
rect 13469 -379 13503 -357
rect 13875 -635 13909 148
rect 14347 2 14421 68
rect 14487 2 14497 68
rect 14347 -128 14487 -122
rect 14347 -188 14409 -128
rect 14475 -188 14487 -128
rect 14347 -194 14487 -188
rect 13961 -492 14087 -486
rect 13961 -594 13973 -492
rect 14075 -594 14087 -492
rect 13961 -600 14087 -594
rect 13602 -636 13909 -635
rect 12459 -641 12775 -636
rect 13489 -641 13909 -636
rect 12459 -652 12842 -641
rect 12459 -679 12791 -652
rect 12459 -826 12493 -679
rect 12775 -686 12791 -679
rect 12825 -686 12842 -652
rect 12775 -692 12842 -686
rect 13422 -652 13909 -641
rect 13422 -686 13439 -652
rect 13473 -679 13909 -652
rect 13473 -686 13489 -679
rect 13602 -680 13909 -679
rect 13422 -692 13489 -686
rect 12600 -719 12656 -707
rect 12600 -753 12606 -719
rect 12640 -720 12656 -719
rect 13713 -720 13769 -708
rect 12640 -736 13107 -720
rect 12640 -753 13057 -736
rect 12600 -769 13057 -753
rect 13041 -770 13057 -769
rect 13091 -770 13107 -736
rect 13041 -777 13107 -770
rect 13159 -735 13729 -720
rect 13159 -769 13175 -735
rect 13209 -754 13729 -735
rect 13763 -754 13769 -720
rect 13209 -769 13769 -754
rect 13159 -779 13226 -769
rect 13713 -770 13769 -769
rect 13875 -826 13909 -680
rect 14527 -634 14561 150
rect 15240 88 15274 150
rect 14829 50 15571 88
rect 14829 -88 14863 50
rect 15065 -92 15099 50
rect 15301 -94 15335 50
rect 15537 -94 15571 50
rect 15797 62 15875 68
rect 15797 8 15809 62
rect 15863 8 15875 62
rect 15797 2 15875 8
rect 14829 -389 14864 -355
rect 15064 -389 15099 -355
rect 15301 -389 15336 -355
rect 15537 -377 15571 -355
rect 15943 -633 15977 150
rect 16029 -490 16155 -484
rect 16029 -592 16041 -490
rect 16143 -592 16155 -490
rect 16029 -598 16155 -592
rect 15670 -634 15977 -633
rect 14527 -639 14843 -634
rect 15557 -639 15977 -634
rect 14527 -650 14910 -639
rect 14527 -677 14859 -650
rect 14527 -824 14561 -677
rect 14843 -684 14859 -677
rect 14893 -684 14910 -650
rect 14843 -690 14910 -684
rect 15490 -650 15977 -639
rect 15490 -684 15507 -650
rect 15541 -677 15977 -650
rect 15541 -684 15557 -677
rect 15670 -678 15977 -677
rect 15490 -690 15557 -684
rect 14668 -717 14724 -705
rect 14668 -751 14674 -717
rect 14708 -718 14724 -717
rect 15781 -718 15837 -706
rect 14708 -734 15175 -718
rect 14708 -751 15125 -734
rect 14668 -767 15125 -751
rect 15109 -768 15125 -767
rect 15159 -768 15175 -734
rect 15109 -775 15175 -768
rect 15227 -733 15797 -718
rect 15227 -767 15243 -733
rect 15277 -752 15797 -733
rect 15831 -752 15837 -718
rect 15277 -767 15837 -752
rect 15227 -777 15294 -767
rect 15781 -768 15837 -767
rect 15943 -824 15977 -678
rect 165 -1304 199 -995
rect 822 -1304 856 -1198
rect 1346 -1304 1379 -982
rect 165 -1336 1379 -1304
rect 2233 -1302 2267 -993
rect 2890 -1302 2924 -1196
rect 3414 -1302 3447 -980
rect 2233 -1334 3447 -1302
rect 4302 -1304 4336 -995
rect 4959 -1304 4993 -1198
rect 5483 -1304 5516 -982
rect 658 -1358 790 -1336
rect 658 -1416 692 -1358
rect 754 -1416 790 -1358
rect 658 -1421 790 -1416
rect 2726 -1356 2858 -1334
rect 4302 -1336 5516 -1304
rect 6370 -1302 6404 -993
rect 7027 -1302 7061 -1196
rect 7551 -1302 7584 -980
rect 6370 -1334 7584 -1302
rect 8439 -1302 8473 -993
rect 9096 -1302 9130 -1196
rect 9620 -1302 9653 -980
rect 8439 -1334 9653 -1302
rect 10507 -1300 10541 -991
rect 11164 -1300 11198 -1194
rect 11688 -1300 11721 -978
rect 10507 -1332 11721 -1300
rect 12576 -1302 12610 -993
rect 13233 -1302 13267 -1196
rect 13757 -1302 13790 -980
rect 2726 -1414 2760 -1356
rect 2822 -1414 2858 -1356
rect 2726 -1419 2858 -1414
rect 4795 -1358 4927 -1336
rect 4795 -1416 4829 -1358
rect 4891 -1416 4927 -1358
rect 4795 -1421 4927 -1416
rect 6863 -1356 6995 -1334
rect 6863 -1414 6897 -1356
rect 6959 -1414 6995 -1356
rect 6863 -1419 6995 -1414
rect 8932 -1356 9064 -1334
rect 8932 -1414 8966 -1356
rect 9028 -1414 9064 -1356
rect 8932 -1419 9064 -1414
rect 11000 -1354 11132 -1332
rect 12576 -1334 13790 -1302
rect 14644 -1300 14678 -991
rect 15301 -1300 15335 -1194
rect 15825 -1300 15858 -978
rect 14644 -1332 15858 -1300
rect 11000 -1412 11034 -1354
rect 11096 -1412 11132 -1354
rect 11000 -1417 11132 -1412
rect 13069 -1356 13201 -1334
rect 13069 -1414 13103 -1356
rect 13165 -1414 13201 -1356
rect 13069 -1419 13201 -1414
rect 15137 -1354 15269 -1332
rect 15137 -1412 15171 -1354
rect 15233 -1412 15269 -1354
rect 15137 -1417 15269 -1412
<< via1 >>
rect 750 858 804 866
rect 750 820 760 858
rect 760 820 798 858
rect 798 820 804 858
rect 2818 860 2872 868
rect 750 812 804 820
rect 2818 822 2828 860
rect 2828 822 2866 860
rect 2866 822 2872 860
rect 2818 814 2872 822
rect 4887 858 4941 866
rect 4887 820 4897 858
rect 4897 820 4935 858
rect 4935 820 4941 858
rect 6955 860 7009 868
rect 4887 812 4941 820
rect 6955 822 6965 860
rect 6965 822 7003 860
rect 7003 822 7009 860
rect 9024 860 9078 868
rect 6955 814 7009 822
rect 9024 822 9034 860
rect 9034 822 9072 860
rect 9072 822 9078 860
rect 11092 862 11146 870
rect 9024 814 9078 822
rect 11092 824 11102 862
rect 11102 824 11140 862
rect 11140 824 11146 862
rect 11092 816 11146 824
rect 13161 860 13215 868
rect 13161 822 13171 860
rect 13171 822 13209 860
rect 13209 822 13215 860
rect 15229 862 15283 870
rect 13161 814 13215 822
rect 15229 824 15239 862
rect 15239 824 15277 862
rect 15277 824 15283 862
rect 15229 816 15283 824
rect -58 -2 8 64
rect 1330 4 1384 58
rect 2010 0 2076 66
rect 3398 6 3452 60
rect 4079 -2 4145 64
rect 5467 4 5521 58
rect 6147 0 6213 66
rect 7535 6 7589 60
rect 8216 0 8282 66
rect 9604 6 9658 60
rect 10284 2 10350 68
rect 11672 8 11726 62
rect 12353 0 12419 66
rect 13741 6 13795 60
rect 14421 2 14487 68
rect 15809 8 15863 62
rect 692 -1364 754 -1358
rect 692 -1406 698 -1364
rect 698 -1406 748 -1364
rect 748 -1406 754 -1364
rect 692 -1416 754 -1406
rect 2760 -1362 2822 -1356
rect 2760 -1404 2766 -1362
rect 2766 -1404 2816 -1362
rect 2816 -1404 2822 -1362
rect 2760 -1414 2822 -1404
rect 4829 -1364 4891 -1358
rect 4829 -1406 4835 -1364
rect 4835 -1406 4885 -1364
rect 4885 -1406 4891 -1364
rect 4829 -1416 4891 -1406
rect 6897 -1362 6959 -1356
rect 6897 -1404 6903 -1362
rect 6903 -1404 6953 -1362
rect 6953 -1404 6959 -1362
rect 6897 -1414 6959 -1404
rect 8966 -1362 9028 -1356
rect 8966 -1404 8972 -1362
rect 8972 -1404 9022 -1362
rect 9022 -1404 9028 -1362
rect 8966 -1414 9028 -1404
rect 11034 -1360 11096 -1354
rect 11034 -1402 11040 -1360
rect 11040 -1402 11090 -1360
rect 11090 -1402 11096 -1360
rect 11034 -1412 11096 -1402
rect 13103 -1362 13165 -1356
rect 13103 -1404 13109 -1362
rect 13109 -1404 13159 -1362
rect 13159 -1404 13165 -1362
rect 13103 -1414 13165 -1404
rect 15171 -1360 15233 -1354
rect 15171 -1402 15177 -1360
rect 15177 -1402 15227 -1360
rect 15227 -1402 15233 -1360
rect 15171 -1412 15233 -1402
<< metal2 >>
rect 738 874 816 884
rect 738 794 816 804
rect 2806 876 2884 886
rect 2806 796 2884 806
rect 4875 874 4953 884
rect 4875 794 4953 804
rect 6943 876 7021 886
rect 6943 796 7021 806
rect 9012 876 9090 886
rect 9012 796 9090 806
rect 11080 878 11158 888
rect 11080 798 11158 808
rect 13149 876 13227 886
rect 13149 796 13227 806
rect 15217 878 15295 888
rect 15217 798 15295 808
rect -64 -2 -58 64
rect 8 58 1384 64
rect 8 4 1330 58
rect 8 -2 1384 4
rect 2004 0 2010 66
rect 2076 60 3452 66
rect 2076 6 3398 60
rect 2076 0 3452 6
rect 4073 -2 4079 64
rect 4145 58 5521 64
rect 4145 4 5467 58
rect 4145 -2 5521 4
rect 6141 0 6147 66
rect 6213 60 7589 66
rect 6213 6 7535 60
rect 6213 0 7589 6
rect 8210 0 8216 66
rect 8282 60 9658 66
rect 8282 6 9604 60
rect 8282 0 9658 6
rect 10278 2 10284 68
rect 10350 62 11726 68
rect 10350 8 11672 62
rect 10350 2 11726 8
rect 12347 0 12353 66
rect 12419 60 13795 66
rect 12419 6 13741 60
rect 12419 0 13795 6
rect 14415 2 14421 68
rect 14487 62 15863 68
rect 14487 8 15809 62
rect 14487 2 15863 8
rect 686 -1356 758 -1346
rect 686 -1436 758 -1426
rect 2754 -1354 2826 -1344
rect 2754 -1434 2826 -1424
rect 4823 -1356 4895 -1346
rect 4823 -1436 4895 -1426
rect 6891 -1354 6963 -1344
rect 6891 -1434 6963 -1424
rect 8960 -1354 9032 -1344
rect 8960 -1434 9032 -1424
rect 11028 -1352 11100 -1342
rect 11028 -1432 11100 -1422
rect 13097 -1354 13169 -1344
rect 13097 -1434 13169 -1424
rect 15165 -1352 15237 -1342
rect 15165 -1432 15237 -1422
<< via2 >>
rect 738 866 816 874
rect 738 812 750 866
rect 750 812 804 866
rect 804 812 816 866
rect 738 804 816 812
rect 2806 868 2884 876
rect 2806 814 2818 868
rect 2818 814 2872 868
rect 2872 814 2884 868
rect 2806 806 2884 814
rect 4875 866 4953 874
rect 4875 812 4887 866
rect 4887 812 4941 866
rect 4941 812 4953 866
rect 4875 804 4953 812
rect 6943 868 7021 876
rect 6943 814 6955 868
rect 6955 814 7009 868
rect 7009 814 7021 868
rect 6943 806 7021 814
rect 9012 868 9090 876
rect 9012 814 9024 868
rect 9024 814 9078 868
rect 9078 814 9090 868
rect 9012 806 9090 814
rect 11080 870 11158 878
rect 11080 816 11092 870
rect 11092 816 11146 870
rect 11146 816 11158 870
rect 11080 808 11158 816
rect 13149 868 13227 876
rect 13149 814 13161 868
rect 13161 814 13215 868
rect 13215 814 13227 868
rect 13149 806 13227 814
rect 15217 870 15295 878
rect 15217 816 15229 870
rect 15229 816 15283 870
rect 15283 816 15295 870
rect 15217 808 15295 816
rect 686 -1358 758 -1356
rect 686 -1416 692 -1358
rect 692 -1416 754 -1358
rect 754 -1416 758 -1358
rect 686 -1426 758 -1416
rect 2754 -1356 2826 -1354
rect 2754 -1414 2760 -1356
rect 2760 -1414 2822 -1356
rect 2822 -1414 2826 -1356
rect 2754 -1424 2826 -1414
rect 4823 -1358 4895 -1356
rect 4823 -1416 4829 -1358
rect 4829 -1416 4891 -1358
rect 4891 -1416 4895 -1358
rect 4823 -1426 4895 -1416
rect 6891 -1356 6963 -1354
rect 6891 -1414 6897 -1356
rect 6897 -1414 6959 -1356
rect 6959 -1414 6963 -1356
rect 6891 -1424 6963 -1414
rect 8960 -1356 9032 -1354
rect 8960 -1414 8966 -1356
rect 8966 -1414 9028 -1356
rect 9028 -1414 9032 -1356
rect 8960 -1424 9032 -1414
rect 11028 -1354 11100 -1352
rect 11028 -1412 11034 -1354
rect 11034 -1412 11096 -1354
rect 11096 -1412 11100 -1354
rect 11028 -1422 11100 -1412
rect 13097 -1356 13169 -1354
rect 13097 -1414 13103 -1356
rect 13103 -1414 13165 -1356
rect 13165 -1414 13169 -1356
rect 13097 -1424 13169 -1414
rect 15165 -1354 15237 -1352
rect 15165 -1412 15171 -1354
rect 15171 -1412 15233 -1354
rect 15233 -1412 15237 -1354
rect 15165 -1422 15237 -1412
<< metal3 >>
rect 668 876 882 880
rect 668 804 738 876
rect 814 874 882 876
rect 816 804 882 874
rect 2736 878 2950 882
rect 2736 806 2806 878
rect 2882 876 2950 878
rect 2884 806 2950 876
rect 2736 804 2950 806
rect 4805 876 5019 880
rect 4805 804 4875 876
rect 4951 874 5019 876
rect 4953 804 5019 874
rect 6873 878 7087 882
rect 6873 806 6943 878
rect 7019 876 7087 878
rect 7021 806 7087 876
rect 6873 804 7087 806
rect 8942 878 9156 882
rect 8942 806 9012 878
rect 9088 876 9156 878
rect 9090 806 9156 876
rect 11010 880 11224 884
rect 11010 808 11080 880
rect 11156 878 11224 880
rect 11158 808 11224 878
rect 11010 806 11224 808
rect 13079 878 13293 882
rect 13079 806 13149 878
rect 13225 876 13293 878
rect 13227 806 13293 876
rect 15147 880 15361 884
rect 15147 808 15217 880
rect 15293 878 15361 880
rect 15295 808 15361 878
rect 15147 806 15361 808
rect 8942 804 9156 806
rect 668 802 882 804
rect 728 799 826 802
rect 2796 801 2894 804
rect 4805 802 5019 804
rect 4865 799 4963 802
rect 6933 801 7031 804
rect 9002 801 9100 804
rect 11070 803 11168 806
rect 13079 804 13293 806
rect 13139 801 13237 804
rect 15207 803 15305 806
rect 10990 -1338 11142 -1336
rect 15127 -1338 15279 -1336
rect 2716 -1340 2868 -1338
rect 6853 -1340 7005 -1338
rect 8922 -1340 9074 -1338
rect 648 -1342 800 -1340
rect 646 -1346 800 -1342
rect 646 -1434 676 -1346
rect 770 -1434 800 -1346
rect 646 -1440 800 -1434
rect 2714 -1344 2868 -1340
rect 4785 -1342 4937 -1340
rect 2714 -1432 2744 -1344
rect 2838 -1432 2868 -1344
rect 2714 -1438 2868 -1432
rect 648 -1450 800 -1440
rect 2716 -1448 2868 -1438
rect 4783 -1346 4937 -1342
rect 4783 -1434 4813 -1346
rect 4907 -1434 4937 -1346
rect 4783 -1440 4937 -1434
rect 6851 -1344 7005 -1340
rect 6851 -1432 6881 -1344
rect 6975 -1432 7005 -1344
rect 6851 -1438 7005 -1432
rect 8920 -1344 9074 -1340
rect 8920 -1432 8950 -1344
rect 9044 -1432 9074 -1344
rect 8920 -1438 9074 -1432
rect 10988 -1342 11142 -1338
rect 13059 -1340 13211 -1338
rect 10988 -1430 11018 -1342
rect 11112 -1430 11142 -1342
rect 10988 -1436 11142 -1430
rect 4785 -1450 4937 -1440
rect 6853 -1448 7005 -1438
rect 8922 -1448 9074 -1438
rect 10990 -1446 11142 -1436
rect 13057 -1344 13211 -1340
rect 13057 -1432 13087 -1344
rect 13181 -1432 13211 -1344
rect 13057 -1438 13211 -1432
rect 15125 -1342 15279 -1338
rect 15125 -1430 15155 -1342
rect 15249 -1430 15279 -1342
rect 15125 -1436 15279 -1430
rect 13059 -1448 13211 -1438
rect 15127 -1446 15279 -1436
<< via3 >>
rect 738 874 814 876
rect 738 810 814 874
rect 2806 876 2882 878
rect 2806 812 2882 876
rect 4875 874 4951 876
rect 4875 810 4951 874
rect 6943 876 7019 878
rect 6943 812 7019 876
rect 9012 876 9088 878
rect 9012 812 9088 876
rect 11080 878 11156 880
rect 11080 814 11156 878
rect 13149 876 13225 878
rect 13149 812 13225 876
rect 15217 878 15293 880
rect 15217 814 15293 878
rect 676 -1356 770 -1346
rect 676 -1426 686 -1356
rect 686 -1426 758 -1356
rect 758 -1426 770 -1356
rect 676 -1434 770 -1426
rect 2744 -1354 2838 -1344
rect 2744 -1424 2754 -1354
rect 2754 -1424 2826 -1354
rect 2826 -1424 2838 -1354
rect 2744 -1432 2838 -1424
rect 4813 -1356 4907 -1346
rect 4813 -1426 4823 -1356
rect 4823 -1426 4895 -1356
rect 4895 -1426 4907 -1356
rect 4813 -1434 4907 -1426
rect 6881 -1354 6975 -1344
rect 6881 -1424 6891 -1354
rect 6891 -1424 6963 -1354
rect 6963 -1424 6975 -1354
rect 6881 -1432 6975 -1424
rect 8950 -1354 9044 -1344
rect 8950 -1424 8960 -1354
rect 8960 -1424 9032 -1354
rect 9032 -1424 9044 -1354
rect 8950 -1432 9044 -1424
rect 11018 -1352 11112 -1342
rect 11018 -1422 11028 -1352
rect 11028 -1422 11100 -1352
rect 11100 -1422 11112 -1352
rect 11018 -1430 11112 -1422
rect 13087 -1354 13181 -1344
rect 13087 -1424 13097 -1354
rect 13097 -1424 13169 -1354
rect 13169 -1424 13181 -1354
rect 13087 -1432 13181 -1424
rect 15155 -1352 15249 -1342
rect 15155 -1422 15165 -1352
rect 15165 -1422 15237 -1352
rect 15237 -1422 15249 -1352
rect 15155 -1430 15249 -1422
<< metal4 >>
rect -106 880 16132 1012
rect -106 878 11080 880
rect -106 876 2806 878
rect -106 810 738 876
rect 814 812 2806 876
rect 2882 876 6943 878
rect 2882 812 4875 876
rect 814 810 4875 812
rect 4951 812 6943 876
rect 7019 812 9012 878
rect 9088 814 11080 878
rect 11156 878 15217 880
rect 11156 814 13149 878
rect 9088 812 13149 814
rect 13225 814 15217 878
rect 15293 814 16132 880
rect 13225 812 16132 814
rect 4951 810 16132 812
rect -106 768 16132 810
rect 2118 -1340 3482 -1338
rect 6255 -1340 7619 -1338
rect 8324 -1340 9688 -1338
rect 10392 -1340 11756 -1336
rect 12461 -1340 13825 -1338
rect 14529 -1340 16080 -1336
rect -10 -1342 16080 -1340
rect -10 -1344 11018 -1342
rect -10 -1346 2744 -1344
rect -10 -1434 676 -1346
rect 770 -1432 2744 -1346
rect 2838 -1346 6881 -1344
rect 2838 -1432 4813 -1346
rect 770 -1434 4813 -1432
rect 4907 -1432 6881 -1346
rect 6975 -1432 8950 -1344
rect 9044 -1430 11018 -1344
rect 11112 -1344 15155 -1342
rect 11112 -1430 13087 -1344
rect 9044 -1432 13087 -1430
rect 13181 -1430 15155 -1344
rect 15249 -1430 16080 -1342
rect 13181 -1432 16080 -1430
rect 4907 -1434 16080 -1432
rect -10 -1530 16080 -1434
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_0
timestamp 1736499154
transform 1 0 2789 0 1 -1008
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_1
timestamp 1736499154
transform 1 0 721 0 1 -1010
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_2
timestamp 1736499154
transform 1 0 6926 0 1 -1008
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_3
timestamp 1736499154
transform 1 0 4858 0 1 -1010
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_4
timestamp 1736499154
transform 1 0 15200 0 1 -1006
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_5
timestamp 1736499154
transform 1 0 13132 0 1 -1008
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_6
timestamp 1736499154
transform 1 0 11063 0 1 -1006
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ALVBQN  sky130_fd_pr__nfet_01v8_ALVBQN_7
timestamp 1736499154
transform 1 0 8995 0 1 -1008
box -265 -226 265 226
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_0
timestamp 1736499154
transform 1 0 3490 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_1
timestamp 1736499154
transform 1 0 2192 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_2
timestamp 1736499154
transform 1 0 124 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_3
timestamp 1736499154
transform 1 0 1422 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_4
timestamp 1736499154
transform 1 0 7627 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_5
timestamp 1736499154
transform 1 0 6329 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_6
timestamp 1736499154
transform 1 0 5559 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_7
timestamp 1736499154
transform 1 0 4261 0 1 -910
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_8
timestamp 1736499154
transform 1 0 15901 0 1 -906
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_9
timestamp 1736499154
transform 1 0 14603 0 1 -906
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_10
timestamp 1736499154
transform 1 0 13833 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_11
timestamp 1736499154
transform 1 0 12535 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_12
timestamp 1736499154
transform 1 0 11764 0 1 -906
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_13
timestamp 1736499154
transform 1 0 10466 0 1 -906
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_14
timestamp 1736499154
transform 1 0 9696 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__nfet_01v8_ZGVMSF  sky130_fd_pr__nfet_01v8_ZGVMSF_15
timestamp 1736499154
transform 1 0 8398 0 1 -908
box -88 -126 88 126
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_0
timestamp 1736499154
transform 1 0 2789 0 1 -276
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_1
timestamp 1736499154
transform 1 0 2846 0 1 417
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_2
timestamp 1736499154
transform 1 0 778 0 1 415
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_3
timestamp 1736499154
transform 1 0 721 0 1 -278
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_4
timestamp 1736499154
transform 1 0 6983 0 1 417
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_5
timestamp 1736499154
transform 1 0 4915 0 1 415
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_6
timestamp 1736499154
transform 1 0 6926 0 1 -276
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_7
timestamp 1736499154
transform 1 0 4858 0 1 -278
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_8
timestamp 1736499154
transform 1 0 15257 0 1 419
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_9
timestamp 1736499154
transform 1 0 13189 0 1 417
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_10
timestamp 1736499154
transform 1 0 11120 0 1 419
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_11
timestamp 1736499154
transform 1 0 9052 0 1 417
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_12
timestamp 1736499154
transform 1 0 15200 0 1 -274
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_13
timestamp 1736499154
transform 1 0 13132 0 1 -276
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_14
timestamp 1736499154
transform 1 0 11063 0 1 -274
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_6C4S85  sky130_fd_pr__pfet_01v8_6C4S85_15
timestamp 1736499154
transform 1 0 8995 0 1 -276
box -419 -262 419 262
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_0
timestamp 1736499154
transform 1 0 3506 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_1
timestamp 1736499154
transform 1 0 2185 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_2
timestamp 1736499154
transform 1 0 117 0 1 315
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_3
timestamp 1736499154
transform 1 0 1438 0 1 315
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_4
timestamp 1736499154
transform 1 0 7643 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_5
timestamp 1736499154
transform 1 0 6322 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_6
timestamp 1736499154
transform 1 0 5575 0 1 315
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_7
timestamp 1736499154
transform 1 0 4254 0 1 315
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_8
timestamp 1736499154
transform 1 0 15917 0 1 319
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_9
timestamp 1736499154
transform 1 0 14596 0 1 319
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_10
timestamp 1736499154
transform 1 0 13849 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_11
timestamp 1736499154
transform 1 0 12528 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_12
timestamp 1736499154
transform 1 0 11780 0 1 319
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_13
timestamp 1736499154
transform 1 0 10459 0 1 319
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_14
timestamp 1736499154
transform 1 0 9712 0 1 317
box -242 -162 242 162
use sky130_fd_pr__pfet_01v8_A6QCZ3  sky130_fd_pr__pfet_01v8_A6QCZ3_15
timestamp 1736499154
transform 1 0 8391 0 1 317
box -242 -162 242 162
<< labels >>
flabel metal4 7782 -1524 8178 -1430 1 FreeSerif 1120 0 0 0 VSS
port 1 n
flabel metal4 7782 776 8182 898 1 FreeSerif 1120 0 0 0 VDD
port 2 n
flabel metal1 -132 -196 -92 -146 1 FreeSerif 480 0 0 0 A[0]
port 3 n
flabel metal1 1938 -192 1978 -142 1 FreeSerif 480 0 0 0 A[1]
port 4 n
flabel metal1 4008 -194 4048 -144 1 FreeSerif 480 0 0 0 A[2]
port 5 n
flabel metal1 6074 -194 6114 -144 1 FreeSerif 480 0 0 0 A[3]
port 6 n
flabel metal1 8144 -194 8184 -144 1 FreeSerif 480 0 0 0 A[4]
port 7 n
flabel metal1 10212 -192 10252 -142 1 FreeSerif 480 0 0 0 A[5]
port 8 n
flabel metal1 12280 -194 12320 -144 1 FreeSerif 480 0 0 0 A[6]
port 9 n
flabel metal1 14348 -194 14388 -144 1 FreeSerif 480 0 0 0 A[7]
port 10 n
flabel metal1 -130 0 -90 50 1 FreeSerif 480 0 0 0 B[0]
port 11 n
flabel metal1 1938 2 1978 52 1 FreeSerif 480 0 0 0 B[1]
port 12 n
flabel metal1 4008 0 4048 50 1 FreeSerif 480 0 0 0 B[2]
port 13 n
flabel metal1 6074 2 6114 52 1 FreeSerif 480 0 0 0 B[3]
port 14 n
flabel metal1 8144 2 8184 52 1 FreeSerif 480 0 0 0 B[4]
port 15 n
flabel metal1 10212 2 10252 52 1 FreeSerif 480 0 0 0 B[5]
port 16 n
flabel metal1 12280 2 12320 52 1 FreeSerif 480 0 0 0 B[6]
port 17 n
flabel metal1 14350 4 14390 54 1 FreeSerif 480 0 0 0 B[7]
port 18 n
flabel metal1 1570 -570 1676 -510 1 FreeSerif 560 0 0 0 Y[0]
port 19 n
flabel metal1 3632 -568 3738 -508 1 FreeSerif 560 0 0 0 Y[1]
port 20 n
flabel metal1 5702 -568 5808 -508 1 FreeSerif 560 0 0 0 Y[2]
port 21 n
flabel metal1 7762 -572 7868 -512 1 FreeSerif 560 0 0 0 Y[3]
port 22 n
flabel metal1 9844 -564 9950 -504 1 FreeSerif 560 0 0 0 Y[4]
port 23 n
flabel metal1 11910 -562 12016 -502 1 FreeSerif 560 0 0 0 Y[5]
port 24 n
flabel metal1 13978 -568 14084 -508 1 FreeSerif 560 0 0 0 Y[6]
port 25 n
flabel metal1 16044 -562 16150 -502 1 FreeSerif 560 0 0 0 Y[7]
port 26 n
<< end >>
