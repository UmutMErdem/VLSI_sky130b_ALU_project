magic
tech sky130B
magscale 1 2
timestamp 1736766762
<< nwell >>
rect 152 3959 1344 4205
rect 1600 3959 2792 4205
rect 3098 3961 4290 4207
rect 4546 3961 5738 4207
rect 152 3947 1345 3959
rect 1600 3947 2793 3959
rect 3098 3949 4291 3961
rect 4546 3949 5739 3961
rect 153 3635 1345 3947
rect 1601 3635 2793 3947
rect 3099 3637 4291 3949
rect 4547 3637 5739 3949
rect 6066 3959 7258 4205
rect 7514 3959 8706 4205
rect 9012 3961 10204 4207
rect 10460 3961 11652 4207
rect 6066 3947 7259 3959
rect 7514 3947 8707 3959
rect 9012 3949 10205 3961
rect 10460 3949 11653 3961
rect 6067 3635 7259 3947
rect 7515 3635 8707 3947
rect 9013 3637 10205 3949
rect 10461 3637 11653 3949
rect 11916 3632 12830 4410
rect 13084 3632 13998 4410
rect 12346 3042 12830 3632
rect 13514 3372 13998 3632
rect 14252 3630 15166 4410
rect 15420 3632 16334 4410
rect 16594 3634 17508 4412
rect 14682 3372 15166 3630
rect 13513 3324 13998 3372
rect 14681 3324 15166 3372
rect 13513 3048 13997 3324
rect 14681 3048 15165 3324
rect 15850 3048 16334 3632
rect 17024 3368 17508 3634
rect 17762 3632 18676 4412
rect 18930 3634 19844 4412
rect 17022 3326 17508 3368
rect 18192 3367 18676 3632
rect 19360 3367 19844 3634
rect 20098 3632 21012 4412
rect 20528 3368 21012 3632
rect 18191 3326 18676 3367
rect 19359 3326 19844 3367
rect 20527 3326 21012 3368
rect 17022 3044 17506 3326
rect 18191 3043 18675 3326
rect 19359 3043 19843 3326
rect 20527 3044 21011 3326
rect 653 2202 2430 2492
rect 3797 2202 5574 2492
rect 6929 2206 8706 2496
rect 10073 2206 11850 2496
rect 653 2002 2431 2202
rect 3797 2002 5575 2202
rect 6929 2006 8707 2206
rect 10073 2006 11851 2206
rect 13275 2202 15052 2492
rect 16419 2202 18196 2492
rect 19551 2206 21328 2496
rect 22695 2206 24472 2496
rect 212 1678 2904 2002
rect 3356 1678 6048 2002
rect 6488 1682 9180 2006
rect 9632 1682 12324 2006
rect 13275 2002 15053 2202
rect 16419 2002 18197 2202
rect 19551 2006 21329 2206
rect 22695 2006 24473 2206
rect 12834 1678 15526 2002
rect 15978 1678 18670 2002
rect 19110 1682 21802 2006
rect 22254 1682 24946 2006
rect 653 -532 2430 -242
rect 3797 -532 5574 -242
rect 6929 -528 8706 -238
rect 10073 -528 11850 -238
rect 653 -732 2431 -532
rect 3797 -732 5575 -532
rect 6929 -728 8707 -528
rect 10073 -728 11851 -528
rect 13275 -532 15052 -242
rect 16419 -532 18196 -242
rect 19551 -528 21328 -238
rect 22695 -528 24472 -238
rect 212 -1056 2904 -732
rect 3356 -1056 6048 -732
rect 6488 -1052 9180 -728
rect 9632 -1052 12324 -728
rect 13275 -732 15053 -532
rect 16419 -732 18197 -532
rect 19551 -728 21329 -528
rect 22695 -728 24473 -528
rect 12834 -1056 15526 -732
rect 15978 -1056 18670 -732
rect 19110 -1052 21802 -728
rect 22254 -1052 24946 -728
rect 643 -3264 2420 -2974
rect 3787 -3264 5564 -2974
rect 6919 -3260 8696 -2970
rect 10063 -3260 11840 -2970
rect 643 -3464 2421 -3264
rect 3787 -3464 5565 -3264
rect 6919 -3460 8697 -3260
rect 10063 -3460 11841 -3260
rect 13265 -3264 15042 -2974
rect 16409 -3264 18186 -2974
rect 19541 -3260 21318 -2970
rect 22685 -3260 24462 -2970
rect 202 -3788 2894 -3464
rect 3346 -3788 6038 -3464
rect 6478 -3784 9170 -3460
rect 9622 -3784 12314 -3460
rect 13265 -3464 15043 -3264
rect 16409 -3464 18187 -3264
rect 19541 -3460 21319 -3260
rect 22685 -3460 24463 -3260
rect 12824 -3788 15516 -3464
rect 15968 -3788 18660 -3464
rect 19100 -3784 21792 -3460
rect 22244 -3784 24936 -3460
rect 610 -6114 1086 -5922
rect 2678 -6112 3154 -5922
rect 420 -6409 1264 -6114
rect 2488 -6407 3332 -6112
rect 4747 -6114 5223 -5922
rect 6815 -6112 7291 -5922
rect 8884 -6112 9360 -5920
rect 10952 -6110 11428 -5920
rect -61 -6733 1744 -6409
rect 2007 -6731 3812 -6407
rect 4557 -6409 5401 -6114
rect 6625 -6407 7469 -6112
rect 8694 -6407 9538 -6112
rect 10762 -6405 11606 -6110
rect 13021 -6112 13497 -5920
rect 15089 -6110 15565 -5920
rect 366 -7426 1204 -6733
rect 2434 -7424 3272 -6731
rect 4076 -6733 5881 -6409
rect 6144 -6731 7949 -6407
rect 8213 -6731 10018 -6407
rect 10281 -6729 12086 -6405
rect 12831 -6407 13675 -6112
rect 14899 -6405 15743 -6110
rect 4503 -7426 5341 -6733
rect 6571 -7424 7409 -6731
rect 8640 -7424 9478 -6731
rect 10708 -7422 11546 -6729
rect 12350 -6731 14155 -6407
rect 14418 -6729 16223 -6405
rect 16671 -6417 17155 -5865
rect 17409 -6413 17893 -5867
rect 18147 -6417 18631 -5867
rect 18889 -6419 19373 -5867
rect 19629 -6419 20113 -5867
rect 20367 -6419 20851 -5867
rect 21105 -6419 21589 -5867
rect 21843 -6419 22327 -5867
rect 12777 -7424 13615 -6731
rect 14845 -7422 15683 -6729
<< nmos >>
rect 484 3060 544 3460
rect 602 3060 662 3460
rect 837 3260 897 3460
rect 1932 3060 1992 3460
rect 2050 3060 2110 3460
rect 2285 3260 2345 3460
rect 3430 3062 3490 3462
rect 3548 3062 3608 3462
rect 3783 3262 3843 3462
rect 4878 3062 4938 3462
rect 4996 3062 5056 3462
rect 5231 3262 5291 3462
rect 6398 3060 6458 3460
rect 6516 3060 6576 3460
rect 6751 3260 6811 3460
rect 7846 3060 7906 3460
rect 7964 3060 8024 3460
rect 8199 3260 8259 3460
rect 9344 3062 9404 3462
rect 9462 3062 9522 3462
rect 9697 3262 9757 3462
rect 10792 3062 10852 3462
rect 10910 3062 10970 3462
rect 11145 3262 11205 3462
rect 11920 3108 11980 3308
rect 12038 3108 12098 3308
rect 12156 3108 12216 3308
rect 13088 3110 13148 3310
rect 13206 3110 13266 3310
rect 13324 3110 13384 3310
rect 14256 3110 14316 3310
rect 14374 3110 14434 3310
rect 14492 3110 14552 3310
rect 15424 3110 15484 3310
rect 15542 3110 15602 3310
rect 15660 3110 15720 3310
rect 16598 3110 16658 3310
rect 16716 3110 16776 3310
rect 16834 3110 16894 3310
rect 17766 3110 17826 3310
rect 17884 3110 17944 3310
rect 18002 3110 18062 3310
rect 18934 3112 18994 3312
rect 19052 3112 19112 3312
rect 19170 3112 19230 3312
rect 20102 3112 20162 3312
rect 20220 3112 20280 3312
rect 20338 3112 20398 3312
rect 1140 607 1200 807
rect 1332 407 1392 807
rect 1450 407 1510 807
rect 1568 407 1628 807
rect 1686 407 1746 807
rect 1882 607 1942 807
rect 4284 607 4344 807
rect 4476 407 4536 807
rect 4594 407 4654 807
rect 4712 407 4772 807
rect 4830 407 4890 807
rect 5026 607 5086 807
rect 7416 611 7476 811
rect 7608 411 7668 811
rect 7726 411 7786 811
rect 7844 411 7904 811
rect 7962 411 8022 811
rect 8158 611 8218 811
rect 10560 611 10620 811
rect 10752 411 10812 811
rect 10870 411 10930 811
rect 10988 411 11048 811
rect 11106 411 11166 811
rect 11302 611 11362 811
rect 13762 607 13822 807
rect 13954 407 14014 807
rect 14072 407 14132 807
rect 14190 407 14250 807
rect 14308 407 14368 807
rect 14504 607 14564 807
rect 16906 607 16966 807
rect 17098 407 17158 807
rect 17216 407 17276 807
rect 17334 407 17394 807
rect 17452 407 17512 807
rect 17648 607 17708 807
rect 20038 611 20098 811
rect 20230 411 20290 811
rect 20348 411 20408 811
rect 20466 411 20526 811
rect 20584 411 20644 811
rect 20780 611 20840 811
rect 23182 611 23242 811
rect 23374 411 23434 811
rect 23492 411 23552 811
rect 23610 411 23670 811
rect 23728 411 23788 811
rect 23924 611 23984 811
rect 1140 -2127 1200 -1927
rect 1332 -2327 1392 -1927
rect 1450 -2327 1510 -1927
rect 1568 -2327 1628 -1927
rect 1686 -2327 1746 -1927
rect 1882 -2127 1942 -1927
rect 4284 -2127 4344 -1927
rect 4476 -2327 4536 -1927
rect 4594 -2327 4654 -1927
rect 4712 -2327 4772 -1927
rect 4830 -2327 4890 -1927
rect 5026 -2127 5086 -1927
rect 7416 -2123 7476 -1923
rect 7608 -2323 7668 -1923
rect 7726 -2323 7786 -1923
rect 7844 -2323 7904 -1923
rect 7962 -2323 8022 -1923
rect 8158 -2123 8218 -1923
rect 10560 -2123 10620 -1923
rect 10752 -2323 10812 -1923
rect 10870 -2323 10930 -1923
rect 10988 -2323 11048 -1923
rect 11106 -2323 11166 -1923
rect 11302 -2123 11362 -1923
rect 13762 -2127 13822 -1927
rect 13954 -2327 14014 -1927
rect 14072 -2327 14132 -1927
rect 14190 -2327 14250 -1927
rect 14308 -2327 14368 -1927
rect 14504 -2127 14564 -1927
rect 16906 -2127 16966 -1927
rect 17098 -2327 17158 -1927
rect 17216 -2327 17276 -1927
rect 17334 -2327 17394 -1927
rect 17452 -2327 17512 -1927
rect 17648 -2127 17708 -1927
rect 20038 -2123 20098 -1923
rect 20230 -2323 20290 -1923
rect 20348 -2323 20408 -1923
rect 20466 -2323 20526 -1923
rect 20584 -2323 20644 -1923
rect 20780 -2123 20840 -1923
rect 23182 -2123 23242 -1923
rect 23374 -2323 23434 -1923
rect 23492 -2323 23552 -1923
rect 23610 -2323 23670 -1923
rect 23728 -2323 23788 -1923
rect 23924 -2123 23984 -1923
rect 1130 -4859 1190 -4659
rect 1322 -5059 1382 -4659
rect 1440 -5059 1500 -4659
rect 1558 -5059 1618 -4659
rect 1676 -5059 1736 -4659
rect 1872 -4859 1932 -4659
rect 4274 -4859 4334 -4659
rect 4466 -5059 4526 -4659
rect 4584 -5059 4644 -4659
rect 4702 -5059 4762 -4659
rect 4820 -5059 4880 -4659
rect 5016 -4859 5076 -4659
rect 7406 -4855 7466 -4655
rect 7598 -5055 7658 -4655
rect 7716 -5055 7776 -4655
rect 7834 -5055 7894 -4655
rect 7952 -5055 8012 -4655
rect 8148 -4855 8208 -4655
rect 10550 -4855 10610 -4655
rect 10742 -5055 10802 -4655
rect 10860 -5055 10920 -4655
rect 10978 -5055 11038 -4655
rect 11096 -5055 11156 -4655
rect 11292 -4855 11352 -4655
rect 13752 -4859 13812 -4659
rect 13944 -5059 14004 -4659
rect 14062 -5059 14122 -4659
rect 14180 -5059 14240 -4659
rect 14298 -5059 14358 -4659
rect 14494 -4859 14554 -4659
rect 16896 -4859 16956 -4659
rect 17088 -5059 17148 -4659
rect 17206 -5059 17266 -4659
rect 17324 -5059 17384 -4659
rect 17442 -5059 17502 -4659
rect 17638 -4859 17698 -4659
rect 20028 -4855 20088 -4655
rect 20220 -5055 20280 -4655
rect 20338 -5055 20398 -4655
rect 20456 -5055 20516 -4655
rect 20574 -5055 20634 -4655
rect 20770 -4855 20830 -4655
rect 23172 -4855 23232 -4655
rect 23364 -5055 23424 -4655
rect 23482 -5055 23542 -4655
rect 23600 -5055 23660 -4655
rect 23718 -5055 23778 -4655
rect 23914 -4855 23974 -4655
rect 158 -7896 218 -7696
rect 578 -8096 638 -7696
rect 696 -8096 756 -7696
rect 814 -8096 874 -7696
rect 932 -8096 992 -7696
rect 1456 -7896 1516 -7696
rect 2226 -7894 2286 -7694
rect 2646 -8094 2706 -7694
rect 2764 -8094 2824 -7694
rect 2882 -8094 2942 -7694
rect 3000 -8094 3060 -7694
rect 3524 -7894 3584 -7694
rect 4295 -7896 4355 -7696
rect 4715 -8096 4775 -7696
rect 4833 -8096 4893 -7696
rect 4951 -8096 5011 -7696
rect 5069 -8096 5129 -7696
rect 5593 -7896 5653 -7696
rect 6363 -7894 6423 -7694
rect 6783 -8094 6843 -7694
rect 6901 -8094 6961 -7694
rect 7019 -8094 7079 -7694
rect 7137 -8094 7197 -7694
rect 7661 -7894 7721 -7694
rect 8432 -7894 8492 -7694
rect 8852 -8094 8912 -7694
rect 8970 -8094 9030 -7694
rect 9088 -8094 9148 -7694
rect 9206 -8094 9266 -7694
rect 9730 -7894 9790 -7694
rect 10500 -7892 10560 -7692
rect 10920 -8092 10980 -7692
rect 11038 -8092 11098 -7692
rect 11156 -8092 11216 -7692
rect 11274 -8092 11334 -7692
rect 11798 -7892 11858 -7692
rect 16883 -6741 16943 -6541
rect 17621 -6739 17681 -6539
rect 18359 -6743 18419 -6543
rect 19101 -6743 19161 -6543
rect 19841 -6743 19901 -6543
rect 20579 -6743 20639 -6543
rect 21317 -6739 21377 -6539
rect 22055 -6739 22115 -6539
rect 12569 -7894 12629 -7694
rect 12989 -8094 13049 -7694
rect 13107 -8094 13167 -7694
rect 13225 -8094 13285 -7694
rect 13343 -8094 13403 -7694
rect 13867 -7894 13927 -7694
rect 14637 -7892 14697 -7692
rect 15057 -8092 15117 -7692
rect 15175 -8092 15235 -7692
rect 15293 -8092 15353 -7692
rect 15411 -8092 15471 -7692
rect 15935 -7892 15995 -7692
<< pmos >>
rect 247 3697 307 3897
rect 365 3697 425 3897
rect 483 3697 543 3897
rect 601 3697 661 3897
rect 719 3697 779 3897
rect 837 3697 897 3897
rect 955 3697 1015 3897
rect 1073 3697 1133 3897
rect 1191 3697 1251 3897
rect 1695 3697 1755 3897
rect 1813 3697 1873 3897
rect 1931 3697 1991 3897
rect 2049 3697 2109 3897
rect 2167 3697 2227 3897
rect 2285 3697 2345 3897
rect 2403 3697 2463 3897
rect 2521 3697 2581 3897
rect 2639 3697 2699 3897
rect 3193 3699 3253 3899
rect 3311 3699 3371 3899
rect 3429 3699 3489 3899
rect 3547 3699 3607 3899
rect 3665 3699 3725 3899
rect 3783 3699 3843 3899
rect 3901 3699 3961 3899
rect 4019 3699 4079 3899
rect 4137 3699 4197 3899
rect 4641 3699 4701 3899
rect 4759 3699 4819 3899
rect 4877 3699 4937 3899
rect 4995 3699 5055 3899
rect 5113 3699 5173 3899
rect 5231 3699 5291 3899
rect 5349 3699 5409 3899
rect 5467 3699 5527 3899
rect 5585 3699 5645 3899
rect 6161 3697 6221 3897
rect 6279 3697 6339 3897
rect 6397 3697 6457 3897
rect 6515 3697 6575 3897
rect 6633 3697 6693 3897
rect 6751 3697 6811 3897
rect 6869 3697 6929 3897
rect 6987 3697 7047 3897
rect 7105 3697 7165 3897
rect 7609 3697 7669 3897
rect 7727 3697 7787 3897
rect 7845 3697 7905 3897
rect 7963 3697 8023 3897
rect 8081 3697 8141 3897
rect 8199 3697 8259 3897
rect 8317 3697 8377 3897
rect 8435 3697 8495 3897
rect 8553 3697 8613 3897
rect 9107 3699 9167 3899
rect 9225 3699 9285 3899
rect 9343 3699 9403 3899
rect 9461 3699 9521 3899
rect 9579 3699 9639 3899
rect 9697 3699 9757 3899
rect 9815 3699 9875 3899
rect 9933 3699 9993 3899
rect 10051 3699 10111 3899
rect 10555 3699 10615 3899
rect 10673 3699 10733 3899
rect 10791 3699 10851 3899
rect 10909 3699 10969 3899
rect 11027 3699 11087 3899
rect 11145 3699 11205 3899
rect 11263 3699 11323 3899
rect 11381 3699 11441 3899
rect 11499 3699 11559 3899
rect 12010 3694 12070 4094
rect 12128 3694 12188 4094
rect 12246 3694 12306 4094
rect 12364 3694 12424 4094
rect 12482 3694 12542 4094
rect 12600 3694 12660 4094
rect 13178 3694 13238 4094
rect 13296 3694 13356 4094
rect 13414 3694 13474 4094
rect 13532 3694 13592 4094
rect 13650 3694 13710 4094
rect 13768 3694 13828 4094
rect 14346 3692 14406 4092
rect 14464 3692 14524 4092
rect 14582 3692 14642 4092
rect 14700 3692 14760 4092
rect 14818 3692 14878 4092
rect 14936 3692 14996 4092
rect 15514 3694 15574 4094
rect 15632 3694 15692 4094
rect 15750 3694 15810 4094
rect 15868 3694 15928 4094
rect 15986 3694 16046 4094
rect 16104 3694 16164 4094
rect 16688 3696 16748 4096
rect 16806 3696 16866 4096
rect 16924 3696 16984 4096
rect 17042 3696 17102 4096
rect 17160 3696 17220 4096
rect 17278 3696 17338 4096
rect 17856 3694 17916 4094
rect 17974 3694 18034 4094
rect 18092 3694 18152 4094
rect 18210 3694 18270 4094
rect 18328 3694 18388 4094
rect 18446 3694 18506 4094
rect 19024 3696 19084 4096
rect 19142 3696 19202 4096
rect 19260 3696 19320 4096
rect 19378 3696 19438 4096
rect 19496 3696 19556 4096
rect 19614 3696 19674 4096
rect 12440 3104 12500 3304
rect 12558 3104 12618 3304
rect 12676 3104 12736 3304
rect 13607 3110 13667 3310
rect 13725 3110 13785 3310
rect 13843 3110 13903 3310
rect 14775 3110 14835 3310
rect 14893 3110 14953 3310
rect 15011 3110 15071 3310
rect 15944 3110 16004 3310
rect 16062 3110 16122 3310
rect 16180 3110 16240 3310
rect 17116 3106 17176 3306
rect 17234 3106 17294 3306
rect 17352 3106 17412 3306
rect 20192 3694 20252 4094
rect 20310 3694 20370 4094
rect 20428 3694 20488 4094
rect 20546 3694 20606 4094
rect 20664 3694 20724 4094
rect 20782 3694 20842 4094
rect 18285 3105 18345 3305
rect 18403 3105 18463 3305
rect 18521 3105 18581 3305
rect 19453 3105 19513 3305
rect 19571 3105 19631 3305
rect 19689 3105 19749 3305
rect 20621 3106 20681 3306
rect 20739 3106 20799 3306
rect 20857 3106 20917 3306
rect 306 1740 366 1940
rect 424 1740 484 1940
rect 542 1740 602 1940
rect 747 1740 807 2140
rect 865 1740 925 2140
rect 983 1740 1043 2140
rect 1214 1740 1274 2140
rect 1332 1740 1392 2140
rect 1450 1740 1510 2140
rect 1568 1740 1628 2140
rect 1686 1740 1746 2140
rect 1804 1740 1864 2140
rect 2041 1740 2101 2140
rect 2159 1740 2219 2140
rect 2277 1740 2337 2140
rect 2514 1740 2574 1940
rect 2632 1740 2692 1940
rect 2750 1740 2810 1940
rect 3450 1740 3510 1940
rect 3568 1740 3628 1940
rect 3686 1740 3746 1940
rect 3891 1740 3951 2140
rect 4009 1740 4069 2140
rect 4127 1740 4187 2140
rect 4358 1740 4418 2140
rect 4476 1740 4536 2140
rect 4594 1740 4654 2140
rect 4712 1740 4772 2140
rect 4830 1740 4890 2140
rect 4948 1740 5008 2140
rect 5185 1740 5245 2140
rect 5303 1740 5363 2140
rect 5421 1740 5481 2140
rect 5658 1740 5718 1940
rect 5776 1740 5836 1940
rect 5894 1740 5954 1940
rect 6582 1744 6642 1944
rect 6700 1744 6760 1944
rect 6818 1744 6878 1944
rect 7023 1744 7083 2144
rect 7141 1744 7201 2144
rect 7259 1744 7319 2144
rect 7490 1744 7550 2144
rect 7608 1744 7668 2144
rect 7726 1744 7786 2144
rect 7844 1744 7904 2144
rect 7962 1744 8022 2144
rect 8080 1744 8140 2144
rect 8317 1744 8377 2144
rect 8435 1744 8495 2144
rect 8553 1744 8613 2144
rect 8790 1744 8850 1944
rect 8908 1744 8968 1944
rect 9026 1744 9086 1944
rect 9726 1744 9786 1944
rect 9844 1744 9904 1944
rect 9962 1744 10022 1944
rect 10167 1744 10227 2144
rect 10285 1744 10345 2144
rect 10403 1744 10463 2144
rect 10634 1744 10694 2144
rect 10752 1744 10812 2144
rect 10870 1744 10930 2144
rect 10988 1744 11048 2144
rect 11106 1744 11166 2144
rect 11224 1744 11284 2144
rect 11461 1744 11521 2144
rect 11579 1744 11639 2144
rect 11697 1744 11757 2144
rect 11934 1744 11994 1944
rect 12052 1744 12112 1944
rect 12170 1744 12230 1944
rect 12928 1740 12988 1940
rect 13046 1740 13106 1940
rect 13164 1740 13224 1940
rect 13369 1740 13429 2140
rect 13487 1740 13547 2140
rect 13605 1740 13665 2140
rect 13836 1740 13896 2140
rect 13954 1740 14014 2140
rect 14072 1740 14132 2140
rect 14190 1740 14250 2140
rect 14308 1740 14368 2140
rect 14426 1740 14486 2140
rect 14663 1740 14723 2140
rect 14781 1740 14841 2140
rect 14899 1740 14959 2140
rect 15136 1740 15196 1940
rect 15254 1740 15314 1940
rect 15372 1740 15432 1940
rect 16072 1740 16132 1940
rect 16190 1740 16250 1940
rect 16308 1740 16368 1940
rect 16513 1740 16573 2140
rect 16631 1740 16691 2140
rect 16749 1740 16809 2140
rect 16980 1740 17040 2140
rect 17098 1740 17158 2140
rect 17216 1740 17276 2140
rect 17334 1740 17394 2140
rect 17452 1740 17512 2140
rect 17570 1740 17630 2140
rect 17807 1740 17867 2140
rect 17925 1740 17985 2140
rect 18043 1740 18103 2140
rect 18280 1740 18340 1940
rect 18398 1740 18458 1940
rect 18516 1740 18576 1940
rect 19204 1744 19264 1944
rect 19322 1744 19382 1944
rect 19440 1744 19500 1944
rect 19645 1744 19705 2144
rect 19763 1744 19823 2144
rect 19881 1744 19941 2144
rect 20112 1744 20172 2144
rect 20230 1744 20290 2144
rect 20348 1744 20408 2144
rect 20466 1744 20526 2144
rect 20584 1744 20644 2144
rect 20702 1744 20762 2144
rect 20939 1744 20999 2144
rect 21057 1744 21117 2144
rect 21175 1744 21235 2144
rect 21412 1744 21472 1944
rect 21530 1744 21590 1944
rect 21648 1744 21708 1944
rect 22348 1744 22408 1944
rect 22466 1744 22526 1944
rect 22584 1744 22644 1944
rect 22789 1744 22849 2144
rect 22907 1744 22967 2144
rect 23025 1744 23085 2144
rect 23256 1744 23316 2144
rect 23374 1744 23434 2144
rect 23492 1744 23552 2144
rect 23610 1744 23670 2144
rect 23728 1744 23788 2144
rect 23846 1744 23906 2144
rect 24083 1744 24143 2144
rect 24201 1744 24261 2144
rect 24319 1744 24379 2144
rect 24556 1744 24616 1944
rect 24674 1744 24734 1944
rect 24792 1744 24852 1944
rect 306 -994 366 -794
rect 424 -994 484 -794
rect 542 -994 602 -794
rect 747 -994 807 -594
rect 865 -994 925 -594
rect 983 -994 1043 -594
rect 1214 -994 1274 -594
rect 1332 -994 1392 -594
rect 1450 -994 1510 -594
rect 1568 -994 1628 -594
rect 1686 -994 1746 -594
rect 1804 -994 1864 -594
rect 2041 -994 2101 -594
rect 2159 -994 2219 -594
rect 2277 -994 2337 -594
rect 2514 -994 2574 -794
rect 2632 -994 2692 -794
rect 2750 -994 2810 -794
rect 3450 -994 3510 -794
rect 3568 -994 3628 -794
rect 3686 -994 3746 -794
rect 3891 -994 3951 -594
rect 4009 -994 4069 -594
rect 4127 -994 4187 -594
rect 4358 -994 4418 -594
rect 4476 -994 4536 -594
rect 4594 -994 4654 -594
rect 4712 -994 4772 -594
rect 4830 -994 4890 -594
rect 4948 -994 5008 -594
rect 5185 -994 5245 -594
rect 5303 -994 5363 -594
rect 5421 -994 5481 -594
rect 5658 -994 5718 -794
rect 5776 -994 5836 -794
rect 5894 -994 5954 -794
rect 6582 -990 6642 -790
rect 6700 -990 6760 -790
rect 6818 -990 6878 -790
rect 7023 -990 7083 -590
rect 7141 -990 7201 -590
rect 7259 -990 7319 -590
rect 7490 -990 7550 -590
rect 7608 -990 7668 -590
rect 7726 -990 7786 -590
rect 7844 -990 7904 -590
rect 7962 -990 8022 -590
rect 8080 -990 8140 -590
rect 8317 -990 8377 -590
rect 8435 -990 8495 -590
rect 8553 -990 8613 -590
rect 8790 -990 8850 -790
rect 8908 -990 8968 -790
rect 9026 -990 9086 -790
rect 9726 -990 9786 -790
rect 9844 -990 9904 -790
rect 9962 -990 10022 -790
rect 10167 -990 10227 -590
rect 10285 -990 10345 -590
rect 10403 -990 10463 -590
rect 10634 -990 10694 -590
rect 10752 -990 10812 -590
rect 10870 -990 10930 -590
rect 10988 -990 11048 -590
rect 11106 -990 11166 -590
rect 11224 -990 11284 -590
rect 11461 -990 11521 -590
rect 11579 -990 11639 -590
rect 11697 -990 11757 -590
rect 11934 -990 11994 -790
rect 12052 -990 12112 -790
rect 12170 -990 12230 -790
rect 12928 -994 12988 -794
rect 13046 -994 13106 -794
rect 13164 -994 13224 -794
rect 13369 -994 13429 -594
rect 13487 -994 13547 -594
rect 13605 -994 13665 -594
rect 13836 -994 13896 -594
rect 13954 -994 14014 -594
rect 14072 -994 14132 -594
rect 14190 -994 14250 -594
rect 14308 -994 14368 -594
rect 14426 -994 14486 -594
rect 14663 -994 14723 -594
rect 14781 -994 14841 -594
rect 14899 -994 14959 -594
rect 15136 -994 15196 -794
rect 15254 -994 15314 -794
rect 15372 -994 15432 -794
rect 16072 -994 16132 -794
rect 16190 -994 16250 -794
rect 16308 -994 16368 -794
rect 16513 -994 16573 -594
rect 16631 -994 16691 -594
rect 16749 -994 16809 -594
rect 16980 -994 17040 -594
rect 17098 -994 17158 -594
rect 17216 -994 17276 -594
rect 17334 -994 17394 -594
rect 17452 -994 17512 -594
rect 17570 -994 17630 -594
rect 17807 -994 17867 -594
rect 17925 -994 17985 -594
rect 18043 -994 18103 -594
rect 18280 -994 18340 -794
rect 18398 -994 18458 -794
rect 18516 -994 18576 -794
rect 19204 -990 19264 -790
rect 19322 -990 19382 -790
rect 19440 -990 19500 -790
rect 19645 -990 19705 -590
rect 19763 -990 19823 -590
rect 19881 -990 19941 -590
rect 20112 -990 20172 -590
rect 20230 -990 20290 -590
rect 20348 -990 20408 -590
rect 20466 -990 20526 -590
rect 20584 -990 20644 -590
rect 20702 -990 20762 -590
rect 20939 -990 20999 -590
rect 21057 -990 21117 -590
rect 21175 -990 21235 -590
rect 21412 -990 21472 -790
rect 21530 -990 21590 -790
rect 21648 -990 21708 -790
rect 22348 -990 22408 -790
rect 22466 -990 22526 -790
rect 22584 -990 22644 -790
rect 22789 -990 22849 -590
rect 22907 -990 22967 -590
rect 23025 -990 23085 -590
rect 23256 -990 23316 -590
rect 23374 -990 23434 -590
rect 23492 -990 23552 -590
rect 23610 -990 23670 -590
rect 23728 -990 23788 -590
rect 23846 -990 23906 -590
rect 24083 -990 24143 -590
rect 24201 -990 24261 -590
rect 24319 -990 24379 -590
rect 24556 -990 24616 -790
rect 24674 -990 24734 -790
rect 24792 -990 24852 -790
rect 296 -3726 356 -3526
rect 414 -3726 474 -3526
rect 532 -3726 592 -3526
rect 737 -3726 797 -3326
rect 855 -3726 915 -3326
rect 973 -3726 1033 -3326
rect 1204 -3726 1264 -3326
rect 1322 -3726 1382 -3326
rect 1440 -3726 1500 -3326
rect 1558 -3726 1618 -3326
rect 1676 -3726 1736 -3326
rect 1794 -3726 1854 -3326
rect 2031 -3726 2091 -3326
rect 2149 -3726 2209 -3326
rect 2267 -3726 2327 -3326
rect 2504 -3726 2564 -3526
rect 2622 -3726 2682 -3526
rect 2740 -3726 2800 -3526
rect 3440 -3726 3500 -3526
rect 3558 -3726 3618 -3526
rect 3676 -3726 3736 -3526
rect 3881 -3726 3941 -3326
rect 3999 -3726 4059 -3326
rect 4117 -3726 4177 -3326
rect 4348 -3726 4408 -3326
rect 4466 -3726 4526 -3326
rect 4584 -3726 4644 -3326
rect 4702 -3726 4762 -3326
rect 4820 -3726 4880 -3326
rect 4938 -3726 4998 -3326
rect 5175 -3726 5235 -3326
rect 5293 -3726 5353 -3326
rect 5411 -3726 5471 -3326
rect 5648 -3726 5708 -3526
rect 5766 -3726 5826 -3526
rect 5884 -3726 5944 -3526
rect 6572 -3722 6632 -3522
rect 6690 -3722 6750 -3522
rect 6808 -3722 6868 -3522
rect 7013 -3722 7073 -3322
rect 7131 -3722 7191 -3322
rect 7249 -3722 7309 -3322
rect 7480 -3722 7540 -3322
rect 7598 -3722 7658 -3322
rect 7716 -3722 7776 -3322
rect 7834 -3722 7894 -3322
rect 7952 -3722 8012 -3322
rect 8070 -3722 8130 -3322
rect 8307 -3722 8367 -3322
rect 8425 -3722 8485 -3322
rect 8543 -3722 8603 -3322
rect 8780 -3722 8840 -3522
rect 8898 -3722 8958 -3522
rect 9016 -3722 9076 -3522
rect 9716 -3722 9776 -3522
rect 9834 -3722 9894 -3522
rect 9952 -3722 10012 -3522
rect 10157 -3722 10217 -3322
rect 10275 -3722 10335 -3322
rect 10393 -3722 10453 -3322
rect 10624 -3722 10684 -3322
rect 10742 -3722 10802 -3322
rect 10860 -3722 10920 -3322
rect 10978 -3722 11038 -3322
rect 11096 -3722 11156 -3322
rect 11214 -3722 11274 -3322
rect 11451 -3722 11511 -3322
rect 11569 -3722 11629 -3322
rect 11687 -3722 11747 -3322
rect 11924 -3722 11984 -3522
rect 12042 -3722 12102 -3522
rect 12160 -3722 12220 -3522
rect 12918 -3726 12978 -3526
rect 13036 -3726 13096 -3526
rect 13154 -3726 13214 -3526
rect 13359 -3726 13419 -3326
rect 13477 -3726 13537 -3326
rect 13595 -3726 13655 -3326
rect 13826 -3726 13886 -3326
rect 13944 -3726 14004 -3326
rect 14062 -3726 14122 -3326
rect 14180 -3726 14240 -3326
rect 14298 -3726 14358 -3326
rect 14416 -3726 14476 -3326
rect 14653 -3726 14713 -3326
rect 14771 -3726 14831 -3326
rect 14889 -3726 14949 -3326
rect 15126 -3726 15186 -3526
rect 15244 -3726 15304 -3526
rect 15362 -3726 15422 -3526
rect 16062 -3726 16122 -3526
rect 16180 -3726 16240 -3526
rect 16298 -3726 16358 -3526
rect 16503 -3726 16563 -3326
rect 16621 -3726 16681 -3326
rect 16739 -3726 16799 -3326
rect 16970 -3726 17030 -3326
rect 17088 -3726 17148 -3326
rect 17206 -3726 17266 -3326
rect 17324 -3726 17384 -3326
rect 17442 -3726 17502 -3326
rect 17560 -3726 17620 -3326
rect 17797 -3726 17857 -3326
rect 17915 -3726 17975 -3326
rect 18033 -3726 18093 -3326
rect 18270 -3726 18330 -3526
rect 18388 -3726 18448 -3526
rect 18506 -3726 18566 -3526
rect 19194 -3722 19254 -3522
rect 19312 -3722 19372 -3522
rect 19430 -3722 19490 -3522
rect 19635 -3722 19695 -3322
rect 19753 -3722 19813 -3322
rect 19871 -3722 19931 -3322
rect 20102 -3722 20162 -3322
rect 20220 -3722 20280 -3322
rect 20338 -3722 20398 -3322
rect 20456 -3722 20516 -3322
rect 20574 -3722 20634 -3322
rect 20692 -3722 20752 -3322
rect 20929 -3722 20989 -3322
rect 21047 -3722 21107 -3322
rect 21165 -3722 21225 -3322
rect 21402 -3722 21462 -3522
rect 21520 -3722 21580 -3522
rect 21638 -3722 21698 -3522
rect 22338 -3722 22398 -3522
rect 22456 -3722 22516 -3522
rect 22574 -3722 22634 -3522
rect 22779 -3722 22839 -3322
rect 22897 -3722 22957 -3322
rect 23015 -3722 23075 -3322
rect 23246 -3722 23306 -3322
rect 23364 -3722 23424 -3322
rect 23482 -3722 23542 -3322
rect 23600 -3722 23660 -3322
rect 23718 -3722 23778 -3322
rect 23836 -3722 23896 -3322
rect 24073 -3722 24133 -3322
rect 24191 -3722 24251 -3322
rect 24309 -3722 24369 -3322
rect 24546 -3722 24606 -3522
rect 24664 -3722 24724 -3522
rect 24782 -3722 24842 -3522
rect 33 -6671 93 -6471
rect 151 -6671 211 -6471
rect 269 -6671 329 -6471
rect 517 -6671 577 -6271
rect 635 -6671 695 -6271
rect 753 -6671 813 -6271
rect 871 -6671 931 -6271
rect 989 -6671 1049 -6271
rect 1107 -6671 1167 -6271
rect 1354 -6671 1414 -6471
rect 1472 -6671 1532 -6471
rect 1590 -6671 1650 -6471
rect 2101 -6669 2161 -6469
rect 2219 -6669 2279 -6469
rect 2337 -6669 2397 -6469
rect 2585 -6669 2645 -6269
rect 2703 -6669 2763 -6269
rect 2821 -6669 2881 -6269
rect 2939 -6669 2999 -6269
rect 3057 -6669 3117 -6269
rect 3175 -6669 3235 -6269
rect 3422 -6669 3482 -6469
rect 3540 -6669 3600 -6469
rect 3658 -6669 3718 -6469
rect 460 -7364 520 -6964
rect 578 -7364 638 -6964
rect 696 -7364 756 -6964
rect 814 -7364 874 -6964
rect 932 -7364 992 -6964
rect 1050 -7364 1110 -6964
rect 4170 -6671 4230 -6471
rect 4288 -6671 4348 -6471
rect 4406 -6671 4466 -6471
rect 4654 -6671 4714 -6271
rect 4772 -6671 4832 -6271
rect 4890 -6671 4950 -6271
rect 5008 -6671 5068 -6271
rect 5126 -6671 5186 -6271
rect 5244 -6671 5304 -6271
rect 5491 -6671 5551 -6471
rect 5609 -6671 5669 -6471
rect 5727 -6671 5787 -6471
rect 6238 -6669 6298 -6469
rect 6356 -6669 6416 -6469
rect 6474 -6669 6534 -6469
rect 6722 -6669 6782 -6269
rect 6840 -6669 6900 -6269
rect 6958 -6669 7018 -6269
rect 7076 -6669 7136 -6269
rect 7194 -6669 7254 -6269
rect 7312 -6669 7372 -6269
rect 7559 -6669 7619 -6469
rect 7677 -6669 7737 -6469
rect 7795 -6669 7855 -6469
rect 8307 -6669 8367 -6469
rect 8425 -6669 8485 -6469
rect 8543 -6669 8603 -6469
rect 8791 -6669 8851 -6269
rect 8909 -6669 8969 -6269
rect 9027 -6669 9087 -6269
rect 9145 -6669 9205 -6269
rect 9263 -6669 9323 -6269
rect 9381 -6669 9441 -6269
rect 9628 -6669 9688 -6469
rect 9746 -6669 9806 -6469
rect 9864 -6669 9924 -6469
rect 10375 -6667 10435 -6467
rect 10493 -6667 10553 -6467
rect 10611 -6667 10671 -6467
rect 10859 -6667 10919 -6267
rect 10977 -6667 11037 -6267
rect 11095 -6667 11155 -6267
rect 11213 -6667 11273 -6267
rect 11331 -6667 11391 -6267
rect 11449 -6667 11509 -6267
rect 11696 -6667 11756 -6467
rect 11814 -6667 11874 -6467
rect 11932 -6667 11992 -6467
rect 2528 -7362 2588 -6962
rect 2646 -7362 2706 -6962
rect 2764 -7362 2824 -6962
rect 2882 -7362 2942 -6962
rect 3000 -7362 3060 -6962
rect 3118 -7362 3178 -6962
rect 4597 -7364 4657 -6964
rect 4715 -7364 4775 -6964
rect 4833 -7364 4893 -6964
rect 4951 -7364 5011 -6964
rect 5069 -7364 5129 -6964
rect 5187 -7364 5247 -6964
rect 6665 -7362 6725 -6962
rect 6783 -7362 6843 -6962
rect 6901 -7362 6961 -6962
rect 7019 -7362 7079 -6962
rect 7137 -7362 7197 -6962
rect 7255 -7362 7315 -6962
rect 8734 -7362 8794 -6962
rect 8852 -7362 8912 -6962
rect 8970 -7362 9030 -6962
rect 9088 -7362 9148 -6962
rect 9206 -7362 9266 -6962
rect 9324 -7362 9384 -6962
rect 12444 -6669 12504 -6469
rect 12562 -6669 12622 -6469
rect 12680 -6669 12740 -6469
rect 12928 -6669 12988 -6269
rect 13046 -6669 13106 -6269
rect 13164 -6669 13224 -6269
rect 13282 -6669 13342 -6269
rect 13400 -6669 13460 -6269
rect 13518 -6669 13578 -6269
rect 13765 -6669 13825 -6469
rect 13883 -6669 13943 -6469
rect 14001 -6669 14061 -6469
rect 14512 -6667 14572 -6467
rect 14630 -6667 14690 -6467
rect 14748 -6667 14808 -6467
rect 14996 -6667 15056 -6267
rect 15114 -6667 15174 -6267
rect 15232 -6667 15292 -6267
rect 15350 -6667 15410 -6267
rect 15468 -6667 15528 -6267
rect 15586 -6667 15646 -6267
rect 16765 -6355 16825 -6155
rect 16883 -6355 16943 -6155
rect 17001 -6355 17061 -6155
rect 17503 -6351 17563 -6151
rect 17621 -6351 17681 -6151
rect 17739 -6351 17799 -6151
rect 18241 -6355 18301 -6155
rect 18359 -6355 18419 -6155
rect 18477 -6355 18537 -6155
rect 18983 -6357 19043 -6157
rect 19101 -6357 19161 -6157
rect 19219 -6357 19279 -6157
rect 19723 -6357 19783 -6157
rect 19841 -6357 19901 -6157
rect 19959 -6357 20019 -6157
rect 20461 -6357 20521 -6157
rect 20579 -6357 20639 -6157
rect 20697 -6357 20757 -6157
rect 21199 -6357 21259 -6157
rect 21317 -6357 21377 -6157
rect 21435 -6357 21495 -6157
rect 21937 -6357 21997 -6157
rect 22055 -6357 22115 -6157
rect 22173 -6357 22233 -6157
rect 15833 -6667 15893 -6467
rect 15951 -6667 16011 -6467
rect 16069 -6667 16129 -6467
rect 10802 -7360 10862 -6960
rect 10920 -7360 10980 -6960
rect 11038 -7360 11098 -6960
rect 11156 -7360 11216 -6960
rect 11274 -7360 11334 -6960
rect 11392 -7360 11452 -6960
rect 12871 -7362 12931 -6962
rect 12989 -7362 13049 -6962
rect 13107 -7362 13167 -6962
rect 13225 -7362 13285 -6962
rect 13343 -7362 13403 -6962
rect 13461 -7362 13521 -6962
rect 14939 -7360 14999 -6960
rect 15057 -7360 15117 -6960
rect 15175 -7360 15235 -6960
rect 15293 -7360 15353 -6960
rect 15411 -7360 15471 -6960
rect 15529 -7360 15589 -6960
<< ndiff >>
rect 426 3448 484 3460
rect 426 3072 438 3448
rect 472 3072 484 3448
rect 426 3060 484 3072
rect 544 3448 602 3460
rect 544 3072 556 3448
rect 590 3072 602 3448
rect 544 3060 602 3072
rect 662 3448 720 3460
rect 662 3072 674 3448
rect 708 3072 720 3448
rect 779 3448 837 3460
rect 779 3272 791 3448
rect 825 3272 837 3448
rect 779 3260 837 3272
rect 897 3448 955 3460
rect 897 3272 909 3448
rect 943 3272 955 3448
rect 897 3260 955 3272
rect 1874 3448 1932 3460
rect 662 3060 720 3072
rect 1874 3072 1886 3448
rect 1920 3072 1932 3448
rect 1874 3060 1932 3072
rect 1992 3448 2050 3460
rect 1992 3072 2004 3448
rect 2038 3072 2050 3448
rect 1992 3060 2050 3072
rect 2110 3448 2168 3460
rect 2110 3072 2122 3448
rect 2156 3072 2168 3448
rect 2227 3448 2285 3460
rect 2227 3272 2239 3448
rect 2273 3272 2285 3448
rect 2227 3260 2285 3272
rect 2345 3448 2403 3460
rect 2345 3272 2357 3448
rect 2391 3272 2403 3448
rect 2345 3260 2403 3272
rect 3372 3450 3430 3462
rect 2110 3060 2168 3072
rect 3372 3074 3384 3450
rect 3418 3074 3430 3450
rect 3372 3062 3430 3074
rect 3490 3450 3548 3462
rect 3490 3074 3502 3450
rect 3536 3074 3548 3450
rect 3490 3062 3548 3074
rect 3608 3450 3666 3462
rect 3608 3074 3620 3450
rect 3654 3074 3666 3450
rect 3725 3450 3783 3462
rect 3725 3274 3737 3450
rect 3771 3274 3783 3450
rect 3725 3262 3783 3274
rect 3843 3450 3901 3462
rect 3843 3274 3855 3450
rect 3889 3274 3901 3450
rect 3843 3262 3901 3274
rect 4820 3450 4878 3462
rect 3608 3062 3666 3074
rect 4820 3074 4832 3450
rect 4866 3074 4878 3450
rect 4820 3062 4878 3074
rect 4938 3450 4996 3462
rect 4938 3074 4950 3450
rect 4984 3074 4996 3450
rect 4938 3062 4996 3074
rect 5056 3450 5114 3462
rect 5056 3074 5068 3450
rect 5102 3074 5114 3450
rect 5173 3450 5231 3462
rect 5173 3274 5185 3450
rect 5219 3274 5231 3450
rect 5173 3262 5231 3274
rect 5291 3450 5349 3462
rect 5291 3274 5303 3450
rect 5337 3274 5349 3450
rect 5291 3262 5349 3274
rect 6340 3448 6398 3460
rect 5056 3062 5114 3074
rect 6340 3072 6352 3448
rect 6386 3072 6398 3448
rect 6340 3060 6398 3072
rect 6458 3448 6516 3460
rect 6458 3072 6470 3448
rect 6504 3072 6516 3448
rect 6458 3060 6516 3072
rect 6576 3448 6634 3460
rect 6576 3072 6588 3448
rect 6622 3072 6634 3448
rect 6693 3448 6751 3460
rect 6693 3272 6705 3448
rect 6739 3272 6751 3448
rect 6693 3260 6751 3272
rect 6811 3448 6869 3460
rect 6811 3272 6823 3448
rect 6857 3272 6869 3448
rect 6811 3260 6869 3272
rect 7788 3448 7846 3460
rect 6576 3060 6634 3072
rect 7788 3072 7800 3448
rect 7834 3072 7846 3448
rect 7788 3060 7846 3072
rect 7906 3448 7964 3460
rect 7906 3072 7918 3448
rect 7952 3072 7964 3448
rect 7906 3060 7964 3072
rect 8024 3448 8082 3460
rect 8024 3072 8036 3448
rect 8070 3072 8082 3448
rect 8141 3448 8199 3460
rect 8141 3272 8153 3448
rect 8187 3272 8199 3448
rect 8141 3260 8199 3272
rect 8259 3448 8317 3460
rect 8259 3272 8271 3448
rect 8305 3272 8317 3448
rect 8259 3260 8317 3272
rect 9286 3450 9344 3462
rect 8024 3060 8082 3072
rect 9286 3074 9298 3450
rect 9332 3074 9344 3450
rect 9286 3062 9344 3074
rect 9404 3450 9462 3462
rect 9404 3074 9416 3450
rect 9450 3074 9462 3450
rect 9404 3062 9462 3074
rect 9522 3450 9580 3462
rect 9522 3074 9534 3450
rect 9568 3074 9580 3450
rect 9639 3450 9697 3462
rect 9639 3274 9651 3450
rect 9685 3274 9697 3450
rect 9639 3262 9697 3274
rect 9757 3450 9815 3462
rect 9757 3274 9769 3450
rect 9803 3274 9815 3450
rect 9757 3262 9815 3274
rect 10734 3450 10792 3462
rect 9522 3062 9580 3074
rect 10734 3074 10746 3450
rect 10780 3074 10792 3450
rect 10734 3062 10792 3074
rect 10852 3450 10910 3462
rect 10852 3074 10864 3450
rect 10898 3074 10910 3450
rect 10852 3062 10910 3074
rect 10970 3450 11028 3462
rect 10970 3074 10982 3450
rect 11016 3074 11028 3450
rect 11087 3450 11145 3462
rect 11087 3274 11099 3450
rect 11133 3274 11145 3450
rect 11087 3262 11145 3274
rect 11205 3450 11263 3462
rect 11205 3274 11217 3450
rect 11251 3274 11263 3450
rect 11205 3262 11263 3274
rect 11862 3296 11920 3308
rect 11862 3120 11874 3296
rect 11908 3120 11920 3296
rect 11862 3108 11920 3120
rect 11980 3296 12038 3308
rect 11980 3120 11992 3296
rect 12026 3120 12038 3296
rect 11980 3108 12038 3120
rect 12098 3296 12156 3308
rect 12098 3120 12110 3296
rect 12144 3120 12156 3296
rect 12098 3108 12156 3120
rect 12216 3296 12274 3308
rect 12216 3120 12228 3296
rect 12262 3120 12274 3296
rect 12216 3108 12274 3120
rect 10970 3062 11028 3074
rect 13030 3298 13088 3310
rect 13030 3122 13042 3298
rect 13076 3122 13088 3298
rect 13030 3110 13088 3122
rect 13148 3298 13206 3310
rect 13148 3122 13160 3298
rect 13194 3122 13206 3298
rect 13148 3110 13206 3122
rect 13266 3298 13324 3310
rect 13266 3122 13278 3298
rect 13312 3122 13324 3298
rect 13266 3110 13324 3122
rect 13384 3298 13442 3310
rect 13384 3122 13396 3298
rect 13430 3122 13442 3298
rect 13384 3110 13442 3122
rect 14198 3298 14256 3310
rect 14198 3122 14210 3298
rect 14244 3122 14256 3298
rect 14198 3110 14256 3122
rect 14316 3298 14374 3310
rect 14316 3122 14328 3298
rect 14362 3122 14374 3298
rect 14316 3110 14374 3122
rect 14434 3298 14492 3310
rect 14434 3122 14446 3298
rect 14480 3122 14492 3298
rect 14434 3110 14492 3122
rect 14552 3298 14610 3310
rect 14552 3122 14564 3298
rect 14598 3122 14610 3298
rect 14552 3110 14610 3122
rect 15366 3298 15424 3310
rect 15366 3122 15378 3298
rect 15412 3122 15424 3298
rect 15366 3110 15424 3122
rect 15484 3298 15542 3310
rect 15484 3122 15496 3298
rect 15530 3122 15542 3298
rect 15484 3110 15542 3122
rect 15602 3298 15660 3310
rect 15602 3122 15614 3298
rect 15648 3122 15660 3298
rect 15602 3110 15660 3122
rect 15720 3298 15778 3310
rect 15720 3122 15732 3298
rect 15766 3122 15778 3298
rect 15720 3110 15778 3122
rect 16540 3298 16598 3310
rect 16540 3122 16552 3298
rect 16586 3122 16598 3298
rect 16540 3110 16598 3122
rect 16658 3298 16716 3310
rect 16658 3122 16670 3298
rect 16704 3122 16716 3298
rect 16658 3110 16716 3122
rect 16776 3298 16834 3310
rect 16776 3122 16788 3298
rect 16822 3122 16834 3298
rect 16776 3110 16834 3122
rect 16894 3298 16952 3310
rect 16894 3122 16906 3298
rect 16940 3122 16952 3298
rect 16894 3110 16952 3122
rect 17708 3298 17766 3310
rect 17708 3122 17720 3298
rect 17754 3122 17766 3298
rect 17708 3110 17766 3122
rect 17826 3298 17884 3310
rect 17826 3122 17838 3298
rect 17872 3122 17884 3298
rect 17826 3110 17884 3122
rect 17944 3298 18002 3310
rect 17944 3122 17956 3298
rect 17990 3122 18002 3298
rect 17944 3110 18002 3122
rect 18062 3298 18120 3310
rect 18062 3122 18074 3298
rect 18108 3122 18120 3298
rect 18062 3110 18120 3122
rect 18876 3300 18934 3312
rect 18876 3124 18888 3300
rect 18922 3124 18934 3300
rect 18876 3112 18934 3124
rect 18994 3300 19052 3312
rect 18994 3124 19006 3300
rect 19040 3124 19052 3300
rect 18994 3112 19052 3124
rect 19112 3300 19170 3312
rect 19112 3124 19124 3300
rect 19158 3124 19170 3300
rect 19112 3112 19170 3124
rect 19230 3300 19288 3312
rect 19230 3124 19242 3300
rect 19276 3124 19288 3300
rect 19230 3112 19288 3124
rect 20044 3300 20102 3312
rect 20044 3124 20056 3300
rect 20090 3124 20102 3300
rect 20044 3112 20102 3124
rect 20162 3300 20220 3312
rect 20162 3124 20174 3300
rect 20208 3124 20220 3300
rect 20162 3112 20220 3124
rect 20280 3300 20338 3312
rect 20280 3124 20292 3300
rect 20326 3124 20338 3300
rect 20280 3112 20338 3124
rect 20398 3300 20456 3312
rect 20398 3124 20410 3300
rect 20444 3124 20456 3300
rect 20398 3112 20456 3124
rect 1082 795 1140 807
rect 1082 619 1094 795
rect 1128 619 1140 795
rect 1082 607 1140 619
rect 1200 795 1332 807
rect 1200 619 1212 795
rect 1246 619 1286 795
rect 1200 607 1286 619
rect 1274 419 1286 607
rect 1320 419 1332 795
rect 1274 407 1332 419
rect 1392 795 1450 807
rect 1392 419 1404 795
rect 1438 419 1450 795
rect 1392 407 1450 419
rect 1510 795 1568 807
rect 1510 419 1522 795
rect 1556 419 1568 795
rect 1510 407 1568 419
rect 1628 795 1686 807
rect 1628 419 1640 795
rect 1674 419 1686 795
rect 1628 407 1686 419
rect 1746 795 1882 807
rect 1746 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1882 795
rect 1792 607 1882 619
rect 1942 795 2000 807
rect 1942 619 1954 795
rect 1988 619 2000 795
rect 1942 607 2000 619
rect 4226 795 4284 807
rect 4226 619 4238 795
rect 4272 619 4284 795
rect 4226 607 4284 619
rect 4344 795 4476 807
rect 4344 619 4356 795
rect 4390 619 4430 795
rect 4344 607 4430 619
rect 1792 419 1804 607
rect 1746 407 1804 419
rect 4418 419 4430 607
rect 4464 419 4476 795
rect 4418 407 4476 419
rect 4536 795 4594 807
rect 4536 419 4548 795
rect 4582 419 4594 795
rect 4536 407 4594 419
rect 4654 795 4712 807
rect 4654 419 4666 795
rect 4700 419 4712 795
rect 4654 407 4712 419
rect 4772 795 4830 807
rect 4772 419 4784 795
rect 4818 419 4830 795
rect 4772 407 4830 419
rect 4890 795 5026 807
rect 4890 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5026 795
rect 4936 607 5026 619
rect 5086 795 5144 807
rect 5086 619 5098 795
rect 5132 619 5144 795
rect 5086 607 5144 619
rect 7358 799 7416 811
rect 7358 623 7370 799
rect 7404 623 7416 799
rect 7358 611 7416 623
rect 7476 799 7608 811
rect 7476 623 7488 799
rect 7522 623 7562 799
rect 7476 611 7562 623
rect 4936 419 4948 607
rect 4890 407 4948 419
rect 7550 423 7562 611
rect 7596 423 7608 799
rect 7550 411 7608 423
rect 7668 799 7726 811
rect 7668 423 7680 799
rect 7714 423 7726 799
rect 7668 411 7726 423
rect 7786 799 7844 811
rect 7786 423 7798 799
rect 7832 423 7844 799
rect 7786 411 7844 423
rect 7904 799 7962 811
rect 7904 423 7916 799
rect 7950 423 7962 799
rect 7904 411 7962 423
rect 8022 799 8158 811
rect 8022 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8158 799
rect 8068 611 8158 623
rect 8218 799 8276 811
rect 8218 623 8230 799
rect 8264 623 8276 799
rect 8218 611 8276 623
rect 10502 799 10560 811
rect 10502 623 10514 799
rect 10548 623 10560 799
rect 10502 611 10560 623
rect 10620 799 10752 811
rect 10620 623 10632 799
rect 10666 623 10706 799
rect 10620 611 10706 623
rect 8068 423 8080 611
rect 8022 411 8080 423
rect 10694 423 10706 611
rect 10740 423 10752 799
rect 10694 411 10752 423
rect 10812 799 10870 811
rect 10812 423 10824 799
rect 10858 423 10870 799
rect 10812 411 10870 423
rect 10930 799 10988 811
rect 10930 423 10942 799
rect 10976 423 10988 799
rect 10930 411 10988 423
rect 11048 799 11106 811
rect 11048 423 11060 799
rect 11094 423 11106 799
rect 11048 411 11106 423
rect 11166 799 11302 811
rect 11166 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11302 799
rect 11212 611 11302 623
rect 11362 799 11420 811
rect 11362 623 11374 799
rect 11408 623 11420 799
rect 11362 611 11420 623
rect 13704 795 13762 807
rect 13704 619 13716 795
rect 13750 619 13762 795
rect 11212 423 11224 611
rect 11166 411 11224 423
rect 13704 607 13762 619
rect 13822 795 13954 807
rect 13822 619 13834 795
rect 13868 619 13908 795
rect 13822 607 13908 619
rect 13896 419 13908 607
rect 13942 419 13954 795
rect 13896 407 13954 419
rect 14014 795 14072 807
rect 14014 419 14026 795
rect 14060 419 14072 795
rect 14014 407 14072 419
rect 14132 795 14190 807
rect 14132 419 14144 795
rect 14178 419 14190 795
rect 14132 407 14190 419
rect 14250 795 14308 807
rect 14250 419 14262 795
rect 14296 419 14308 795
rect 14250 407 14308 419
rect 14368 795 14504 807
rect 14368 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14504 795
rect 14414 607 14504 619
rect 14564 795 14622 807
rect 14564 619 14576 795
rect 14610 619 14622 795
rect 14564 607 14622 619
rect 16848 795 16906 807
rect 16848 619 16860 795
rect 16894 619 16906 795
rect 16848 607 16906 619
rect 16966 795 17098 807
rect 16966 619 16978 795
rect 17012 619 17052 795
rect 16966 607 17052 619
rect 14414 419 14426 607
rect 14368 407 14426 419
rect 17040 419 17052 607
rect 17086 419 17098 795
rect 17040 407 17098 419
rect 17158 795 17216 807
rect 17158 419 17170 795
rect 17204 419 17216 795
rect 17158 407 17216 419
rect 17276 795 17334 807
rect 17276 419 17288 795
rect 17322 419 17334 795
rect 17276 407 17334 419
rect 17394 795 17452 807
rect 17394 419 17406 795
rect 17440 419 17452 795
rect 17394 407 17452 419
rect 17512 795 17648 807
rect 17512 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17648 795
rect 17558 607 17648 619
rect 17708 795 17766 807
rect 17708 619 17720 795
rect 17754 619 17766 795
rect 17708 607 17766 619
rect 19980 799 20038 811
rect 19980 623 19992 799
rect 20026 623 20038 799
rect 19980 611 20038 623
rect 20098 799 20230 811
rect 20098 623 20110 799
rect 20144 623 20184 799
rect 20098 611 20184 623
rect 17558 419 17570 607
rect 17512 407 17570 419
rect 20172 423 20184 611
rect 20218 423 20230 799
rect 20172 411 20230 423
rect 20290 799 20348 811
rect 20290 423 20302 799
rect 20336 423 20348 799
rect 20290 411 20348 423
rect 20408 799 20466 811
rect 20408 423 20420 799
rect 20454 423 20466 799
rect 20408 411 20466 423
rect 20526 799 20584 811
rect 20526 423 20538 799
rect 20572 423 20584 799
rect 20526 411 20584 423
rect 20644 799 20780 811
rect 20644 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20780 799
rect 20690 611 20780 623
rect 20840 799 20898 811
rect 20840 623 20852 799
rect 20886 623 20898 799
rect 20840 611 20898 623
rect 23124 799 23182 811
rect 23124 623 23136 799
rect 23170 623 23182 799
rect 23124 611 23182 623
rect 23242 799 23374 811
rect 23242 623 23254 799
rect 23288 623 23328 799
rect 23242 611 23328 623
rect 20690 423 20702 611
rect 20644 411 20702 423
rect 23316 423 23328 611
rect 23362 423 23374 799
rect 23316 411 23374 423
rect 23434 799 23492 811
rect 23434 423 23446 799
rect 23480 423 23492 799
rect 23434 411 23492 423
rect 23552 799 23610 811
rect 23552 423 23564 799
rect 23598 423 23610 799
rect 23552 411 23610 423
rect 23670 799 23728 811
rect 23670 423 23682 799
rect 23716 423 23728 799
rect 23670 411 23728 423
rect 23788 799 23924 811
rect 23788 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23924 799
rect 23834 611 23924 623
rect 23984 799 24042 811
rect 23984 623 23996 799
rect 24030 623 24042 799
rect 23984 611 24042 623
rect 23834 423 23846 611
rect 23788 411 23846 423
rect 1082 -1939 1140 -1927
rect 1082 -2115 1094 -1939
rect 1128 -2115 1140 -1939
rect 1082 -2127 1140 -2115
rect 1200 -1939 1332 -1927
rect 1200 -2115 1212 -1939
rect 1246 -2115 1286 -1939
rect 1200 -2127 1286 -2115
rect 1274 -2315 1286 -2127
rect 1320 -2315 1332 -1939
rect 1274 -2327 1332 -2315
rect 1392 -1939 1450 -1927
rect 1392 -2315 1404 -1939
rect 1438 -2315 1450 -1939
rect 1392 -2327 1450 -2315
rect 1510 -1939 1568 -1927
rect 1510 -2315 1522 -1939
rect 1556 -2315 1568 -1939
rect 1510 -2327 1568 -2315
rect 1628 -1939 1686 -1927
rect 1628 -2315 1640 -1939
rect 1674 -2315 1686 -1939
rect 1628 -2327 1686 -2315
rect 1746 -1939 1882 -1927
rect 1746 -2315 1758 -1939
rect 1792 -2115 1836 -1939
rect 1870 -2115 1882 -1939
rect 1792 -2127 1882 -2115
rect 1942 -1939 2000 -1927
rect 1942 -2115 1954 -1939
rect 1988 -2115 2000 -1939
rect 1942 -2127 2000 -2115
rect 4226 -1939 4284 -1927
rect 4226 -2115 4238 -1939
rect 4272 -2115 4284 -1939
rect 4226 -2127 4284 -2115
rect 4344 -1939 4476 -1927
rect 4344 -2115 4356 -1939
rect 4390 -2115 4430 -1939
rect 4344 -2127 4430 -2115
rect 1792 -2315 1804 -2127
rect 1746 -2327 1804 -2315
rect 4418 -2315 4430 -2127
rect 4464 -2315 4476 -1939
rect 4418 -2327 4476 -2315
rect 4536 -1939 4594 -1927
rect 4536 -2315 4548 -1939
rect 4582 -2315 4594 -1939
rect 4536 -2327 4594 -2315
rect 4654 -1939 4712 -1927
rect 4654 -2315 4666 -1939
rect 4700 -2315 4712 -1939
rect 4654 -2327 4712 -2315
rect 4772 -1939 4830 -1927
rect 4772 -2315 4784 -1939
rect 4818 -2315 4830 -1939
rect 4772 -2327 4830 -2315
rect 4890 -1939 5026 -1927
rect 4890 -2315 4902 -1939
rect 4936 -2115 4980 -1939
rect 5014 -2115 5026 -1939
rect 4936 -2127 5026 -2115
rect 5086 -1939 5144 -1927
rect 5086 -2115 5098 -1939
rect 5132 -2115 5144 -1939
rect 5086 -2127 5144 -2115
rect 7358 -1935 7416 -1923
rect 7358 -2111 7370 -1935
rect 7404 -2111 7416 -1935
rect 7358 -2123 7416 -2111
rect 7476 -1935 7608 -1923
rect 7476 -2111 7488 -1935
rect 7522 -2111 7562 -1935
rect 7476 -2123 7562 -2111
rect 4936 -2315 4948 -2127
rect 4890 -2327 4948 -2315
rect 7550 -2311 7562 -2123
rect 7596 -2311 7608 -1935
rect 7550 -2323 7608 -2311
rect 7668 -1935 7726 -1923
rect 7668 -2311 7680 -1935
rect 7714 -2311 7726 -1935
rect 7668 -2323 7726 -2311
rect 7786 -1935 7844 -1923
rect 7786 -2311 7798 -1935
rect 7832 -2311 7844 -1935
rect 7786 -2323 7844 -2311
rect 7904 -1935 7962 -1923
rect 7904 -2311 7916 -1935
rect 7950 -2311 7962 -1935
rect 7904 -2323 7962 -2311
rect 8022 -1935 8158 -1923
rect 8022 -2311 8034 -1935
rect 8068 -2111 8112 -1935
rect 8146 -2111 8158 -1935
rect 8068 -2123 8158 -2111
rect 8218 -1935 8276 -1923
rect 8218 -2111 8230 -1935
rect 8264 -2111 8276 -1935
rect 8218 -2123 8276 -2111
rect 10502 -1935 10560 -1923
rect 10502 -2111 10514 -1935
rect 10548 -2111 10560 -1935
rect 10502 -2123 10560 -2111
rect 10620 -1935 10752 -1923
rect 10620 -2111 10632 -1935
rect 10666 -2111 10706 -1935
rect 10620 -2123 10706 -2111
rect 8068 -2311 8080 -2123
rect 8022 -2323 8080 -2311
rect 10694 -2311 10706 -2123
rect 10740 -2311 10752 -1935
rect 10694 -2323 10752 -2311
rect 10812 -1935 10870 -1923
rect 10812 -2311 10824 -1935
rect 10858 -2311 10870 -1935
rect 10812 -2323 10870 -2311
rect 10930 -1935 10988 -1923
rect 10930 -2311 10942 -1935
rect 10976 -2311 10988 -1935
rect 10930 -2323 10988 -2311
rect 11048 -1935 11106 -1923
rect 11048 -2311 11060 -1935
rect 11094 -2311 11106 -1935
rect 11048 -2323 11106 -2311
rect 11166 -1935 11302 -1923
rect 11166 -2311 11178 -1935
rect 11212 -2111 11256 -1935
rect 11290 -2111 11302 -1935
rect 11212 -2123 11302 -2111
rect 11362 -1935 11420 -1923
rect 11362 -2111 11374 -1935
rect 11408 -2111 11420 -1935
rect 11362 -2123 11420 -2111
rect 13704 -1939 13762 -1927
rect 13704 -2115 13716 -1939
rect 13750 -2115 13762 -1939
rect 11212 -2311 11224 -2123
rect 11166 -2323 11224 -2311
rect 13704 -2127 13762 -2115
rect 13822 -1939 13954 -1927
rect 13822 -2115 13834 -1939
rect 13868 -2115 13908 -1939
rect 13822 -2127 13908 -2115
rect 13896 -2315 13908 -2127
rect 13942 -2315 13954 -1939
rect 13896 -2327 13954 -2315
rect 14014 -1939 14072 -1927
rect 14014 -2315 14026 -1939
rect 14060 -2315 14072 -1939
rect 14014 -2327 14072 -2315
rect 14132 -1939 14190 -1927
rect 14132 -2315 14144 -1939
rect 14178 -2315 14190 -1939
rect 14132 -2327 14190 -2315
rect 14250 -1939 14308 -1927
rect 14250 -2315 14262 -1939
rect 14296 -2315 14308 -1939
rect 14250 -2327 14308 -2315
rect 14368 -1939 14504 -1927
rect 14368 -2315 14380 -1939
rect 14414 -2115 14458 -1939
rect 14492 -2115 14504 -1939
rect 14414 -2127 14504 -2115
rect 14564 -1939 14622 -1927
rect 14564 -2115 14576 -1939
rect 14610 -2115 14622 -1939
rect 14564 -2127 14622 -2115
rect 16848 -1939 16906 -1927
rect 16848 -2115 16860 -1939
rect 16894 -2115 16906 -1939
rect 16848 -2127 16906 -2115
rect 16966 -1939 17098 -1927
rect 16966 -2115 16978 -1939
rect 17012 -2115 17052 -1939
rect 16966 -2127 17052 -2115
rect 14414 -2315 14426 -2127
rect 14368 -2327 14426 -2315
rect 17040 -2315 17052 -2127
rect 17086 -2315 17098 -1939
rect 17040 -2327 17098 -2315
rect 17158 -1939 17216 -1927
rect 17158 -2315 17170 -1939
rect 17204 -2315 17216 -1939
rect 17158 -2327 17216 -2315
rect 17276 -1939 17334 -1927
rect 17276 -2315 17288 -1939
rect 17322 -2315 17334 -1939
rect 17276 -2327 17334 -2315
rect 17394 -1939 17452 -1927
rect 17394 -2315 17406 -1939
rect 17440 -2315 17452 -1939
rect 17394 -2327 17452 -2315
rect 17512 -1939 17648 -1927
rect 17512 -2315 17524 -1939
rect 17558 -2115 17602 -1939
rect 17636 -2115 17648 -1939
rect 17558 -2127 17648 -2115
rect 17708 -1939 17766 -1927
rect 17708 -2115 17720 -1939
rect 17754 -2115 17766 -1939
rect 17708 -2127 17766 -2115
rect 19980 -1935 20038 -1923
rect 19980 -2111 19992 -1935
rect 20026 -2111 20038 -1935
rect 19980 -2123 20038 -2111
rect 20098 -1935 20230 -1923
rect 20098 -2111 20110 -1935
rect 20144 -2111 20184 -1935
rect 20098 -2123 20184 -2111
rect 17558 -2315 17570 -2127
rect 17512 -2327 17570 -2315
rect 20172 -2311 20184 -2123
rect 20218 -2311 20230 -1935
rect 20172 -2323 20230 -2311
rect 20290 -1935 20348 -1923
rect 20290 -2311 20302 -1935
rect 20336 -2311 20348 -1935
rect 20290 -2323 20348 -2311
rect 20408 -1935 20466 -1923
rect 20408 -2311 20420 -1935
rect 20454 -2311 20466 -1935
rect 20408 -2323 20466 -2311
rect 20526 -1935 20584 -1923
rect 20526 -2311 20538 -1935
rect 20572 -2311 20584 -1935
rect 20526 -2323 20584 -2311
rect 20644 -1935 20780 -1923
rect 20644 -2311 20656 -1935
rect 20690 -2111 20734 -1935
rect 20768 -2111 20780 -1935
rect 20690 -2123 20780 -2111
rect 20840 -1935 20898 -1923
rect 20840 -2111 20852 -1935
rect 20886 -2111 20898 -1935
rect 20840 -2123 20898 -2111
rect 23124 -1935 23182 -1923
rect 23124 -2111 23136 -1935
rect 23170 -2111 23182 -1935
rect 23124 -2123 23182 -2111
rect 23242 -1935 23374 -1923
rect 23242 -2111 23254 -1935
rect 23288 -2111 23328 -1935
rect 23242 -2123 23328 -2111
rect 20690 -2311 20702 -2123
rect 20644 -2323 20702 -2311
rect 23316 -2311 23328 -2123
rect 23362 -2311 23374 -1935
rect 23316 -2323 23374 -2311
rect 23434 -1935 23492 -1923
rect 23434 -2311 23446 -1935
rect 23480 -2311 23492 -1935
rect 23434 -2323 23492 -2311
rect 23552 -1935 23610 -1923
rect 23552 -2311 23564 -1935
rect 23598 -2311 23610 -1935
rect 23552 -2323 23610 -2311
rect 23670 -1935 23728 -1923
rect 23670 -2311 23682 -1935
rect 23716 -2311 23728 -1935
rect 23670 -2323 23728 -2311
rect 23788 -1935 23924 -1923
rect 23788 -2311 23800 -1935
rect 23834 -2111 23878 -1935
rect 23912 -2111 23924 -1935
rect 23834 -2123 23924 -2111
rect 23984 -1935 24042 -1923
rect 23984 -2111 23996 -1935
rect 24030 -2111 24042 -1935
rect 23984 -2123 24042 -2111
rect 23834 -2311 23846 -2123
rect 23788 -2323 23846 -2311
rect 1072 -4671 1130 -4659
rect 1072 -4847 1084 -4671
rect 1118 -4847 1130 -4671
rect 1072 -4859 1130 -4847
rect 1190 -4671 1322 -4659
rect 1190 -4847 1202 -4671
rect 1236 -4847 1276 -4671
rect 1190 -4859 1276 -4847
rect 1264 -5047 1276 -4859
rect 1310 -5047 1322 -4671
rect 1264 -5059 1322 -5047
rect 1382 -4671 1440 -4659
rect 1382 -5047 1394 -4671
rect 1428 -5047 1440 -4671
rect 1382 -5059 1440 -5047
rect 1500 -4671 1558 -4659
rect 1500 -5047 1512 -4671
rect 1546 -5047 1558 -4671
rect 1500 -5059 1558 -5047
rect 1618 -4671 1676 -4659
rect 1618 -5047 1630 -4671
rect 1664 -5047 1676 -4671
rect 1618 -5059 1676 -5047
rect 1736 -4671 1872 -4659
rect 1736 -5047 1748 -4671
rect 1782 -4847 1826 -4671
rect 1860 -4847 1872 -4671
rect 1782 -4859 1872 -4847
rect 1932 -4671 1990 -4659
rect 1932 -4847 1944 -4671
rect 1978 -4847 1990 -4671
rect 1932 -4859 1990 -4847
rect 4216 -4671 4274 -4659
rect 4216 -4847 4228 -4671
rect 4262 -4847 4274 -4671
rect 4216 -4859 4274 -4847
rect 4334 -4671 4466 -4659
rect 4334 -4847 4346 -4671
rect 4380 -4847 4420 -4671
rect 4334 -4859 4420 -4847
rect 1782 -5047 1794 -4859
rect 1736 -5059 1794 -5047
rect 4408 -5047 4420 -4859
rect 4454 -5047 4466 -4671
rect 4408 -5059 4466 -5047
rect 4526 -4671 4584 -4659
rect 4526 -5047 4538 -4671
rect 4572 -5047 4584 -4671
rect 4526 -5059 4584 -5047
rect 4644 -4671 4702 -4659
rect 4644 -5047 4656 -4671
rect 4690 -5047 4702 -4671
rect 4644 -5059 4702 -5047
rect 4762 -4671 4820 -4659
rect 4762 -5047 4774 -4671
rect 4808 -5047 4820 -4671
rect 4762 -5059 4820 -5047
rect 4880 -4671 5016 -4659
rect 4880 -5047 4892 -4671
rect 4926 -4847 4970 -4671
rect 5004 -4847 5016 -4671
rect 4926 -4859 5016 -4847
rect 5076 -4671 5134 -4659
rect 5076 -4847 5088 -4671
rect 5122 -4847 5134 -4671
rect 5076 -4859 5134 -4847
rect 7348 -4667 7406 -4655
rect 7348 -4843 7360 -4667
rect 7394 -4843 7406 -4667
rect 7348 -4855 7406 -4843
rect 7466 -4667 7598 -4655
rect 7466 -4843 7478 -4667
rect 7512 -4843 7552 -4667
rect 7466 -4855 7552 -4843
rect 4926 -5047 4938 -4859
rect 4880 -5059 4938 -5047
rect 7540 -5043 7552 -4855
rect 7586 -5043 7598 -4667
rect 7540 -5055 7598 -5043
rect 7658 -4667 7716 -4655
rect 7658 -5043 7670 -4667
rect 7704 -5043 7716 -4667
rect 7658 -5055 7716 -5043
rect 7776 -4667 7834 -4655
rect 7776 -5043 7788 -4667
rect 7822 -5043 7834 -4667
rect 7776 -5055 7834 -5043
rect 7894 -4667 7952 -4655
rect 7894 -5043 7906 -4667
rect 7940 -5043 7952 -4667
rect 7894 -5055 7952 -5043
rect 8012 -4667 8148 -4655
rect 8012 -5043 8024 -4667
rect 8058 -4843 8102 -4667
rect 8136 -4843 8148 -4667
rect 8058 -4855 8148 -4843
rect 8208 -4667 8266 -4655
rect 8208 -4843 8220 -4667
rect 8254 -4843 8266 -4667
rect 8208 -4855 8266 -4843
rect 10492 -4667 10550 -4655
rect 10492 -4843 10504 -4667
rect 10538 -4843 10550 -4667
rect 10492 -4855 10550 -4843
rect 10610 -4667 10742 -4655
rect 10610 -4843 10622 -4667
rect 10656 -4843 10696 -4667
rect 10610 -4855 10696 -4843
rect 8058 -5043 8070 -4855
rect 8012 -5055 8070 -5043
rect 10684 -5043 10696 -4855
rect 10730 -5043 10742 -4667
rect 10684 -5055 10742 -5043
rect 10802 -4667 10860 -4655
rect 10802 -5043 10814 -4667
rect 10848 -5043 10860 -4667
rect 10802 -5055 10860 -5043
rect 10920 -4667 10978 -4655
rect 10920 -5043 10932 -4667
rect 10966 -5043 10978 -4667
rect 10920 -5055 10978 -5043
rect 11038 -4667 11096 -4655
rect 11038 -5043 11050 -4667
rect 11084 -5043 11096 -4667
rect 11038 -5055 11096 -5043
rect 11156 -4667 11292 -4655
rect 11156 -5043 11168 -4667
rect 11202 -4843 11246 -4667
rect 11280 -4843 11292 -4667
rect 11202 -4855 11292 -4843
rect 11352 -4667 11410 -4655
rect 11352 -4843 11364 -4667
rect 11398 -4843 11410 -4667
rect 11352 -4855 11410 -4843
rect 13694 -4671 13752 -4659
rect 13694 -4847 13706 -4671
rect 13740 -4847 13752 -4671
rect 11202 -5043 11214 -4855
rect 11156 -5055 11214 -5043
rect 13694 -4859 13752 -4847
rect 13812 -4671 13944 -4659
rect 13812 -4847 13824 -4671
rect 13858 -4847 13898 -4671
rect 13812 -4859 13898 -4847
rect 13886 -5047 13898 -4859
rect 13932 -5047 13944 -4671
rect 13886 -5059 13944 -5047
rect 14004 -4671 14062 -4659
rect 14004 -5047 14016 -4671
rect 14050 -5047 14062 -4671
rect 14004 -5059 14062 -5047
rect 14122 -4671 14180 -4659
rect 14122 -5047 14134 -4671
rect 14168 -5047 14180 -4671
rect 14122 -5059 14180 -5047
rect 14240 -4671 14298 -4659
rect 14240 -5047 14252 -4671
rect 14286 -5047 14298 -4671
rect 14240 -5059 14298 -5047
rect 14358 -4671 14494 -4659
rect 14358 -5047 14370 -4671
rect 14404 -4847 14448 -4671
rect 14482 -4847 14494 -4671
rect 14404 -4859 14494 -4847
rect 14554 -4671 14612 -4659
rect 14554 -4847 14566 -4671
rect 14600 -4847 14612 -4671
rect 14554 -4859 14612 -4847
rect 16838 -4671 16896 -4659
rect 16838 -4847 16850 -4671
rect 16884 -4847 16896 -4671
rect 16838 -4859 16896 -4847
rect 16956 -4671 17088 -4659
rect 16956 -4847 16968 -4671
rect 17002 -4847 17042 -4671
rect 16956 -4859 17042 -4847
rect 14404 -5047 14416 -4859
rect 14358 -5059 14416 -5047
rect 17030 -5047 17042 -4859
rect 17076 -5047 17088 -4671
rect 17030 -5059 17088 -5047
rect 17148 -4671 17206 -4659
rect 17148 -5047 17160 -4671
rect 17194 -5047 17206 -4671
rect 17148 -5059 17206 -5047
rect 17266 -4671 17324 -4659
rect 17266 -5047 17278 -4671
rect 17312 -5047 17324 -4671
rect 17266 -5059 17324 -5047
rect 17384 -4671 17442 -4659
rect 17384 -5047 17396 -4671
rect 17430 -5047 17442 -4671
rect 17384 -5059 17442 -5047
rect 17502 -4671 17638 -4659
rect 17502 -5047 17514 -4671
rect 17548 -4847 17592 -4671
rect 17626 -4847 17638 -4671
rect 17548 -4859 17638 -4847
rect 17698 -4671 17756 -4659
rect 17698 -4847 17710 -4671
rect 17744 -4847 17756 -4671
rect 17698 -4859 17756 -4847
rect 19970 -4667 20028 -4655
rect 19970 -4843 19982 -4667
rect 20016 -4843 20028 -4667
rect 19970 -4855 20028 -4843
rect 20088 -4667 20220 -4655
rect 20088 -4843 20100 -4667
rect 20134 -4843 20174 -4667
rect 20088 -4855 20174 -4843
rect 17548 -5047 17560 -4859
rect 17502 -5059 17560 -5047
rect 20162 -5043 20174 -4855
rect 20208 -5043 20220 -4667
rect 20162 -5055 20220 -5043
rect 20280 -4667 20338 -4655
rect 20280 -5043 20292 -4667
rect 20326 -5043 20338 -4667
rect 20280 -5055 20338 -5043
rect 20398 -4667 20456 -4655
rect 20398 -5043 20410 -4667
rect 20444 -5043 20456 -4667
rect 20398 -5055 20456 -5043
rect 20516 -4667 20574 -4655
rect 20516 -5043 20528 -4667
rect 20562 -5043 20574 -4667
rect 20516 -5055 20574 -5043
rect 20634 -4667 20770 -4655
rect 20634 -5043 20646 -4667
rect 20680 -4843 20724 -4667
rect 20758 -4843 20770 -4667
rect 20680 -4855 20770 -4843
rect 20830 -4667 20888 -4655
rect 20830 -4843 20842 -4667
rect 20876 -4843 20888 -4667
rect 20830 -4855 20888 -4843
rect 23114 -4667 23172 -4655
rect 23114 -4843 23126 -4667
rect 23160 -4843 23172 -4667
rect 23114 -4855 23172 -4843
rect 23232 -4667 23364 -4655
rect 23232 -4843 23244 -4667
rect 23278 -4843 23318 -4667
rect 23232 -4855 23318 -4843
rect 20680 -5043 20692 -4855
rect 20634 -5055 20692 -5043
rect 23306 -5043 23318 -4855
rect 23352 -5043 23364 -4667
rect 23306 -5055 23364 -5043
rect 23424 -4667 23482 -4655
rect 23424 -5043 23436 -4667
rect 23470 -5043 23482 -4667
rect 23424 -5055 23482 -5043
rect 23542 -4667 23600 -4655
rect 23542 -5043 23554 -4667
rect 23588 -5043 23600 -4667
rect 23542 -5055 23600 -5043
rect 23660 -4667 23718 -4655
rect 23660 -5043 23672 -4667
rect 23706 -5043 23718 -4667
rect 23660 -5055 23718 -5043
rect 23778 -4667 23914 -4655
rect 23778 -5043 23790 -4667
rect 23824 -4843 23868 -4667
rect 23902 -4843 23914 -4667
rect 23824 -4855 23914 -4843
rect 23974 -4667 24032 -4655
rect 23974 -4843 23986 -4667
rect 24020 -4843 24032 -4667
rect 23974 -4855 24032 -4843
rect 23824 -5043 23836 -4855
rect 23778 -5055 23836 -5043
rect 100 -7708 158 -7696
rect 100 -7884 112 -7708
rect 146 -7884 158 -7708
rect 100 -7896 158 -7884
rect 218 -7708 276 -7696
rect 218 -7884 230 -7708
rect 264 -7884 276 -7708
rect 218 -7896 276 -7884
rect 520 -7708 578 -7696
rect 520 -8084 532 -7708
rect 566 -8084 578 -7708
rect 520 -8096 578 -8084
rect 638 -7708 696 -7696
rect 638 -8084 650 -7708
rect 684 -8084 696 -7708
rect 638 -8096 696 -8084
rect 756 -7708 814 -7696
rect 756 -8084 768 -7708
rect 802 -8084 814 -7708
rect 756 -8096 814 -8084
rect 874 -7708 932 -7696
rect 874 -8084 886 -7708
rect 920 -8084 932 -7708
rect 874 -8096 932 -8084
rect 992 -7708 1050 -7696
rect 992 -8084 1004 -7708
rect 1038 -8084 1050 -7708
rect 1398 -7708 1456 -7696
rect 1398 -7884 1410 -7708
rect 1444 -7884 1456 -7708
rect 1398 -7896 1456 -7884
rect 1516 -7708 1574 -7696
rect 1516 -7884 1528 -7708
rect 1562 -7884 1574 -7708
rect 1516 -7896 1574 -7884
rect 2168 -7706 2226 -7694
rect 2168 -7882 2180 -7706
rect 2214 -7882 2226 -7706
rect 2168 -7894 2226 -7882
rect 2286 -7706 2344 -7694
rect 2286 -7882 2298 -7706
rect 2332 -7882 2344 -7706
rect 2286 -7894 2344 -7882
rect 2588 -7706 2646 -7694
rect 992 -8096 1050 -8084
rect 2588 -8082 2600 -7706
rect 2634 -8082 2646 -7706
rect 2588 -8094 2646 -8082
rect 2706 -7706 2764 -7694
rect 2706 -8082 2718 -7706
rect 2752 -8082 2764 -7706
rect 2706 -8094 2764 -8082
rect 2824 -7706 2882 -7694
rect 2824 -8082 2836 -7706
rect 2870 -8082 2882 -7706
rect 2824 -8094 2882 -8082
rect 2942 -7706 3000 -7694
rect 2942 -8082 2954 -7706
rect 2988 -8082 3000 -7706
rect 2942 -8094 3000 -8082
rect 3060 -7706 3118 -7694
rect 3060 -8082 3072 -7706
rect 3106 -8082 3118 -7706
rect 3466 -7706 3524 -7694
rect 3466 -7882 3478 -7706
rect 3512 -7882 3524 -7706
rect 3466 -7894 3524 -7882
rect 3584 -7706 3642 -7694
rect 16825 -6553 16883 -6541
rect 3584 -7882 3596 -7706
rect 3630 -7882 3642 -7706
rect 3584 -7894 3642 -7882
rect 4237 -7708 4295 -7696
rect 4237 -7884 4249 -7708
rect 4283 -7884 4295 -7708
rect 4237 -7896 4295 -7884
rect 4355 -7708 4413 -7696
rect 4355 -7884 4367 -7708
rect 4401 -7884 4413 -7708
rect 4355 -7896 4413 -7884
rect 4657 -7708 4715 -7696
rect 3060 -8094 3118 -8082
rect 4657 -8084 4669 -7708
rect 4703 -8084 4715 -7708
rect 4657 -8096 4715 -8084
rect 4775 -7708 4833 -7696
rect 4775 -8084 4787 -7708
rect 4821 -8084 4833 -7708
rect 4775 -8096 4833 -8084
rect 4893 -7708 4951 -7696
rect 4893 -8084 4905 -7708
rect 4939 -8084 4951 -7708
rect 4893 -8096 4951 -8084
rect 5011 -7708 5069 -7696
rect 5011 -8084 5023 -7708
rect 5057 -8084 5069 -7708
rect 5011 -8096 5069 -8084
rect 5129 -7708 5187 -7696
rect 5129 -8084 5141 -7708
rect 5175 -8084 5187 -7708
rect 5535 -7708 5593 -7696
rect 5535 -7884 5547 -7708
rect 5581 -7884 5593 -7708
rect 5535 -7896 5593 -7884
rect 5653 -7708 5711 -7696
rect 5653 -7884 5665 -7708
rect 5699 -7884 5711 -7708
rect 5653 -7896 5711 -7884
rect 6305 -7706 6363 -7694
rect 6305 -7882 6317 -7706
rect 6351 -7882 6363 -7706
rect 6305 -7894 6363 -7882
rect 6423 -7706 6481 -7694
rect 6423 -7882 6435 -7706
rect 6469 -7882 6481 -7706
rect 6423 -7894 6481 -7882
rect 6725 -7706 6783 -7694
rect 5129 -8096 5187 -8084
rect 6725 -8082 6737 -7706
rect 6771 -8082 6783 -7706
rect 6725 -8094 6783 -8082
rect 6843 -7706 6901 -7694
rect 6843 -8082 6855 -7706
rect 6889 -8082 6901 -7706
rect 6843 -8094 6901 -8082
rect 6961 -7706 7019 -7694
rect 6961 -8082 6973 -7706
rect 7007 -8082 7019 -7706
rect 6961 -8094 7019 -8082
rect 7079 -7706 7137 -7694
rect 7079 -8082 7091 -7706
rect 7125 -8082 7137 -7706
rect 7079 -8094 7137 -8082
rect 7197 -7706 7255 -7694
rect 7197 -8082 7209 -7706
rect 7243 -8082 7255 -7706
rect 7603 -7706 7661 -7694
rect 7603 -7882 7615 -7706
rect 7649 -7882 7661 -7706
rect 7603 -7894 7661 -7882
rect 7721 -7706 7779 -7694
rect 7721 -7882 7733 -7706
rect 7767 -7882 7779 -7706
rect 7721 -7894 7779 -7882
rect 8374 -7706 8432 -7694
rect 8374 -7882 8386 -7706
rect 8420 -7882 8432 -7706
rect 8374 -7894 8432 -7882
rect 8492 -7706 8550 -7694
rect 8492 -7882 8504 -7706
rect 8538 -7882 8550 -7706
rect 8492 -7894 8550 -7882
rect 8794 -7706 8852 -7694
rect 7197 -8094 7255 -8082
rect 8794 -8082 8806 -7706
rect 8840 -8082 8852 -7706
rect 8794 -8094 8852 -8082
rect 8912 -7706 8970 -7694
rect 8912 -8082 8924 -7706
rect 8958 -8082 8970 -7706
rect 8912 -8094 8970 -8082
rect 9030 -7706 9088 -7694
rect 9030 -8082 9042 -7706
rect 9076 -8082 9088 -7706
rect 9030 -8094 9088 -8082
rect 9148 -7706 9206 -7694
rect 9148 -8082 9160 -7706
rect 9194 -8082 9206 -7706
rect 9148 -8094 9206 -8082
rect 9266 -7706 9324 -7694
rect 9266 -8082 9278 -7706
rect 9312 -8082 9324 -7706
rect 9672 -7706 9730 -7694
rect 9672 -7882 9684 -7706
rect 9718 -7882 9730 -7706
rect 9672 -7894 9730 -7882
rect 9790 -7706 9848 -7694
rect 9790 -7882 9802 -7706
rect 9836 -7882 9848 -7706
rect 9790 -7894 9848 -7882
rect 10442 -7704 10500 -7692
rect 10442 -7880 10454 -7704
rect 10488 -7880 10500 -7704
rect 10442 -7892 10500 -7880
rect 10560 -7704 10618 -7692
rect 10560 -7880 10572 -7704
rect 10606 -7880 10618 -7704
rect 10560 -7892 10618 -7880
rect 10862 -7704 10920 -7692
rect 9266 -8094 9324 -8082
rect 10862 -8080 10874 -7704
rect 10908 -8080 10920 -7704
rect 10862 -8092 10920 -8080
rect 10980 -7704 11038 -7692
rect 10980 -8080 10992 -7704
rect 11026 -8080 11038 -7704
rect 10980 -8092 11038 -8080
rect 11098 -7704 11156 -7692
rect 11098 -8080 11110 -7704
rect 11144 -8080 11156 -7704
rect 11098 -8092 11156 -8080
rect 11216 -7704 11274 -7692
rect 11216 -8080 11228 -7704
rect 11262 -8080 11274 -7704
rect 11216 -8092 11274 -8080
rect 11334 -7704 11392 -7692
rect 11334 -8080 11346 -7704
rect 11380 -8080 11392 -7704
rect 11740 -7704 11798 -7692
rect 11740 -7880 11752 -7704
rect 11786 -7880 11798 -7704
rect 11740 -7892 11798 -7880
rect 11858 -7704 11916 -7692
rect 16825 -6729 16837 -6553
rect 16871 -6729 16883 -6553
rect 16825 -6741 16883 -6729
rect 16943 -6553 17001 -6541
rect 16943 -6729 16955 -6553
rect 16989 -6729 17001 -6553
rect 16943 -6741 17001 -6729
rect 17563 -6551 17621 -6539
rect 17563 -6727 17575 -6551
rect 17609 -6727 17621 -6551
rect 17563 -6739 17621 -6727
rect 17681 -6551 17739 -6539
rect 17681 -6727 17693 -6551
rect 17727 -6727 17739 -6551
rect 17681 -6739 17739 -6727
rect 18301 -6555 18359 -6543
rect 18301 -6731 18313 -6555
rect 18347 -6731 18359 -6555
rect 18301 -6743 18359 -6731
rect 18419 -6555 18477 -6543
rect 18419 -6731 18431 -6555
rect 18465 -6731 18477 -6555
rect 18419 -6743 18477 -6731
rect 19043 -6555 19101 -6543
rect 19043 -6731 19055 -6555
rect 19089 -6731 19101 -6555
rect 19043 -6743 19101 -6731
rect 19161 -6555 19219 -6543
rect 19161 -6731 19173 -6555
rect 19207 -6731 19219 -6555
rect 19161 -6743 19219 -6731
rect 19783 -6555 19841 -6543
rect 19783 -6731 19795 -6555
rect 19829 -6731 19841 -6555
rect 19783 -6743 19841 -6731
rect 19901 -6555 19959 -6543
rect 19901 -6731 19913 -6555
rect 19947 -6731 19959 -6555
rect 19901 -6743 19959 -6731
rect 20521 -6555 20579 -6543
rect 20521 -6731 20533 -6555
rect 20567 -6731 20579 -6555
rect 20521 -6743 20579 -6731
rect 20639 -6555 20697 -6543
rect 20639 -6731 20651 -6555
rect 20685 -6731 20697 -6555
rect 20639 -6743 20697 -6731
rect 21259 -6551 21317 -6539
rect 21259 -6727 21271 -6551
rect 21305 -6727 21317 -6551
rect 21259 -6739 21317 -6727
rect 21377 -6551 21435 -6539
rect 21377 -6727 21389 -6551
rect 21423 -6727 21435 -6551
rect 21377 -6739 21435 -6727
rect 21997 -6551 22055 -6539
rect 21997 -6727 22009 -6551
rect 22043 -6727 22055 -6551
rect 21997 -6739 22055 -6727
rect 22115 -6551 22173 -6539
rect 22115 -6727 22127 -6551
rect 22161 -6727 22173 -6551
rect 22115 -6739 22173 -6727
rect 11858 -7880 11870 -7704
rect 11904 -7880 11916 -7704
rect 11858 -7892 11916 -7880
rect 12511 -7706 12569 -7694
rect 12511 -7882 12523 -7706
rect 12557 -7882 12569 -7706
rect 12511 -7894 12569 -7882
rect 12629 -7706 12687 -7694
rect 12629 -7882 12641 -7706
rect 12675 -7882 12687 -7706
rect 12629 -7894 12687 -7882
rect 12931 -7706 12989 -7694
rect 11334 -8092 11392 -8080
rect 12931 -8082 12943 -7706
rect 12977 -8082 12989 -7706
rect 12931 -8094 12989 -8082
rect 13049 -7706 13107 -7694
rect 13049 -8082 13061 -7706
rect 13095 -8082 13107 -7706
rect 13049 -8094 13107 -8082
rect 13167 -7706 13225 -7694
rect 13167 -8082 13179 -7706
rect 13213 -8082 13225 -7706
rect 13167 -8094 13225 -8082
rect 13285 -7706 13343 -7694
rect 13285 -8082 13297 -7706
rect 13331 -8082 13343 -7706
rect 13285 -8094 13343 -8082
rect 13403 -7706 13461 -7694
rect 13403 -8082 13415 -7706
rect 13449 -8082 13461 -7706
rect 13809 -7706 13867 -7694
rect 13809 -7882 13821 -7706
rect 13855 -7882 13867 -7706
rect 13809 -7894 13867 -7882
rect 13927 -7706 13985 -7694
rect 13927 -7882 13939 -7706
rect 13973 -7882 13985 -7706
rect 13927 -7894 13985 -7882
rect 14579 -7704 14637 -7692
rect 14579 -7880 14591 -7704
rect 14625 -7880 14637 -7704
rect 14579 -7892 14637 -7880
rect 14697 -7704 14755 -7692
rect 14697 -7880 14709 -7704
rect 14743 -7880 14755 -7704
rect 14697 -7892 14755 -7880
rect 14999 -7704 15057 -7692
rect 13403 -8094 13461 -8082
rect 14999 -8080 15011 -7704
rect 15045 -8080 15057 -7704
rect 14999 -8092 15057 -8080
rect 15117 -7704 15175 -7692
rect 15117 -8080 15129 -7704
rect 15163 -8080 15175 -7704
rect 15117 -8092 15175 -8080
rect 15235 -7704 15293 -7692
rect 15235 -8080 15247 -7704
rect 15281 -8080 15293 -7704
rect 15235 -8092 15293 -8080
rect 15353 -7704 15411 -7692
rect 15353 -8080 15365 -7704
rect 15399 -8080 15411 -7704
rect 15353 -8092 15411 -8080
rect 15471 -7704 15529 -7692
rect 15471 -8080 15483 -7704
rect 15517 -8080 15529 -7704
rect 15877 -7704 15935 -7692
rect 15877 -7880 15889 -7704
rect 15923 -7880 15935 -7704
rect 15877 -7892 15935 -7880
rect 15995 -7704 16053 -7692
rect 15995 -7880 16007 -7704
rect 16041 -7880 16053 -7704
rect 15995 -7892 16053 -7880
rect 15471 -8092 15529 -8080
<< pdiff >>
rect 11952 4082 12010 4094
rect 189 3885 247 3897
rect 189 3709 201 3885
rect 235 3709 247 3885
rect 189 3697 247 3709
rect 307 3885 365 3897
rect 307 3709 319 3885
rect 353 3709 365 3885
rect 307 3697 365 3709
rect 425 3885 483 3897
rect 425 3709 437 3885
rect 471 3709 483 3885
rect 425 3697 483 3709
rect 543 3885 601 3897
rect 543 3709 555 3885
rect 589 3709 601 3885
rect 543 3697 601 3709
rect 661 3885 719 3897
rect 661 3709 673 3885
rect 707 3709 719 3885
rect 661 3697 719 3709
rect 779 3885 837 3897
rect 779 3709 791 3885
rect 825 3709 837 3885
rect 779 3697 837 3709
rect 897 3885 955 3897
rect 897 3709 909 3885
rect 943 3709 955 3885
rect 897 3697 955 3709
rect 1015 3885 1073 3897
rect 1015 3709 1027 3885
rect 1061 3709 1073 3885
rect 1015 3697 1073 3709
rect 1133 3885 1191 3897
rect 1133 3709 1145 3885
rect 1179 3709 1191 3885
rect 1133 3697 1191 3709
rect 1251 3885 1309 3897
rect 1251 3709 1263 3885
rect 1297 3709 1309 3885
rect 1251 3697 1309 3709
rect 1637 3885 1695 3897
rect 1637 3709 1649 3885
rect 1683 3709 1695 3885
rect 1637 3697 1695 3709
rect 1755 3885 1813 3897
rect 1755 3709 1767 3885
rect 1801 3709 1813 3885
rect 1755 3697 1813 3709
rect 1873 3885 1931 3897
rect 1873 3709 1885 3885
rect 1919 3709 1931 3885
rect 1873 3697 1931 3709
rect 1991 3885 2049 3897
rect 1991 3709 2003 3885
rect 2037 3709 2049 3885
rect 1991 3697 2049 3709
rect 2109 3885 2167 3897
rect 2109 3709 2121 3885
rect 2155 3709 2167 3885
rect 2109 3697 2167 3709
rect 2227 3885 2285 3897
rect 2227 3709 2239 3885
rect 2273 3709 2285 3885
rect 2227 3697 2285 3709
rect 2345 3885 2403 3897
rect 2345 3709 2357 3885
rect 2391 3709 2403 3885
rect 2345 3697 2403 3709
rect 2463 3885 2521 3897
rect 2463 3709 2475 3885
rect 2509 3709 2521 3885
rect 2463 3697 2521 3709
rect 2581 3885 2639 3897
rect 2581 3709 2593 3885
rect 2627 3709 2639 3885
rect 2581 3697 2639 3709
rect 2699 3885 2757 3897
rect 2699 3709 2711 3885
rect 2745 3709 2757 3885
rect 2699 3697 2757 3709
rect 3135 3887 3193 3899
rect 3135 3711 3147 3887
rect 3181 3711 3193 3887
rect 3135 3699 3193 3711
rect 3253 3887 3311 3899
rect 3253 3711 3265 3887
rect 3299 3711 3311 3887
rect 3253 3699 3311 3711
rect 3371 3887 3429 3899
rect 3371 3711 3383 3887
rect 3417 3711 3429 3887
rect 3371 3699 3429 3711
rect 3489 3887 3547 3899
rect 3489 3711 3501 3887
rect 3535 3711 3547 3887
rect 3489 3699 3547 3711
rect 3607 3887 3665 3899
rect 3607 3711 3619 3887
rect 3653 3711 3665 3887
rect 3607 3699 3665 3711
rect 3725 3887 3783 3899
rect 3725 3711 3737 3887
rect 3771 3711 3783 3887
rect 3725 3699 3783 3711
rect 3843 3887 3901 3899
rect 3843 3711 3855 3887
rect 3889 3711 3901 3887
rect 3843 3699 3901 3711
rect 3961 3887 4019 3899
rect 3961 3711 3973 3887
rect 4007 3711 4019 3887
rect 3961 3699 4019 3711
rect 4079 3887 4137 3899
rect 4079 3711 4091 3887
rect 4125 3711 4137 3887
rect 4079 3699 4137 3711
rect 4197 3887 4255 3899
rect 4197 3711 4209 3887
rect 4243 3711 4255 3887
rect 4197 3699 4255 3711
rect 4583 3887 4641 3899
rect 4583 3711 4595 3887
rect 4629 3711 4641 3887
rect 4583 3699 4641 3711
rect 4701 3887 4759 3899
rect 4701 3711 4713 3887
rect 4747 3711 4759 3887
rect 4701 3699 4759 3711
rect 4819 3887 4877 3899
rect 4819 3711 4831 3887
rect 4865 3711 4877 3887
rect 4819 3699 4877 3711
rect 4937 3887 4995 3899
rect 4937 3711 4949 3887
rect 4983 3711 4995 3887
rect 4937 3699 4995 3711
rect 5055 3887 5113 3899
rect 5055 3711 5067 3887
rect 5101 3711 5113 3887
rect 5055 3699 5113 3711
rect 5173 3887 5231 3899
rect 5173 3711 5185 3887
rect 5219 3711 5231 3887
rect 5173 3699 5231 3711
rect 5291 3887 5349 3899
rect 5291 3711 5303 3887
rect 5337 3711 5349 3887
rect 5291 3699 5349 3711
rect 5409 3887 5467 3899
rect 5409 3711 5421 3887
rect 5455 3711 5467 3887
rect 5409 3699 5467 3711
rect 5527 3887 5585 3899
rect 5527 3711 5539 3887
rect 5573 3711 5585 3887
rect 5527 3699 5585 3711
rect 5645 3887 5703 3899
rect 5645 3711 5657 3887
rect 5691 3711 5703 3887
rect 5645 3699 5703 3711
rect 6103 3885 6161 3897
rect 6103 3709 6115 3885
rect 6149 3709 6161 3885
rect 6103 3697 6161 3709
rect 6221 3885 6279 3897
rect 6221 3709 6233 3885
rect 6267 3709 6279 3885
rect 6221 3697 6279 3709
rect 6339 3885 6397 3897
rect 6339 3709 6351 3885
rect 6385 3709 6397 3885
rect 6339 3697 6397 3709
rect 6457 3885 6515 3897
rect 6457 3709 6469 3885
rect 6503 3709 6515 3885
rect 6457 3697 6515 3709
rect 6575 3885 6633 3897
rect 6575 3709 6587 3885
rect 6621 3709 6633 3885
rect 6575 3697 6633 3709
rect 6693 3885 6751 3897
rect 6693 3709 6705 3885
rect 6739 3709 6751 3885
rect 6693 3697 6751 3709
rect 6811 3885 6869 3897
rect 6811 3709 6823 3885
rect 6857 3709 6869 3885
rect 6811 3697 6869 3709
rect 6929 3885 6987 3897
rect 6929 3709 6941 3885
rect 6975 3709 6987 3885
rect 6929 3697 6987 3709
rect 7047 3885 7105 3897
rect 7047 3709 7059 3885
rect 7093 3709 7105 3885
rect 7047 3697 7105 3709
rect 7165 3885 7223 3897
rect 7165 3709 7177 3885
rect 7211 3709 7223 3885
rect 7165 3697 7223 3709
rect 7551 3885 7609 3897
rect 7551 3709 7563 3885
rect 7597 3709 7609 3885
rect 7551 3697 7609 3709
rect 7669 3885 7727 3897
rect 7669 3709 7681 3885
rect 7715 3709 7727 3885
rect 7669 3697 7727 3709
rect 7787 3885 7845 3897
rect 7787 3709 7799 3885
rect 7833 3709 7845 3885
rect 7787 3697 7845 3709
rect 7905 3885 7963 3897
rect 7905 3709 7917 3885
rect 7951 3709 7963 3885
rect 7905 3697 7963 3709
rect 8023 3885 8081 3897
rect 8023 3709 8035 3885
rect 8069 3709 8081 3885
rect 8023 3697 8081 3709
rect 8141 3885 8199 3897
rect 8141 3709 8153 3885
rect 8187 3709 8199 3885
rect 8141 3697 8199 3709
rect 8259 3885 8317 3897
rect 8259 3709 8271 3885
rect 8305 3709 8317 3885
rect 8259 3697 8317 3709
rect 8377 3885 8435 3897
rect 8377 3709 8389 3885
rect 8423 3709 8435 3885
rect 8377 3697 8435 3709
rect 8495 3885 8553 3897
rect 8495 3709 8507 3885
rect 8541 3709 8553 3885
rect 8495 3697 8553 3709
rect 8613 3885 8671 3897
rect 8613 3709 8625 3885
rect 8659 3709 8671 3885
rect 8613 3697 8671 3709
rect 9049 3887 9107 3899
rect 9049 3711 9061 3887
rect 9095 3711 9107 3887
rect 9049 3699 9107 3711
rect 9167 3887 9225 3899
rect 9167 3711 9179 3887
rect 9213 3711 9225 3887
rect 9167 3699 9225 3711
rect 9285 3887 9343 3899
rect 9285 3711 9297 3887
rect 9331 3711 9343 3887
rect 9285 3699 9343 3711
rect 9403 3887 9461 3899
rect 9403 3711 9415 3887
rect 9449 3711 9461 3887
rect 9403 3699 9461 3711
rect 9521 3887 9579 3899
rect 9521 3711 9533 3887
rect 9567 3711 9579 3887
rect 9521 3699 9579 3711
rect 9639 3887 9697 3899
rect 9639 3711 9651 3887
rect 9685 3711 9697 3887
rect 9639 3699 9697 3711
rect 9757 3887 9815 3899
rect 9757 3711 9769 3887
rect 9803 3711 9815 3887
rect 9757 3699 9815 3711
rect 9875 3887 9933 3899
rect 9875 3711 9887 3887
rect 9921 3711 9933 3887
rect 9875 3699 9933 3711
rect 9993 3887 10051 3899
rect 9993 3711 10005 3887
rect 10039 3711 10051 3887
rect 9993 3699 10051 3711
rect 10111 3887 10169 3899
rect 10111 3711 10123 3887
rect 10157 3711 10169 3887
rect 10111 3699 10169 3711
rect 10497 3887 10555 3899
rect 10497 3711 10509 3887
rect 10543 3711 10555 3887
rect 10497 3699 10555 3711
rect 10615 3887 10673 3899
rect 10615 3711 10627 3887
rect 10661 3711 10673 3887
rect 10615 3699 10673 3711
rect 10733 3887 10791 3899
rect 10733 3711 10745 3887
rect 10779 3711 10791 3887
rect 10733 3699 10791 3711
rect 10851 3887 10909 3899
rect 10851 3711 10863 3887
rect 10897 3711 10909 3887
rect 10851 3699 10909 3711
rect 10969 3887 11027 3899
rect 10969 3711 10981 3887
rect 11015 3711 11027 3887
rect 10969 3699 11027 3711
rect 11087 3887 11145 3899
rect 11087 3711 11099 3887
rect 11133 3711 11145 3887
rect 11087 3699 11145 3711
rect 11205 3887 11263 3899
rect 11205 3711 11217 3887
rect 11251 3711 11263 3887
rect 11205 3699 11263 3711
rect 11323 3887 11381 3899
rect 11323 3711 11335 3887
rect 11369 3711 11381 3887
rect 11323 3699 11381 3711
rect 11441 3887 11499 3899
rect 11441 3711 11453 3887
rect 11487 3711 11499 3887
rect 11441 3699 11499 3711
rect 11559 3887 11617 3899
rect 11559 3711 11571 3887
rect 11605 3711 11617 3887
rect 11559 3699 11617 3711
rect 11952 3706 11964 4082
rect 11998 3706 12010 4082
rect 11952 3694 12010 3706
rect 12070 4082 12128 4094
rect 12070 3706 12082 4082
rect 12116 3706 12128 4082
rect 12070 3694 12128 3706
rect 12188 4082 12246 4094
rect 12188 3706 12200 4082
rect 12234 3706 12246 4082
rect 12188 3694 12246 3706
rect 12306 4082 12364 4094
rect 12306 3706 12318 4082
rect 12352 3706 12364 4082
rect 12306 3694 12364 3706
rect 12424 4082 12482 4094
rect 12424 3706 12436 4082
rect 12470 3706 12482 4082
rect 12424 3694 12482 3706
rect 12542 4082 12600 4094
rect 12542 3706 12554 4082
rect 12588 3706 12600 4082
rect 12542 3694 12600 3706
rect 12660 4082 12718 4094
rect 12660 3706 12672 4082
rect 12706 3706 12718 4082
rect 12660 3694 12718 3706
rect 13120 4082 13178 4094
rect 13120 3706 13132 4082
rect 13166 3706 13178 4082
rect 13120 3694 13178 3706
rect 13238 4082 13296 4094
rect 13238 3706 13250 4082
rect 13284 3706 13296 4082
rect 13238 3694 13296 3706
rect 13356 4082 13414 4094
rect 13356 3706 13368 4082
rect 13402 3706 13414 4082
rect 13356 3694 13414 3706
rect 13474 4082 13532 4094
rect 13474 3706 13486 4082
rect 13520 3706 13532 4082
rect 13474 3694 13532 3706
rect 13592 4082 13650 4094
rect 13592 3706 13604 4082
rect 13638 3706 13650 4082
rect 13592 3694 13650 3706
rect 13710 4082 13768 4094
rect 13710 3706 13722 4082
rect 13756 3706 13768 4082
rect 13710 3694 13768 3706
rect 13828 4082 13886 4094
rect 13828 3706 13840 4082
rect 13874 3706 13886 4082
rect 13828 3694 13886 3706
rect 14288 4080 14346 4092
rect 14288 3704 14300 4080
rect 14334 3704 14346 4080
rect 14288 3692 14346 3704
rect 14406 4080 14464 4092
rect 14406 3704 14418 4080
rect 14452 3704 14464 4080
rect 14406 3692 14464 3704
rect 14524 4080 14582 4092
rect 14524 3704 14536 4080
rect 14570 3704 14582 4080
rect 14524 3692 14582 3704
rect 14642 4080 14700 4092
rect 14642 3704 14654 4080
rect 14688 3704 14700 4080
rect 14642 3692 14700 3704
rect 14760 4080 14818 4092
rect 14760 3704 14772 4080
rect 14806 3704 14818 4080
rect 14760 3692 14818 3704
rect 14878 4080 14936 4092
rect 14878 3704 14890 4080
rect 14924 3704 14936 4080
rect 14878 3692 14936 3704
rect 14996 4080 15054 4092
rect 14996 3704 15008 4080
rect 15042 3704 15054 4080
rect 14996 3692 15054 3704
rect 15456 4082 15514 4094
rect 15456 3706 15468 4082
rect 15502 3706 15514 4082
rect 15456 3694 15514 3706
rect 15574 4082 15632 4094
rect 15574 3706 15586 4082
rect 15620 3706 15632 4082
rect 15574 3694 15632 3706
rect 15692 4082 15750 4094
rect 15692 3706 15704 4082
rect 15738 3706 15750 4082
rect 15692 3694 15750 3706
rect 15810 4082 15868 4094
rect 15810 3706 15822 4082
rect 15856 3706 15868 4082
rect 15810 3694 15868 3706
rect 15928 4082 15986 4094
rect 15928 3706 15940 4082
rect 15974 3706 15986 4082
rect 15928 3694 15986 3706
rect 16046 4082 16104 4094
rect 16046 3706 16058 4082
rect 16092 3706 16104 4082
rect 16046 3694 16104 3706
rect 16164 4082 16222 4094
rect 16164 3706 16176 4082
rect 16210 3706 16222 4082
rect 16164 3694 16222 3706
rect 16630 4084 16688 4096
rect 16630 3708 16642 4084
rect 16676 3708 16688 4084
rect 16630 3696 16688 3708
rect 16748 4084 16806 4096
rect 16748 3708 16760 4084
rect 16794 3708 16806 4084
rect 16748 3696 16806 3708
rect 16866 4084 16924 4096
rect 16866 3708 16878 4084
rect 16912 3708 16924 4084
rect 16866 3696 16924 3708
rect 16984 4084 17042 4096
rect 16984 3708 16996 4084
rect 17030 3708 17042 4084
rect 16984 3696 17042 3708
rect 17102 4084 17160 4096
rect 17102 3708 17114 4084
rect 17148 3708 17160 4084
rect 17102 3696 17160 3708
rect 17220 4084 17278 4096
rect 17220 3708 17232 4084
rect 17266 3708 17278 4084
rect 17220 3696 17278 3708
rect 17338 4084 17396 4096
rect 17338 3708 17350 4084
rect 17384 3708 17396 4084
rect 17338 3696 17396 3708
rect 17798 4082 17856 4094
rect 17798 3706 17810 4082
rect 17844 3706 17856 4082
rect 17798 3694 17856 3706
rect 17916 4082 17974 4094
rect 17916 3706 17928 4082
rect 17962 3706 17974 4082
rect 17916 3694 17974 3706
rect 18034 4082 18092 4094
rect 18034 3706 18046 4082
rect 18080 3706 18092 4082
rect 18034 3694 18092 3706
rect 18152 4082 18210 4094
rect 18152 3706 18164 4082
rect 18198 3706 18210 4082
rect 18152 3694 18210 3706
rect 18270 4082 18328 4094
rect 18270 3706 18282 4082
rect 18316 3706 18328 4082
rect 18270 3694 18328 3706
rect 18388 4082 18446 4094
rect 18388 3706 18400 4082
rect 18434 3706 18446 4082
rect 18388 3694 18446 3706
rect 18506 4082 18564 4094
rect 18506 3706 18518 4082
rect 18552 3706 18564 4082
rect 18506 3694 18564 3706
rect 18966 4084 19024 4096
rect 18966 3708 18978 4084
rect 19012 3708 19024 4084
rect 18966 3696 19024 3708
rect 19084 4084 19142 4096
rect 19084 3708 19096 4084
rect 19130 3708 19142 4084
rect 19084 3696 19142 3708
rect 19202 4084 19260 4096
rect 19202 3708 19214 4084
rect 19248 3708 19260 4084
rect 19202 3696 19260 3708
rect 19320 4084 19378 4096
rect 19320 3708 19332 4084
rect 19366 3708 19378 4084
rect 19320 3696 19378 3708
rect 19438 4084 19496 4096
rect 19438 3708 19450 4084
rect 19484 3708 19496 4084
rect 19438 3696 19496 3708
rect 19556 4084 19614 4096
rect 19556 3708 19568 4084
rect 19602 3708 19614 4084
rect 19556 3696 19614 3708
rect 19674 4084 19732 4096
rect 19674 3708 19686 4084
rect 19720 3708 19732 4084
rect 19674 3696 19732 3708
rect 20134 4082 20192 4094
rect 20134 3706 20146 4082
rect 20180 3706 20192 4082
rect 12382 3292 12440 3304
rect 12382 3116 12394 3292
rect 12428 3116 12440 3292
rect 12382 3104 12440 3116
rect 12500 3292 12558 3304
rect 12500 3116 12512 3292
rect 12546 3116 12558 3292
rect 12500 3104 12558 3116
rect 12618 3292 12676 3304
rect 12618 3116 12630 3292
rect 12664 3116 12676 3292
rect 12618 3104 12676 3116
rect 12736 3292 12794 3304
rect 12736 3116 12748 3292
rect 12782 3116 12794 3292
rect 12736 3104 12794 3116
rect 13549 3298 13607 3310
rect 13549 3122 13561 3298
rect 13595 3122 13607 3298
rect 13549 3110 13607 3122
rect 13667 3298 13725 3310
rect 13667 3122 13679 3298
rect 13713 3122 13725 3298
rect 13667 3110 13725 3122
rect 13785 3298 13843 3310
rect 13785 3122 13797 3298
rect 13831 3122 13843 3298
rect 13785 3110 13843 3122
rect 13903 3298 13961 3310
rect 13903 3122 13915 3298
rect 13949 3122 13961 3298
rect 13903 3110 13961 3122
rect 14717 3298 14775 3310
rect 14717 3122 14729 3298
rect 14763 3122 14775 3298
rect 14717 3110 14775 3122
rect 14835 3298 14893 3310
rect 14835 3122 14847 3298
rect 14881 3122 14893 3298
rect 14835 3110 14893 3122
rect 14953 3298 15011 3310
rect 14953 3122 14965 3298
rect 14999 3122 15011 3298
rect 14953 3110 15011 3122
rect 15071 3298 15129 3310
rect 15071 3122 15083 3298
rect 15117 3122 15129 3298
rect 15071 3110 15129 3122
rect 15886 3298 15944 3310
rect 15886 3122 15898 3298
rect 15932 3122 15944 3298
rect 15886 3110 15944 3122
rect 16004 3298 16062 3310
rect 16004 3122 16016 3298
rect 16050 3122 16062 3298
rect 16004 3110 16062 3122
rect 16122 3298 16180 3310
rect 16122 3122 16134 3298
rect 16168 3122 16180 3298
rect 16122 3110 16180 3122
rect 16240 3298 16298 3310
rect 16240 3122 16252 3298
rect 16286 3122 16298 3298
rect 16240 3110 16298 3122
rect 17058 3294 17116 3306
rect 17058 3118 17070 3294
rect 17104 3118 17116 3294
rect 17058 3106 17116 3118
rect 17176 3294 17234 3306
rect 17176 3118 17188 3294
rect 17222 3118 17234 3294
rect 17176 3106 17234 3118
rect 17294 3294 17352 3306
rect 17294 3118 17306 3294
rect 17340 3118 17352 3294
rect 17294 3106 17352 3118
rect 17412 3294 17470 3306
rect 17412 3118 17424 3294
rect 17458 3118 17470 3294
rect 17412 3106 17470 3118
rect 20134 3694 20192 3706
rect 20252 4082 20310 4094
rect 20252 3706 20264 4082
rect 20298 3706 20310 4082
rect 20252 3694 20310 3706
rect 20370 4082 20428 4094
rect 20370 3706 20382 4082
rect 20416 3706 20428 4082
rect 20370 3694 20428 3706
rect 20488 4082 20546 4094
rect 20488 3706 20500 4082
rect 20534 3706 20546 4082
rect 20488 3694 20546 3706
rect 20606 4082 20664 4094
rect 20606 3706 20618 4082
rect 20652 3706 20664 4082
rect 20606 3694 20664 3706
rect 20724 4082 20782 4094
rect 20724 3706 20736 4082
rect 20770 3706 20782 4082
rect 20724 3694 20782 3706
rect 20842 4082 20900 4094
rect 20842 3706 20854 4082
rect 20888 3706 20900 4082
rect 20842 3694 20900 3706
rect 18227 3293 18285 3305
rect 18227 3117 18239 3293
rect 18273 3117 18285 3293
rect 18227 3105 18285 3117
rect 18345 3293 18403 3305
rect 18345 3117 18357 3293
rect 18391 3117 18403 3293
rect 18345 3105 18403 3117
rect 18463 3293 18521 3305
rect 18463 3117 18475 3293
rect 18509 3117 18521 3293
rect 18463 3105 18521 3117
rect 18581 3293 18639 3305
rect 18581 3117 18593 3293
rect 18627 3117 18639 3293
rect 18581 3105 18639 3117
rect 19395 3293 19453 3305
rect 19395 3117 19407 3293
rect 19441 3117 19453 3293
rect 19395 3105 19453 3117
rect 19513 3293 19571 3305
rect 19513 3117 19525 3293
rect 19559 3117 19571 3293
rect 19513 3105 19571 3117
rect 19631 3293 19689 3305
rect 19631 3117 19643 3293
rect 19677 3117 19689 3293
rect 19631 3105 19689 3117
rect 19749 3293 19807 3305
rect 19749 3117 19761 3293
rect 19795 3117 19807 3293
rect 19749 3105 19807 3117
rect 20563 3294 20621 3306
rect 20563 3118 20575 3294
rect 20609 3118 20621 3294
rect 20563 3106 20621 3118
rect 20681 3294 20739 3306
rect 20681 3118 20693 3294
rect 20727 3118 20739 3294
rect 20681 3106 20739 3118
rect 20799 3294 20857 3306
rect 20799 3118 20811 3294
rect 20845 3118 20857 3294
rect 20799 3106 20857 3118
rect 20917 3294 20975 3306
rect 20917 3118 20929 3294
rect 20963 3118 20975 3294
rect 20917 3106 20975 3118
rect 689 2128 747 2140
rect 689 1940 701 2128
rect 248 1928 306 1940
rect 248 1752 260 1928
rect 294 1752 306 1928
rect 248 1740 306 1752
rect 366 1928 424 1940
rect 366 1752 378 1928
rect 412 1752 424 1928
rect 366 1740 424 1752
rect 484 1928 542 1940
rect 484 1752 496 1928
rect 530 1752 542 1928
rect 484 1740 542 1752
rect 602 1928 701 1940
rect 602 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 747 2128
rect 602 1740 747 1752
rect 807 2128 865 2140
rect 807 1752 819 2128
rect 853 1752 865 2128
rect 807 1740 865 1752
rect 925 2128 983 2140
rect 925 1752 937 2128
rect 971 1752 983 2128
rect 925 1740 983 1752
rect 1043 2128 1101 2140
rect 1043 1752 1055 2128
rect 1089 1752 1101 2128
rect 1043 1740 1101 1752
rect 1156 2128 1214 2140
rect 1156 1752 1168 2128
rect 1202 1752 1214 2128
rect 1156 1740 1214 1752
rect 1274 2128 1332 2140
rect 1274 1752 1286 2128
rect 1320 1752 1332 2128
rect 1274 1740 1332 1752
rect 1392 2128 1450 2140
rect 1392 1752 1404 2128
rect 1438 1752 1450 2128
rect 1392 1740 1450 1752
rect 1510 2128 1568 2140
rect 1510 1752 1522 2128
rect 1556 1752 1568 2128
rect 1510 1740 1568 1752
rect 1628 2128 1686 2140
rect 1628 1752 1640 2128
rect 1674 1752 1686 2128
rect 1628 1740 1686 1752
rect 1746 2128 1804 2140
rect 1746 1752 1758 2128
rect 1792 1752 1804 2128
rect 1746 1740 1804 1752
rect 1864 2128 1922 2140
rect 1864 1752 1876 2128
rect 1910 1752 1922 2128
rect 1864 1740 1922 1752
rect 1983 2128 2041 2140
rect 1983 1752 1995 2128
rect 2029 1752 2041 2128
rect 1983 1740 2041 1752
rect 2101 2128 2159 2140
rect 2101 1752 2113 2128
rect 2147 1752 2159 2128
rect 2101 1740 2159 1752
rect 2219 2128 2277 2140
rect 2219 1752 2231 2128
rect 2265 1752 2277 2128
rect 2219 1740 2277 1752
rect 2337 2128 2395 2140
rect 2337 1752 2349 2128
rect 2383 1752 2395 2128
rect 3833 2128 3891 2140
rect 3833 1940 3845 2128
rect 2337 1740 2395 1752
rect 2456 1928 2514 1940
rect 2456 1752 2468 1928
rect 2502 1752 2514 1928
rect 2456 1740 2514 1752
rect 2574 1928 2632 1940
rect 2574 1752 2586 1928
rect 2620 1752 2632 1928
rect 2574 1740 2632 1752
rect 2692 1928 2750 1940
rect 2692 1752 2704 1928
rect 2738 1752 2750 1928
rect 2692 1740 2750 1752
rect 2810 1928 2868 1940
rect 2810 1752 2822 1928
rect 2856 1752 2868 1928
rect 2810 1740 2868 1752
rect 3392 1928 3450 1940
rect 3392 1752 3404 1928
rect 3438 1752 3450 1928
rect 3392 1740 3450 1752
rect 3510 1928 3568 1940
rect 3510 1752 3522 1928
rect 3556 1752 3568 1928
rect 3510 1740 3568 1752
rect 3628 1928 3686 1940
rect 3628 1752 3640 1928
rect 3674 1752 3686 1928
rect 3628 1740 3686 1752
rect 3746 1928 3845 1940
rect 3746 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3891 2128
rect 3746 1740 3891 1752
rect 3951 2128 4009 2140
rect 3951 1752 3963 2128
rect 3997 1752 4009 2128
rect 3951 1740 4009 1752
rect 4069 2128 4127 2140
rect 4069 1752 4081 2128
rect 4115 1752 4127 2128
rect 4069 1740 4127 1752
rect 4187 2128 4245 2140
rect 4187 1752 4199 2128
rect 4233 1752 4245 2128
rect 4187 1740 4245 1752
rect 4300 2128 4358 2140
rect 4300 1752 4312 2128
rect 4346 1752 4358 2128
rect 4300 1740 4358 1752
rect 4418 2128 4476 2140
rect 4418 1752 4430 2128
rect 4464 1752 4476 2128
rect 4418 1740 4476 1752
rect 4536 2128 4594 2140
rect 4536 1752 4548 2128
rect 4582 1752 4594 2128
rect 4536 1740 4594 1752
rect 4654 2128 4712 2140
rect 4654 1752 4666 2128
rect 4700 1752 4712 2128
rect 4654 1740 4712 1752
rect 4772 2128 4830 2140
rect 4772 1752 4784 2128
rect 4818 1752 4830 2128
rect 4772 1740 4830 1752
rect 4890 2128 4948 2140
rect 4890 1752 4902 2128
rect 4936 1752 4948 2128
rect 4890 1740 4948 1752
rect 5008 2128 5066 2140
rect 5008 1752 5020 2128
rect 5054 1752 5066 2128
rect 5008 1740 5066 1752
rect 5127 2128 5185 2140
rect 5127 1752 5139 2128
rect 5173 1752 5185 2128
rect 5127 1740 5185 1752
rect 5245 2128 5303 2140
rect 5245 1752 5257 2128
rect 5291 1752 5303 2128
rect 5245 1740 5303 1752
rect 5363 2128 5421 2140
rect 5363 1752 5375 2128
rect 5409 1752 5421 2128
rect 5363 1740 5421 1752
rect 5481 2128 5539 2140
rect 5481 1752 5493 2128
rect 5527 1752 5539 2128
rect 6965 2132 7023 2144
rect 6965 1944 6977 2132
rect 5481 1740 5539 1752
rect 5600 1928 5658 1940
rect 5600 1752 5612 1928
rect 5646 1752 5658 1928
rect 5600 1740 5658 1752
rect 5718 1928 5776 1940
rect 5718 1752 5730 1928
rect 5764 1752 5776 1928
rect 5718 1740 5776 1752
rect 5836 1928 5894 1940
rect 5836 1752 5848 1928
rect 5882 1752 5894 1928
rect 5836 1740 5894 1752
rect 5954 1928 6012 1940
rect 5954 1752 5966 1928
rect 6000 1752 6012 1928
rect 5954 1740 6012 1752
rect 6524 1932 6582 1944
rect 6524 1756 6536 1932
rect 6570 1756 6582 1932
rect 6524 1744 6582 1756
rect 6642 1932 6700 1944
rect 6642 1756 6654 1932
rect 6688 1756 6700 1932
rect 6642 1744 6700 1756
rect 6760 1932 6818 1944
rect 6760 1756 6772 1932
rect 6806 1756 6818 1932
rect 6760 1744 6818 1756
rect 6878 1932 6977 1944
rect 6878 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7023 2132
rect 6878 1744 7023 1756
rect 7083 2132 7141 2144
rect 7083 1756 7095 2132
rect 7129 1756 7141 2132
rect 7083 1744 7141 1756
rect 7201 2132 7259 2144
rect 7201 1756 7213 2132
rect 7247 1756 7259 2132
rect 7201 1744 7259 1756
rect 7319 2132 7377 2144
rect 7319 1756 7331 2132
rect 7365 1756 7377 2132
rect 7319 1744 7377 1756
rect 7432 2132 7490 2144
rect 7432 1756 7444 2132
rect 7478 1756 7490 2132
rect 7432 1744 7490 1756
rect 7550 2132 7608 2144
rect 7550 1756 7562 2132
rect 7596 1756 7608 2132
rect 7550 1744 7608 1756
rect 7668 2132 7726 2144
rect 7668 1756 7680 2132
rect 7714 1756 7726 2132
rect 7668 1744 7726 1756
rect 7786 2132 7844 2144
rect 7786 1756 7798 2132
rect 7832 1756 7844 2132
rect 7786 1744 7844 1756
rect 7904 2132 7962 2144
rect 7904 1756 7916 2132
rect 7950 1756 7962 2132
rect 7904 1744 7962 1756
rect 8022 2132 8080 2144
rect 8022 1756 8034 2132
rect 8068 1756 8080 2132
rect 8022 1744 8080 1756
rect 8140 2132 8198 2144
rect 8140 1756 8152 2132
rect 8186 1756 8198 2132
rect 8140 1744 8198 1756
rect 8259 2132 8317 2144
rect 8259 1756 8271 2132
rect 8305 1756 8317 2132
rect 8259 1744 8317 1756
rect 8377 2132 8435 2144
rect 8377 1756 8389 2132
rect 8423 1756 8435 2132
rect 8377 1744 8435 1756
rect 8495 2132 8553 2144
rect 8495 1756 8507 2132
rect 8541 1756 8553 2132
rect 8495 1744 8553 1756
rect 8613 2132 8671 2144
rect 8613 1756 8625 2132
rect 8659 1756 8671 2132
rect 10109 2132 10167 2144
rect 10109 1944 10121 2132
rect 8613 1744 8671 1756
rect 8732 1932 8790 1944
rect 8732 1756 8744 1932
rect 8778 1756 8790 1932
rect 8732 1744 8790 1756
rect 8850 1932 8908 1944
rect 8850 1756 8862 1932
rect 8896 1756 8908 1932
rect 8850 1744 8908 1756
rect 8968 1932 9026 1944
rect 8968 1756 8980 1932
rect 9014 1756 9026 1932
rect 8968 1744 9026 1756
rect 9086 1932 9144 1944
rect 9086 1756 9098 1932
rect 9132 1756 9144 1932
rect 9086 1744 9144 1756
rect 9668 1932 9726 1944
rect 9668 1756 9680 1932
rect 9714 1756 9726 1932
rect 9668 1744 9726 1756
rect 9786 1932 9844 1944
rect 9786 1756 9798 1932
rect 9832 1756 9844 1932
rect 9786 1744 9844 1756
rect 9904 1932 9962 1944
rect 9904 1756 9916 1932
rect 9950 1756 9962 1932
rect 9904 1744 9962 1756
rect 10022 1932 10121 1944
rect 10022 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10167 2132
rect 10022 1744 10167 1756
rect 10227 2132 10285 2144
rect 10227 1756 10239 2132
rect 10273 1756 10285 2132
rect 10227 1744 10285 1756
rect 10345 2132 10403 2144
rect 10345 1756 10357 2132
rect 10391 1756 10403 2132
rect 10345 1744 10403 1756
rect 10463 2132 10521 2144
rect 10463 1756 10475 2132
rect 10509 1756 10521 2132
rect 10463 1744 10521 1756
rect 10576 2132 10634 2144
rect 10576 1756 10588 2132
rect 10622 1756 10634 2132
rect 10576 1744 10634 1756
rect 10694 2132 10752 2144
rect 10694 1756 10706 2132
rect 10740 1756 10752 2132
rect 10694 1744 10752 1756
rect 10812 2132 10870 2144
rect 10812 1756 10824 2132
rect 10858 1756 10870 2132
rect 10812 1744 10870 1756
rect 10930 2132 10988 2144
rect 10930 1756 10942 2132
rect 10976 1756 10988 2132
rect 10930 1744 10988 1756
rect 11048 2132 11106 2144
rect 11048 1756 11060 2132
rect 11094 1756 11106 2132
rect 11048 1744 11106 1756
rect 11166 2132 11224 2144
rect 11166 1756 11178 2132
rect 11212 1756 11224 2132
rect 11166 1744 11224 1756
rect 11284 2132 11342 2144
rect 11284 1756 11296 2132
rect 11330 1756 11342 2132
rect 11284 1744 11342 1756
rect 11403 2132 11461 2144
rect 11403 1756 11415 2132
rect 11449 1756 11461 2132
rect 11403 1744 11461 1756
rect 11521 2132 11579 2144
rect 11521 1756 11533 2132
rect 11567 1756 11579 2132
rect 11521 1744 11579 1756
rect 11639 2132 11697 2144
rect 11639 1756 11651 2132
rect 11685 1756 11697 2132
rect 11639 1744 11697 1756
rect 11757 2132 11815 2144
rect 11757 1756 11769 2132
rect 11803 1756 11815 2132
rect 13311 2128 13369 2140
rect 11757 1744 11815 1756
rect 11876 1932 11934 1944
rect 11876 1756 11888 1932
rect 11922 1756 11934 1932
rect 11876 1744 11934 1756
rect 11994 1932 12052 1944
rect 11994 1756 12006 1932
rect 12040 1756 12052 1932
rect 11994 1744 12052 1756
rect 12112 1932 12170 1944
rect 12112 1756 12124 1932
rect 12158 1756 12170 1932
rect 12112 1744 12170 1756
rect 12230 1932 12288 1944
rect 13311 1940 13323 2128
rect 12230 1756 12242 1932
rect 12276 1756 12288 1932
rect 12230 1744 12288 1756
rect 12870 1928 12928 1940
rect 12870 1752 12882 1928
rect 12916 1752 12928 1928
rect 12870 1740 12928 1752
rect 12988 1928 13046 1940
rect 12988 1752 13000 1928
rect 13034 1752 13046 1928
rect 12988 1740 13046 1752
rect 13106 1928 13164 1940
rect 13106 1752 13118 1928
rect 13152 1752 13164 1928
rect 13106 1740 13164 1752
rect 13224 1928 13323 1940
rect 13224 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13369 2128
rect 13224 1740 13369 1752
rect 13429 2128 13487 2140
rect 13429 1752 13441 2128
rect 13475 1752 13487 2128
rect 13429 1740 13487 1752
rect 13547 2128 13605 2140
rect 13547 1752 13559 2128
rect 13593 1752 13605 2128
rect 13547 1740 13605 1752
rect 13665 2128 13723 2140
rect 13665 1752 13677 2128
rect 13711 1752 13723 2128
rect 13665 1740 13723 1752
rect 13778 2128 13836 2140
rect 13778 1752 13790 2128
rect 13824 1752 13836 2128
rect 13778 1740 13836 1752
rect 13896 2128 13954 2140
rect 13896 1752 13908 2128
rect 13942 1752 13954 2128
rect 13896 1740 13954 1752
rect 14014 2128 14072 2140
rect 14014 1752 14026 2128
rect 14060 1752 14072 2128
rect 14014 1740 14072 1752
rect 14132 2128 14190 2140
rect 14132 1752 14144 2128
rect 14178 1752 14190 2128
rect 14132 1740 14190 1752
rect 14250 2128 14308 2140
rect 14250 1752 14262 2128
rect 14296 1752 14308 2128
rect 14250 1740 14308 1752
rect 14368 2128 14426 2140
rect 14368 1752 14380 2128
rect 14414 1752 14426 2128
rect 14368 1740 14426 1752
rect 14486 2128 14544 2140
rect 14486 1752 14498 2128
rect 14532 1752 14544 2128
rect 14486 1740 14544 1752
rect 14605 2128 14663 2140
rect 14605 1752 14617 2128
rect 14651 1752 14663 2128
rect 14605 1740 14663 1752
rect 14723 2128 14781 2140
rect 14723 1752 14735 2128
rect 14769 1752 14781 2128
rect 14723 1740 14781 1752
rect 14841 2128 14899 2140
rect 14841 1752 14853 2128
rect 14887 1752 14899 2128
rect 14841 1740 14899 1752
rect 14959 2128 15017 2140
rect 14959 1752 14971 2128
rect 15005 1752 15017 2128
rect 16455 2128 16513 2140
rect 16455 1940 16467 2128
rect 14959 1740 15017 1752
rect 15078 1928 15136 1940
rect 15078 1752 15090 1928
rect 15124 1752 15136 1928
rect 15078 1740 15136 1752
rect 15196 1928 15254 1940
rect 15196 1752 15208 1928
rect 15242 1752 15254 1928
rect 15196 1740 15254 1752
rect 15314 1928 15372 1940
rect 15314 1752 15326 1928
rect 15360 1752 15372 1928
rect 15314 1740 15372 1752
rect 15432 1928 15490 1940
rect 15432 1752 15444 1928
rect 15478 1752 15490 1928
rect 15432 1740 15490 1752
rect 16014 1928 16072 1940
rect 16014 1752 16026 1928
rect 16060 1752 16072 1928
rect 16014 1740 16072 1752
rect 16132 1928 16190 1940
rect 16132 1752 16144 1928
rect 16178 1752 16190 1928
rect 16132 1740 16190 1752
rect 16250 1928 16308 1940
rect 16250 1752 16262 1928
rect 16296 1752 16308 1928
rect 16250 1740 16308 1752
rect 16368 1928 16467 1940
rect 16368 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16513 2128
rect 16368 1740 16513 1752
rect 16573 2128 16631 2140
rect 16573 1752 16585 2128
rect 16619 1752 16631 2128
rect 16573 1740 16631 1752
rect 16691 2128 16749 2140
rect 16691 1752 16703 2128
rect 16737 1752 16749 2128
rect 16691 1740 16749 1752
rect 16809 2128 16867 2140
rect 16809 1752 16821 2128
rect 16855 1752 16867 2128
rect 16809 1740 16867 1752
rect 16922 2128 16980 2140
rect 16922 1752 16934 2128
rect 16968 1752 16980 2128
rect 16922 1740 16980 1752
rect 17040 2128 17098 2140
rect 17040 1752 17052 2128
rect 17086 1752 17098 2128
rect 17040 1740 17098 1752
rect 17158 2128 17216 2140
rect 17158 1752 17170 2128
rect 17204 1752 17216 2128
rect 17158 1740 17216 1752
rect 17276 2128 17334 2140
rect 17276 1752 17288 2128
rect 17322 1752 17334 2128
rect 17276 1740 17334 1752
rect 17394 2128 17452 2140
rect 17394 1752 17406 2128
rect 17440 1752 17452 2128
rect 17394 1740 17452 1752
rect 17512 2128 17570 2140
rect 17512 1752 17524 2128
rect 17558 1752 17570 2128
rect 17512 1740 17570 1752
rect 17630 2128 17688 2140
rect 17630 1752 17642 2128
rect 17676 1752 17688 2128
rect 17630 1740 17688 1752
rect 17749 2128 17807 2140
rect 17749 1752 17761 2128
rect 17795 1752 17807 2128
rect 17749 1740 17807 1752
rect 17867 2128 17925 2140
rect 17867 1752 17879 2128
rect 17913 1752 17925 2128
rect 17867 1740 17925 1752
rect 17985 2128 18043 2140
rect 17985 1752 17997 2128
rect 18031 1752 18043 2128
rect 17985 1740 18043 1752
rect 18103 2128 18161 2140
rect 18103 1752 18115 2128
rect 18149 1752 18161 2128
rect 19587 2132 19645 2144
rect 19587 1944 19599 2132
rect 18103 1740 18161 1752
rect 18222 1928 18280 1940
rect 18222 1752 18234 1928
rect 18268 1752 18280 1928
rect 18222 1740 18280 1752
rect 18340 1928 18398 1940
rect 18340 1752 18352 1928
rect 18386 1752 18398 1928
rect 18340 1740 18398 1752
rect 18458 1928 18516 1940
rect 18458 1752 18470 1928
rect 18504 1752 18516 1928
rect 18458 1740 18516 1752
rect 18576 1928 18634 1940
rect 18576 1752 18588 1928
rect 18622 1752 18634 1928
rect 18576 1740 18634 1752
rect 19146 1932 19204 1944
rect 19146 1756 19158 1932
rect 19192 1756 19204 1932
rect 19146 1744 19204 1756
rect 19264 1932 19322 1944
rect 19264 1756 19276 1932
rect 19310 1756 19322 1932
rect 19264 1744 19322 1756
rect 19382 1932 19440 1944
rect 19382 1756 19394 1932
rect 19428 1756 19440 1932
rect 19382 1744 19440 1756
rect 19500 1932 19599 1944
rect 19500 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19645 2132
rect 19500 1744 19645 1756
rect 19705 2132 19763 2144
rect 19705 1756 19717 2132
rect 19751 1756 19763 2132
rect 19705 1744 19763 1756
rect 19823 2132 19881 2144
rect 19823 1756 19835 2132
rect 19869 1756 19881 2132
rect 19823 1744 19881 1756
rect 19941 2132 19999 2144
rect 19941 1756 19953 2132
rect 19987 1756 19999 2132
rect 19941 1744 19999 1756
rect 20054 2132 20112 2144
rect 20054 1756 20066 2132
rect 20100 1756 20112 2132
rect 20054 1744 20112 1756
rect 20172 2132 20230 2144
rect 20172 1756 20184 2132
rect 20218 1756 20230 2132
rect 20172 1744 20230 1756
rect 20290 2132 20348 2144
rect 20290 1756 20302 2132
rect 20336 1756 20348 2132
rect 20290 1744 20348 1756
rect 20408 2132 20466 2144
rect 20408 1756 20420 2132
rect 20454 1756 20466 2132
rect 20408 1744 20466 1756
rect 20526 2132 20584 2144
rect 20526 1756 20538 2132
rect 20572 1756 20584 2132
rect 20526 1744 20584 1756
rect 20644 2132 20702 2144
rect 20644 1756 20656 2132
rect 20690 1756 20702 2132
rect 20644 1744 20702 1756
rect 20762 2132 20820 2144
rect 20762 1756 20774 2132
rect 20808 1756 20820 2132
rect 20762 1744 20820 1756
rect 20881 2132 20939 2144
rect 20881 1756 20893 2132
rect 20927 1756 20939 2132
rect 20881 1744 20939 1756
rect 20999 2132 21057 2144
rect 20999 1756 21011 2132
rect 21045 1756 21057 2132
rect 20999 1744 21057 1756
rect 21117 2132 21175 2144
rect 21117 1756 21129 2132
rect 21163 1756 21175 2132
rect 21117 1744 21175 1756
rect 21235 2132 21293 2144
rect 21235 1756 21247 2132
rect 21281 1756 21293 2132
rect 22731 2132 22789 2144
rect 22731 1944 22743 2132
rect 21235 1744 21293 1756
rect 21354 1932 21412 1944
rect 21354 1756 21366 1932
rect 21400 1756 21412 1932
rect 21354 1744 21412 1756
rect 21472 1932 21530 1944
rect 21472 1756 21484 1932
rect 21518 1756 21530 1932
rect 21472 1744 21530 1756
rect 21590 1932 21648 1944
rect 21590 1756 21602 1932
rect 21636 1756 21648 1932
rect 21590 1744 21648 1756
rect 21708 1932 21766 1944
rect 21708 1756 21720 1932
rect 21754 1756 21766 1932
rect 21708 1744 21766 1756
rect 22290 1932 22348 1944
rect 22290 1756 22302 1932
rect 22336 1756 22348 1932
rect 22290 1744 22348 1756
rect 22408 1932 22466 1944
rect 22408 1756 22420 1932
rect 22454 1756 22466 1932
rect 22408 1744 22466 1756
rect 22526 1932 22584 1944
rect 22526 1756 22538 1932
rect 22572 1756 22584 1932
rect 22526 1744 22584 1756
rect 22644 1932 22743 1944
rect 22644 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22789 2132
rect 22644 1744 22789 1756
rect 22849 2132 22907 2144
rect 22849 1756 22861 2132
rect 22895 1756 22907 2132
rect 22849 1744 22907 1756
rect 22967 2132 23025 2144
rect 22967 1756 22979 2132
rect 23013 1756 23025 2132
rect 22967 1744 23025 1756
rect 23085 2132 23143 2144
rect 23085 1756 23097 2132
rect 23131 1756 23143 2132
rect 23085 1744 23143 1756
rect 23198 2132 23256 2144
rect 23198 1756 23210 2132
rect 23244 1756 23256 2132
rect 23198 1744 23256 1756
rect 23316 2132 23374 2144
rect 23316 1756 23328 2132
rect 23362 1756 23374 2132
rect 23316 1744 23374 1756
rect 23434 2132 23492 2144
rect 23434 1756 23446 2132
rect 23480 1756 23492 2132
rect 23434 1744 23492 1756
rect 23552 2132 23610 2144
rect 23552 1756 23564 2132
rect 23598 1756 23610 2132
rect 23552 1744 23610 1756
rect 23670 2132 23728 2144
rect 23670 1756 23682 2132
rect 23716 1756 23728 2132
rect 23670 1744 23728 1756
rect 23788 2132 23846 2144
rect 23788 1756 23800 2132
rect 23834 1756 23846 2132
rect 23788 1744 23846 1756
rect 23906 2132 23964 2144
rect 23906 1756 23918 2132
rect 23952 1756 23964 2132
rect 23906 1744 23964 1756
rect 24025 2132 24083 2144
rect 24025 1756 24037 2132
rect 24071 1756 24083 2132
rect 24025 1744 24083 1756
rect 24143 2132 24201 2144
rect 24143 1756 24155 2132
rect 24189 1756 24201 2132
rect 24143 1744 24201 1756
rect 24261 2132 24319 2144
rect 24261 1756 24273 2132
rect 24307 1756 24319 2132
rect 24261 1744 24319 1756
rect 24379 2132 24437 2144
rect 24379 1756 24391 2132
rect 24425 1756 24437 2132
rect 24379 1744 24437 1756
rect 24498 1932 24556 1944
rect 24498 1756 24510 1932
rect 24544 1756 24556 1932
rect 24498 1744 24556 1756
rect 24616 1932 24674 1944
rect 24616 1756 24628 1932
rect 24662 1756 24674 1932
rect 24616 1744 24674 1756
rect 24734 1932 24792 1944
rect 24734 1756 24746 1932
rect 24780 1756 24792 1932
rect 24734 1744 24792 1756
rect 24852 1932 24910 1944
rect 24852 1756 24864 1932
rect 24898 1756 24910 1932
rect 24852 1744 24910 1756
rect 689 -606 747 -594
rect 689 -794 701 -606
rect 248 -806 306 -794
rect 248 -982 260 -806
rect 294 -982 306 -806
rect 248 -994 306 -982
rect 366 -806 424 -794
rect 366 -982 378 -806
rect 412 -982 424 -806
rect 366 -994 424 -982
rect 484 -806 542 -794
rect 484 -982 496 -806
rect 530 -982 542 -806
rect 484 -994 542 -982
rect 602 -806 701 -794
rect 602 -982 614 -806
rect 648 -982 701 -806
rect 735 -982 747 -606
rect 602 -994 747 -982
rect 807 -606 865 -594
rect 807 -982 819 -606
rect 853 -982 865 -606
rect 807 -994 865 -982
rect 925 -606 983 -594
rect 925 -982 937 -606
rect 971 -982 983 -606
rect 925 -994 983 -982
rect 1043 -606 1101 -594
rect 1043 -982 1055 -606
rect 1089 -982 1101 -606
rect 1043 -994 1101 -982
rect 1156 -606 1214 -594
rect 1156 -982 1168 -606
rect 1202 -982 1214 -606
rect 1156 -994 1214 -982
rect 1274 -606 1332 -594
rect 1274 -982 1286 -606
rect 1320 -982 1332 -606
rect 1274 -994 1332 -982
rect 1392 -606 1450 -594
rect 1392 -982 1404 -606
rect 1438 -982 1450 -606
rect 1392 -994 1450 -982
rect 1510 -606 1568 -594
rect 1510 -982 1522 -606
rect 1556 -982 1568 -606
rect 1510 -994 1568 -982
rect 1628 -606 1686 -594
rect 1628 -982 1640 -606
rect 1674 -982 1686 -606
rect 1628 -994 1686 -982
rect 1746 -606 1804 -594
rect 1746 -982 1758 -606
rect 1792 -982 1804 -606
rect 1746 -994 1804 -982
rect 1864 -606 1922 -594
rect 1864 -982 1876 -606
rect 1910 -982 1922 -606
rect 1864 -994 1922 -982
rect 1983 -606 2041 -594
rect 1983 -982 1995 -606
rect 2029 -982 2041 -606
rect 1983 -994 2041 -982
rect 2101 -606 2159 -594
rect 2101 -982 2113 -606
rect 2147 -982 2159 -606
rect 2101 -994 2159 -982
rect 2219 -606 2277 -594
rect 2219 -982 2231 -606
rect 2265 -982 2277 -606
rect 2219 -994 2277 -982
rect 2337 -606 2395 -594
rect 2337 -982 2349 -606
rect 2383 -982 2395 -606
rect 3833 -606 3891 -594
rect 3833 -794 3845 -606
rect 2337 -994 2395 -982
rect 2456 -806 2514 -794
rect 2456 -982 2468 -806
rect 2502 -982 2514 -806
rect 2456 -994 2514 -982
rect 2574 -806 2632 -794
rect 2574 -982 2586 -806
rect 2620 -982 2632 -806
rect 2574 -994 2632 -982
rect 2692 -806 2750 -794
rect 2692 -982 2704 -806
rect 2738 -982 2750 -806
rect 2692 -994 2750 -982
rect 2810 -806 2868 -794
rect 2810 -982 2822 -806
rect 2856 -982 2868 -806
rect 2810 -994 2868 -982
rect 3392 -806 3450 -794
rect 3392 -982 3404 -806
rect 3438 -982 3450 -806
rect 3392 -994 3450 -982
rect 3510 -806 3568 -794
rect 3510 -982 3522 -806
rect 3556 -982 3568 -806
rect 3510 -994 3568 -982
rect 3628 -806 3686 -794
rect 3628 -982 3640 -806
rect 3674 -982 3686 -806
rect 3628 -994 3686 -982
rect 3746 -806 3845 -794
rect 3746 -982 3758 -806
rect 3792 -982 3845 -806
rect 3879 -982 3891 -606
rect 3746 -994 3891 -982
rect 3951 -606 4009 -594
rect 3951 -982 3963 -606
rect 3997 -982 4009 -606
rect 3951 -994 4009 -982
rect 4069 -606 4127 -594
rect 4069 -982 4081 -606
rect 4115 -982 4127 -606
rect 4069 -994 4127 -982
rect 4187 -606 4245 -594
rect 4187 -982 4199 -606
rect 4233 -982 4245 -606
rect 4187 -994 4245 -982
rect 4300 -606 4358 -594
rect 4300 -982 4312 -606
rect 4346 -982 4358 -606
rect 4300 -994 4358 -982
rect 4418 -606 4476 -594
rect 4418 -982 4430 -606
rect 4464 -982 4476 -606
rect 4418 -994 4476 -982
rect 4536 -606 4594 -594
rect 4536 -982 4548 -606
rect 4582 -982 4594 -606
rect 4536 -994 4594 -982
rect 4654 -606 4712 -594
rect 4654 -982 4666 -606
rect 4700 -982 4712 -606
rect 4654 -994 4712 -982
rect 4772 -606 4830 -594
rect 4772 -982 4784 -606
rect 4818 -982 4830 -606
rect 4772 -994 4830 -982
rect 4890 -606 4948 -594
rect 4890 -982 4902 -606
rect 4936 -982 4948 -606
rect 4890 -994 4948 -982
rect 5008 -606 5066 -594
rect 5008 -982 5020 -606
rect 5054 -982 5066 -606
rect 5008 -994 5066 -982
rect 5127 -606 5185 -594
rect 5127 -982 5139 -606
rect 5173 -982 5185 -606
rect 5127 -994 5185 -982
rect 5245 -606 5303 -594
rect 5245 -982 5257 -606
rect 5291 -982 5303 -606
rect 5245 -994 5303 -982
rect 5363 -606 5421 -594
rect 5363 -982 5375 -606
rect 5409 -982 5421 -606
rect 5363 -994 5421 -982
rect 5481 -606 5539 -594
rect 5481 -982 5493 -606
rect 5527 -982 5539 -606
rect 6965 -602 7023 -590
rect 6965 -790 6977 -602
rect 5481 -994 5539 -982
rect 5600 -806 5658 -794
rect 5600 -982 5612 -806
rect 5646 -982 5658 -806
rect 5600 -994 5658 -982
rect 5718 -806 5776 -794
rect 5718 -982 5730 -806
rect 5764 -982 5776 -806
rect 5718 -994 5776 -982
rect 5836 -806 5894 -794
rect 5836 -982 5848 -806
rect 5882 -982 5894 -806
rect 5836 -994 5894 -982
rect 5954 -806 6012 -794
rect 5954 -982 5966 -806
rect 6000 -982 6012 -806
rect 5954 -994 6012 -982
rect 6524 -802 6582 -790
rect 6524 -978 6536 -802
rect 6570 -978 6582 -802
rect 6524 -990 6582 -978
rect 6642 -802 6700 -790
rect 6642 -978 6654 -802
rect 6688 -978 6700 -802
rect 6642 -990 6700 -978
rect 6760 -802 6818 -790
rect 6760 -978 6772 -802
rect 6806 -978 6818 -802
rect 6760 -990 6818 -978
rect 6878 -802 6977 -790
rect 6878 -978 6890 -802
rect 6924 -978 6977 -802
rect 7011 -978 7023 -602
rect 6878 -990 7023 -978
rect 7083 -602 7141 -590
rect 7083 -978 7095 -602
rect 7129 -978 7141 -602
rect 7083 -990 7141 -978
rect 7201 -602 7259 -590
rect 7201 -978 7213 -602
rect 7247 -978 7259 -602
rect 7201 -990 7259 -978
rect 7319 -602 7377 -590
rect 7319 -978 7331 -602
rect 7365 -978 7377 -602
rect 7319 -990 7377 -978
rect 7432 -602 7490 -590
rect 7432 -978 7444 -602
rect 7478 -978 7490 -602
rect 7432 -990 7490 -978
rect 7550 -602 7608 -590
rect 7550 -978 7562 -602
rect 7596 -978 7608 -602
rect 7550 -990 7608 -978
rect 7668 -602 7726 -590
rect 7668 -978 7680 -602
rect 7714 -978 7726 -602
rect 7668 -990 7726 -978
rect 7786 -602 7844 -590
rect 7786 -978 7798 -602
rect 7832 -978 7844 -602
rect 7786 -990 7844 -978
rect 7904 -602 7962 -590
rect 7904 -978 7916 -602
rect 7950 -978 7962 -602
rect 7904 -990 7962 -978
rect 8022 -602 8080 -590
rect 8022 -978 8034 -602
rect 8068 -978 8080 -602
rect 8022 -990 8080 -978
rect 8140 -602 8198 -590
rect 8140 -978 8152 -602
rect 8186 -978 8198 -602
rect 8140 -990 8198 -978
rect 8259 -602 8317 -590
rect 8259 -978 8271 -602
rect 8305 -978 8317 -602
rect 8259 -990 8317 -978
rect 8377 -602 8435 -590
rect 8377 -978 8389 -602
rect 8423 -978 8435 -602
rect 8377 -990 8435 -978
rect 8495 -602 8553 -590
rect 8495 -978 8507 -602
rect 8541 -978 8553 -602
rect 8495 -990 8553 -978
rect 8613 -602 8671 -590
rect 8613 -978 8625 -602
rect 8659 -978 8671 -602
rect 10109 -602 10167 -590
rect 10109 -790 10121 -602
rect 8613 -990 8671 -978
rect 8732 -802 8790 -790
rect 8732 -978 8744 -802
rect 8778 -978 8790 -802
rect 8732 -990 8790 -978
rect 8850 -802 8908 -790
rect 8850 -978 8862 -802
rect 8896 -978 8908 -802
rect 8850 -990 8908 -978
rect 8968 -802 9026 -790
rect 8968 -978 8980 -802
rect 9014 -978 9026 -802
rect 8968 -990 9026 -978
rect 9086 -802 9144 -790
rect 9086 -978 9098 -802
rect 9132 -978 9144 -802
rect 9086 -990 9144 -978
rect 9668 -802 9726 -790
rect 9668 -978 9680 -802
rect 9714 -978 9726 -802
rect 9668 -990 9726 -978
rect 9786 -802 9844 -790
rect 9786 -978 9798 -802
rect 9832 -978 9844 -802
rect 9786 -990 9844 -978
rect 9904 -802 9962 -790
rect 9904 -978 9916 -802
rect 9950 -978 9962 -802
rect 9904 -990 9962 -978
rect 10022 -802 10121 -790
rect 10022 -978 10034 -802
rect 10068 -978 10121 -802
rect 10155 -978 10167 -602
rect 10022 -990 10167 -978
rect 10227 -602 10285 -590
rect 10227 -978 10239 -602
rect 10273 -978 10285 -602
rect 10227 -990 10285 -978
rect 10345 -602 10403 -590
rect 10345 -978 10357 -602
rect 10391 -978 10403 -602
rect 10345 -990 10403 -978
rect 10463 -602 10521 -590
rect 10463 -978 10475 -602
rect 10509 -978 10521 -602
rect 10463 -990 10521 -978
rect 10576 -602 10634 -590
rect 10576 -978 10588 -602
rect 10622 -978 10634 -602
rect 10576 -990 10634 -978
rect 10694 -602 10752 -590
rect 10694 -978 10706 -602
rect 10740 -978 10752 -602
rect 10694 -990 10752 -978
rect 10812 -602 10870 -590
rect 10812 -978 10824 -602
rect 10858 -978 10870 -602
rect 10812 -990 10870 -978
rect 10930 -602 10988 -590
rect 10930 -978 10942 -602
rect 10976 -978 10988 -602
rect 10930 -990 10988 -978
rect 11048 -602 11106 -590
rect 11048 -978 11060 -602
rect 11094 -978 11106 -602
rect 11048 -990 11106 -978
rect 11166 -602 11224 -590
rect 11166 -978 11178 -602
rect 11212 -978 11224 -602
rect 11166 -990 11224 -978
rect 11284 -602 11342 -590
rect 11284 -978 11296 -602
rect 11330 -978 11342 -602
rect 11284 -990 11342 -978
rect 11403 -602 11461 -590
rect 11403 -978 11415 -602
rect 11449 -978 11461 -602
rect 11403 -990 11461 -978
rect 11521 -602 11579 -590
rect 11521 -978 11533 -602
rect 11567 -978 11579 -602
rect 11521 -990 11579 -978
rect 11639 -602 11697 -590
rect 11639 -978 11651 -602
rect 11685 -978 11697 -602
rect 11639 -990 11697 -978
rect 11757 -602 11815 -590
rect 11757 -978 11769 -602
rect 11803 -978 11815 -602
rect 13311 -606 13369 -594
rect 11757 -990 11815 -978
rect 11876 -802 11934 -790
rect 11876 -978 11888 -802
rect 11922 -978 11934 -802
rect 11876 -990 11934 -978
rect 11994 -802 12052 -790
rect 11994 -978 12006 -802
rect 12040 -978 12052 -802
rect 11994 -990 12052 -978
rect 12112 -802 12170 -790
rect 12112 -978 12124 -802
rect 12158 -978 12170 -802
rect 12112 -990 12170 -978
rect 12230 -802 12288 -790
rect 13311 -794 13323 -606
rect 12230 -978 12242 -802
rect 12276 -978 12288 -802
rect 12230 -990 12288 -978
rect 12870 -806 12928 -794
rect 12870 -982 12882 -806
rect 12916 -982 12928 -806
rect 12870 -994 12928 -982
rect 12988 -806 13046 -794
rect 12988 -982 13000 -806
rect 13034 -982 13046 -806
rect 12988 -994 13046 -982
rect 13106 -806 13164 -794
rect 13106 -982 13118 -806
rect 13152 -982 13164 -806
rect 13106 -994 13164 -982
rect 13224 -806 13323 -794
rect 13224 -982 13236 -806
rect 13270 -982 13323 -806
rect 13357 -982 13369 -606
rect 13224 -994 13369 -982
rect 13429 -606 13487 -594
rect 13429 -982 13441 -606
rect 13475 -982 13487 -606
rect 13429 -994 13487 -982
rect 13547 -606 13605 -594
rect 13547 -982 13559 -606
rect 13593 -982 13605 -606
rect 13547 -994 13605 -982
rect 13665 -606 13723 -594
rect 13665 -982 13677 -606
rect 13711 -982 13723 -606
rect 13665 -994 13723 -982
rect 13778 -606 13836 -594
rect 13778 -982 13790 -606
rect 13824 -982 13836 -606
rect 13778 -994 13836 -982
rect 13896 -606 13954 -594
rect 13896 -982 13908 -606
rect 13942 -982 13954 -606
rect 13896 -994 13954 -982
rect 14014 -606 14072 -594
rect 14014 -982 14026 -606
rect 14060 -982 14072 -606
rect 14014 -994 14072 -982
rect 14132 -606 14190 -594
rect 14132 -982 14144 -606
rect 14178 -982 14190 -606
rect 14132 -994 14190 -982
rect 14250 -606 14308 -594
rect 14250 -982 14262 -606
rect 14296 -982 14308 -606
rect 14250 -994 14308 -982
rect 14368 -606 14426 -594
rect 14368 -982 14380 -606
rect 14414 -982 14426 -606
rect 14368 -994 14426 -982
rect 14486 -606 14544 -594
rect 14486 -982 14498 -606
rect 14532 -982 14544 -606
rect 14486 -994 14544 -982
rect 14605 -606 14663 -594
rect 14605 -982 14617 -606
rect 14651 -982 14663 -606
rect 14605 -994 14663 -982
rect 14723 -606 14781 -594
rect 14723 -982 14735 -606
rect 14769 -982 14781 -606
rect 14723 -994 14781 -982
rect 14841 -606 14899 -594
rect 14841 -982 14853 -606
rect 14887 -982 14899 -606
rect 14841 -994 14899 -982
rect 14959 -606 15017 -594
rect 14959 -982 14971 -606
rect 15005 -982 15017 -606
rect 16455 -606 16513 -594
rect 16455 -794 16467 -606
rect 14959 -994 15017 -982
rect 15078 -806 15136 -794
rect 15078 -982 15090 -806
rect 15124 -982 15136 -806
rect 15078 -994 15136 -982
rect 15196 -806 15254 -794
rect 15196 -982 15208 -806
rect 15242 -982 15254 -806
rect 15196 -994 15254 -982
rect 15314 -806 15372 -794
rect 15314 -982 15326 -806
rect 15360 -982 15372 -806
rect 15314 -994 15372 -982
rect 15432 -806 15490 -794
rect 15432 -982 15444 -806
rect 15478 -982 15490 -806
rect 15432 -994 15490 -982
rect 16014 -806 16072 -794
rect 16014 -982 16026 -806
rect 16060 -982 16072 -806
rect 16014 -994 16072 -982
rect 16132 -806 16190 -794
rect 16132 -982 16144 -806
rect 16178 -982 16190 -806
rect 16132 -994 16190 -982
rect 16250 -806 16308 -794
rect 16250 -982 16262 -806
rect 16296 -982 16308 -806
rect 16250 -994 16308 -982
rect 16368 -806 16467 -794
rect 16368 -982 16380 -806
rect 16414 -982 16467 -806
rect 16501 -982 16513 -606
rect 16368 -994 16513 -982
rect 16573 -606 16631 -594
rect 16573 -982 16585 -606
rect 16619 -982 16631 -606
rect 16573 -994 16631 -982
rect 16691 -606 16749 -594
rect 16691 -982 16703 -606
rect 16737 -982 16749 -606
rect 16691 -994 16749 -982
rect 16809 -606 16867 -594
rect 16809 -982 16821 -606
rect 16855 -982 16867 -606
rect 16809 -994 16867 -982
rect 16922 -606 16980 -594
rect 16922 -982 16934 -606
rect 16968 -982 16980 -606
rect 16922 -994 16980 -982
rect 17040 -606 17098 -594
rect 17040 -982 17052 -606
rect 17086 -982 17098 -606
rect 17040 -994 17098 -982
rect 17158 -606 17216 -594
rect 17158 -982 17170 -606
rect 17204 -982 17216 -606
rect 17158 -994 17216 -982
rect 17276 -606 17334 -594
rect 17276 -982 17288 -606
rect 17322 -982 17334 -606
rect 17276 -994 17334 -982
rect 17394 -606 17452 -594
rect 17394 -982 17406 -606
rect 17440 -982 17452 -606
rect 17394 -994 17452 -982
rect 17512 -606 17570 -594
rect 17512 -982 17524 -606
rect 17558 -982 17570 -606
rect 17512 -994 17570 -982
rect 17630 -606 17688 -594
rect 17630 -982 17642 -606
rect 17676 -982 17688 -606
rect 17630 -994 17688 -982
rect 17749 -606 17807 -594
rect 17749 -982 17761 -606
rect 17795 -982 17807 -606
rect 17749 -994 17807 -982
rect 17867 -606 17925 -594
rect 17867 -982 17879 -606
rect 17913 -982 17925 -606
rect 17867 -994 17925 -982
rect 17985 -606 18043 -594
rect 17985 -982 17997 -606
rect 18031 -982 18043 -606
rect 17985 -994 18043 -982
rect 18103 -606 18161 -594
rect 18103 -982 18115 -606
rect 18149 -982 18161 -606
rect 19587 -602 19645 -590
rect 19587 -790 19599 -602
rect 18103 -994 18161 -982
rect 18222 -806 18280 -794
rect 18222 -982 18234 -806
rect 18268 -982 18280 -806
rect 18222 -994 18280 -982
rect 18340 -806 18398 -794
rect 18340 -982 18352 -806
rect 18386 -982 18398 -806
rect 18340 -994 18398 -982
rect 18458 -806 18516 -794
rect 18458 -982 18470 -806
rect 18504 -982 18516 -806
rect 18458 -994 18516 -982
rect 18576 -806 18634 -794
rect 18576 -982 18588 -806
rect 18622 -982 18634 -806
rect 18576 -994 18634 -982
rect 19146 -802 19204 -790
rect 19146 -978 19158 -802
rect 19192 -978 19204 -802
rect 19146 -990 19204 -978
rect 19264 -802 19322 -790
rect 19264 -978 19276 -802
rect 19310 -978 19322 -802
rect 19264 -990 19322 -978
rect 19382 -802 19440 -790
rect 19382 -978 19394 -802
rect 19428 -978 19440 -802
rect 19382 -990 19440 -978
rect 19500 -802 19599 -790
rect 19500 -978 19512 -802
rect 19546 -978 19599 -802
rect 19633 -978 19645 -602
rect 19500 -990 19645 -978
rect 19705 -602 19763 -590
rect 19705 -978 19717 -602
rect 19751 -978 19763 -602
rect 19705 -990 19763 -978
rect 19823 -602 19881 -590
rect 19823 -978 19835 -602
rect 19869 -978 19881 -602
rect 19823 -990 19881 -978
rect 19941 -602 19999 -590
rect 19941 -978 19953 -602
rect 19987 -978 19999 -602
rect 19941 -990 19999 -978
rect 20054 -602 20112 -590
rect 20054 -978 20066 -602
rect 20100 -978 20112 -602
rect 20054 -990 20112 -978
rect 20172 -602 20230 -590
rect 20172 -978 20184 -602
rect 20218 -978 20230 -602
rect 20172 -990 20230 -978
rect 20290 -602 20348 -590
rect 20290 -978 20302 -602
rect 20336 -978 20348 -602
rect 20290 -990 20348 -978
rect 20408 -602 20466 -590
rect 20408 -978 20420 -602
rect 20454 -978 20466 -602
rect 20408 -990 20466 -978
rect 20526 -602 20584 -590
rect 20526 -978 20538 -602
rect 20572 -978 20584 -602
rect 20526 -990 20584 -978
rect 20644 -602 20702 -590
rect 20644 -978 20656 -602
rect 20690 -978 20702 -602
rect 20644 -990 20702 -978
rect 20762 -602 20820 -590
rect 20762 -978 20774 -602
rect 20808 -978 20820 -602
rect 20762 -990 20820 -978
rect 20881 -602 20939 -590
rect 20881 -978 20893 -602
rect 20927 -978 20939 -602
rect 20881 -990 20939 -978
rect 20999 -602 21057 -590
rect 20999 -978 21011 -602
rect 21045 -978 21057 -602
rect 20999 -990 21057 -978
rect 21117 -602 21175 -590
rect 21117 -978 21129 -602
rect 21163 -978 21175 -602
rect 21117 -990 21175 -978
rect 21235 -602 21293 -590
rect 21235 -978 21247 -602
rect 21281 -978 21293 -602
rect 22731 -602 22789 -590
rect 22731 -790 22743 -602
rect 21235 -990 21293 -978
rect 21354 -802 21412 -790
rect 21354 -978 21366 -802
rect 21400 -978 21412 -802
rect 21354 -990 21412 -978
rect 21472 -802 21530 -790
rect 21472 -978 21484 -802
rect 21518 -978 21530 -802
rect 21472 -990 21530 -978
rect 21590 -802 21648 -790
rect 21590 -978 21602 -802
rect 21636 -978 21648 -802
rect 21590 -990 21648 -978
rect 21708 -802 21766 -790
rect 21708 -978 21720 -802
rect 21754 -978 21766 -802
rect 21708 -990 21766 -978
rect 22290 -802 22348 -790
rect 22290 -978 22302 -802
rect 22336 -978 22348 -802
rect 22290 -990 22348 -978
rect 22408 -802 22466 -790
rect 22408 -978 22420 -802
rect 22454 -978 22466 -802
rect 22408 -990 22466 -978
rect 22526 -802 22584 -790
rect 22526 -978 22538 -802
rect 22572 -978 22584 -802
rect 22526 -990 22584 -978
rect 22644 -802 22743 -790
rect 22644 -978 22656 -802
rect 22690 -978 22743 -802
rect 22777 -978 22789 -602
rect 22644 -990 22789 -978
rect 22849 -602 22907 -590
rect 22849 -978 22861 -602
rect 22895 -978 22907 -602
rect 22849 -990 22907 -978
rect 22967 -602 23025 -590
rect 22967 -978 22979 -602
rect 23013 -978 23025 -602
rect 22967 -990 23025 -978
rect 23085 -602 23143 -590
rect 23085 -978 23097 -602
rect 23131 -978 23143 -602
rect 23085 -990 23143 -978
rect 23198 -602 23256 -590
rect 23198 -978 23210 -602
rect 23244 -978 23256 -602
rect 23198 -990 23256 -978
rect 23316 -602 23374 -590
rect 23316 -978 23328 -602
rect 23362 -978 23374 -602
rect 23316 -990 23374 -978
rect 23434 -602 23492 -590
rect 23434 -978 23446 -602
rect 23480 -978 23492 -602
rect 23434 -990 23492 -978
rect 23552 -602 23610 -590
rect 23552 -978 23564 -602
rect 23598 -978 23610 -602
rect 23552 -990 23610 -978
rect 23670 -602 23728 -590
rect 23670 -978 23682 -602
rect 23716 -978 23728 -602
rect 23670 -990 23728 -978
rect 23788 -602 23846 -590
rect 23788 -978 23800 -602
rect 23834 -978 23846 -602
rect 23788 -990 23846 -978
rect 23906 -602 23964 -590
rect 23906 -978 23918 -602
rect 23952 -978 23964 -602
rect 23906 -990 23964 -978
rect 24025 -602 24083 -590
rect 24025 -978 24037 -602
rect 24071 -978 24083 -602
rect 24025 -990 24083 -978
rect 24143 -602 24201 -590
rect 24143 -978 24155 -602
rect 24189 -978 24201 -602
rect 24143 -990 24201 -978
rect 24261 -602 24319 -590
rect 24261 -978 24273 -602
rect 24307 -978 24319 -602
rect 24261 -990 24319 -978
rect 24379 -602 24437 -590
rect 24379 -978 24391 -602
rect 24425 -978 24437 -602
rect 24379 -990 24437 -978
rect 24498 -802 24556 -790
rect 24498 -978 24510 -802
rect 24544 -978 24556 -802
rect 24498 -990 24556 -978
rect 24616 -802 24674 -790
rect 24616 -978 24628 -802
rect 24662 -978 24674 -802
rect 24616 -990 24674 -978
rect 24734 -802 24792 -790
rect 24734 -978 24746 -802
rect 24780 -978 24792 -802
rect 24734 -990 24792 -978
rect 24852 -802 24910 -790
rect 24852 -978 24864 -802
rect 24898 -978 24910 -802
rect 24852 -990 24910 -978
rect 679 -3338 737 -3326
rect 679 -3526 691 -3338
rect 238 -3538 296 -3526
rect 238 -3714 250 -3538
rect 284 -3714 296 -3538
rect 238 -3726 296 -3714
rect 356 -3538 414 -3526
rect 356 -3714 368 -3538
rect 402 -3714 414 -3538
rect 356 -3726 414 -3714
rect 474 -3538 532 -3526
rect 474 -3714 486 -3538
rect 520 -3714 532 -3538
rect 474 -3726 532 -3714
rect 592 -3538 691 -3526
rect 592 -3714 604 -3538
rect 638 -3714 691 -3538
rect 725 -3714 737 -3338
rect 592 -3726 737 -3714
rect 797 -3338 855 -3326
rect 797 -3714 809 -3338
rect 843 -3714 855 -3338
rect 797 -3726 855 -3714
rect 915 -3338 973 -3326
rect 915 -3714 927 -3338
rect 961 -3714 973 -3338
rect 915 -3726 973 -3714
rect 1033 -3338 1091 -3326
rect 1033 -3714 1045 -3338
rect 1079 -3714 1091 -3338
rect 1033 -3726 1091 -3714
rect 1146 -3338 1204 -3326
rect 1146 -3714 1158 -3338
rect 1192 -3714 1204 -3338
rect 1146 -3726 1204 -3714
rect 1264 -3338 1322 -3326
rect 1264 -3714 1276 -3338
rect 1310 -3714 1322 -3338
rect 1264 -3726 1322 -3714
rect 1382 -3338 1440 -3326
rect 1382 -3714 1394 -3338
rect 1428 -3714 1440 -3338
rect 1382 -3726 1440 -3714
rect 1500 -3338 1558 -3326
rect 1500 -3714 1512 -3338
rect 1546 -3714 1558 -3338
rect 1500 -3726 1558 -3714
rect 1618 -3338 1676 -3326
rect 1618 -3714 1630 -3338
rect 1664 -3714 1676 -3338
rect 1618 -3726 1676 -3714
rect 1736 -3338 1794 -3326
rect 1736 -3714 1748 -3338
rect 1782 -3714 1794 -3338
rect 1736 -3726 1794 -3714
rect 1854 -3338 1912 -3326
rect 1854 -3714 1866 -3338
rect 1900 -3714 1912 -3338
rect 1854 -3726 1912 -3714
rect 1973 -3338 2031 -3326
rect 1973 -3714 1985 -3338
rect 2019 -3714 2031 -3338
rect 1973 -3726 2031 -3714
rect 2091 -3338 2149 -3326
rect 2091 -3714 2103 -3338
rect 2137 -3714 2149 -3338
rect 2091 -3726 2149 -3714
rect 2209 -3338 2267 -3326
rect 2209 -3714 2221 -3338
rect 2255 -3714 2267 -3338
rect 2209 -3726 2267 -3714
rect 2327 -3338 2385 -3326
rect 2327 -3714 2339 -3338
rect 2373 -3714 2385 -3338
rect 3823 -3338 3881 -3326
rect 3823 -3526 3835 -3338
rect 2327 -3726 2385 -3714
rect 2446 -3538 2504 -3526
rect 2446 -3714 2458 -3538
rect 2492 -3714 2504 -3538
rect 2446 -3726 2504 -3714
rect 2564 -3538 2622 -3526
rect 2564 -3714 2576 -3538
rect 2610 -3714 2622 -3538
rect 2564 -3726 2622 -3714
rect 2682 -3538 2740 -3526
rect 2682 -3714 2694 -3538
rect 2728 -3714 2740 -3538
rect 2682 -3726 2740 -3714
rect 2800 -3538 2858 -3526
rect 2800 -3714 2812 -3538
rect 2846 -3714 2858 -3538
rect 2800 -3726 2858 -3714
rect 3382 -3538 3440 -3526
rect 3382 -3714 3394 -3538
rect 3428 -3714 3440 -3538
rect 3382 -3726 3440 -3714
rect 3500 -3538 3558 -3526
rect 3500 -3714 3512 -3538
rect 3546 -3714 3558 -3538
rect 3500 -3726 3558 -3714
rect 3618 -3538 3676 -3526
rect 3618 -3714 3630 -3538
rect 3664 -3714 3676 -3538
rect 3618 -3726 3676 -3714
rect 3736 -3538 3835 -3526
rect 3736 -3714 3748 -3538
rect 3782 -3714 3835 -3538
rect 3869 -3714 3881 -3338
rect 3736 -3726 3881 -3714
rect 3941 -3338 3999 -3326
rect 3941 -3714 3953 -3338
rect 3987 -3714 3999 -3338
rect 3941 -3726 3999 -3714
rect 4059 -3338 4117 -3326
rect 4059 -3714 4071 -3338
rect 4105 -3714 4117 -3338
rect 4059 -3726 4117 -3714
rect 4177 -3338 4235 -3326
rect 4177 -3714 4189 -3338
rect 4223 -3714 4235 -3338
rect 4177 -3726 4235 -3714
rect 4290 -3338 4348 -3326
rect 4290 -3714 4302 -3338
rect 4336 -3714 4348 -3338
rect 4290 -3726 4348 -3714
rect 4408 -3338 4466 -3326
rect 4408 -3714 4420 -3338
rect 4454 -3714 4466 -3338
rect 4408 -3726 4466 -3714
rect 4526 -3338 4584 -3326
rect 4526 -3714 4538 -3338
rect 4572 -3714 4584 -3338
rect 4526 -3726 4584 -3714
rect 4644 -3338 4702 -3326
rect 4644 -3714 4656 -3338
rect 4690 -3714 4702 -3338
rect 4644 -3726 4702 -3714
rect 4762 -3338 4820 -3326
rect 4762 -3714 4774 -3338
rect 4808 -3714 4820 -3338
rect 4762 -3726 4820 -3714
rect 4880 -3338 4938 -3326
rect 4880 -3714 4892 -3338
rect 4926 -3714 4938 -3338
rect 4880 -3726 4938 -3714
rect 4998 -3338 5056 -3326
rect 4998 -3714 5010 -3338
rect 5044 -3714 5056 -3338
rect 4998 -3726 5056 -3714
rect 5117 -3338 5175 -3326
rect 5117 -3714 5129 -3338
rect 5163 -3714 5175 -3338
rect 5117 -3726 5175 -3714
rect 5235 -3338 5293 -3326
rect 5235 -3714 5247 -3338
rect 5281 -3714 5293 -3338
rect 5235 -3726 5293 -3714
rect 5353 -3338 5411 -3326
rect 5353 -3714 5365 -3338
rect 5399 -3714 5411 -3338
rect 5353 -3726 5411 -3714
rect 5471 -3338 5529 -3326
rect 5471 -3714 5483 -3338
rect 5517 -3714 5529 -3338
rect 6955 -3334 7013 -3322
rect 6955 -3522 6967 -3334
rect 5471 -3726 5529 -3714
rect 5590 -3538 5648 -3526
rect 5590 -3714 5602 -3538
rect 5636 -3714 5648 -3538
rect 5590 -3726 5648 -3714
rect 5708 -3538 5766 -3526
rect 5708 -3714 5720 -3538
rect 5754 -3714 5766 -3538
rect 5708 -3726 5766 -3714
rect 5826 -3538 5884 -3526
rect 5826 -3714 5838 -3538
rect 5872 -3714 5884 -3538
rect 5826 -3726 5884 -3714
rect 5944 -3538 6002 -3526
rect 5944 -3714 5956 -3538
rect 5990 -3714 6002 -3538
rect 5944 -3726 6002 -3714
rect 6514 -3534 6572 -3522
rect 6514 -3710 6526 -3534
rect 6560 -3710 6572 -3534
rect 6514 -3722 6572 -3710
rect 6632 -3534 6690 -3522
rect 6632 -3710 6644 -3534
rect 6678 -3710 6690 -3534
rect 6632 -3722 6690 -3710
rect 6750 -3534 6808 -3522
rect 6750 -3710 6762 -3534
rect 6796 -3710 6808 -3534
rect 6750 -3722 6808 -3710
rect 6868 -3534 6967 -3522
rect 6868 -3710 6880 -3534
rect 6914 -3710 6967 -3534
rect 7001 -3710 7013 -3334
rect 6868 -3722 7013 -3710
rect 7073 -3334 7131 -3322
rect 7073 -3710 7085 -3334
rect 7119 -3710 7131 -3334
rect 7073 -3722 7131 -3710
rect 7191 -3334 7249 -3322
rect 7191 -3710 7203 -3334
rect 7237 -3710 7249 -3334
rect 7191 -3722 7249 -3710
rect 7309 -3334 7367 -3322
rect 7309 -3710 7321 -3334
rect 7355 -3710 7367 -3334
rect 7309 -3722 7367 -3710
rect 7422 -3334 7480 -3322
rect 7422 -3710 7434 -3334
rect 7468 -3710 7480 -3334
rect 7422 -3722 7480 -3710
rect 7540 -3334 7598 -3322
rect 7540 -3710 7552 -3334
rect 7586 -3710 7598 -3334
rect 7540 -3722 7598 -3710
rect 7658 -3334 7716 -3322
rect 7658 -3710 7670 -3334
rect 7704 -3710 7716 -3334
rect 7658 -3722 7716 -3710
rect 7776 -3334 7834 -3322
rect 7776 -3710 7788 -3334
rect 7822 -3710 7834 -3334
rect 7776 -3722 7834 -3710
rect 7894 -3334 7952 -3322
rect 7894 -3710 7906 -3334
rect 7940 -3710 7952 -3334
rect 7894 -3722 7952 -3710
rect 8012 -3334 8070 -3322
rect 8012 -3710 8024 -3334
rect 8058 -3710 8070 -3334
rect 8012 -3722 8070 -3710
rect 8130 -3334 8188 -3322
rect 8130 -3710 8142 -3334
rect 8176 -3710 8188 -3334
rect 8130 -3722 8188 -3710
rect 8249 -3334 8307 -3322
rect 8249 -3710 8261 -3334
rect 8295 -3710 8307 -3334
rect 8249 -3722 8307 -3710
rect 8367 -3334 8425 -3322
rect 8367 -3710 8379 -3334
rect 8413 -3710 8425 -3334
rect 8367 -3722 8425 -3710
rect 8485 -3334 8543 -3322
rect 8485 -3710 8497 -3334
rect 8531 -3710 8543 -3334
rect 8485 -3722 8543 -3710
rect 8603 -3334 8661 -3322
rect 8603 -3710 8615 -3334
rect 8649 -3710 8661 -3334
rect 10099 -3334 10157 -3322
rect 10099 -3522 10111 -3334
rect 8603 -3722 8661 -3710
rect 8722 -3534 8780 -3522
rect 8722 -3710 8734 -3534
rect 8768 -3710 8780 -3534
rect 8722 -3722 8780 -3710
rect 8840 -3534 8898 -3522
rect 8840 -3710 8852 -3534
rect 8886 -3710 8898 -3534
rect 8840 -3722 8898 -3710
rect 8958 -3534 9016 -3522
rect 8958 -3710 8970 -3534
rect 9004 -3710 9016 -3534
rect 8958 -3722 9016 -3710
rect 9076 -3534 9134 -3522
rect 9076 -3710 9088 -3534
rect 9122 -3710 9134 -3534
rect 9076 -3722 9134 -3710
rect 9658 -3534 9716 -3522
rect 9658 -3710 9670 -3534
rect 9704 -3710 9716 -3534
rect 9658 -3722 9716 -3710
rect 9776 -3534 9834 -3522
rect 9776 -3710 9788 -3534
rect 9822 -3710 9834 -3534
rect 9776 -3722 9834 -3710
rect 9894 -3534 9952 -3522
rect 9894 -3710 9906 -3534
rect 9940 -3710 9952 -3534
rect 9894 -3722 9952 -3710
rect 10012 -3534 10111 -3522
rect 10012 -3710 10024 -3534
rect 10058 -3710 10111 -3534
rect 10145 -3710 10157 -3334
rect 10012 -3722 10157 -3710
rect 10217 -3334 10275 -3322
rect 10217 -3710 10229 -3334
rect 10263 -3710 10275 -3334
rect 10217 -3722 10275 -3710
rect 10335 -3334 10393 -3322
rect 10335 -3710 10347 -3334
rect 10381 -3710 10393 -3334
rect 10335 -3722 10393 -3710
rect 10453 -3334 10511 -3322
rect 10453 -3710 10465 -3334
rect 10499 -3710 10511 -3334
rect 10453 -3722 10511 -3710
rect 10566 -3334 10624 -3322
rect 10566 -3710 10578 -3334
rect 10612 -3710 10624 -3334
rect 10566 -3722 10624 -3710
rect 10684 -3334 10742 -3322
rect 10684 -3710 10696 -3334
rect 10730 -3710 10742 -3334
rect 10684 -3722 10742 -3710
rect 10802 -3334 10860 -3322
rect 10802 -3710 10814 -3334
rect 10848 -3710 10860 -3334
rect 10802 -3722 10860 -3710
rect 10920 -3334 10978 -3322
rect 10920 -3710 10932 -3334
rect 10966 -3710 10978 -3334
rect 10920 -3722 10978 -3710
rect 11038 -3334 11096 -3322
rect 11038 -3710 11050 -3334
rect 11084 -3710 11096 -3334
rect 11038 -3722 11096 -3710
rect 11156 -3334 11214 -3322
rect 11156 -3710 11168 -3334
rect 11202 -3710 11214 -3334
rect 11156 -3722 11214 -3710
rect 11274 -3334 11332 -3322
rect 11274 -3710 11286 -3334
rect 11320 -3710 11332 -3334
rect 11274 -3722 11332 -3710
rect 11393 -3334 11451 -3322
rect 11393 -3710 11405 -3334
rect 11439 -3710 11451 -3334
rect 11393 -3722 11451 -3710
rect 11511 -3334 11569 -3322
rect 11511 -3710 11523 -3334
rect 11557 -3710 11569 -3334
rect 11511 -3722 11569 -3710
rect 11629 -3334 11687 -3322
rect 11629 -3710 11641 -3334
rect 11675 -3710 11687 -3334
rect 11629 -3722 11687 -3710
rect 11747 -3334 11805 -3322
rect 11747 -3710 11759 -3334
rect 11793 -3710 11805 -3334
rect 13301 -3338 13359 -3326
rect 11747 -3722 11805 -3710
rect 11866 -3534 11924 -3522
rect 11866 -3710 11878 -3534
rect 11912 -3710 11924 -3534
rect 11866 -3722 11924 -3710
rect 11984 -3534 12042 -3522
rect 11984 -3710 11996 -3534
rect 12030 -3710 12042 -3534
rect 11984 -3722 12042 -3710
rect 12102 -3534 12160 -3522
rect 12102 -3710 12114 -3534
rect 12148 -3710 12160 -3534
rect 12102 -3722 12160 -3710
rect 12220 -3534 12278 -3522
rect 13301 -3526 13313 -3338
rect 12220 -3710 12232 -3534
rect 12266 -3710 12278 -3534
rect 12220 -3722 12278 -3710
rect 12860 -3538 12918 -3526
rect 12860 -3714 12872 -3538
rect 12906 -3714 12918 -3538
rect 12860 -3726 12918 -3714
rect 12978 -3538 13036 -3526
rect 12978 -3714 12990 -3538
rect 13024 -3714 13036 -3538
rect 12978 -3726 13036 -3714
rect 13096 -3538 13154 -3526
rect 13096 -3714 13108 -3538
rect 13142 -3714 13154 -3538
rect 13096 -3726 13154 -3714
rect 13214 -3538 13313 -3526
rect 13214 -3714 13226 -3538
rect 13260 -3714 13313 -3538
rect 13347 -3714 13359 -3338
rect 13214 -3726 13359 -3714
rect 13419 -3338 13477 -3326
rect 13419 -3714 13431 -3338
rect 13465 -3714 13477 -3338
rect 13419 -3726 13477 -3714
rect 13537 -3338 13595 -3326
rect 13537 -3714 13549 -3338
rect 13583 -3714 13595 -3338
rect 13537 -3726 13595 -3714
rect 13655 -3338 13713 -3326
rect 13655 -3714 13667 -3338
rect 13701 -3714 13713 -3338
rect 13655 -3726 13713 -3714
rect 13768 -3338 13826 -3326
rect 13768 -3714 13780 -3338
rect 13814 -3714 13826 -3338
rect 13768 -3726 13826 -3714
rect 13886 -3338 13944 -3326
rect 13886 -3714 13898 -3338
rect 13932 -3714 13944 -3338
rect 13886 -3726 13944 -3714
rect 14004 -3338 14062 -3326
rect 14004 -3714 14016 -3338
rect 14050 -3714 14062 -3338
rect 14004 -3726 14062 -3714
rect 14122 -3338 14180 -3326
rect 14122 -3714 14134 -3338
rect 14168 -3714 14180 -3338
rect 14122 -3726 14180 -3714
rect 14240 -3338 14298 -3326
rect 14240 -3714 14252 -3338
rect 14286 -3714 14298 -3338
rect 14240 -3726 14298 -3714
rect 14358 -3338 14416 -3326
rect 14358 -3714 14370 -3338
rect 14404 -3714 14416 -3338
rect 14358 -3726 14416 -3714
rect 14476 -3338 14534 -3326
rect 14476 -3714 14488 -3338
rect 14522 -3714 14534 -3338
rect 14476 -3726 14534 -3714
rect 14595 -3338 14653 -3326
rect 14595 -3714 14607 -3338
rect 14641 -3714 14653 -3338
rect 14595 -3726 14653 -3714
rect 14713 -3338 14771 -3326
rect 14713 -3714 14725 -3338
rect 14759 -3714 14771 -3338
rect 14713 -3726 14771 -3714
rect 14831 -3338 14889 -3326
rect 14831 -3714 14843 -3338
rect 14877 -3714 14889 -3338
rect 14831 -3726 14889 -3714
rect 14949 -3338 15007 -3326
rect 14949 -3714 14961 -3338
rect 14995 -3714 15007 -3338
rect 16445 -3338 16503 -3326
rect 16445 -3526 16457 -3338
rect 14949 -3726 15007 -3714
rect 15068 -3538 15126 -3526
rect 15068 -3714 15080 -3538
rect 15114 -3714 15126 -3538
rect 15068 -3726 15126 -3714
rect 15186 -3538 15244 -3526
rect 15186 -3714 15198 -3538
rect 15232 -3714 15244 -3538
rect 15186 -3726 15244 -3714
rect 15304 -3538 15362 -3526
rect 15304 -3714 15316 -3538
rect 15350 -3714 15362 -3538
rect 15304 -3726 15362 -3714
rect 15422 -3538 15480 -3526
rect 15422 -3714 15434 -3538
rect 15468 -3714 15480 -3538
rect 15422 -3726 15480 -3714
rect 16004 -3538 16062 -3526
rect 16004 -3714 16016 -3538
rect 16050 -3714 16062 -3538
rect 16004 -3726 16062 -3714
rect 16122 -3538 16180 -3526
rect 16122 -3714 16134 -3538
rect 16168 -3714 16180 -3538
rect 16122 -3726 16180 -3714
rect 16240 -3538 16298 -3526
rect 16240 -3714 16252 -3538
rect 16286 -3714 16298 -3538
rect 16240 -3726 16298 -3714
rect 16358 -3538 16457 -3526
rect 16358 -3714 16370 -3538
rect 16404 -3714 16457 -3538
rect 16491 -3714 16503 -3338
rect 16358 -3726 16503 -3714
rect 16563 -3338 16621 -3326
rect 16563 -3714 16575 -3338
rect 16609 -3714 16621 -3338
rect 16563 -3726 16621 -3714
rect 16681 -3338 16739 -3326
rect 16681 -3714 16693 -3338
rect 16727 -3714 16739 -3338
rect 16681 -3726 16739 -3714
rect 16799 -3338 16857 -3326
rect 16799 -3714 16811 -3338
rect 16845 -3714 16857 -3338
rect 16799 -3726 16857 -3714
rect 16912 -3338 16970 -3326
rect 16912 -3714 16924 -3338
rect 16958 -3714 16970 -3338
rect 16912 -3726 16970 -3714
rect 17030 -3338 17088 -3326
rect 17030 -3714 17042 -3338
rect 17076 -3714 17088 -3338
rect 17030 -3726 17088 -3714
rect 17148 -3338 17206 -3326
rect 17148 -3714 17160 -3338
rect 17194 -3714 17206 -3338
rect 17148 -3726 17206 -3714
rect 17266 -3338 17324 -3326
rect 17266 -3714 17278 -3338
rect 17312 -3714 17324 -3338
rect 17266 -3726 17324 -3714
rect 17384 -3338 17442 -3326
rect 17384 -3714 17396 -3338
rect 17430 -3714 17442 -3338
rect 17384 -3726 17442 -3714
rect 17502 -3338 17560 -3326
rect 17502 -3714 17514 -3338
rect 17548 -3714 17560 -3338
rect 17502 -3726 17560 -3714
rect 17620 -3338 17678 -3326
rect 17620 -3714 17632 -3338
rect 17666 -3714 17678 -3338
rect 17620 -3726 17678 -3714
rect 17739 -3338 17797 -3326
rect 17739 -3714 17751 -3338
rect 17785 -3714 17797 -3338
rect 17739 -3726 17797 -3714
rect 17857 -3338 17915 -3326
rect 17857 -3714 17869 -3338
rect 17903 -3714 17915 -3338
rect 17857 -3726 17915 -3714
rect 17975 -3338 18033 -3326
rect 17975 -3714 17987 -3338
rect 18021 -3714 18033 -3338
rect 17975 -3726 18033 -3714
rect 18093 -3338 18151 -3326
rect 18093 -3714 18105 -3338
rect 18139 -3714 18151 -3338
rect 19577 -3334 19635 -3322
rect 19577 -3522 19589 -3334
rect 18093 -3726 18151 -3714
rect 18212 -3538 18270 -3526
rect 18212 -3714 18224 -3538
rect 18258 -3714 18270 -3538
rect 18212 -3726 18270 -3714
rect 18330 -3538 18388 -3526
rect 18330 -3714 18342 -3538
rect 18376 -3714 18388 -3538
rect 18330 -3726 18388 -3714
rect 18448 -3538 18506 -3526
rect 18448 -3714 18460 -3538
rect 18494 -3714 18506 -3538
rect 18448 -3726 18506 -3714
rect 18566 -3538 18624 -3526
rect 18566 -3714 18578 -3538
rect 18612 -3714 18624 -3538
rect 18566 -3726 18624 -3714
rect 19136 -3534 19194 -3522
rect 19136 -3710 19148 -3534
rect 19182 -3710 19194 -3534
rect 19136 -3722 19194 -3710
rect 19254 -3534 19312 -3522
rect 19254 -3710 19266 -3534
rect 19300 -3710 19312 -3534
rect 19254 -3722 19312 -3710
rect 19372 -3534 19430 -3522
rect 19372 -3710 19384 -3534
rect 19418 -3710 19430 -3534
rect 19372 -3722 19430 -3710
rect 19490 -3534 19589 -3522
rect 19490 -3710 19502 -3534
rect 19536 -3710 19589 -3534
rect 19623 -3710 19635 -3334
rect 19490 -3722 19635 -3710
rect 19695 -3334 19753 -3322
rect 19695 -3710 19707 -3334
rect 19741 -3710 19753 -3334
rect 19695 -3722 19753 -3710
rect 19813 -3334 19871 -3322
rect 19813 -3710 19825 -3334
rect 19859 -3710 19871 -3334
rect 19813 -3722 19871 -3710
rect 19931 -3334 19989 -3322
rect 19931 -3710 19943 -3334
rect 19977 -3710 19989 -3334
rect 19931 -3722 19989 -3710
rect 20044 -3334 20102 -3322
rect 20044 -3710 20056 -3334
rect 20090 -3710 20102 -3334
rect 20044 -3722 20102 -3710
rect 20162 -3334 20220 -3322
rect 20162 -3710 20174 -3334
rect 20208 -3710 20220 -3334
rect 20162 -3722 20220 -3710
rect 20280 -3334 20338 -3322
rect 20280 -3710 20292 -3334
rect 20326 -3710 20338 -3334
rect 20280 -3722 20338 -3710
rect 20398 -3334 20456 -3322
rect 20398 -3710 20410 -3334
rect 20444 -3710 20456 -3334
rect 20398 -3722 20456 -3710
rect 20516 -3334 20574 -3322
rect 20516 -3710 20528 -3334
rect 20562 -3710 20574 -3334
rect 20516 -3722 20574 -3710
rect 20634 -3334 20692 -3322
rect 20634 -3710 20646 -3334
rect 20680 -3710 20692 -3334
rect 20634 -3722 20692 -3710
rect 20752 -3334 20810 -3322
rect 20752 -3710 20764 -3334
rect 20798 -3710 20810 -3334
rect 20752 -3722 20810 -3710
rect 20871 -3334 20929 -3322
rect 20871 -3710 20883 -3334
rect 20917 -3710 20929 -3334
rect 20871 -3722 20929 -3710
rect 20989 -3334 21047 -3322
rect 20989 -3710 21001 -3334
rect 21035 -3710 21047 -3334
rect 20989 -3722 21047 -3710
rect 21107 -3334 21165 -3322
rect 21107 -3710 21119 -3334
rect 21153 -3710 21165 -3334
rect 21107 -3722 21165 -3710
rect 21225 -3334 21283 -3322
rect 21225 -3710 21237 -3334
rect 21271 -3710 21283 -3334
rect 22721 -3334 22779 -3322
rect 22721 -3522 22733 -3334
rect 21225 -3722 21283 -3710
rect 21344 -3534 21402 -3522
rect 21344 -3710 21356 -3534
rect 21390 -3710 21402 -3534
rect 21344 -3722 21402 -3710
rect 21462 -3534 21520 -3522
rect 21462 -3710 21474 -3534
rect 21508 -3710 21520 -3534
rect 21462 -3722 21520 -3710
rect 21580 -3534 21638 -3522
rect 21580 -3710 21592 -3534
rect 21626 -3710 21638 -3534
rect 21580 -3722 21638 -3710
rect 21698 -3534 21756 -3522
rect 21698 -3710 21710 -3534
rect 21744 -3710 21756 -3534
rect 21698 -3722 21756 -3710
rect 22280 -3534 22338 -3522
rect 22280 -3710 22292 -3534
rect 22326 -3710 22338 -3534
rect 22280 -3722 22338 -3710
rect 22398 -3534 22456 -3522
rect 22398 -3710 22410 -3534
rect 22444 -3710 22456 -3534
rect 22398 -3722 22456 -3710
rect 22516 -3534 22574 -3522
rect 22516 -3710 22528 -3534
rect 22562 -3710 22574 -3534
rect 22516 -3722 22574 -3710
rect 22634 -3534 22733 -3522
rect 22634 -3710 22646 -3534
rect 22680 -3710 22733 -3534
rect 22767 -3710 22779 -3334
rect 22634 -3722 22779 -3710
rect 22839 -3334 22897 -3322
rect 22839 -3710 22851 -3334
rect 22885 -3710 22897 -3334
rect 22839 -3722 22897 -3710
rect 22957 -3334 23015 -3322
rect 22957 -3710 22969 -3334
rect 23003 -3710 23015 -3334
rect 22957 -3722 23015 -3710
rect 23075 -3334 23133 -3322
rect 23075 -3710 23087 -3334
rect 23121 -3710 23133 -3334
rect 23075 -3722 23133 -3710
rect 23188 -3334 23246 -3322
rect 23188 -3710 23200 -3334
rect 23234 -3710 23246 -3334
rect 23188 -3722 23246 -3710
rect 23306 -3334 23364 -3322
rect 23306 -3710 23318 -3334
rect 23352 -3710 23364 -3334
rect 23306 -3722 23364 -3710
rect 23424 -3334 23482 -3322
rect 23424 -3710 23436 -3334
rect 23470 -3710 23482 -3334
rect 23424 -3722 23482 -3710
rect 23542 -3334 23600 -3322
rect 23542 -3710 23554 -3334
rect 23588 -3710 23600 -3334
rect 23542 -3722 23600 -3710
rect 23660 -3334 23718 -3322
rect 23660 -3710 23672 -3334
rect 23706 -3710 23718 -3334
rect 23660 -3722 23718 -3710
rect 23778 -3334 23836 -3322
rect 23778 -3710 23790 -3334
rect 23824 -3710 23836 -3334
rect 23778 -3722 23836 -3710
rect 23896 -3334 23954 -3322
rect 23896 -3710 23908 -3334
rect 23942 -3710 23954 -3334
rect 23896 -3722 23954 -3710
rect 24015 -3334 24073 -3322
rect 24015 -3710 24027 -3334
rect 24061 -3710 24073 -3334
rect 24015 -3722 24073 -3710
rect 24133 -3334 24191 -3322
rect 24133 -3710 24145 -3334
rect 24179 -3710 24191 -3334
rect 24133 -3722 24191 -3710
rect 24251 -3334 24309 -3322
rect 24251 -3710 24263 -3334
rect 24297 -3710 24309 -3334
rect 24251 -3722 24309 -3710
rect 24369 -3334 24427 -3322
rect 24369 -3710 24381 -3334
rect 24415 -3710 24427 -3334
rect 24369 -3722 24427 -3710
rect 24488 -3534 24546 -3522
rect 24488 -3710 24500 -3534
rect 24534 -3710 24546 -3534
rect 24488 -3722 24546 -3710
rect 24606 -3534 24664 -3522
rect 24606 -3710 24618 -3534
rect 24652 -3710 24664 -3534
rect 24606 -3722 24664 -3710
rect 24724 -3534 24782 -3522
rect 24724 -3710 24736 -3534
rect 24770 -3710 24782 -3534
rect 24724 -3722 24782 -3710
rect 24842 -3534 24900 -3522
rect 24842 -3710 24854 -3534
rect 24888 -3710 24900 -3534
rect 24842 -3722 24900 -3710
rect 16707 -6167 16765 -6155
rect 459 -6283 517 -6271
rect -25 -6483 33 -6471
rect -25 -6659 -13 -6483
rect 21 -6659 33 -6483
rect -25 -6671 33 -6659
rect 93 -6483 151 -6471
rect 93 -6659 105 -6483
rect 139 -6659 151 -6483
rect 93 -6671 151 -6659
rect 211 -6483 269 -6471
rect 211 -6659 223 -6483
rect 257 -6659 269 -6483
rect 211 -6671 269 -6659
rect 329 -6483 387 -6471
rect 329 -6659 341 -6483
rect 375 -6659 387 -6483
rect 329 -6671 387 -6659
rect 459 -6659 471 -6283
rect 505 -6659 517 -6283
rect 459 -6671 517 -6659
rect 577 -6283 635 -6271
rect 577 -6659 589 -6283
rect 623 -6659 635 -6283
rect 577 -6671 635 -6659
rect 695 -6283 753 -6271
rect 695 -6659 707 -6283
rect 741 -6659 753 -6283
rect 695 -6671 753 -6659
rect 813 -6283 871 -6271
rect 813 -6659 825 -6283
rect 859 -6659 871 -6283
rect 813 -6671 871 -6659
rect 931 -6283 989 -6271
rect 931 -6659 943 -6283
rect 977 -6659 989 -6283
rect 931 -6671 989 -6659
rect 1049 -6283 1107 -6271
rect 1049 -6659 1061 -6283
rect 1095 -6659 1107 -6283
rect 1049 -6671 1107 -6659
rect 1167 -6283 1225 -6271
rect 1167 -6659 1179 -6283
rect 1213 -6659 1225 -6283
rect 2527 -6281 2585 -6269
rect 1167 -6671 1225 -6659
rect 1296 -6483 1354 -6471
rect 1296 -6659 1308 -6483
rect 1342 -6659 1354 -6483
rect 1296 -6671 1354 -6659
rect 1414 -6483 1472 -6471
rect 1414 -6659 1426 -6483
rect 1460 -6659 1472 -6483
rect 1414 -6671 1472 -6659
rect 1532 -6483 1590 -6471
rect 1532 -6659 1544 -6483
rect 1578 -6659 1590 -6483
rect 1532 -6671 1590 -6659
rect 1650 -6483 1708 -6471
rect 1650 -6659 1662 -6483
rect 1696 -6659 1708 -6483
rect 1650 -6671 1708 -6659
rect 2043 -6481 2101 -6469
rect 2043 -6657 2055 -6481
rect 2089 -6657 2101 -6481
rect 2043 -6669 2101 -6657
rect 2161 -6481 2219 -6469
rect 2161 -6657 2173 -6481
rect 2207 -6657 2219 -6481
rect 2161 -6669 2219 -6657
rect 2279 -6481 2337 -6469
rect 2279 -6657 2291 -6481
rect 2325 -6657 2337 -6481
rect 2279 -6669 2337 -6657
rect 2397 -6481 2455 -6469
rect 2397 -6657 2409 -6481
rect 2443 -6657 2455 -6481
rect 2397 -6669 2455 -6657
rect 2527 -6657 2539 -6281
rect 2573 -6657 2585 -6281
rect 2527 -6669 2585 -6657
rect 2645 -6281 2703 -6269
rect 2645 -6657 2657 -6281
rect 2691 -6657 2703 -6281
rect 2645 -6669 2703 -6657
rect 2763 -6281 2821 -6269
rect 2763 -6657 2775 -6281
rect 2809 -6657 2821 -6281
rect 2763 -6669 2821 -6657
rect 2881 -6281 2939 -6269
rect 2881 -6657 2893 -6281
rect 2927 -6657 2939 -6281
rect 2881 -6669 2939 -6657
rect 2999 -6281 3057 -6269
rect 2999 -6657 3011 -6281
rect 3045 -6657 3057 -6281
rect 2999 -6669 3057 -6657
rect 3117 -6281 3175 -6269
rect 3117 -6657 3129 -6281
rect 3163 -6657 3175 -6281
rect 3117 -6669 3175 -6657
rect 3235 -6281 3293 -6269
rect 3235 -6657 3247 -6281
rect 3281 -6657 3293 -6281
rect 4596 -6283 4654 -6271
rect 3235 -6669 3293 -6657
rect 3364 -6481 3422 -6469
rect 3364 -6657 3376 -6481
rect 3410 -6657 3422 -6481
rect 3364 -6669 3422 -6657
rect 3482 -6481 3540 -6469
rect 3482 -6657 3494 -6481
rect 3528 -6657 3540 -6481
rect 3482 -6669 3540 -6657
rect 3600 -6481 3658 -6469
rect 3600 -6657 3612 -6481
rect 3646 -6657 3658 -6481
rect 3600 -6669 3658 -6657
rect 3718 -6481 3776 -6469
rect 3718 -6657 3730 -6481
rect 3764 -6657 3776 -6481
rect 3718 -6669 3776 -6657
rect 4112 -6483 4170 -6471
rect 4112 -6659 4124 -6483
rect 4158 -6659 4170 -6483
rect 402 -6976 460 -6964
rect 402 -7352 414 -6976
rect 448 -7352 460 -6976
rect 402 -7364 460 -7352
rect 520 -6976 578 -6964
rect 520 -7352 532 -6976
rect 566 -7352 578 -6976
rect 520 -7364 578 -7352
rect 638 -6976 696 -6964
rect 638 -7352 650 -6976
rect 684 -7352 696 -6976
rect 638 -7364 696 -7352
rect 756 -6976 814 -6964
rect 756 -7352 768 -6976
rect 802 -7352 814 -6976
rect 756 -7364 814 -7352
rect 874 -6976 932 -6964
rect 874 -7352 886 -6976
rect 920 -7352 932 -6976
rect 874 -7364 932 -7352
rect 992 -6976 1050 -6964
rect 992 -7352 1004 -6976
rect 1038 -7352 1050 -6976
rect 992 -7364 1050 -7352
rect 1110 -6976 1168 -6964
rect 1110 -7352 1122 -6976
rect 1156 -7352 1168 -6976
rect 1110 -7364 1168 -7352
rect 4112 -6671 4170 -6659
rect 4230 -6483 4288 -6471
rect 4230 -6659 4242 -6483
rect 4276 -6659 4288 -6483
rect 4230 -6671 4288 -6659
rect 4348 -6483 4406 -6471
rect 4348 -6659 4360 -6483
rect 4394 -6659 4406 -6483
rect 4348 -6671 4406 -6659
rect 4466 -6483 4524 -6471
rect 4466 -6659 4478 -6483
rect 4512 -6659 4524 -6483
rect 4466 -6671 4524 -6659
rect 4596 -6659 4608 -6283
rect 4642 -6659 4654 -6283
rect 4596 -6671 4654 -6659
rect 4714 -6283 4772 -6271
rect 4714 -6659 4726 -6283
rect 4760 -6659 4772 -6283
rect 4714 -6671 4772 -6659
rect 4832 -6283 4890 -6271
rect 4832 -6659 4844 -6283
rect 4878 -6659 4890 -6283
rect 4832 -6671 4890 -6659
rect 4950 -6283 5008 -6271
rect 4950 -6659 4962 -6283
rect 4996 -6659 5008 -6283
rect 4950 -6671 5008 -6659
rect 5068 -6283 5126 -6271
rect 5068 -6659 5080 -6283
rect 5114 -6659 5126 -6283
rect 5068 -6671 5126 -6659
rect 5186 -6283 5244 -6271
rect 5186 -6659 5198 -6283
rect 5232 -6659 5244 -6283
rect 5186 -6671 5244 -6659
rect 5304 -6283 5362 -6271
rect 5304 -6659 5316 -6283
rect 5350 -6659 5362 -6283
rect 6664 -6281 6722 -6269
rect 5304 -6671 5362 -6659
rect 5433 -6483 5491 -6471
rect 5433 -6659 5445 -6483
rect 5479 -6659 5491 -6483
rect 5433 -6671 5491 -6659
rect 5551 -6483 5609 -6471
rect 5551 -6659 5563 -6483
rect 5597 -6659 5609 -6483
rect 5551 -6671 5609 -6659
rect 5669 -6483 5727 -6471
rect 5669 -6659 5681 -6483
rect 5715 -6659 5727 -6483
rect 5669 -6671 5727 -6659
rect 5787 -6483 5845 -6471
rect 5787 -6659 5799 -6483
rect 5833 -6659 5845 -6483
rect 5787 -6671 5845 -6659
rect 6180 -6481 6238 -6469
rect 6180 -6657 6192 -6481
rect 6226 -6657 6238 -6481
rect 6180 -6669 6238 -6657
rect 6298 -6481 6356 -6469
rect 6298 -6657 6310 -6481
rect 6344 -6657 6356 -6481
rect 6298 -6669 6356 -6657
rect 6416 -6481 6474 -6469
rect 6416 -6657 6428 -6481
rect 6462 -6657 6474 -6481
rect 6416 -6669 6474 -6657
rect 6534 -6481 6592 -6469
rect 6534 -6657 6546 -6481
rect 6580 -6657 6592 -6481
rect 6534 -6669 6592 -6657
rect 6664 -6657 6676 -6281
rect 6710 -6657 6722 -6281
rect 6664 -6669 6722 -6657
rect 6782 -6281 6840 -6269
rect 6782 -6657 6794 -6281
rect 6828 -6657 6840 -6281
rect 6782 -6669 6840 -6657
rect 6900 -6281 6958 -6269
rect 6900 -6657 6912 -6281
rect 6946 -6657 6958 -6281
rect 6900 -6669 6958 -6657
rect 7018 -6281 7076 -6269
rect 7018 -6657 7030 -6281
rect 7064 -6657 7076 -6281
rect 7018 -6669 7076 -6657
rect 7136 -6281 7194 -6269
rect 7136 -6657 7148 -6281
rect 7182 -6657 7194 -6281
rect 7136 -6669 7194 -6657
rect 7254 -6281 7312 -6269
rect 7254 -6657 7266 -6281
rect 7300 -6657 7312 -6281
rect 7254 -6669 7312 -6657
rect 7372 -6281 7430 -6269
rect 7372 -6657 7384 -6281
rect 7418 -6657 7430 -6281
rect 8733 -6281 8791 -6269
rect 7372 -6669 7430 -6657
rect 7501 -6481 7559 -6469
rect 7501 -6657 7513 -6481
rect 7547 -6657 7559 -6481
rect 7501 -6669 7559 -6657
rect 7619 -6481 7677 -6469
rect 7619 -6657 7631 -6481
rect 7665 -6657 7677 -6481
rect 7619 -6669 7677 -6657
rect 7737 -6481 7795 -6469
rect 7737 -6657 7749 -6481
rect 7783 -6657 7795 -6481
rect 7737 -6669 7795 -6657
rect 7855 -6481 7913 -6469
rect 7855 -6657 7867 -6481
rect 7901 -6657 7913 -6481
rect 7855 -6669 7913 -6657
rect 8249 -6481 8307 -6469
rect 8249 -6657 8261 -6481
rect 8295 -6657 8307 -6481
rect 8249 -6669 8307 -6657
rect 8367 -6481 8425 -6469
rect 8367 -6657 8379 -6481
rect 8413 -6657 8425 -6481
rect 8367 -6669 8425 -6657
rect 8485 -6481 8543 -6469
rect 8485 -6657 8497 -6481
rect 8531 -6657 8543 -6481
rect 8485 -6669 8543 -6657
rect 8603 -6481 8661 -6469
rect 8603 -6657 8615 -6481
rect 8649 -6657 8661 -6481
rect 8603 -6669 8661 -6657
rect 8733 -6657 8745 -6281
rect 8779 -6657 8791 -6281
rect 8733 -6669 8791 -6657
rect 8851 -6281 8909 -6269
rect 8851 -6657 8863 -6281
rect 8897 -6657 8909 -6281
rect 8851 -6669 8909 -6657
rect 8969 -6281 9027 -6269
rect 8969 -6657 8981 -6281
rect 9015 -6657 9027 -6281
rect 8969 -6669 9027 -6657
rect 9087 -6281 9145 -6269
rect 9087 -6657 9099 -6281
rect 9133 -6657 9145 -6281
rect 9087 -6669 9145 -6657
rect 9205 -6281 9263 -6269
rect 9205 -6657 9217 -6281
rect 9251 -6657 9263 -6281
rect 9205 -6669 9263 -6657
rect 9323 -6281 9381 -6269
rect 9323 -6657 9335 -6281
rect 9369 -6657 9381 -6281
rect 9323 -6669 9381 -6657
rect 9441 -6281 9499 -6269
rect 9441 -6657 9453 -6281
rect 9487 -6657 9499 -6281
rect 10801 -6279 10859 -6267
rect 9441 -6669 9499 -6657
rect 9570 -6481 9628 -6469
rect 9570 -6657 9582 -6481
rect 9616 -6657 9628 -6481
rect 9570 -6669 9628 -6657
rect 9688 -6481 9746 -6469
rect 9688 -6657 9700 -6481
rect 9734 -6657 9746 -6481
rect 9688 -6669 9746 -6657
rect 9806 -6481 9864 -6469
rect 9806 -6657 9818 -6481
rect 9852 -6657 9864 -6481
rect 9806 -6669 9864 -6657
rect 9924 -6481 9982 -6469
rect 9924 -6657 9936 -6481
rect 9970 -6657 9982 -6481
rect 9924 -6669 9982 -6657
rect 10317 -6479 10375 -6467
rect 10317 -6655 10329 -6479
rect 10363 -6655 10375 -6479
rect 10317 -6667 10375 -6655
rect 10435 -6479 10493 -6467
rect 10435 -6655 10447 -6479
rect 10481 -6655 10493 -6479
rect 10435 -6667 10493 -6655
rect 10553 -6479 10611 -6467
rect 10553 -6655 10565 -6479
rect 10599 -6655 10611 -6479
rect 10553 -6667 10611 -6655
rect 10671 -6479 10729 -6467
rect 10671 -6655 10683 -6479
rect 10717 -6655 10729 -6479
rect 10671 -6667 10729 -6655
rect 10801 -6655 10813 -6279
rect 10847 -6655 10859 -6279
rect 10801 -6667 10859 -6655
rect 10919 -6279 10977 -6267
rect 10919 -6655 10931 -6279
rect 10965 -6655 10977 -6279
rect 10919 -6667 10977 -6655
rect 11037 -6279 11095 -6267
rect 11037 -6655 11049 -6279
rect 11083 -6655 11095 -6279
rect 11037 -6667 11095 -6655
rect 11155 -6279 11213 -6267
rect 11155 -6655 11167 -6279
rect 11201 -6655 11213 -6279
rect 11155 -6667 11213 -6655
rect 11273 -6279 11331 -6267
rect 11273 -6655 11285 -6279
rect 11319 -6655 11331 -6279
rect 11273 -6667 11331 -6655
rect 11391 -6279 11449 -6267
rect 11391 -6655 11403 -6279
rect 11437 -6655 11449 -6279
rect 11391 -6667 11449 -6655
rect 11509 -6279 11567 -6267
rect 11509 -6655 11521 -6279
rect 11555 -6655 11567 -6279
rect 12870 -6281 12928 -6269
rect 11509 -6667 11567 -6655
rect 11638 -6479 11696 -6467
rect 11638 -6655 11650 -6479
rect 11684 -6655 11696 -6479
rect 11638 -6667 11696 -6655
rect 11756 -6479 11814 -6467
rect 11756 -6655 11768 -6479
rect 11802 -6655 11814 -6479
rect 11756 -6667 11814 -6655
rect 11874 -6479 11932 -6467
rect 11874 -6655 11886 -6479
rect 11920 -6655 11932 -6479
rect 11874 -6667 11932 -6655
rect 11992 -6479 12050 -6467
rect 11992 -6655 12004 -6479
rect 12038 -6655 12050 -6479
rect 11992 -6667 12050 -6655
rect 12386 -6481 12444 -6469
rect 12386 -6657 12398 -6481
rect 12432 -6657 12444 -6481
rect 2470 -6974 2528 -6962
rect 2470 -7350 2482 -6974
rect 2516 -7350 2528 -6974
rect 2470 -7362 2528 -7350
rect 2588 -6974 2646 -6962
rect 2588 -7350 2600 -6974
rect 2634 -7350 2646 -6974
rect 2588 -7362 2646 -7350
rect 2706 -6974 2764 -6962
rect 2706 -7350 2718 -6974
rect 2752 -7350 2764 -6974
rect 2706 -7362 2764 -7350
rect 2824 -6974 2882 -6962
rect 2824 -7350 2836 -6974
rect 2870 -7350 2882 -6974
rect 2824 -7362 2882 -7350
rect 2942 -6974 3000 -6962
rect 2942 -7350 2954 -6974
rect 2988 -7350 3000 -6974
rect 2942 -7362 3000 -7350
rect 3060 -6974 3118 -6962
rect 3060 -7350 3072 -6974
rect 3106 -7350 3118 -6974
rect 3060 -7362 3118 -7350
rect 3178 -6974 3236 -6962
rect 3178 -7350 3190 -6974
rect 3224 -7350 3236 -6974
rect 3178 -7362 3236 -7350
rect 4539 -6976 4597 -6964
rect 4539 -7352 4551 -6976
rect 4585 -7352 4597 -6976
rect 4539 -7364 4597 -7352
rect 4657 -6976 4715 -6964
rect 4657 -7352 4669 -6976
rect 4703 -7352 4715 -6976
rect 4657 -7364 4715 -7352
rect 4775 -6976 4833 -6964
rect 4775 -7352 4787 -6976
rect 4821 -7352 4833 -6976
rect 4775 -7364 4833 -7352
rect 4893 -6976 4951 -6964
rect 4893 -7352 4905 -6976
rect 4939 -7352 4951 -6976
rect 4893 -7364 4951 -7352
rect 5011 -6976 5069 -6964
rect 5011 -7352 5023 -6976
rect 5057 -7352 5069 -6976
rect 5011 -7364 5069 -7352
rect 5129 -6976 5187 -6964
rect 5129 -7352 5141 -6976
rect 5175 -7352 5187 -6976
rect 5129 -7364 5187 -7352
rect 5247 -6976 5305 -6964
rect 5247 -7352 5259 -6976
rect 5293 -7352 5305 -6976
rect 5247 -7364 5305 -7352
rect 6607 -6974 6665 -6962
rect 6607 -7350 6619 -6974
rect 6653 -7350 6665 -6974
rect 6607 -7362 6665 -7350
rect 6725 -6974 6783 -6962
rect 6725 -7350 6737 -6974
rect 6771 -7350 6783 -6974
rect 6725 -7362 6783 -7350
rect 6843 -6974 6901 -6962
rect 6843 -7350 6855 -6974
rect 6889 -7350 6901 -6974
rect 6843 -7362 6901 -7350
rect 6961 -6974 7019 -6962
rect 6961 -7350 6973 -6974
rect 7007 -7350 7019 -6974
rect 6961 -7362 7019 -7350
rect 7079 -6974 7137 -6962
rect 7079 -7350 7091 -6974
rect 7125 -7350 7137 -6974
rect 7079 -7362 7137 -7350
rect 7197 -6974 7255 -6962
rect 7197 -7350 7209 -6974
rect 7243 -7350 7255 -6974
rect 7197 -7362 7255 -7350
rect 7315 -6974 7373 -6962
rect 7315 -7350 7327 -6974
rect 7361 -7350 7373 -6974
rect 7315 -7362 7373 -7350
rect 8676 -6974 8734 -6962
rect 8676 -7350 8688 -6974
rect 8722 -7350 8734 -6974
rect 8676 -7362 8734 -7350
rect 8794 -6974 8852 -6962
rect 8794 -7350 8806 -6974
rect 8840 -7350 8852 -6974
rect 8794 -7362 8852 -7350
rect 8912 -6974 8970 -6962
rect 8912 -7350 8924 -6974
rect 8958 -7350 8970 -6974
rect 8912 -7362 8970 -7350
rect 9030 -6974 9088 -6962
rect 9030 -7350 9042 -6974
rect 9076 -7350 9088 -6974
rect 9030 -7362 9088 -7350
rect 9148 -6974 9206 -6962
rect 9148 -7350 9160 -6974
rect 9194 -7350 9206 -6974
rect 9148 -7362 9206 -7350
rect 9266 -6974 9324 -6962
rect 9266 -7350 9278 -6974
rect 9312 -7350 9324 -6974
rect 9266 -7362 9324 -7350
rect 9384 -6974 9442 -6962
rect 9384 -7350 9396 -6974
rect 9430 -7350 9442 -6974
rect 9384 -7362 9442 -7350
rect 12386 -6669 12444 -6657
rect 12504 -6481 12562 -6469
rect 12504 -6657 12516 -6481
rect 12550 -6657 12562 -6481
rect 12504 -6669 12562 -6657
rect 12622 -6481 12680 -6469
rect 12622 -6657 12634 -6481
rect 12668 -6657 12680 -6481
rect 12622 -6669 12680 -6657
rect 12740 -6481 12798 -6469
rect 12740 -6657 12752 -6481
rect 12786 -6657 12798 -6481
rect 12740 -6669 12798 -6657
rect 12870 -6657 12882 -6281
rect 12916 -6657 12928 -6281
rect 12870 -6669 12928 -6657
rect 12988 -6281 13046 -6269
rect 12988 -6657 13000 -6281
rect 13034 -6657 13046 -6281
rect 12988 -6669 13046 -6657
rect 13106 -6281 13164 -6269
rect 13106 -6657 13118 -6281
rect 13152 -6657 13164 -6281
rect 13106 -6669 13164 -6657
rect 13224 -6281 13282 -6269
rect 13224 -6657 13236 -6281
rect 13270 -6657 13282 -6281
rect 13224 -6669 13282 -6657
rect 13342 -6281 13400 -6269
rect 13342 -6657 13354 -6281
rect 13388 -6657 13400 -6281
rect 13342 -6669 13400 -6657
rect 13460 -6281 13518 -6269
rect 13460 -6657 13472 -6281
rect 13506 -6657 13518 -6281
rect 13460 -6669 13518 -6657
rect 13578 -6281 13636 -6269
rect 13578 -6657 13590 -6281
rect 13624 -6657 13636 -6281
rect 14938 -6279 14996 -6267
rect 13578 -6669 13636 -6657
rect 13707 -6481 13765 -6469
rect 13707 -6657 13719 -6481
rect 13753 -6657 13765 -6481
rect 13707 -6669 13765 -6657
rect 13825 -6481 13883 -6469
rect 13825 -6657 13837 -6481
rect 13871 -6657 13883 -6481
rect 13825 -6669 13883 -6657
rect 13943 -6481 14001 -6469
rect 13943 -6657 13955 -6481
rect 13989 -6657 14001 -6481
rect 13943 -6669 14001 -6657
rect 14061 -6481 14119 -6469
rect 14061 -6657 14073 -6481
rect 14107 -6657 14119 -6481
rect 14061 -6669 14119 -6657
rect 14454 -6479 14512 -6467
rect 14454 -6655 14466 -6479
rect 14500 -6655 14512 -6479
rect 14454 -6667 14512 -6655
rect 14572 -6479 14630 -6467
rect 14572 -6655 14584 -6479
rect 14618 -6655 14630 -6479
rect 14572 -6667 14630 -6655
rect 14690 -6479 14748 -6467
rect 14690 -6655 14702 -6479
rect 14736 -6655 14748 -6479
rect 14690 -6667 14748 -6655
rect 14808 -6479 14866 -6467
rect 14808 -6655 14820 -6479
rect 14854 -6655 14866 -6479
rect 14808 -6667 14866 -6655
rect 14938 -6655 14950 -6279
rect 14984 -6655 14996 -6279
rect 14938 -6667 14996 -6655
rect 15056 -6279 15114 -6267
rect 15056 -6655 15068 -6279
rect 15102 -6655 15114 -6279
rect 15056 -6667 15114 -6655
rect 15174 -6279 15232 -6267
rect 15174 -6655 15186 -6279
rect 15220 -6655 15232 -6279
rect 15174 -6667 15232 -6655
rect 15292 -6279 15350 -6267
rect 15292 -6655 15304 -6279
rect 15338 -6655 15350 -6279
rect 15292 -6667 15350 -6655
rect 15410 -6279 15468 -6267
rect 15410 -6655 15422 -6279
rect 15456 -6655 15468 -6279
rect 15410 -6667 15468 -6655
rect 15528 -6279 15586 -6267
rect 15528 -6655 15540 -6279
rect 15574 -6655 15586 -6279
rect 15528 -6667 15586 -6655
rect 15646 -6279 15704 -6267
rect 15646 -6655 15658 -6279
rect 15692 -6655 15704 -6279
rect 16707 -6343 16719 -6167
rect 16753 -6343 16765 -6167
rect 16707 -6355 16765 -6343
rect 16825 -6167 16883 -6155
rect 16825 -6343 16837 -6167
rect 16871 -6343 16883 -6167
rect 16825 -6355 16883 -6343
rect 16943 -6167 17001 -6155
rect 16943 -6343 16955 -6167
rect 16989 -6343 17001 -6167
rect 16943 -6355 17001 -6343
rect 17061 -6167 17119 -6155
rect 17061 -6343 17073 -6167
rect 17107 -6343 17119 -6167
rect 17061 -6355 17119 -6343
rect 17445 -6163 17503 -6151
rect 17445 -6339 17457 -6163
rect 17491 -6339 17503 -6163
rect 17445 -6351 17503 -6339
rect 17563 -6163 17621 -6151
rect 17563 -6339 17575 -6163
rect 17609 -6339 17621 -6163
rect 17563 -6351 17621 -6339
rect 17681 -6163 17739 -6151
rect 17681 -6339 17693 -6163
rect 17727 -6339 17739 -6163
rect 17681 -6351 17739 -6339
rect 17799 -6163 17857 -6151
rect 17799 -6339 17811 -6163
rect 17845 -6339 17857 -6163
rect 17799 -6351 17857 -6339
rect 18183 -6167 18241 -6155
rect 18183 -6343 18195 -6167
rect 18229 -6343 18241 -6167
rect 18183 -6355 18241 -6343
rect 18301 -6167 18359 -6155
rect 18301 -6343 18313 -6167
rect 18347 -6343 18359 -6167
rect 18301 -6355 18359 -6343
rect 18419 -6167 18477 -6155
rect 18419 -6343 18431 -6167
rect 18465 -6343 18477 -6167
rect 18419 -6355 18477 -6343
rect 18537 -6167 18595 -6155
rect 18537 -6343 18549 -6167
rect 18583 -6343 18595 -6167
rect 18537 -6355 18595 -6343
rect 18925 -6169 18983 -6157
rect 18925 -6345 18937 -6169
rect 18971 -6345 18983 -6169
rect 18925 -6357 18983 -6345
rect 19043 -6169 19101 -6157
rect 19043 -6345 19055 -6169
rect 19089 -6345 19101 -6169
rect 19043 -6357 19101 -6345
rect 19161 -6169 19219 -6157
rect 19161 -6345 19173 -6169
rect 19207 -6345 19219 -6169
rect 19161 -6357 19219 -6345
rect 19279 -6169 19337 -6157
rect 19279 -6345 19291 -6169
rect 19325 -6345 19337 -6169
rect 19279 -6357 19337 -6345
rect 19665 -6169 19723 -6157
rect 19665 -6345 19677 -6169
rect 19711 -6345 19723 -6169
rect 19665 -6357 19723 -6345
rect 19783 -6169 19841 -6157
rect 19783 -6345 19795 -6169
rect 19829 -6345 19841 -6169
rect 19783 -6357 19841 -6345
rect 19901 -6169 19959 -6157
rect 19901 -6345 19913 -6169
rect 19947 -6345 19959 -6169
rect 19901 -6357 19959 -6345
rect 20019 -6169 20077 -6157
rect 20019 -6345 20031 -6169
rect 20065 -6345 20077 -6169
rect 20019 -6357 20077 -6345
rect 20403 -6169 20461 -6157
rect 20403 -6345 20415 -6169
rect 20449 -6345 20461 -6169
rect 20403 -6357 20461 -6345
rect 20521 -6169 20579 -6157
rect 20521 -6345 20533 -6169
rect 20567 -6345 20579 -6169
rect 20521 -6357 20579 -6345
rect 20639 -6169 20697 -6157
rect 20639 -6345 20651 -6169
rect 20685 -6345 20697 -6169
rect 20639 -6357 20697 -6345
rect 20757 -6169 20815 -6157
rect 20757 -6345 20769 -6169
rect 20803 -6345 20815 -6169
rect 20757 -6357 20815 -6345
rect 21141 -6169 21199 -6157
rect 21141 -6345 21153 -6169
rect 21187 -6345 21199 -6169
rect 21141 -6357 21199 -6345
rect 21259 -6169 21317 -6157
rect 21259 -6345 21271 -6169
rect 21305 -6345 21317 -6169
rect 21259 -6357 21317 -6345
rect 21377 -6169 21435 -6157
rect 21377 -6345 21389 -6169
rect 21423 -6345 21435 -6169
rect 21377 -6357 21435 -6345
rect 21495 -6169 21553 -6157
rect 21495 -6345 21507 -6169
rect 21541 -6345 21553 -6169
rect 21495 -6357 21553 -6345
rect 21879 -6169 21937 -6157
rect 21879 -6345 21891 -6169
rect 21925 -6345 21937 -6169
rect 21879 -6357 21937 -6345
rect 21997 -6169 22055 -6157
rect 21997 -6345 22009 -6169
rect 22043 -6345 22055 -6169
rect 21997 -6357 22055 -6345
rect 22115 -6169 22173 -6157
rect 22115 -6345 22127 -6169
rect 22161 -6345 22173 -6169
rect 22115 -6357 22173 -6345
rect 22233 -6169 22291 -6157
rect 22233 -6345 22245 -6169
rect 22279 -6345 22291 -6169
rect 22233 -6357 22291 -6345
rect 15646 -6667 15704 -6655
rect 15775 -6479 15833 -6467
rect 15775 -6655 15787 -6479
rect 15821 -6655 15833 -6479
rect 15775 -6667 15833 -6655
rect 15893 -6479 15951 -6467
rect 15893 -6655 15905 -6479
rect 15939 -6655 15951 -6479
rect 15893 -6667 15951 -6655
rect 16011 -6479 16069 -6467
rect 16011 -6655 16023 -6479
rect 16057 -6655 16069 -6479
rect 16011 -6667 16069 -6655
rect 16129 -6479 16187 -6467
rect 16129 -6655 16141 -6479
rect 16175 -6655 16187 -6479
rect 16129 -6667 16187 -6655
rect 10744 -6972 10802 -6960
rect 10744 -7348 10756 -6972
rect 10790 -7348 10802 -6972
rect 10744 -7360 10802 -7348
rect 10862 -6972 10920 -6960
rect 10862 -7348 10874 -6972
rect 10908 -7348 10920 -6972
rect 10862 -7360 10920 -7348
rect 10980 -6972 11038 -6960
rect 10980 -7348 10992 -6972
rect 11026 -7348 11038 -6972
rect 10980 -7360 11038 -7348
rect 11098 -6972 11156 -6960
rect 11098 -7348 11110 -6972
rect 11144 -7348 11156 -6972
rect 11098 -7360 11156 -7348
rect 11216 -6972 11274 -6960
rect 11216 -7348 11228 -6972
rect 11262 -7348 11274 -6972
rect 11216 -7360 11274 -7348
rect 11334 -6972 11392 -6960
rect 11334 -7348 11346 -6972
rect 11380 -7348 11392 -6972
rect 11334 -7360 11392 -7348
rect 11452 -6972 11510 -6960
rect 11452 -7348 11464 -6972
rect 11498 -7348 11510 -6972
rect 11452 -7360 11510 -7348
rect 12813 -6974 12871 -6962
rect 12813 -7350 12825 -6974
rect 12859 -7350 12871 -6974
rect 12813 -7362 12871 -7350
rect 12931 -6974 12989 -6962
rect 12931 -7350 12943 -6974
rect 12977 -7350 12989 -6974
rect 12931 -7362 12989 -7350
rect 13049 -6974 13107 -6962
rect 13049 -7350 13061 -6974
rect 13095 -7350 13107 -6974
rect 13049 -7362 13107 -7350
rect 13167 -6974 13225 -6962
rect 13167 -7350 13179 -6974
rect 13213 -7350 13225 -6974
rect 13167 -7362 13225 -7350
rect 13285 -6974 13343 -6962
rect 13285 -7350 13297 -6974
rect 13331 -7350 13343 -6974
rect 13285 -7362 13343 -7350
rect 13403 -6974 13461 -6962
rect 13403 -7350 13415 -6974
rect 13449 -7350 13461 -6974
rect 13403 -7362 13461 -7350
rect 13521 -6974 13579 -6962
rect 13521 -7350 13533 -6974
rect 13567 -7350 13579 -6974
rect 13521 -7362 13579 -7350
rect 14881 -6972 14939 -6960
rect 14881 -7348 14893 -6972
rect 14927 -7348 14939 -6972
rect 14881 -7360 14939 -7348
rect 14999 -6972 15057 -6960
rect 14999 -7348 15011 -6972
rect 15045 -7348 15057 -6972
rect 14999 -7360 15057 -7348
rect 15117 -6972 15175 -6960
rect 15117 -7348 15129 -6972
rect 15163 -7348 15175 -6972
rect 15117 -7360 15175 -7348
rect 15235 -6972 15293 -6960
rect 15235 -7348 15247 -6972
rect 15281 -7348 15293 -6972
rect 15235 -7360 15293 -7348
rect 15353 -6972 15411 -6960
rect 15353 -7348 15365 -6972
rect 15399 -7348 15411 -6972
rect 15353 -7360 15411 -7348
rect 15471 -6972 15529 -6960
rect 15471 -7348 15483 -6972
rect 15517 -7348 15529 -6972
rect 15471 -7360 15529 -7348
rect 15589 -6972 15647 -6960
rect 15589 -7348 15601 -6972
rect 15635 -7348 15647 -6972
rect 15589 -7360 15647 -7348
<< ndiffc >>
rect 438 3072 472 3448
rect 556 3072 590 3448
rect 674 3072 708 3448
rect 791 3272 825 3448
rect 909 3272 943 3448
rect 1886 3072 1920 3448
rect 2004 3072 2038 3448
rect 2122 3072 2156 3448
rect 2239 3272 2273 3448
rect 2357 3272 2391 3448
rect 3384 3074 3418 3450
rect 3502 3074 3536 3450
rect 3620 3074 3654 3450
rect 3737 3274 3771 3450
rect 3855 3274 3889 3450
rect 4832 3074 4866 3450
rect 4950 3074 4984 3450
rect 5068 3074 5102 3450
rect 5185 3274 5219 3450
rect 5303 3274 5337 3450
rect 6352 3072 6386 3448
rect 6470 3072 6504 3448
rect 6588 3072 6622 3448
rect 6705 3272 6739 3448
rect 6823 3272 6857 3448
rect 7800 3072 7834 3448
rect 7918 3072 7952 3448
rect 8036 3072 8070 3448
rect 8153 3272 8187 3448
rect 8271 3272 8305 3448
rect 9298 3074 9332 3450
rect 9416 3074 9450 3450
rect 9534 3074 9568 3450
rect 9651 3274 9685 3450
rect 9769 3274 9803 3450
rect 10746 3074 10780 3450
rect 10864 3074 10898 3450
rect 10982 3074 11016 3450
rect 11099 3274 11133 3450
rect 11217 3274 11251 3450
rect 11874 3120 11908 3296
rect 11992 3120 12026 3296
rect 12110 3120 12144 3296
rect 12228 3120 12262 3296
rect 13042 3122 13076 3298
rect 13160 3122 13194 3298
rect 13278 3122 13312 3298
rect 13396 3122 13430 3298
rect 14210 3122 14244 3298
rect 14328 3122 14362 3298
rect 14446 3122 14480 3298
rect 14564 3122 14598 3298
rect 15378 3122 15412 3298
rect 15496 3122 15530 3298
rect 15614 3122 15648 3298
rect 15732 3122 15766 3298
rect 16552 3122 16586 3298
rect 16670 3122 16704 3298
rect 16788 3122 16822 3298
rect 16906 3122 16940 3298
rect 17720 3122 17754 3298
rect 17838 3122 17872 3298
rect 17956 3122 17990 3298
rect 18074 3122 18108 3298
rect 18888 3124 18922 3300
rect 19006 3124 19040 3300
rect 19124 3124 19158 3300
rect 19242 3124 19276 3300
rect 20056 3124 20090 3300
rect 20174 3124 20208 3300
rect 20292 3124 20326 3300
rect 20410 3124 20444 3300
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 1094 -2115 1128 -1939
rect 1212 -2115 1246 -1939
rect 1286 -2315 1320 -1939
rect 1404 -2315 1438 -1939
rect 1522 -2315 1556 -1939
rect 1640 -2315 1674 -1939
rect 1758 -2315 1792 -1939
rect 1836 -2115 1870 -1939
rect 1954 -2115 1988 -1939
rect 4238 -2115 4272 -1939
rect 4356 -2115 4390 -1939
rect 4430 -2315 4464 -1939
rect 4548 -2315 4582 -1939
rect 4666 -2315 4700 -1939
rect 4784 -2315 4818 -1939
rect 4902 -2315 4936 -1939
rect 4980 -2115 5014 -1939
rect 5098 -2115 5132 -1939
rect 7370 -2111 7404 -1935
rect 7488 -2111 7522 -1935
rect 7562 -2311 7596 -1935
rect 7680 -2311 7714 -1935
rect 7798 -2311 7832 -1935
rect 7916 -2311 7950 -1935
rect 8034 -2311 8068 -1935
rect 8112 -2111 8146 -1935
rect 8230 -2111 8264 -1935
rect 10514 -2111 10548 -1935
rect 10632 -2111 10666 -1935
rect 10706 -2311 10740 -1935
rect 10824 -2311 10858 -1935
rect 10942 -2311 10976 -1935
rect 11060 -2311 11094 -1935
rect 11178 -2311 11212 -1935
rect 11256 -2111 11290 -1935
rect 11374 -2111 11408 -1935
rect 13716 -2115 13750 -1939
rect 13834 -2115 13868 -1939
rect 13908 -2315 13942 -1939
rect 14026 -2315 14060 -1939
rect 14144 -2315 14178 -1939
rect 14262 -2315 14296 -1939
rect 14380 -2315 14414 -1939
rect 14458 -2115 14492 -1939
rect 14576 -2115 14610 -1939
rect 16860 -2115 16894 -1939
rect 16978 -2115 17012 -1939
rect 17052 -2315 17086 -1939
rect 17170 -2315 17204 -1939
rect 17288 -2315 17322 -1939
rect 17406 -2315 17440 -1939
rect 17524 -2315 17558 -1939
rect 17602 -2115 17636 -1939
rect 17720 -2115 17754 -1939
rect 19992 -2111 20026 -1935
rect 20110 -2111 20144 -1935
rect 20184 -2311 20218 -1935
rect 20302 -2311 20336 -1935
rect 20420 -2311 20454 -1935
rect 20538 -2311 20572 -1935
rect 20656 -2311 20690 -1935
rect 20734 -2111 20768 -1935
rect 20852 -2111 20886 -1935
rect 23136 -2111 23170 -1935
rect 23254 -2111 23288 -1935
rect 23328 -2311 23362 -1935
rect 23446 -2311 23480 -1935
rect 23564 -2311 23598 -1935
rect 23682 -2311 23716 -1935
rect 23800 -2311 23834 -1935
rect 23878 -2111 23912 -1935
rect 23996 -2111 24030 -1935
rect 1084 -4847 1118 -4671
rect 1202 -4847 1236 -4671
rect 1276 -5047 1310 -4671
rect 1394 -5047 1428 -4671
rect 1512 -5047 1546 -4671
rect 1630 -5047 1664 -4671
rect 1748 -5047 1782 -4671
rect 1826 -4847 1860 -4671
rect 1944 -4847 1978 -4671
rect 4228 -4847 4262 -4671
rect 4346 -4847 4380 -4671
rect 4420 -5047 4454 -4671
rect 4538 -5047 4572 -4671
rect 4656 -5047 4690 -4671
rect 4774 -5047 4808 -4671
rect 4892 -5047 4926 -4671
rect 4970 -4847 5004 -4671
rect 5088 -4847 5122 -4671
rect 7360 -4843 7394 -4667
rect 7478 -4843 7512 -4667
rect 7552 -5043 7586 -4667
rect 7670 -5043 7704 -4667
rect 7788 -5043 7822 -4667
rect 7906 -5043 7940 -4667
rect 8024 -5043 8058 -4667
rect 8102 -4843 8136 -4667
rect 8220 -4843 8254 -4667
rect 10504 -4843 10538 -4667
rect 10622 -4843 10656 -4667
rect 10696 -5043 10730 -4667
rect 10814 -5043 10848 -4667
rect 10932 -5043 10966 -4667
rect 11050 -5043 11084 -4667
rect 11168 -5043 11202 -4667
rect 11246 -4843 11280 -4667
rect 11364 -4843 11398 -4667
rect 13706 -4847 13740 -4671
rect 13824 -4847 13858 -4671
rect 13898 -5047 13932 -4671
rect 14016 -5047 14050 -4671
rect 14134 -5047 14168 -4671
rect 14252 -5047 14286 -4671
rect 14370 -5047 14404 -4671
rect 14448 -4847 14482 -4671
rect 14566 -4847 14600 -4671
rect 16850 -4847 16884 -4671
rect 16968 -4847 17002 -4671
rect 17042 -5047 17076 -4671
rect 17160 -5047 17194 -4671
rect 17278 -5047 17312 -4671
rect 17396 -5047 17430 -4671
rect 17514 -5047 17548 -4671
rect 17592 -4847 17626 -4671
rect 17710 -4847 17744 -4671
rect 19982 -4843 20016 -4667
rect 20100 -4843 20134 -4667
rect 20174 -5043 20208 -4667
rect 20292 -5043 20326 -4667
rect 20410 -5043 20444 -4667
rect 20528 -5043 20562 -4667
rect 20646 -5043 20680 -4667
rect 20724 -4843 20758 -4667
rect 20842 -4843 20876 -4667
rect 23126 -4843 23160 -4667
rect 23244 -4843 23278 -4667
rect 23318 -5043 23352 -4667
rect 23436 -5043 23470 -4667
rect 23554 -5043 23588 -4667
rect 23672 -5043 23706 -4667
rect 23790 -5043 23824 -4667
rect 23868 -4843 23902 -4667
rect 23986 -4843 24020 -4667
rect 112 -7884 146 -7708
rect 230 -7884 264 -7708
rect 532 -8084 566 -7708
rect 650 -8084 684 -7708
rect 768 -8084 802 -7708
rect 886 -8084 920 -7708
rect 1004 -8084 1038 -7708
rect 1410 -7884 1444 -7708
rect 1528 -7884 1562 -7708
rect 2180 -7882 2214 -7706
rect 2298 -7882 2332 -7706
rect 2600 -8082 2634 -7706
rect 2718 -8082 2752 -7706
rect 2836 -8082 2870 -7706
rect 2954 -8082 2988 -7706
rect 3072 -8082 3106 -7706
rect 3478 -7882 3512 -7706
rect 3596 -7882 3630 -7706
rect 4249 -7884 4283 -7708
rect 4367 -7884 4401 -7708
rect 4669 -8084 4703 -7708
rect 4787 -8084 4821 -7708
rect 4905 -8084 4939 -7708
rect 5023 -8084 5057 -7708
rect 5141 -8084 5175 -7708
rect 5547 -7884 5581 -7708
rect 5665 -7884 5699 -7708
rect 6317 -7882 6351 -7706
rect 6435 -7882 6469 -7706
rect 6737 -8082 6771 -7706
rect 6855 -8082 6889 -7706
rect 6973 -8082 7007 -7706
rect 7091 -8082 7125 -7706
rect 7209 -8082 7243 -7706
rect 7615 -7882 7649 -7706
rect 7733 -7882 7767 -7706
rect 8386 -7882 8420 -7706
rect 8504 -7882 8538 -7706
rect 8806 -8082 8840 -7706
rect 8924 -8082 8958 -7706
rect 9042 -8082 9076 -7706
rect 9160 -8082 9194 -7706
rect 9278 -8082 9312 -7706
rect 9684 -7882 9718 -7706
rect 9802 -7882 9836 -7706
rect 10454 -7880 10488 -7704
rect 10572 -7880 10606 -7704
rect 10874 -8080 10908 -7704
rect 10992 -8080 11026 -7704
rect 11110 -8080 11144 -7704
rect 11228 -8080 11262 -7704
rect 11346 -8080 11380 -7704
rect 11752 -7880 11786 -7704
rect 16837 -6729 16871 -6553
rect 16955 -6729 16989 -6553
rect 17575 -6727 17609 -6551
rect 17693 -6727 17727 -6551
rect 18313 -6731 18347 -6555
rect 18431 -6731 18465 -6555
rect 19055 -6731 19089 -6555
rect 19173 -6731 19207 -6555
rect 19795 -6731 19829 -6555
rect 19913 -6731 19947 -6555
rect 20533 -6731 20567 -6555
rect 20651 -6731 20685 -6555
rect 21271 -6727 21305 -6551
rect 21389 -6727 21423 -6551
rect 22009 -6727 22043 -6551
rect 22127 -6727 22161 -6551
rect 11870 -7880 11904 -7704
rect 12523 -7882 12557 -7706
rect 12641 -7882 12675 -7706
rect 12943 -8082 12977 -7706
rect 13061 -8082 13095 -7706
rect 13179 -8082 13213 -7706
rect 13297 -8082 13331 -7706
rect 13415 -8082 13449 -7706
rect 13821 -7882 13855 -7706
rect 13939 -7882 13973 -7706
rect 14591 -7880 14625 -7704
rect 14709 -7880 14743 -7704
rect 15011 -8080 15045 -7704
rect 15129 -8080 15163 -7704
rect 15247 -8080 15281 -7704
rect 15365 -8080 15399 -7704
rect 15483 -8080 15517 -7704
rect 15889 -7880 15923 -7704
rect 16007 -7880 16041 -7704
<< pdiffc >>
rect 201 3709 235 3885
rect 319 3709 353 3885
rect 437 3709 471 3885
rect 555 3709 589 3885
rect 673 3709 707 3885
rect 791 3709 825 3885
rect 909 3709 943 3885
rect 1027 3709 1061 3885
rect 1145 3709 1179 3885
rect 1263 3709 1297 3885
rect 1649 3709 1683 3885
rect 1767 3709 1801 3885
rect 1885 3709 1919 3885
rect 2003 3709 2037 3885
rect 2121 3709 2155 3885
rect 2239 3709 2273 3885
rect 2357 3709 2391 3885
rect 2475 3709 2509 3885
rect 2593 3709 2627 3885
rect 2711 3709 2745 3885
rect 3147 3711 3181 3887
rect 3265 3711 3299 3887
rect 3383 3711 3417 3887
rect 3501 3711 3535 3887
rect 3619 3711 3653 3887
rect 3737 3711 3771 3887
rect 3855 3711 3889 3887
rect 3973 3711 4007 3887
rect 4091 3711 4125 3887
rect 4209 3711 4243 3887
rect 4595 3711 4629 3887
rect 4713 3711 4747 3887
rect 4831 3711 4865 3887
rect 4949 3711 4983 3887
rect 5067 3711 5101 3887
rect 5185 3711 5219 3887
rect 5303 3711 5337 3887
rect 5421 3711 5455 3887
rect 5539 3711 5573 3887
rect 5657 3711 5691 3887
rect 6115 3709 6149 3885
rect 6233 3709 6267 3885
rect 6351 3709 6385 3885
rect 6469 3709 6503 3885
rect 6587 3709 6621 3885
rect 6705 3709 6739 3885
rect 6823 3709 6857 3885
rect 6941 3709 6975 3885
rect 7059 3709 7093 3885
rect 7177 3709 7211 3885
rect 7563 3709 7597 3885
rect 7681 3709 7715 3885
rect 7799 3709 7833 3885
rect 7917 3709 7951 3885
rect 8035 3709 8069 3885
rect 8153 3709 8187 3885
rect 8271 3709 8305 3885
rect 8389 3709 8423 3885
rect 8507 3709 8541 3885
rect 8625 3709 8659 3885
rect 9061 3711 9095 3887
rect 9179 3711 9213 3887
rect 9297 3711 9331 3887
rect 9415 3711 9449 3887
rect 9533 3711 9567 3887
rect 9651 3711 9685 3887
rect 9769 3711 9803 3887
rect 9887 3711 9921 3887
rect 10005 3711 10039 3887
rect 10123 3711 10157 3887
rect 10509 3711 10543 3887
rect 10627 3711 10661 3887
rect 10745 3711 10779 3887
rect 10863 3711 10897 3887
rect 10981 3711 11015 3887
rect 11099 3711 11133 3887
rect 11217 3711 11251 3887
rect 11335 3711 11369 3887
rect 11453 3711 11487 3887
rect 11571 3711 11605 3887
rect 11964 3706 11998 4082
rect 12082 3706 12116 4082
rect 12200 3706 12234 4082
rect 12318 3706 12352 4082
rect 12436 3706 12470 4082
rect 12554 3706 12588 4082
rect 12672 3706 12706 4082
rect 13132 3706 13166 4082
rect 13250 3706 13284 4082
rect 13368 3706 13402 4082
rect 13486 3706 13520 4082
rect 13604 3706 13638 4082
rect 13722 3706 13756 4082
rect 13840 3706 13874 4082
rect 14300 3704 14334 4080
rect 14418 3704 14452 4080
rect 14536 3704 14570 4080
rect 14654 3704 14688 4080
rect 14772 3704 14806 4080
rect 14890 3704 14924 4080
rect 15008 3704 15042 4080
rect 15468 3706 15502 4082
rect 15586 3706 15620 4082
rect 15704 3706 15738 4082
rect 15822 3706 15856 4082
rect 15940 3706 15974 4082
rect 16058 3706 16092 4082
rect 16176 3706 16210 4082
rect 16642 3708 16676 4084
rect 16760 3708 16794 4084
rect 16878 3708 16912 4084
rect 16996 3708 17030 4084
rect 17114 3708 17148 4084
rect 17232 3708 17266 4084
rect 17350 3708 17384 4084
rect 17810 3706 17844 4082
rect 17928 3706 17962 4082
rect 18046 3706 18080 4082
rect 18164 3706 18198 4082
rect 18282 3706 18316 4082
rect 18400 3706 18434 4082
rect 18518 3706 18552 4082
rect 18978 3708 19012 4084
rect 19096 3708 19130 4084
rect 19214 3708 19248 4084
rect 19332 3708 19366 4084
rect 19450 3708 19484 4084
rect 19568 3708 19602 4084
rect 19686 3708 19720 4084
rect 20146 3706 20180 4082
rect 12394 3116 12428 3292
rect 12512 3116 12546 3292
rect 12630 3116 12664 3292
rect 12748 3116 12782 3292
rect 13561 3122 13595 3298
rect 13679 3122 13713 3298
rect 13797 3122 13831 3298
rect 13915 3122 13949 3298
rect 14729 3122 14763 3298
rect 14847 3122 14881 3298
rect 14965 3122 14999 3298
rect 15083 3122 15117 3298
rect 15898 3122 15932 3298
rect 16016 3122 16050 3298
rect 16134 3122 16168 3298
rect 16252 3122 16286 3298
rect 17070 3118 17104 3294
rect 17188 3118 17222 3294
rect 17306 3118 17340 3294
rect 17424 3118 17458 3294
rect 20264 3706 20298 4082
rect 20382 3706 20416 4082
rect 20500 3706 20534 4082
rect 20618 3706 20652 4082
rect 20736 3706 20770 4082
rect 20854 3706 20888 4082
rect 18239 3117 18273 3293
rect 18357 3117 18391 3293
rect 18475 3117 18509 3293
rect 18593 3117 18627 3293
rect 19407 3117 19441 3293
rect 19525 3117 19559 3293
rect 19643 3117 19677 3293
rect 19761 3117 19795 3293
rect 20575 3118 20609 3294
rect 20693 3118 20727 3294
rect 20811 3118 20845 3294
rect 20929 3118 20963 3294
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 260 -982 294 -806
rect 378 -982 412 -806
rect 496 -982 530 -806
rect 614 -982 648 -806
rect 701 -982 735 -606
rect 819 -982 853 -606
rect 937 -982 971 -606
rect 1055 -982 1089 -606
rect 1168 -982 1202 -606
rect 1286 -982 1320 -606
rect 1404 -982 1438 -606
rect 1522 -982 1556 -606
rect 1640 -982 1674 -606
rect 1758 -982 1792 -606
rect 1876 -982 1910 -606
rect 1995 -982 2029 -606
rect 2113 -982 2147 -606
rect 2231 -982 2265 -606
rect 2349 -982 2383 -606
rect 2468 -982 2502 -806
rect 2586 -982 2620 -806
rect 2704 -982 2738 -806
rect 2822 -982 2856 -806
rect 3404 -982 3438 -806
rect 3522 -982 3556 -806
rect 3640 -982 3674 -806
rect 3758 -982 3792 -806
rect 3845 -982 3879 -606
rect 3963 -982 3997 -606
rect 4081 -982 4115 -606
rect 4199 -982 4233 -606
rect 4312 -982 4346 -606
rect 4430 -982 4464 -606
rect 4548 -982 4582 -606
rect 4666 -982 4700 -606
rect 4784 -982 4818 -606
rect 4902 -982 4936 -606
rect 5020 -982 5054 -606
rect 5139 -982 5173 -606
rect 5257 -982 5291 -606
rect 5375 -982 5409 -606
rect 5493 -982 5527 -606
rect 5612 -982 5646 -806
rect 5730 -982 5764 -806
rect 5848 -982 5882 -806
rect 5966 -982 6000 -806
rect 6536 -978 6570 -802
rect 6654 -978 6688 -802
rect 6772 -978 6806 -802
rect 6890 -978 6924 -802
rect 6977 -978 7011 -602
rect 7095 -978 7129 -602
rect 7213 -978 7247 -602
rect 7331 -978 7365 -602
rect 7444 -978 7478 -602
rect 7562 -978 7596 -602
rect 7680 -978 7714 -602
rect 7798 -978 7832 -602
rect 7916 -978 7950 -602
rect 8034 -978 8068 -602
rect 8152 -978 8186 -602
rect 8271 -978 8305 -602
rect 8389 -978 8423 -602
rect 8507 -978 8541 -602
rect 8625 -978 8659 -602
rect 8744 -978 8778 -802
rect 8862 -978 8896 -802
rect 8980 -978 9014 -802
rect 9098 -978 9132 -802
rect 9680 -978 9714 -802
rect 9798 -978 9832 -802
rect 9916 -978 9950 -802
rect 10034 -978 10068 -802
rect 10121 -978 10155 -602
rect 10239 -978 10273 -602
rect 10357 -978 10391 -602
rect 10475 -978 10509 -602
rect 10588 -978 10622 -602
rect 10706 -978 10740 -602
rect 10824 -978 10858 -602
rect 10942 -978 10976 -602
rect 11060 -978 11094 -602
rect 11178 -978 11212 -602
rect 11296 -978 11330 -602
rect 11415 -978 11449 -602
rect 11533 -978 11567 -602
rect 11651 -978 11685 -602
rect 11769 -978 11803 -602
rect 11888 -978 11922 -802
rect 12006 -978 12040 -802
rect 12124 -978 12158 -802
rect 12242 -978 12276 -802
rect 12882 -982 12916 -806
rect 13000 -982 13034 -806
rect 13118 -982 13152 -806
rect 13236 -982 13270 -806
rect 13323 -982 13357 -606
rect 13441 -982 13475 -606
rect 13559 -982 13593 -606
rect 13677 -982 13711 -606
rect 13790 -982 13824 -606
rect 13908 -982 13942 -606
rect 14026 -982 14060 -606
rect 14144 -982 14178 -606
rect 14262 -982 14296 -606
rect 14380 -982 14414 -606
rect 14498 -982 14532 -606
rect 14617 -982 14651 -606
rect 14735 -982 14769 -606
rect 14853 -982 14887 -606
rect 14971 -982 15005 -606
rect 15090 -982 15124 -806
rect 15208 -982 15242 -806
rect 15326 -982 15360 -806
rect 15444 -982 15478 -806
rect 16026 -982 16060 -806
rect 16144 -982 16178 -806
rect 16262 -982 16296 -806
rect 16380 -982 16414 -806
rect 16467 -982 16501 -606
rect 16585 -982 16619 -606
rect 16703 -982 16737 -606
rect 16821 -982 16855 -606
rect 16934 -982 16968 -606
rect 17052 -982 17086 -606
rect 17170 -982 17204 -606
rect 17288 -982 17322 -606
rect 17406 -982 17440 -606
rect 17524 -982 17558 -606
rect 17642 -982 17676 -606
rect 17761 -982 17795 -606
rect 17879 -982 17913 -606
rect 17997 -982 18031 -606
rect 18115 -982 18149 -606
rect 18234 -982 18268 -806
rect 18352 -982 18386 -806
rect 18470 -982 18504 -806
rect 18588 -982 18622 -806
rect 19158 -978 19192 -802
rect 19276 -978 19310 -802
rect 19394 -978 19428 -802
rect 19512 -978 19546 -802
rect 19599 -978 19633 -602
rect 19717 -978 19751 -602
rect 19835 -978 19869 -602
rect 19953 -978 19987 -602
rect 20066 -978 20100 -602
rect 20184 -978 20218 -602
rect 20302 -978 20336 -602
rect 20420 -978 20454 -602
rect 20538 -978 20572 -602
rect 20656 -978 20690 -602
rect 20774 -978 20808 -602
rect 20893 -978 20927 -602
rect 21011 -978 21045 -602
rect 21129 -978 21163 -602
rect 21247 -978 21281 -602
rect 21366 -978 21400 -802
rect 21484 -978 21518 -802
rect 21602 -978 21636 -802
rect 21720 -978 21754 -802
rect 22302 -978 22336 -802
rect 22420 -978 22454 -802
rect 22538 -978 22572 -802
rect 22656 -978 22690 -802
rect 22743 -978 22777 -602
rect 22861 -978 22895 -602
rect 22979 -978 23013 -602
rect 23097 -978 23131 -602
rect 23210 -978 23244 -602
rect 23328 -978 23362 -602
rect 23446 -978 23480 -602
rect 23564 -978 23598 -602
rect 23682 -978 23716 -602
rect 23800 -978 23834 -602
rect 23918 -978 23952 -602
rect 24037 -978 24071 -602
rect 24155 -978 24189 -602
rect 24273 -978 24307 -602
rect 24391 -978 24425 -602
rect 24510 -978 24544 -802
rect 24628 -978 24662 -802
rect 24746 -978 24780 -802
rect 24864 -978 24898 -802
rect 250 -3714 284 -3538
rect 368 -3714 402 -3538
rect 486 -3714 520 -3538
rect 604 -3714 638 -3538
rect 691 -3714 725 -3338
rect 809 -3714 843 -3338
rect 927 -3714 961 -3338
rect 1045 -3714 1079 -3338
rect 1158 -3714 1192 -3338
rect 1276 -3714 1310 -3338
rect 1394 -3714 1428 -3338
rect 1512 -3714 1546 -3338
rect 1630 -3714 1664 -3338
rect 1748 -3714 1782 -3338
rect 1866 -3714 1900 -3338
rect 1985 -3714 2019 -3338
rect 2103 -3714 2137 -3338
rect 2221 -3714 2255 -3338
rect 2339 -3714 2373 -3338
rect 2458 -3714 2492 -3538
rect 2576 -3714 2610 -3538
rect 2694 -3714 2728 -3538
rect 2812 -3714 2846 -3538
rect 3394 -3714 3428 -3538
rect 3512 -3714 3546 -3538
rect 3630 -3714 3664 -3538
rect 3748 -3714 3782 -3538
rect 3835 -3714 3869 -3338
rect 3953 -3714 3987 -3338
rect 4071 -3714 4105 -3338
rect 4189 -3714 4223 -3338
rect 4302 -3714 4336 -3338
rect 4420 -3714 4454 -3338
rect 4538 -3714 4572 -3338
rect 4656 -3714 4690 -3338
rect 4774 -3714 4808 -3338
rect 4892 -3714 4926 -3338
rect 5010 -3714 5044 -3338
rect 5129 -3714 5163 -3338
rect 5247 -3714 5281 -3338
rect 5365 -3714 5399 -3338
rect 5483 -3714 5517 -3338
rect 5602 -3714 5636 -3538
rect 5720 -3714 5754 -3538
rect 5838 -3714 5872 -3538
rect 5956 -3714 5990 -3538
rect 6526 -3710 6560 -3534
rect 6644 -3710 6678 -3534
rect 6762 -3710 6796 -3534
rect 6880 -3710 6914 -3534
rect 6967 -3710 7001 -3334
rect 7085 -3710 7119 -3334
rect 7203 -3710 7237 -3334
rect 7321 -3710 7355 -3334
rect 7434 -3710 7468 -3334
rect 7552 -3710 7586 -3334
rect 7670 -3710 7704 -3334
rect 7788 -3710 7822 -3334
rect 7906 -3710 7940 -3334
rect 8024 -3710 8058 -3334
rect 8142 -3710 8176 -3334
rect 8261 -3710 8295 -3334
rect 8379 -3710 8413 -3334
rect 8497 -3710 8531 -3334
rect 8615 -3710 8649 -3334
rect 8734 -3710 8768 -3534
rect 8852 -3710 8886 -3534
rect 8970 -3710 9004 -3534
rect 9088 -3710 9122 -3534
rect 9670 -3710 9704 -3534
rect 9788 -3710 9822 -3534
rect 9906 -3710 9940 -3534
rect 10024 -3710 10058 -3534
rect 10111 -3710 10145 -3334
rect 10229 -3710 10263 -3334
rect 10347 -3710 10381 -3334
rect 10465 -3710 10499 -3334
rect 10578 -3710 10612 -3334
rect 10696 -3710 10730 -3334
rect 10814 -3710 10848 -3334
rect 10932 -3710 10966 -3334
rect 11050 -3710 11084 -3334
rect 11168 -3710 11202 -3334
rect 11286 -3710 11320 -3334
rect 11405 -3710 11439 -3334
rect 11523 -3710 11557 -3334
rect 11641 -3710 11675 -3334
rect 11759 -3710 11793 -3334
rect 11878 -3710 11912 -3534
rect 11996 -3710 12030 -3534
rect 12114 -3710 12148 -3534
rect 12232 -3710 12266 -3534
rect 12872 -3714 12906 -3538
rect 12990 -3714 13024 -3538
rect 13108 -3714 13142 -3538
rect 13226 -3714 13260 -3538
rect 13313 -3714 13347 -3338
rect 13431 -3714 13465 -3338
rect 13549 -3714 13583 -3338
rect 13667 -3714 13701 -3338
rect 13780 -3714 13814 -3338
rect 13898 -3714 13932 -3338
rect 14016 -3714 14050 -3338
rect 14134 -3714 14168 -3338
rect 14252 -3714 14286 -3338
rect 14370 -3714 14404 -3338
rect 14488 -3714 14522 -3338
rect 14607 -3714 14641 -3338
rect 14725 -3714 14759 -3338
rect 14843 -3714 14877 -3338
rect 14961 -3714 14995 -3338
rect 15080 -3714 15114 -3538
rect 15198 -3714 15232 -3538
rect 15316 -3714 15350 -3538
rect 15434 -3714 15468 -3538
rect 16016 -3714 16050 -3538
rect 16134 -3714 16168 -3538
rect 16252 -3714 16286 -3538
rect 16370 -3714 16404 -3538
rect 16457 -3714 16491 -3338
rect 16575 -3714 16609 -3338
rect 16693 -3714 16727 -3338
rect 16811 -3714 16845 -3338
rect 16924 -3714 16958 -3338
rect 17042 -3714 17076 -3338
rect 17160 -3714 17194 -3338
rect 17278 -3714 17312 -3338
rect 17396 -3714 17430 -3338
rect 17514 -3714 17548 -3338
rect 17632 -3714 17666 -3338
rect 17751 -3714 17785 -3338
rect 17869 -3714 17903 -3338
rect 17987 -3714 18021 -3338
rect 18105 -3714 18139 -3338
rect 18224 -3714 18258 -3538
rect 18342 -3714 18376 -3538
rect 18460 -3714 18494 -3538
rect 18578 -3714 18612 -3538
rect 19148 -3710 19182 -3534
rect 19266 -3710 19300 -3534
rect 19384 -3710 19418 -3534
rect 19502 -3710 19536 -3534
rect 19589 -3710 19623 -3334
rect 19707 -3710 19741 -3334
rect 19825 -3710 19859 -3334
rect 19943 -3710 19977 -3334
rect 20056 -3710 20090 -3334
rect 20174 -3710 20208 -3334
rect 20292 -3710 20326 -3334
rect 20410 -3710 20444 -3334
rect 20528 -3710 20562 -3334
rect 20646 -3710 20680 -3334
rect 20764 -3710 20798 -3334
rect 20883 -3710 20917 -3334
rect 21001 -3710 21035 -3334
rect 21119 -3710 21153 -3334
rect 21237 -3710 21271 -3334
rect 21356 -3710 21390 -3534
rect 21474 -3710 21508 -3534
rect 21592 -3710 21626 -3534
rect 21710 -3710 21744 -3534
rect 22292 -3710 22326 -3534
rect 22410 -3710 22444 -3534
rect 22528 -3710 22562 -3534
rect 22646 -3710 22680 -3534
rect 22733 -3710 22767 -3334
rect 22851 -3710 22885 -3334
rect 22969 -3710 23003 -3334
rect 23087 -3710 23121 -3334
rect 23200 -3710 23234 -3334
rect 23318 -3710 23352 -3334
rect 23436 -3710 23470 -3334
rect 23554 -3710 23588 -3334
rect 23672 -3710 23706 -3334
rect 23790 -3710 23824 -3334
rect 23908 -3710 23942 -3334
rect 24027 -3710 24061 -3334
rect 24145 -3710 24179 -3334
rect 24263 -3710 24297 -3334
rect 24381 -3710 24415 -3334
rect 24500 -3710 24534 -3534
rect 24618 -3710 24652 -3534
rect 24736 -3710 24770 -3534
rect 24854 -3710 24888 -3534
rect -13 -6659 21 -6483
rect 105 -6659 139 -6483
rect 223 -6659 257 -6483
rect 341 -6659 375 -6483
rect 471 -6659 505 -6283
rect 589 -6659 623 -6283
rect 707 -6659 741 -6283
rect 825 -6659 859 -6283
rect 943 -6659 977 -6283
rect 1061 -6659 1095 -6283
rect 1179 -6659 1213 -6283
rect 1308 -6659 1342 -6483
rect 1426 -6659 1460 -6483
rect 1544 -6659 1578 -6483
rect 1662 -6659 1696 -6483
rect 2055 -6657 2089 -6481
rect 2173 -6657 2207 -6481
rect 2291 -6657 2325 -6481
rect 2409 -6657 2443 -6481
rect 2539 -6657 2573 -6281
rect 2657 -6657 2691 -6281
rect 2775 -6657 2809 -6281
rect 2893 -6657 2927 -6281
rect 3011 -6657 3045 -6281
rect 3129 -6657 3163 -6281
rect 3247 -6657 3281 -6281
rect 3376 -6657 3410 -6481
rect 3494 -6657 3528 -6481
rect 3612 -6657 3646 -6481
rect 3730 -6657 3764 -6481
rect 4124 -6659 4158 -6483
rect 414 -7352 448 -6976
rect 532 -7352 566 -6976
rect 650 -7352 684 -6976
rect 768 -7352 802 -6976
rect 886 -7352 920 -6976
rect 1004 -7352 1038 -6976
rect 1122 -7352 1156 -6976
rect 4242 -6659 4276 -6483
rect 4360 -6659 4394 -6483
rect 4478 -6659 4512 -6483
rect 4608 -6659 4642 -6283
rect 4726 -6659 4760 -6283
rect 4844 -6659 4878 -6283
rect 4962 -6659 4996 -6283
rect 5080 -6659 5114 -6283
rect 5198 -6659 5232 -6283
rect 5316 -6659 5350 -6283
rect 5445 -6659 5479 -6483
rect 5563 -6659 5597 -6483
rect 5681 -6659 5715 -6483
rect 5799 -6659 5833 -6483
rect 6192 -6657 6226 -6481
rect 6310 -6657 6344 -6481
rect 6428 -6657 6462 -6481
rect 6546 -6657 6580 -6481
rect 6676 -6657 6710 -6281
rect 6794 -6657 6828 -6281
rect 6912 -6657 6946 -6281
rect 7030 -6657 7064 -6281
rect 7148 -6657 7182 -6281
rect 7266 -6657 7300 -6281
rect 7384 -6657 7418 -6281
rect 7513 -6657 7547 -6481
rect 7631 -6657 7665 -6481
rect 7749 -6657 7783 -6481
rect 7867 -6657 7901 -6481
rect 8261 -6657 8295 -6481
rect 8379 -6657 8413 -6481
rect 8497 -6657 8531 -6481
rect 8615 -6657 8649 -6481
rect 8745 -6657 8779 -6281
rect 8863 -6657 8897 -6281
rect 8981 -6657 9015 -6281
rect 9099 -6657 9133 -6281
rect 9217 -6657 9251 -6281
rect 9335 -6657 9369 -6281
rect 9453 -6657 9487 -6281
rect 9582 -6657 9616 -6481
rect 9700 -6657 9734 -6481
rect 9818 -6657 9852 -6481
rect 9936 -6657 9970 -6481
rect 10329 -6655 10363 -6479
rect 10447 -6655 10481 -6479
rect 10565 -6655 10599 -6479
rect 10683 -6655 10717 -6479
rect 10813 -6655 10847 -6279
rect 10931 -6655 10965 -6279
rect 11049 -6655 11083 -6279
rect 11167 -6655 11201 -6279
rect 11285 -6655 11319 -6279
rect 11403 -6655 11437 -6279
rect 11521 -6655 11555 -6279
rect 11650 -6655 11684 -6479
rect 11768 -6655 11802 -6479
rect 11886 -6655 11920 -6479
rect 12004 -6655 12038 -6479
rect 12398 -6657 12432 -6481
rect 2482 -7350 2516 -6974
rect 2600 -7350 2634 -6974
rect 2718 -7350 2752 -6974
rect 2836 -7350 2870 -6974
rect 2954 -7350 2988 -6974
rect 3072 -7350 3106 -6974
rect 3190 -7350 3224 -6974
rect 4551 -7352 4585 -6976
rect 4669 -7352 4703 -6976
rect 4787 -7352 4821 -6976
rect 4905 -7352 4939 -6976
rect 5023 -7352 5057 -6976
rect 5141 -7352 5175 -6976
rect 5259 -7352 5293 -6976
rect 6619 -7350 6653 -6974
rect 6737 -7350 6771 -6974
rect 6855 -7350 6889 -6974
rect 6973 -7350 7007 -6974
rect 7091 -7350 7125 -6974
rect 7209 -7350 7243 -6974
rect 7327 -7350 7361 -6974
rect 8688 -7350 8722 -6974
rect 8806 -7350 8840 -6974
rect 8924 -7350 8958 -6974
rect 9042 -7350 9076 -6974
rect 9160 -7350 9194 -6974
rect 9278 -7350 9312 -6974
rect 9396 -7350 9430 -6974
rect 12516 -6657 12550 -6481
rect 12634 -6657 12668 -6481
rect 12752 -6657 12786 -6481
rect 12882 -6657 12916 -6281
rect 13000 -6657 13034 -6281
rect 13118 -6657 13152 -6281
rect 13236 -6657 13270 -6281
rect 13354 -6657 13388 -6281
rect 13472 -6657 13506 -6281
rect 13590 -6657 13624 -6281
rect 13719 -6657 13753 -6481
rect 13837 -6657 13871 -6481
rect 13955 -6657 13989 -6481
rect 14073 -6657 14107 -6481
rect 14466 -6655 14500 -6479
rect 14584 -6655 14618 -6479
rect 14702 -6655 14736 -6479
rect 14820 -6655 14854 -6479
rect 14950 -6655 14984 -6279
rect 15068 -6655 15102 -6279
rect 15186 -6655 15220 -6279
rect 15304 -6655 15338 -6279
rect 15422 -6655 15456 -6279
rect 15540 -6655 15574 -6279
rect 15658 -6655 15692 -6279
rect 16719 -6343 16753 -6167
rect 16837 -6343 16871 -6167
rect 16955 -6343 16989 -6167
rect 17073 -6343 17107 -6167
rect 17457 -6339 17491 -6163
rect 17575 -6339 17609 -6163
rect 17693 -6339 17727 -6163
rect 17811 -6339 17845 -6163
rect 18195 -6343 18229 -6167
rect 18313 -6343 18347 -6167
rect 18431 -6343 18465 -6167
rect 18549 -6343 18583 -6167
rect 18937 -6345 18971 -6169
rect 19055 -6345 19089 -6169
rect 19173 -6345 19207 -6169
rect 19291 -6345 19325 -6169
rect 19677 -6345 19711 -6169
rect 19795 -6345 19829 -6169
rect 19913 -6345 19947 -6169
rect 20031 -6345 20065 -6169
rect 20415 -6345 20449 -6169
rect 20533 -6345 20567 -6169
rect 20651 -6345 20685 -6169
rect 20769 -6345 20803 -6169
rect 21153 -6345 21187 -6169
rect 21271 -6345 21305 -6169
rect 21389 -6345 21423 -6169
rect 21507 -6345 21541 -6169
rect 21891 -6345 21925 -6169
rect 22009 -6345 22043 -6169
rect 22127 -6345 22161 -6169
rect 22245 -6345 22279 -6169
rect 15787 -6655 15821 -6479
rect 15905 -6655 15939 -6479
rect 16023 -6655 16057 -6479
rect 16141 -6655 16175 -6479
rect 10756 -7348 10790 -6972
rect 10874 -7348 10908 -6972
rect 10992 -7348 11026 -6972
rect 11110 -7348 11144 -6972
rect 11228 -7348 11262 -6972
rect 11346 -7348 11380 -6972
rect 11464 -7348 11498 -6972
rect 12825 -7350 12859 -6974
rect 12943 -7350 12977 -6974
rect 13061 -7350 13095 -6974
rect 13179 -7350 13213 -6974
rect 13297 -7350 13331 -6974
rect 13415 -7350 13449 -6974
rect 13533 -7350 13567 -6974
rect 14893 -7348 14927 -6972
rect 15011 -7348 15045 -6972
rect 15129 -7348 15163 -6972
rect 15247 -7348 15281 -6972
rect 15365 -7348 15399 -6972
rect 15483 -7348 15517 -6972
rect 15601 -7348 15635 -6972
<< psubdiff >>
rect 11996 2988 12192 3018
rect 690 2917 902 2947
rect 690 2861 730 2917
rect 864 2861 902 2917
rect 690 2839 902 2861
rect 2138 2917 2350 2947
rect 2138 2861 2178 2917
rect 2312 2861 2350 2917
rect 2138 2839 2350 2861
rect 3636 2919 3848 2949
rect 3636 2863 3676 2919
rect 3810 2863 3848 2919
rect 3636 2841 3848 2863
rect 5084 2919 5296 2949
rect 5084 2863 5124 2919
rect 5258 2863 5296 2919
rect 5084 2841 5296 2863
rect 6604 2917 6816 2947
rect 6604 2861 6644 2917
rect 6778 2861 6816 2917
rect 6604 2839 6816 2861
rect 8052 2917 8264 2947
rect 8052 2861 8092 2917
rect 8226 2861 8264 2917
rect 8052 2839 8264 2861
rect 9550 2919 9762 2949
rect 9550 2863 9590 2919
rect 9724 2863 9762 2919
rect 9550 2841 9762 2863
rect 10998 2919 11210 2949
rect 10998 2863 11038 2919
rect 11172 2863 11210 2919
rect 11996 2922 12036 2988
rect 12154 2922 12192 2988
rect 11996 2874 12192 2922
rect 13164 2988 13360 3018
rect 13164 2922 13204 2988
rect 13322 2922 13360 2988
rect 13164 2874 13360 2922
rect 14332 2988 14528 3018
rect 14332 2922 14372 2988
rect 14490 2922 14528 2988
rect 14332 2874 14528 2922
rect 15500 2988 15696 3018
rect 15500 2922 15540 2988
rect 15658 2922 15696 2988
rect 15500 2874 15696 2922
rect 16674 2990 16870 3020
rect 16674 2924 16714 2990
rect 16832 2924 16870 2990
rect 16674 2876 16870 2924
rect 17842 2990 18038 3020
rect 17842 2924 17882 2990
rect 18000 2924 18038 2990
rect 17842 2876 18038 2924
rect 19010 2990 19206 3020
rect 19010 2924 19050 2990
rect 19168 2924 19206 2990
rect 19010 2876 19206 2924
rect 20178 2990 20374 3020
rect 20178 2924 20218 2990
rect 20336 2924 20374 2990
rect 20178 2876 20374 2924
rect 10998 2841 11210 2863
rect 1462 152 1648 176
rect 1462 106 1504 152
rect 1608 106 1648 152
rect 1462 70 1648 106
rect 4606 152 4792 176
rect 4606 106 4648 152
rect 4752 106 4792 152
rect 4606 70 4792 106
rect 7738 156 7924 180
rect 7738 110 7780 156
rect 7884 110 7924 156
rect 7738 74 7924 110
rect 10882 156 11068 180
rect 10882 110 10924 156
rect 11028 110 11068 156
rect 10882 74 11068 110
rect 14084 152 14270 176
rect 14084 106 14126 152
rect 14230 106 14270 152
rect 14084 70 14270 106
rect 17228 152 17414 176
rect 17228 106 17270 152
rect 17374 106 17414 152
rect 17228 70 17414 106
rect 20360 156 20546 180
rect 20360 110 20402 156
rect 20506 110 20546 156
rect 20360 74 20546 110
rect 23504 156 23690 180
rect 23504 110 23546 156
rect 23650 110 23690 156
rect 23504 74 23690 110
rect 1462 -2582 1648 -2558
rect 1462 -2628 1504 -2582
rect 1608 -2628 1648 -2582
rect 1462 -2664 1648 -2628
rect 4606 -2582 4792 -2558
rect 4606 -2628 4648 -2582
rect 4752 -2628 4792 -2582
rect 4606 -2664 4792 -2628
rect 7738 -2578 7924 -2554
rect 7738 -2624 7780 -2578
rect 7884 -2624 7924 -2578
rect 7738 -2660 7924 -2624
rect 10882 -2578 11068 -2554
rect 10882 -2624 10924 -2578
rect 11028 -2624 11068 -2578
rect 10882 -2660 11068 -2624
rect 14084 -2582 14270 -2558
rect 14084 -2628 14126 -2582
rect 14230 -2628 14270 -2582
rect 14084 -2664 14270 -2628
rect 17228 -2582 17414 -2558
rect 17228 -2628 17270 -2582
rect 17374 -2628 17414 -2582
rect 17228 -2664 17414 -2628
rect 20360 -2578 20546 -2554
rect 20360 -2624 20402 -2578
rect 20506 -2624 20546 -2578
rect 20360 -2660 20546 -2624
rect 23504 -2578 23690 -2554
rect 23504 -2624 23546 -2578
rect 23650 -2624 23690 -2578
rect 23504 -2660 23690 -2624
rect 1452 -5314 1638 -5290
rect 1452 -5360 1494 -5314
rect 1598 -5360 1638 -5314
rect 1452 -5396 1638 -5360
rect 4596 -5314 4782 -5290
rect 4596 -5360 4638 -5314
rect 4742 -5360 4782 -5314
rect 4596 -5396 4782 -5360
rect 7728 -5310 7914 -5286
rect 7728 -5356 7770 -5310
rect 7874 -5356 7914 -5310
rect 7728 -5392 7914 -5356
rect 10872 -5310 11058 -5286
rect 10872 -5356 10914 -5310
rect 11018 -5356 11058 -5310
rect 10872 -5392 11058 -5356
rect 14074 -5314 14260 -5290
rect 14074 -5360 14116 -5314
rect 14220 -5360 14260 -5314
rect 14074 -5396 14260 -5360
rect 17218 -5314 17404 -5290
rect 17218 -5360 17260 -5314
rect 17364 -5360 17404 -5314
rect 17218 -5396 17404 -5360
rect 20350 -5310 20536 -5286
rect 20350 -5356 20392 -5310
rect 20496 -5356 20536 -5310
rect 20350 -5392 20536 -5356
rect 23494 -5310 23680 -5286
rect 23494 -5356 23536 -5310
rect 23640 -5356 23680 -5310
rect 23494 -5392 23680 -5356
rect 16715 -6841 16975 -6795
rect 16715 -6911 16777 -6841
rect 16921 -6911 16975 -6841
rect 16715 -6945 16975 -6911
rect 17453 -6843 17713 -6797
rect 17453 -6913 17515 -6843
rect 17659 -6913 17713 -6843
rect 17453 -6947 17713 -6913
rect 18191 -6843 18451 -6797
rect 18191 -6913 18253 -6843
rect 18397 -6913 18451 -6843
rect 18191 -6947 18451 -6913
rect 18933 -6843 19193 -6797
rect 18933 -6913 18995 -6843
rect 19139 -6913 19193 -6843
rect 18933 -6947 19193 -6913
rect 19673 -6843 19933 -6797
rect 19673 -6913 19735 -6843
rect 19879 -6913 19933 -6843
rect 19673 -6947 19933 -6913
rect 20411 -6843 20671 -6797
rect 20411 -6913 20473 -6843
rect 20617 -6913 20671 -6843
rect 20411 -6947 20671 -6913
rect 21149 -6843 21409 -6797
rect 21149 -6913 21211 -6843
rect 21355 -6913 21409 -6843
rect 21149 -6947 21409 -6913
rect 21887 -6843 22147 -6797
rect 21887 -6913 21949 -6843
rect 22093 -6913 22147 -6843
rect 21887 -6947 22147 -6913
rect 664 -8272 916 -8252
rect 664 -8328 722 -8272
rect 854 -8328 916 -8272
rect 664 -8350 916 -8328
rect 2732 -8270 2984 -8250
rect 2732 -8326 2790 -8270
rect 2922 -8326 2984 -8270
rect 2732 -8348 2984 -8326
rect 4801 -8272 5053 -8252
rect 4801 -8328 4859 -8272
rect 4991 -8328 5053 -8272
rect 4801 -8350 5053 -8328
rect 6869 -8270 7121 -8250
rect 6869 -8326 6927 -8270
rect 7059 -8326 7121 -8270
rect 6869 -8348 7121 -8326
rect 8938 -8270 9190 -8250
rect 8938 -8326 8996 -8270
rect 9128 -8326 9190 -8270
rect 8938 -8348 9190 -8326
rect 11006 -8268 11258 -8248
rect 11006 -8324 11064 -8268
rect 11196 -8324 11258 -8268
rect 11006 -8346 11258 -8324
rect 13075 -8270 13327 -8250
rect 13075 -8326 13133 -8270
rect 13265 -8326 13327 -8270
rect 13075 -8348 13327 -8326
rect 15143 -8268 15395 -8248
rect 15143 -8324 15201 -8268
rect 15333 -8324 15395 -8268
rect 15143 -8346 15395 -8324
<< nsubdiff >>
rect 12436 4332 12702 4370
rect 12436 4260 12492 4332
rect 12636 4260 12702 4332
rect 13604 4332 13870 4370
rect 12436 4230 12702 4260
rect 450 4125 694 4163
rect 450 4055 506 4125
rect 642 4055 694 4125
rect 450 4033 694 4055
rect 1898 4125 2142 4163
rect 1898 4055 1954 4125
rect 2090 4055 2142 4125
rect 1898 4033 2142 4055
rect 3396 4127 3640 4165
rect 3396 4057 3452 4127
rect 3588 4057 3640 4127
rect 3396 4035 3640 4057
rect 4844 4127 5088 4165
rect 4844 4057 4900 4127
rect 5036 4057 5088 4127
rect 4844 4035 5088 4057
rect 6364 4125 6608 4163
rect 6364 4055 6420 4125
rect 6556 4055 6608 4125
rect 6364 4033 6608 4055
rect 7812 4125 8056 4163
rect 7812 4055 7868 4125
rect 8004 4055 8056 4125
rect 7812 4033 8056 4055
rect 9310 4127 9554 4165
rect 9310 4057 9366 4127
rect 9502 4057 9554 4127
rect 9310 4035 9554 4057
rect 10758 4127 11002 4165
rect 10758 4057 10814 4127
rect 10950 4057 11002 4127
rect 13604 4260 13660 4332
rect 13804 4260 13870 4332
rect 14772 4332 15038 4370
rect 13604 4230 13870 4260
rect 14772 4260 14828 4332
rect 14972 4260 15038 4332
rect 15940 4332 16206 4370
rect 14772 4230 15038 4260
rect 15940 4260 15996 4332
rect 16140 4260 16206 4332
rect 17114 4334 17380 4372
rect 15940 4230 16206 4260
rect 17114 4262 17170 4334
rect 17314 4262 17380 4334
rect 18282 4334 18548 4372
rect 17114 4232 17380 4262
rect 18282 4262 18338 4334
rect 18482 4262 18548 4334
rect 19450 4334 19716 4372
rect 18282 4232 18548 4262
rect 19450 4262 19506 4334
rect 19650 4262 19716 4334
rect 20618 4334 20884 4372
rect 19450 4232 19716 4262
rect 20618 4262 20674 4334
rect 20818 4262 20884 4334
rect 20618 4232 20884 4262
rect 10758 4035 11002 4057
rect 1392 2398 1696 2454
rect 1392 2322 1446 2398
rect 1642 2322 1696 2398
rect 1392 2308 1696 2322
rect 4536 2398 4840 2454
rect 4536 2322 4590 2398
rect 4786 2322 4840 2398
rect 4536 2308 4840 2322
rect 7668 2402 7972 2458
rect 7668 2326 7722 2402
rect 7918 2326 7972 2402
rect 7668 2312 7972 2326
rect 10812 2402 11116 2458
rect 10812 2326 10866 2402
rect 11062 2326 11116 2402
rect 10812 2312 11116 2326
rect 14014 2398 14318 2454
rect 14014 2322 14068 2398
rect 14264 2322 14318 2398
rect 14014 2308 14318 2322
rect 17158 2398 17462 2454
rect 17158 2322 17212 2398
rect 17408 2322 17462 2398
rect 17158 2308 17462 2322
rect 20290 2402 20594 2458
rect 20290 2326 20344 2402
rect 20540 2326 20594 2402
rect 20290 2312 20594 2326
rect 23434 2402 23738 2458
rect 23434 2326 23488 2402
rect 23684 2326 23738 2402
rect 23434 2312 23738 2326
rect 1392 -336 1696 -280
rect 1392 -412 1446 -336
rect 1642 -412 1696 -336
rect 1392 -426 1696 -412
rect 4536 -336 4840 -280
rect 4536 -412 4590 -336
rect 4786 -412 4840 -336
rect 4536 -426 4840 -412
rect 7668 -332 7972 -276
rect 7668 -408 7722 -332
rect 7918 -408 7972 -332
rect 7668 -422 7972 -408
rect 10812 -332 11116 -276
rect 10812 -408 10866 -332
rect 11062 -408 11116 -332
rect 10812 -422 11116 -408
rect 14014 -336 14318 -280
rect 14014 -412 14068 -336
rect 14264 -412 14318 -336
rect 14014 -426 14318 -412
rect 17158 -336 17462 -280
rect 17158 -412 17212 -336
rect 17408 -412 17462 -336
rect 17158 -426 17462 -412
rect 20290 -332 20594 -276
rect 20290 -408 20344 -332
rect 20540 -408 20594 -332
rect 20290 -422 20594 -408
rect 23434 -332 23738 -276
rect 23434 -408 23488 -332
rect 23684 -408 23738 -332
rect 23434 -422 23738 -408
rect 1382 -3068 1686 -3012
rect 1382 -3144 1436 -3068
rect 1632 -3144 1686 -3068
rect 1382 -3158 1686 -3144
rect 4526 -3068 4830 -3012
rect 4526 -3144 4580 -3068
rect 4776 -3144 4830 -3068
rect 4526 -3158 4830 -3144
rect 7658 -3064 7962 -3008
rect 7658 -3140 7712 -3064
rect 7908 -3140 7962 -3064
rect 7658 -3154 7962 -3140
rect 10802 -3064 11106 -3008
rect 10802 -3140 10856 -3064
rect 11052 -3140 11106 -3064
rect 10802 -3154 11106 -3140
rect 14004 -3068 14308 -3012
rect 14004 -3144 14058 -3068
rect 14254 -3144 14308 -3068
rect 14004 -3158 14308 -3144
rect 17148 -3068 17452 -3012
rect 17148 -3144 17202 -3068
rect 17398 -3144 17452 -3068
rect 17148 -3158 17452 -3144
rect 20280 -3064 20584 -3008
rect 20280 -3140 20334 -3064
rect 20530 -3140 20584 -3064
rect 20280 -3154 20584 -3140
rect 23424 -3064 23728 -3008
rect 23424 -3140 23478 -3064
rect 23674 -3140 23728 -3064
rect 23424 -3154 23728 -3140
rect 648 -6012 1048 -5960
rect 648 -6056 772 -6012
rect 894 -6056 1048 -6012
rect 648 -6104 1048 -6056
rect 2716 -6010 3116 -5958
rect 2716 -6054 2840 -6010
rect 2962 -6054 3116 -6010
rect 2716 -6102 3116 -6054
rect 4785 -6012 5185 -5960
rect 4785 -6056 4909 -6012
rect 5031 -6056 5185 -6012
rect 4785 -6104 5185 -6056
rect 6853 -6010 7253 -5958
rect 6853 -6054 6977 -6010
rect 7099 -6054 7253 -6010
rect 6853 -6102 7253 -6054
rect 8922 -6010 9322 -5958
rect 8922 -6054 9046 -6010
rect 9168 -6054 9322 -6010
rect 8922 -6102 9322 -6054
rect 10990 -6008 11390 -5956
rect 10990 -6052 11114 -6008
rect 11236 -6052 11390 -6008
rect 10990 -6100 11390 -6052
rect 13059 -6010 13459 -5958
rect 13059 -6054 13183 -6010
rect 13305 -6054 13459 -6010
rect 13059 -6102 13459 -6054
rect 15127 -6008 15527 -5956
rect 15127 -6052 15251 -6008
rect 15373 -6052 15527 -6008
rect 15127 -6100 15527 -6052
rect 16765 -5961 17061 -5947
rect 16765 -6023 16843 -5961
rect 16983 -6023 17061 -5961
rect 16765 -6079 17061 -6023
rect 17503 -5963 17799 -5949
rect 17503 -6025 17581 -5963
rect 17721 -6025 17799 -5963
rect 17503 -6081 17799 -6025
rect 18241 -5963 18537 -5949
rect 18241 -6025 18319 -5963
rect 18459 -6025 18537 -5963
rect 18241 -6081 18537 -6025
rect 18983 -5963 19279 -5949
rect 18983 -6025 19061 -5963
rect 19201 -6025 19279 -5963
rect 18983 -6081 19279 -6025
rect 19723 -5963 20019 -5949
rect 19723 -6025 19801 -5963
rect 19941 -6025 20019 -5963
rect 19723 -6081 20019 -6025
rect 20461 -5963 20757 -5949
rect 20461 -6025 20539 -5963
rect 20679 -6025 20757 -5963
rect 20461 -6081 20757 -6025
rect 21199 -5963 21495 -5949
rect 21199 -6025 21277 -5963
rect 21417 -6025 21495 -5963
rect 21199 -6081 21495 -6025
rect 21937 -5963 22233 -5949
rect 21937 -6025 22015 -5963
rect 22155 -6025 22233 -5963
rect 21937 -6081 22233 -6025
<< psubdiffcont >>
rect 730 2861 864 2917
rect 2178 2861 2312 2917
rect 3676 2863 3810 2919
rect 5124 2863 5258 2919
rect 6644 2861 6778 2917
rect 8092 2861 8226 2917
rect 9590 2863 9724 2919
rect 11038 2863 11172 2919
rect 12036 2922 12154 2988
rect 13204 2922 13322 2988
rect 14372 2922 14490 2988
rect 15540 2922 15658 2988
rect 16714 2924 16832 2990
rect 17882 2924 18000 2990
rect 19050 2924 19168 2990
rect 20218 2924 20336 2990
rect 1504 106 1608 152
rect 4648 106 4752 152
rect 7780 110 7884 156
rect 10924 110 11028 156
rect 14126 106 14230 152
rect 17270 106 17374 152
rect 20402 110 20506 156
rect 23546 110 23650 156
rect 1504 -2628 1608 -2582
rect 4648 -2628 4752 -2582
rect 7780 -2624 7884 -2578
rect 10924 -2624 11028 -2578
rect 14126 -2628 14230 -2582
rect 17270 -2628 17374 -2582
rect 20402 -2624 20506 -2578
rect 23546 -2624 23650 -2578
rect 1494 -5360 1598 -5314
rect 4638 -5360 4742 -5314
rect 7770 -5356 7874 -5310
rect 10914 -5356 11018 -5310
rect 14116 -5360 14220 -5314
rect 17260 -5360 17364 -5314
rect 20392 -5356 20496 -5310
rect 23536 -5356 23640 -5310
rect 16777 -6911 16921 -6841
rect 17515 -6913 17659 -6843
rect 18253 -6913 18397 -6843
rect 18995 -6913 19139 -6843
rect 19735 -6913 19879 -6843
rect 20473 -6913 20617 -6843
rect 21211 -6913 21355 -6843
rect 21949 -6913 22093 -6843
rect 722 -8328 854 -8272
rect 2790 -8326 2922 -8270
rect 4859 -8328 4991 -8272
rect 6927 -8326 7059 -8270
rect 8996 -8326 9128 -8270
rect 11064 -8324 11196 -8268
rect 13133 -8326 13265 -8270
rect 15201 -8324 15333 -8268
<< nsubdiffcont >>
rect 12492 4260 12636 4332
rect 506 4055 642 4125
rect 1954 4055 2090 4125
rect 3452 4057 3588 4127
rect 4900 4057 5036 4127
rect 6420 4055 6556 4125
rect 7868 4055 8004 4125
rect 9366 4057 9502 4127
rect 10814 4057 10950 4127
rect 13660 4260 13804 4332
rect 14828 4260 14972 4332
rect 15996 4260 16140 4332
rect 17170 4262 17314 4334
rect 18338 4262 18482 4334
rect 19506 4262 19650 4334
rect 20674 4262 20818 4334
rect 1446 2322 1642 2398
rect 4590 2322 4786 2398
rect 7722 2326 7918 2402
rect 10866 2326 11062 2402
rect 14068 2322 14264 2398
rect 17212 2322 17408 2398
rect 20344 2326 20540 2402
rect 23488 2326 23684 2402
rect 1446 -412 1642 -336
rect 4590 -412 4786 -336
rect 7722 -408 7918 -332
rect 10866 -408 11062 -332
rect 14068 -412 14264 -336
rect 17212 -412 17408 -336
rect 20344 -408 20540 -332
rect 23488 -408 23684 -332
rect 1436 -3144 1632 -3068
rect 4580 -3144 4776 -3068
rect 7712 -3140 7908 -3064
rect 10856 -3140 11052 -3064
rect 14058 -3144 14254 -3068
rect 17202 -3144 17398 -3068
rect 20334 -3140 20530 -3064
rect 23478 -3140 23674 -3064
rect 772 -6056 894 -6012
rect 2840 -6054 2962 -6010
rect 4909 -6056 5031 -6012
rect 6977 -6054 7099 -6010
rect 9046 -6054 9168 -6010
rect 11114 -6052 11236 -6008
rect 13183 -6054 13305 -6010
rect 15251 -6052 15373 -6008
rect 16843 -6023 16983 -5961
rect 17581 -6025 17721 -5963
rect 18319 -6025 18459 -5963
rect 19061 -6025 19201 -5963
rect 19801 -6025 19941 -5963
rect 20539 -6025 20679 -5963
rect 21277 -6025 21417 -5963
rect 22015 -6025 22155 -5963
<< poly >>
rect 11858 4254 11924 4270
rect 11858 4220 11874 4254
rect 11908 4250 11924 4254
rect 11908 4220 12408 4250
rect 13026 4254 13092 4270
rect 11858 4207 12408 4220
rect 11858 4204 11924 4207
rect 11858 4155 11924 4162
rect 12364 4155 12408 4207
rect 13026 4220 13042 4254
rect 13076 4250 13092 4254
rect 13076 4220 13576 4250
rect 14194 4254 14260 4270
rect 13026 4207 13576 4220
rect 13026 4204 13092 4207
rect 13026 4155 13092 4162
rect 13532 4155 13576 4207
rect 14194 4220 14210 4254
rect 14244 4250 14260 4254
rect 14244 4220 14744 4250
rect 15362 4254 15428 4270
rect 14194 4207 14744 4220
rect 14194 4204 14260 4207
rect 14194 4155 14260 4162
rect 14700 4155 14744 4207
rect 15362 4220 15378 4254
rect 15412 4250 15428 4254
rect 15412 4220 15912 4250
rect 16536 4256 16602 4272
rect 15362 4207 15912 4220
rect 15362 4204 15428 4207
rect 15362 4155 15428 4162
rect 15868 4155 15912 4207
rect 16536 4222 16552 4256
rect 16586 4252 16602 4256
rect 16586 4222 17086 4252
rect 17704 4256 17770 4272
rect 16536 4209 17086 4222
rect 16536 4206 16602 4209
rect 16536 4157 16602 4164
rect 17042 4157 17086 4209
rect 17704 4222 17720 4256
rect 17754 4252 17770 4256
rect 17754 4222 18254 4252
rect 18872 4256 18938 4272
rect 17704 4209 18254 4222
rect 17704 4206 17770 4209
rect 17704 4157 17770 4164
rect 18210 4157 18254 4209
rect 18872 4222 18888 4256
rect 18922 4252 18938 4256
rect 18922 4222 19422 4252
rect 20040 4256 20106 4272
rect 18872 4209 19422 4222
rect 18872 4206 18938 4209
rect 18872 4157 18938 4164
rect 19378 4157 19422 4209
rect 20040 4222 20056 4256
rect 20090 4252 20106 4256
rect 20090 4222 20590 4252
rect 20040 4209 20590 4222
rect 20040 4206 20106 4209
rect 20040 4157 20106 4164
rect 20546 4157 20590 4209
rect 11858 4146 12306 4155
rect 11858 4112 11874 4146
rect 11908 4114 12306 4146
rect 11908 4113 12070 4114
rect 11908 4112 11924 4113
rect 11858 4096 11924 4112
rect 12010 4094 12070 4113
rect 12128 4094 12188 4114
rect 12246 4094 12306 4114
rect 12364 4114 12660 4155
rect 12364 4094 12424 4114
rect 12482 4094 12542 4114
rect 12600 4094 12660 4114
rect 13026 4146 13474 4155
rect 13026 4112 13042 4146
rect 13076 4114 13474 4146
rect 13076 4113 13238 4114
rect 13076 4112 13092 4113
rect 13026 4096 13092 4112
rect 13178 4094 13238 4113
rect 13296 4094 13356 4114
rect 13414 4094 13474 4114
rect 13532 4114 13828 4155
rect 13532 4094 13592 4114
rect 13650 4094 13710 4114
rect 13768 4094 13828 4114
rect 14194 4146 14642 4155
rect 14194 4112 14210 4146
rect 14244 4114 14642 4146
rect 14244 4113 14406 4114
rect 14244 4112 14260 4113
rect 14194 4096 14260 4112
rect 247 3918 543 3954
rect 247 3897 307 3918
rect 365 3897 425 3918
rect 483 3897 543 3918
rect 601 3917 897 3953
rect 601 3897 661 3917
rect 719 3897 779 3917
rect 837 3897 897 3917
rect 955 3917 1251 3953
rect 955 3897 1015 3917
rect 1073 3897 1133 3917
rect 1191 3897 1251 3917
rect 1695 3918 1991 3954
rect 1695 3897 1755 3918
rect 1813 3897 1873 3918
rect 1931 3897 1991 3918
rect 2049 3917 2345 3953
rect 2049 3897 2109 3917
rect 2167 3897 2227 3917
rect 2285 3897 2345 3917
rect 2403 3917 2699 3953
rect 2403 3897 2463 3917
rect 2521 3897 2581 3917
rect 2639 3897 2699 3917
rect 3193 3920 3489 3956
rect 3193 3899 3253 3920
rect 3311 3899 3371 3920
rect 3429 3899 3489 3920
rect 3547 3919 3843 3955
rect 3547 3899 3607 3919
rect 3665 3899 3725 3919
rect 3783 3899 3843 3919
rect 3901 3919 4197 3955
rect 3901 3899 3961 3919
rect 4019 3899 4079 3919
rect 4137 3899 4197 3919
rect 4641 3920 4937 3956
rect 4641 3899 4701 3920
rect 4759 3899 4819 3920
rect 4877 3899 4937 3920
rect 4995 3919 5291 3955
rect 4995 3899 5055 3919
rect 5113 3899 5173 3919
rect 5231 3899 5291 3919
rect 5349 3919 5645 3955
rect 5349 3899 5409 3919
rect 5467 3899 5527 3919
rect 5585 3899 5645 3919
rect 6161 3918 6457 3954
rect 6161 3897 6221 3918
rect 6279 3897 6339 3918
rect 6397 3897 6457 3918
rect 6515 3917 6811 3953
rect 6515 3897 6575 3917
rect 6633 3897 6693 3917
rect 6751 3897 6811 3917
rect 6869 3917 7165 3953
rect 6869 3897 6929 3917
rect 6987 3897 7047 3917
rect 7105 3897 7165 3917
rect 7609 3918 7905 3954
rect 7609 3897 7669 3918
rect 7727 3897 7787 3918
rect 7845 3897 7905 3918
rect 7963 3917 8259 3953
rect 7963 3897 8023 3917
rect 8081 3897 8141 3917
rect 8199 3897 8259 3917
rect 8317 3917 8613 3953
rect 8317 3897 8377 3917
rect 8435 3897 8495 3917
rect 8553 3897 8613 3917
rect 9107 3920 9403 3956
rect 9107 3899 9167 3920
rect 9225 3899 9285 3920
rect 9343 3899 9403 3920
rect 9461 3919 9757 3955
rect 9461 3899 9521 3919
rect 9579 3899 9639 3919
rect 9697 3899 9757 3919
rect 9815 3919 10111 3955
rect 9815 3899 9875 3919
rect 9933 3899 9993 3919
rect 10051 3899 10111 3919
rect 10555 3920 10851 3956
rect 10555 3899 10615 3920
rect 10673 3899 10733 3920
rect 10791 3899 10851 3920
rect 10909 3919 11205 3955
rect 10909 3899 10969 3919
rect 11027 3899 11087 3919
rect 11145 3899 11205 3919
rect 11263 3919 11559 3955
rect 11263 3899 11323 3919
rect 11381 3899 11441 3919
rect 11499 3899 11559 3919
rect 247 3671 307 3697
rect 365 3671 425 3697
rect 483 3671 543 3697
rect 601 3677 661 3697
rect 601 3671 662 3677
rect 719 3671 779 3697
rect 837 3671 897 3697
rect 484 3486 542 3671
rect 484 3460 544 3486
rect 602 3460 662 3671
rect 955 3665 1015 3697
rect 1073 3671 1133 3697
rect 1191 3671 1251 3697
rect 1695 3671 1755 3697
rect 1813 3671 1873 3697
rect 1931 3671 1991 3697
rect 2049 3677 2109 3697
rect 2049 3671 2110 3677
rect 2167 3671 2227 3697
rect 2285 3671 2345 3697
rect 952 3649 1018 3665
rect 952 3615 968 3649
rect 1002 3615 1018 3649
rect 952 3599 1018 3615
rect 834 3532 900 3548
rect 834 3498 850 3532
rect 884 3498 900 3532
rect 834 3482 900 3498
rect 1932 3486 1990 3671
rect 837 3460 897 3482
rect 1932 3460 1992 3486
rect 2050 3460 2110 3671
rect 2403 3665 2463 3697
rect 2521 3671 2581 3697
rect 2639 3671 2699 3697
rect 3193 3673 3253 3699
rect 3311 3673 3371 3699
rect 3429 3673 3489 3699
rect 3547 3679 3607 3699
rect 3547 3673 3608 3679
rect 3665 3673 3725 3699
rect 3783 3673 3843 3699
rect 2400 3649 2466 3665
rect 2400 3615 2416 3649
rect 2450 3615 2466 3649
rect 2400 3599 2466 3615
rect 2282 3532 2348 3548
rect 2282 3498 2298 3532
rect 2332 3498 2348 3532
rect 2282 3482 2348 3498
rect 3430 3488 3488 3673
rect 2285 3460 2345 3482
rect 3430 3462 3490 3488
rect 3548 3462 3608 3673
rect 3901 3667 3961 3699
rect 4019 3673 4079 3699
rect 4137 3673 4197 3699
rect 4641 3673 4701 3699
rect 4759 3673 4819 3699
rect 4877 3673 4937 3699
rect 4995 3679 5055 3699
rect 4995 3673 5056 3679
rect 5113 3673 5173 3699
rect 5231 3673 5291 3699
rect 3898 3651 3964 3667
rect 3898 3617 3914 3651
rect 3948 3617 3964 3651
rect 3898 3601 3964 3617
rect 3780 3534 3846 3550
rect 3780 3500 3796 3534
rect 3830 3500 3846 3534
rect 3780 3484 3846 3500
rect 4878 3488 4936 3673
rect 3783 3462 3843 3484
rect 4878 3462 4938 3488
rect 4996 3462 5056 3673
rect 5349 3667 5409 3699
rect 5467 3673 5527 3699
rect 5585 3673 5645 3699
rect 6161 3671 6221 3697
rect 6279 3671 6339 3697
rect 6397 3671 6457 3697
rect 6515 3677 6575 3697
rect 6515 3671 6576 3677
rect 6633 3671 6693 3697
rect 6751 3671 6811 3697
rect 5346 3651 5412 3667
rect 5346 3617 5362 3651
rect 5396 3617 5412 3651
rect 5346 3601 5412 3617
rect 5228 3534 5294 3550
rect 5228 3500 5244 3534
rect 5278 3500 5294 3534
rect 5228 3484 5294 3500
rect 6398 3486 6456 3671
rect 5231 3462 5291 3484
rect 837 3234 897 3260
rect 2285 3234 2345 3260
rect 3783 3236 3843 3262
rect 6398 3460 6458 3486
rect 6516 3460 6576 3671
rect 6869 3665 6929 3697
rect 6987 3671 7047 3697
rect 7105 3671 7165 3697
rect 7609 3671 7669 3697
rect 7727 3671 7787 3697
rect 7845 3671 7905 3697
rect 7963 3677 8023 3697
rect 7963 3671 8024 3677
rect 8081 3671 8141 3697
rect 8199 3671 8259 3697
rect 6866 3649 6932 3665
rect 6866 3615 6882 3649
rect 6916 3615 6932 3649
rect 6866 3599 6932 3615
rect 6748 3532 6814 3548
rect 6748 3498 6764 3532
rect 6798 3498 6814 3532
rect 6748 3482 6814 3498
rect 7846 3486 7904 3671
rect 6751 3460 6811 3482
rect 7846 3460 7906 3486
rect 7964 3460 8024 3671
rect 8317 3665 8377 3697
rect 8435 3671 8495 3697
rect 8553 3671 8613 3697
rect 9107 3673 9167 3699
rect 9225 3673 9285 3699
rect 9343 3673 9403 3699
rect 9461 3679 9521 3699
rect 9461 3673 9522 3679
rect 9579 3673 9639 3699
rect 9697 3673 9757 3699
rect 8314 3649 8380 3665
rect 8314 3615 8330 3649
rect 8364 3615 8380 3649
rect 8314 3599 8380 3615
rect 8196 3532 8262 3548
rect 8196 3498 8212 3532
rect 8246 3498 8262 3532
rect 8196 3482 8262 3498
rect 9344 3488 9402 3673
rect 8199 3460 8259 3482
rect 9344 3462 9404 3488
rect 9462 3462 9522 3673
rect 9815 3667 9875 3699
rect 9933 3673 9993 3699
rect 10051 3673 10111 3699
rect 10555 3673 10615 3699
rect 10673 3673 10733 3699
rect 10791 3673 10851 3699
rect 10909 3679 10969 3699
rect 10909 3673 10970 3679
rect 11027 3673 11087 3699
rect 11145 3673 11205 3699
rect 9812 3651 9878 3667
rect 9812 3617 9828 3651
rect 9862 3617 9878 3651
rect 9812 3601 9878 3617
rect 9694 3534 9760 3550
rect 9694 3500 9710 3534
rect 9744 3500 9760 3534
rect 9694 3484 9760 3500
rect 10792 3488 10850 3673
rect 9697 3462 9757 3484
rect 10792 3462 10852 3488
rect 10910 3462 10970 3673
rect 11263 3667 11323 3699
rect 11381 3673 11441 3699
rect 11499 3673 11559 3699
rect 14346 4092 14406 4113
rect 14464 4092 14524 4114
rect 14582 4092 14642 4114
rect 14700 4114 14996 4155
rect 14700 4092 14760 4114
rect 14818 4092 14878 4114
rect 14936 4092 14996 4114
rect 15362 4146 15810 4155
rect 15362 4112 15378 4146
rect 15412 4114 15810 4146
rect 15412 4113 15574 4114
rect 15412 4112 15428 4113
rect 15362 4096 15428 4112
rect 15514 4094 15574 4113
rect 15632 4094 15692 4114
rect 15750 4094 15810 4114
rect 15868 4114 16164 4155
rect 15868 4094 15928 4114
rect 15986 4094 16046 4114
rect 16104 4094 16164 4114
rect 16536 4148 16984 4157
rect 16536 4114 16552 4148
rect 16586 4116 16984 4148
rect 16586 4115 16748 4116
rect 16586 4114 16602 4115
rect 16536 4098 16602 4114
rect 16688 4096 16748 4115
rect 16806 4096 16866 4116
rect 16924 4096 16984 4116
rect 17042 4116 17338 4157
rect 17042 4096 17102 4116
rect 17160 4096 17220 4116
rect 17278 4096 17338 4116
rect 17704 4148 18152 4157
rect 17704 4114 17720 4148
rect 17754 4116 18152 4148
rect 17754 4115 17916 4116
rect 17754 4114 17770 4115
rect 17704 4098 17770 4114
rect 12010 3676 12070 3694
rect 11260 3651 11326 3667
rect 11260 3617 11276 3651
rect 11310 3617 11326 3651
rect 11260 3601 11326 3617
rect 12010 3587 12071 3676
rect 12128 3668 12188 3694
rect 12246 3668 12306 3694
rect 11142 3534 11208 3550
rect 11142 3500 11158 3534
rect 11192 3500 11208 3534
rect 11142 3484 11208 3500
rect 11920 3534 12071 3587
rect 11145 3462 11205 3484
rect 5231 3236 5291 3262
rect 484 3038 544 3060
rect 602 3038 662 3060
rect 1932 3038 1992 3060
rect 2050 3038 2110 3060
rect 3430 3040 3490 3062
rect 3548 3040 3608 3062
rect 4878 3040 4938 3062
rect 4996 3040 5056 3062
rect 6751 3234 6811 3260
rect 8199 3234 8259 3260
rect 9697 3236 9757 3262
rect 11920 3308 11980 3534
rect 12364 3492 12424 3694
rect 12482 3668 12542 3694
rect 12600 3668 12660 3694
rect 13178 3676 13238 3694
rect 13178 3587 13239 3676
rect 13296 3668 13356 3694
rect 13414 3668 13474 3694
rect 12038 3441 12424 3492
rect 13088 3534 13239 3587
rect 12038 3308 12098 3441
rect 12153 3383 12219 3399
rect 12153 3349 12169 3383
rect 12203 3349 12219 3383
rect 12153 3333 12219 3349
rect 12156 3308 12216 3333
rect 11145 3236 11205 3262
rect 12440 3304 12500 3330
rect 12558 3304 12618 3330
rect 12676 3304 12736 3330
rect 13088 3310 13148 3534
rect 13532 3492 13592 3694
rect 13650 3668 13710 3694
rect 13768 3668 13828 3694
rect 17856 4094 17916 4115
rect 17974 4094 18034 4116
rect 18092 4094 18152 4116
rect 18210 4116 18506 4157
rect 18210 4094 18270 4116
rect 18328 4094 18388 4116
rect 18446 4094 18506 4116
rect 18872 4148 19320 4157
rect 18872 4114 18888 4148
rect 18922 4116 19320 4148
rect 18922 4115 19084 4116
rect 18922 4114 18938 4115
rect 18872 4098 18938 4114
rect 19024 4096 19084 4115
rect 19142 4096 19202 4116
rect 19260 4096 19320 4116
rect 19378 4116 19674 4157
rect 19378 4096 19438 4116
rect 19496 4096 19556 4116
rect 19614 4096 19674 4116
rect 20040 4148 20488 4157
rect 20040 4114 20056 4148
rect 20090 4116 20488 4148
rect 20090 4115 20252 4116
rect 20090 4114 20106 4115
rect 20040 4098 20106 4114
rect 14346 3676 14406 3692
rect 14346 3587 14407 3676
rect 14464 3666 14524 3692
rect 14582 3666 14642 3692
rect 13206 3441 13592 3492
rect 14256 3534 14407 3587
rect 13206 3310 13266 3441
rect 13321 3383 13387 3399
rect 13321 3349 13337 3383
rect 13371 3349 13387 3383
rect 13321 3333 13387 3349
rect 13324 3310 13384 3333
rect 13607 3310 13667 3336
rect 13725 3310 13785 3336
rect 13843 3310 13903 3336
rect 14256 3310 14316 3534
rect 14700 3492 14760 3692
rect 14818 3666 14878 3692
rect 14936 3666 14996 3692
rect 15514 3676 15574 3694
rect 15514 3587 15575 3676
rect 15632 3668 15692 3694
rect 15750 3668 15810 3694
rect 14374 3441 14760 3492
rect 15424 3534 15575 3587
rect 14374 3310 14434 3441
rect 14489 3383 14555 3399
rect 14489 3349 14505 3383
rect 14539 3349 14555 3383
rect 14489 3333 14555 3349
rect 14492 3310 14552 3333
rect 14775 3310 14835 3336
rect 14893 3310 14953 3336
rect 15011 3310 15071 3336
rect 15424 3310 15484 3534
rect 15868 3492 15928 3694
rect 15986 3668 16046 3694
rect 16104 3668 16164 3694
rect 16688 3678 16748 3696
rect 16688 3589 16749 3678
rect 16806 3670 16866 3696
rect 16924 3670 16984 3696
rect 15542 3441 15928 3492
rect 16598 3536 16749 3589
rect 15542 3310 15602 3441
rect 15657 3383 15723 3399
rect 15657 3349 15673 3383
rect 15707 3349 15723 3383
rect 15657 3333 15723 3349
rect 15660 3310 15720 3333
rect 15944 3310 16004 3336
rect 16062 3310 16122 3336
rect 16180 3310 16240 3336
rect 16598 3310 16658 3536
rect 17042 3494 17102 3696
rect 17160 3670 17220 3696
rect 17278 3670 17338 3696
rect 20192 4094 20252 4115
rect 20310 4094 20370 4116
rect 20428 4094 20488 4116
rect 20546 4116 20842 4157
rect 20546 4094 20606 4116
rect 20664 4094 20724 4116
rect 20782 4094 20842 4116
rect 17856 3678 17916 3694
rect 17856 3589 17917 3678
rect 17974 3668 18034 3694
rect 18092 3668 18152 3694
rect 16716 3443 17102 3494
rect 17766 3536 17917 3589
rect 16716 3310 16776 3443
rect 16831 3385 16897 3401
rect 16831 3351 16847 3385
rect 16881 3351 16897 3385
rect 16831 3335 16897 3351
rect 16834 3310 16894 3335
rect 11920 3082 11980 3108
rect 12038 3082 12098 3108
rect 12156 3078 12216 3108
rect 17116 3306 17176 3332
rect 17234 3306 17294 3332
rect 17352 3306 17412 3332
rect 17766 3310 17826 3536
rect 18210 3494 18270 3694
rect 18328 3668 18388 3694
rect 18446 3668 18506 3694
rect 19024 3678 19084 3696
rect 19024 3589 19085 3678
rect 19142 3670 19202 3696
rect 19260 3670 19320 3696
rect 17884 3443 18270 3494
rect 18934 3536 19085 3589
rect 17884 3310 17944 3443
rect 17999 3385 18065 3401
rect 17999 3351 18015 3385
rect 18049 3351 18065 3385
rect 17999 3335 18065 3351
rect 18002 3310 18062 3335
rect 12440 3078 12500 3104
rect 12558 3078 12618 3104
rect 12676 3078 12736 3104
rect 13088 3084 13148 3110
rect 13206 3084 13266 3110
rect 13324 3078 13384 3110
rect 13607 3078 13667 3110
rect 13725 3078 13785 3110
rect 13843 3078 13903 3110
rect 14256 3084 14316 3110
rect 14374 3084 14434 3110
rect 481 3022 547 3038
rect 481 2988 497 3022
rect 531 2988 547 3022
rect 481 2972 547 2988
rect 599 3022 665 3038
rect 599 2988 615 3022
rect 649 2988 665 3022
rect 599 2972 665 2988
rect 1929 3022 1995 3038
rect 1929 2988 1945 3022
rect 1979 2988 1995 3022
rect 1929 2972 1995 2988
rect 2047 3022 2113 3038
rect 2047 2988 2063 3022
rect 2097 2988 2113 3022
rect 2047 2972 2113 2988
rect 3427 3024 3493 3040
rect 3427 2990 3443 3024
rect 3477 2990 3493 3024
rect 3427 2974 3493 2990
rect 3545 3024 3611 3040
rect 3545 2990 3561 3024
rect 3595 2990 3611 3024
rect 3545 2974 3611 2990
rect 4875 3024 4941 3040
rect 4875 2990 4891 3024
rect 4925 2990 4941 3024
rect 4875 2974 4941 2990
rect 4993 3024 5059 3040
rect 6398 3038 6458 3060
rect 6516 3038 6576 3060
rect 7846 3038 7906 3060
rect 7964 3038 8024 3060
rect 9344 3040 9404 3062
rect 9462 3040 9522 3062
rect 10792 3040 10852 3062
rect 10910 3040 10970 3062
rect 4993 2990 5009 3024
rect 5043 2990 5059 3024
rect 4993 2974 5059 2990
rect 6395 3022 6461 3038
rect 6395 2988 6411 3022
rect 6445 2988 6461 3022
rect 6395 2972 6461 2988
rect 6513 3022 6579 3038
rect 6513 2988 6529 3022
rect 6563 2988 6579 3022
rect 6513 2972 6579 2988
rect 7843 3022 7909 3038
rect 7843 2988 7859 3022
rect 7893 2988 7909 3022
rect 7843 2972 7909 2988
rect 7961 3022 8027 3038
rect 7961 2988 7977 3022
rect 8011 2988 8027 3022
rect 7961 2972 8027 2988
rect 9341 3024 9407 3040
rect 9341 2990 9357 3024
rect 9391 2990 9407 3024
rect 9341 2974 9407 2990
rect 9459 3024 9525 3040
rect 9459 2990 9475 3024
rect 9509 2990 9525 3024
rect 9459 2974 9525 2990
rect 10789 3024 10855 3040
rect 10789 2990 10805 3024
rect 10839 2990 10855 3024
rect 10789 2974 10855 2990
rect 10907 3024 10973 3040
rect 12156 3037 12735 3078
rect 13324 3037 13903 3078
rect 14492 3078 14552 3110
rect 14775 3078 14835 3110
rect 14893 3078 14953 3110
rect 15011 3078 15071 3110
rect 15424 3084 15484 3110
rect 15542 3084 15602 3110
rect 14492 3037 15071 3078
rect 15660 3078 15720 3110
rect 15944 3078 16004 3110
rect 16062 3078 16122 3110
rect 16180 3084 16240 3110
rect 16598 3084 16658 3110
rect 16716 3084 16776 3110
rect 16180 3078 16239 3084
rect 15660 3037 16239 3078
rect 16834 3080 16894 3110
rect 18285 3305 18345 3331
rect 18403 3305 18463 3331
rect 18521 3305 18581 3331
rect 18934 3312 18994 3536
rect 19378 3494 19438 3696
rect 19496 3670 19556 3696
rect 19614 3670 19674 3696
rect 20192 3678 20252 3694
rect 20192 3589 20253 3678
rect 20310 3668 20370 3694
rect 20428 3668 20488 3694
rect 19052 3443 19438 3494
rect 20102 3536 20253 3589
rect 19052 3312 19112 3443
rect 19167 3385 19233 3401
rect 19167 3351 19183 3385
rect 19217 3351 19233 3385
rect 19167 3335 19233 3351
rect 19170 3312 19230 3335
rect 17116 3080 17176 3106
rect 17234 3080 17294 3106
rect 17352 3080 17412 3106
rect 17766 3084 17826 3110
rect 17884 3084 17944 3110
rect 16834 3074 17412 3080
rect 18002 3080 18062 3110
rect 19453 3305 19513 3331
rect 19571 3305 19631 3331
rect 19689 3305 19749 3331
rect 20102 3312 20162 3536
rect 20546 3494 20606 3694
rect 20664 3668 20724 3694
rect 20782 3668 20842 3694
rect 20220 3443 20606 3494
rect 20220 3312 20280 3443
rect 20335 3385 20401 3401
rect 20335 3351 20351 3385
rect 20385 3351 20401 3385
rect 20335 3335 20401 3351
rect 20338 3312 20398 3335
rect 18285 3080 18345 3105
rect 18403 3080 18463 3105
rect 18521 3080 18581 3105
rect 18934 3086 18994 3112
rect 19052 3086 19112 3112
rect 16834 3039 17413 3074
rect 18002 3039 18581 3080
rect 19170 3080 19230 3112
rect 20621 3306 20681 3332
rect 20739 3306 20799 3332
rect 20857 3306 20917 3332
rect 19453 3080 19513 3105
rect 19571 3080 19631 3105
rect 19689 3080 19749 3105
rect 20102 3086 20162 3112
rect 20220 3086 20280 3112
rect 19170 3039 19749 3080
rect 20338 3080 20398 3112
rect 20621 3080 20681 3106
rect 20739 3080 20799 3106
rect 20857 3080 20917 3106
rect 20338 3039 20917 3080
rect 10907 2990 10923 3024
rect 10957 2990 10973 3024
rect 10907 2974 10973 2990
rect 747 2155 1043 2194
rect 747 2140 807 2155
rect 865 2140 925 2155
rect 983 2140 1043 2155
rect 1214 2155 1510 2194
rect 1214 2140 1274 2155
rect 1332 2140 1392 2155
rect 1450 2140 1510 2155
rect 1568 2155 1864 2194
rect 1568 2140 1628 2155
rect 1686 2140 1746 2155
rect 1804 2140 1864 2155
rect 2041 2155 2337 2194
rect 2041 2140 2101 2155
rect 2159 2140 2219 2155
rect 2277 2140 2337 2155
rect 3891 2155 4187 2194
rect 3891 2140 3951 2155
rect 4009 2140 4069 2155
rect 4127 2140 4187 2155
rect 4358 2155 4654 2194
rect 4358 2140 4418 2155
rect 4476 2140 4536 2155
rect 4594 2140 4654 2155
rect 4712 2155 5008 2194
rect 4712 2140 4772 2155
rect 4830 2140 4890 2155
rect 4948 2140 5008 2155
rect 5185 2155 5481 2194
rect 5185 2140 5245 2155
rect 5303 2140 5363 2155
rect 5421 2140 5481 2155
rect 7023 2159 7319 2198
rect 7023 2144 7083 2159
rect 7141 2144 7201 2159
rect 7259 2144 7319 2159
rect 7490 2159 7786 2198
rect 7490 2144 7550 2159
rect 7608 2144 7668 2159
rect 7726 2144 7786 2159
rect 7844 2159 8140 2198
rect 7844 2144 7904 2159
rect 7962 2144 8022 2159
rect 8080 2144 8140 2159
rect 8317 2159 8613 2198
rect 8317 2144 8377 2159
rect 8435 2144 8495 2159
rect 8553 2144 8613 2159
rect 10167 2159 10463 2198
rect 10167 2144 10227 2159
rect 10285 2144 10345 2159
rect 10403 2144 10463 2159
rect 10634 2159 10930 2198
rect 10634 2144 10694 2159
rect 10752 2144 10812 2159
rect 10870 2144 10930 2159
rect 10988 2159 11284 2198
rect 10988 2144 11048 2159
rect 11106 2144 11166 2159
rect 11224 2144 11284 2159
rect 11461 2159 11757 2198
rect 11461 2144 11521 2159
rect 11579 2144 11639 2159
rect 11697 2144 11757 2159
rect 13369 2155 13665 2194
rect 306 1956 602 1995
rect 306 1940 366 1956
rect 424 1940 484 1956
rect 542 1940 602 1956
rect 2514 1956 2810 1995
rect 2514 1940 2574 1956
rect 2632 1940 2692 1956
rect 2750 1940 2810 1956
rect 3450 1956 3746 1995
rect 3450 1940 3510 1956
rect 3568 1940 3628 1956
rect 3686 1940 3746 1956
rect 5658 1956 5954 1995
rect 5658 1940 5718 1956
rect 5776 1940 5836 1956
rect 5894 1940 5954 1956
rect 6582 1960 6878 1999
rect 6582 1944 6642 1960
rect 6700 1944 6760 1960
rect 6818 1944 6878 1960
rect 8790 1960 9086 1999
rect 8790 1944 8850 1960
rect 8908 1944 8968 1960
rect 9026 1944 9086 1960
rect 9726 1960 10022 1999
rect 9726 1944 9786 1960
rect 9844 1944 9904 1960
rect 9962 1944 10022 1960
rect 13369 2140 13429 2155
rect 13487 2140 13547 2155
rect 13605 2140 13665 2155
rect 13836 2155 14132 2194
rect 13836 2140 13896 2155
rect 13954 2140 14014 2155
rect 14072 2140 14132 2155
rect 14190 2155 14486 2194
rect 14190 2140 14250 2155
rect 14308 2140 14368 2155
rect 14426 2140 14486 2155
rect 14663 2155 14959 2194
rect 14663 2140 14723 2155
rect 14781 2140 14841 2155
rect 14899 2140 14959 2155
rect 16513 2155 16809 2194
rect 16513 2140 16573 2155
rect 16631 2140 16691 2155
rect 16749 2140 16809 2155
rect 16980 2155 17276 2194
rect 16980 2140 17040 2155
rect 17098 2140 17158 2155
rect 17216 2140 17276 2155
rect 17334 2155 17630 2194
rect 17334 2140 17394 2155
rect 17452 2140 17512 2155
rect 17570 2140 17630 2155
rect 17807 2155 18103 2194
rect 17807 2140 17867 2155
rect 17925 2140 17985 2155
rect 18043 2140 18103 2155
rect 19645 2159 19941 2198
rect 19645 2144 19705 2159
rect 19763 2144 19823 2159
rect 19881 2144 19941 2159
rect 20112 2159 20408 2198
rect 20112 2144 20172 2159
rect 20230 2144 20290 2159
rect 20348 2144 20408 2159
rect 20466 2159 20762 2198
rect 20466 2144 20526 2159
rect 20584 2144 20644 2159
rect 20702 2144 20762 2159
rect 20939 2159 21235 2198
rect 20939 2144 20999 2159
rect 21057 2144 21117 2159
rect 21175 2144 21235 2159
rect 22789 2159 23085 2198
rect 22789 2144 22849 2159
rect 22907 2144 22967 2159
rect 23025 2144 23085 2159
rect 23256 2159 23552 2198
rect 23256 2144 23316 2159
rect 23374 2144 23434 2159
rect 23492 2144 23552 2159
rect 23610 2159 23906 2198
rect 23610 2144 23670 2159
rect 23728 2144 23788 2159
rect 23846 2144 23906 2159
rect 24083 2159 24379 2198
rect 24083 2144 24143 2159
rect 24201 2144 24261 2159
rect 24319 2144 24379 2159
rect 11934 1960 12230 1999
rect 11934 1944 11994 1960
rect 12052 1944 12112 1960
rect 12170 1944 12230 1960
rect 12928 1956 13224 1995
rect 12928 1940 12988 1956
rect 13046 1940 13106 1956
rect 13164 1940 13224 1956
rect 306 1454 366 1740
rect 424 1714 484 1740
rect 542 1714 602 1740
rect 747 1714 807 1740
rect 306 1437 442 1454
rect 306 1382 365 1437
rect 423 1382 442 1437
rect 306 1367 442 1382
rect 306 1055 366 1367
rect 865 1322 925 1740
rect 983 1714 1043 1740
rect 1214 1714 1274 1740
rect 1332 1714 1392 1740
rect 1450 1714 1510 1740
rect 1568 1714 1628 1740
rect 1333 1554 1392 1714
rect 1333 1553 1396 1554
rect 1330 1537 1396 1553
rect 1330 1503 1346 1537
rect 1380 1503 1396 1537
rect 1330 1487 1396 1503
rect 1433 1438 1528 1453
rect 1433 1383 1452 1438
rect 1510 1415 1528 1438
rect 1686 1415 1746 1740
rect 1804 1714 1864 1740
rect 2041 1714 2101 1740
rect 1510 1383 1746 1415
rect 1433 1366 1746 1383
rect 865 1265 1392 1322
rect 1332 1166 1392 1265
rect 1321 1153 1402 1166
rect 1321 1098 1334 1153
rect 1392 1098 1402 1153
rect 1321 1087 1402 1098
rect 306 1010 1200 1055
rect 1140 807 1200 1010
rect 1332 807 1392 1087
rect 1450 807 1510 1366
rect 2159 1324 2219 1740
rect 2277 1714 2337 1740
rect 2514 1714 2574 1740
rect 2632 1714 2692 1740
rect 2640 1591 2706 1594
rect 2750 1591 2810 1740
rect 2640 1578 2810 1591
rect 2640 1544 2656 1578
rect 2690 1544 2810 1578
rect 2640 1531 2810 1544
rect 2640 1528 2706 1531
rect 1681 1307 2219 1324
rect 1681 1273 1700 1307
rect 1734 1273 2219 1307
rect 1681 1267 2219 1273
rect 1681 1257 1750 1267
rect 1681 1255 1746 1257
rect 1565 917 1631 933
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1568 807 1628 867
rect 1686 807 1746 1255
rect 2750 1055 2810 1531
rect 1882 1010 2810 1055
rect 3450 1454 3510 1740
rect 3568 1714 3628 1740
rect 3686 1714 3746 1740
rect 3891 1714 3951 1740
rect 3450 1437 3586 1454
rect 3450 1382 3509 1437
rect 3567 1382 3586 1437
rect 3450 1367 3586 1382
rect 3450 1055 3510 1367
rect 4009 1322 4069 1740
rect 4127 1714 4187 1740
rect 4358 1714 4418 1740
rect 4476 1714 4536 1740
rect 4594 1714 4654 1740
rect 4712 1714 4772 1740
rect 4477 1554 4536 1714
rect 4477 1553 4540 1554
rect 4474 1537 4540 1553
rect 4474 1503 4490 1537
rect 4524 1503 4540 1537
rect 4474 1487 4540 1503
rect 4577 1438 4672 1453
rect 4577 1383 4596 1438
rect 4654 1415 4672 1438
rect 4830 1415 4890 1740
rect 4948 1714 5008 1740
rect 5185 1714 5245 1740
rect 4654 1383 4890 1415
rect 4577 1366 4890 1383
rect 4009 1265 4536 1322
rect 4476 1166 4536 1265
rect 4465 1153 4546 1166
rect 4465 1098 4478 1153
rect 4536 1098 4546 1153
rect 4465 1087 4546 1098
rect 3450 1010 4344 1055
rect 1882 807 1942 1010
rect 4284 807 4344 1010
rect 4476 807 4536 1087
rect 4594 807 4654 1366
rect 5303 1324 5363 1740
rect 5421 1714 5481 1740
rect 5658 1714 5718 1740
rect 5776 1714 5836 1740
rect 5784 1591 5850 1594
rect 5894 1591 5954 1740
rect 5784 1578 5954 1591
rect 5784 1544 5800 1578
rect 5834 1544 5954 1578
rect 5784 1531 5954 1544
rect 5784 1528 5850 1531
rect 4825 1307 5363 1324
rect 4825 1273 4844 1307
rect 4878 1273 5363 1307
rect 4825 1267 5363 1273
rect 4825 1257 4894 1267
rect 4825 1255 4890 1257
rect 4709 917 4775 933
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 4712 807 4772 867
rect 4830 807 4890 1255
rect 5894 1055 5954 1531
rect 5026 1010 5954 1055
rect 6582 1458 6642 1744
rect 6700 1718 6760 1744
rect 6818 1718 6878 1744
rect 7023 1718 7083 1744
rect 6582 1441 6718 1458
rect 6582 1386 6641 1441
rect 6699 1386 6718 1441
rect 6582 1371 6718 1386
rect 6582 1059 6642 1371
rect 7141 1326 7201 1744
rect 7259 1718 7319 1744
rect 7490 1718 7550 1744
rect 7608 1718 7668 1744
rect 7726 1718 7786 1744
rect 7844 1718 7904 1744
rect 7609 1558 7668 1718
rect 7609 1557 7672 1558
rect 7606 1541 7672 1557
rect 7606 1507 7622 1541
rect 7656 1507 7672 1541
rect 7606 1491 7672 1507
rect 7709 1442 7804 1457
rect 7709 1387 7728 1442
rect 7786 1419 7804 1442
rect 7962 1419 8022 1744
rect 8080 1718 8140 1744
rect 8317 1718 8377 1744
rect 7786 1387 8022 1419
rect 7709 1370 8022 1387
rect 7141 1269 7668 1326
rect 7608 1170 7668 1269
rect 7597 1157 7678 1170
rect 7597 1102 7610 1157
rect 7668 1102 7678 1157
rect 7597 1091 7678 1102
rect 6582 1014 7476 1059
rect 5026 807 5086 1010
rect 7416 811 7476 1014
rect 7608 811 7668 1091
rect 7726 811 7786 1370
rect 8435 1328 8495 1744
rect 8553 1718 8613 1744
rect 8790 1718 8850 1744
rect 8908 1718 8968 1744
rect 8916 1595 8982 1598
rect 9026 1595 9086 1744
rect 8916 1582 9086 1595
rect 8916 1548 8932 1582
rect 8966 1548 9086 1582
rect 8916 1535 9086 1548
rect 8916 1532 8982 1535
rect 7957 1311 8495 1328
rect 7957 1277 7976 1311
rect 8010 1277 8495 1311
rect 7957 1271 8495 1277
rect 7957 1261 8026 1271
rect 7957 1259 8022 1261
rect 7841 921 7907 937
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 7844 811 7904 871
rect 7962 811 8022 1259
rect 9026 1059 9086 1535
rect 8158 1014 9086 1059
rect 9726 1458 9786 1744
rect 9844 1718 9904 1744
rect 9962 1718 10022 1744
rect 10167 1718 10227 1744
rect 9726 1441 9862 1458
rect 9726 1386 9785 1441
rect 9843 1386 9862 1441
rect 9726 1371 9862 1386
rect 9726 1059 9786 1371
rect 10285 1326 10345 1744
rect 10403 1718 10463 1744
rect 10634 1718 10694 1744
rect 10752 1718 10812 1744
rect 10870 1718 10930 1744
rect 10988 1718 11048 1744
rect 10753 1558 10812 1718
rect 10753 1557 10816 1558
rect 10750 1541 10816 1557
rect 10750 1507 10766 1541
rect 10800 1507 10816 1541
rect 10750 1491 10816 1507
rect 10853 1442 10948 1457
rect 10853 1387 10872 1442
rect 10930 1419 10948 1442
rect 11106 1419 11166 1744
rect 11224 1718 11284 1744
rect 11461 1718 11521 1744
rect 10930 1387 11166 1419
rect 10853 1370 11166 1387
rect 10285 1269 10812 1326
rect 10752 1170 10812 1269
rect 10741 1157 10822 1170
rect 10741 1102 10754 1157
rect 10812 1102 10822 1157
rect 10741 1091 10822 1102
rect 9726 1014 10620 1059
rect 8158 811 8218 1014
rect 10560 811 10620 1014
rect 10752 811 10812 1091
rect 10870 811 10930 1370
rect 11579 1328 11639 1744
rect 11697 1718 11757 1744
rect 11934 1718 11994 1744
rect 12052 1718 12112 1744
rect 12060 1595 12126 1598
rect 12170 1595 12230 1744
rect 15136 1956 15432 1995
rect 15136 1940 15196 1956
rect 15254 1940 15314 1956
rect 15372 1940 15432 1956
rect 16072 1956 16368 1995
rect 16072 1940 16132 1956
rect 16190 1940 16250 1956
rect 16308 1940 16368 1956
rect 18280 1956 18576 1995
rect 18280 1940 18340 1956
rect 18398 1940 18458 1956
rect 18516 1940 18576 1956
rect 19204 1960 19500 1999
rect 19204 1944 19264 1960
rect 19322 1944 19382 1960
rect 19440 1944 19500 1960
rect 21412 1960 21708 1999
rect 21412 1944 21472 1960
rect 21530 1944 21590 1960
rect 21648 1944 21708 1960
rect 22348 1960 22644 1999
rect 22348 1944 22408 1960
rect 22466 1944 22526 1960
rect 22584 1944 22644 1960
rect 24556 1960 24852 1999
rect 24556 1944 24616 1960
rect 24674 1944 24734 1960
rect 24792 1944 24852 1960
rect 12060 1582 12230 1595
rect 12060 1548 12076 1582
rect 12110 1548 12230 1582
rect 12060 1535 12230 1548
rect 12060 1532 12126 1535
rect 11101 1311 11639 1328
rect 11101 1277 11120 1311
rect 11154 1277 11639 1311
rect 11101 1271 11639 1277
rect 11101 1261 11170 1271
rect 11101 1259 11166 1261
rect 10985 921 11051 937
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 10988 811 11048 871
rect 11106 811 11166 1259
rect 12170 1059 12230 1535
rect 11302 1014 12230 1059
rect 12928 1454 12988 1740
rect 13046 1714 13106 1740
rect 13164 1714 13224 1740
rect 13369 1714 13429 1740
rect 12928 1437 13064 1454
rect 12928 1382 12987 1437
rect 13045 1382 13064 1437
rect 12928 1367 13064 1382
rect 12928 1055 12988 1367
rect 13487 1322 13547 1740
rect 13605 1714 13665 1740
rect 13836 1714 13896 1740
rect 13954 1714 14014 1740
rect 14072 1714 14132 1740
rect 14190 1714 14250 1740
rect 13955 1554 14014 1714
rect 13955 1553 14018 1554
rect 13952 1537 14018 1553
rect 13952 1503 13968 1537
rect 14002 1503 14018 1537
rect 13952 1487 14018 1503
rect 14055 1438 14150 1453
rect 14055 1383 14074 1438
rect 14132 1415 14150 1438
rect 14308 1415 14368 1740
rect 14426 1714 14486 1740
rect 14663 1714 14723 1740
rect 14132 1383 14368 1415
rect 14055 1366 14368 1383
rect 13487 1265 14014 1322
rect 13954 1166 14014 1265
rect 13943 1153 14024 1166
rect 13943 1098 13956 1153
rect 14014 1098 14024 1153
rect 13943 1087 14024 1098
rect 11302 811 11362 1014
rect 12928 1010 13822 1055
rect 1140 581 1200 607
rect 1332 381 1392 407
rect 1450 381 1510 407
rect 1568 381 1628 407
rect 1686 381 1746 407
rect 1507 326 1573 334
rect 1882 326 1942 607
rect 4284 581 4344 607
rect 4476 381 4536 407
rect 4594 381 4654 407
rect 4712 381 4772 407
rect 4830 381 4890 407
rect 1507 318 1942 326
rect 1507 284 1523 318
rect 1557 284 1942 318
rect 1507 275 1942 284
rect 4651 326 4717 334
rect 5026 326 5086 607
rect 7416 585 7476 611
rect 7608 385 7668 411
rect 7726 385 7786 411
rect 7844 385 7904 411
rect 7962 385 8022 411
rect 4651 318 5086 326
rect 4651 284 4667 318
rect 4701 284 5086 318
rect 4651 275 5086 284
rect 7783 330 7849 338
rect 8158 330 8218 611
rect 10560 585 10620 611
rect 13762 807 13822 1010
rect 13954 807 14014 1087
rect 14072 807 14132 1366
rect 14781 1324 14841 1740
rect 14899 1714 14959 1740
rect 15136 1714 15196 1740
rect 15254 1714 15314 1740
rect 15262 1591 15328 1594
rect 15372 1591 15432 1740
rect 15262 1578 15432 1591
rect 15262 1544 15278 1578
rect 15312 1544 15432 1578
rect 15262 1531 15432 1544
rect 15262 1528 15328 1531
rect 14303 1307 14841 1324
rect 14303 1273 14322 1307
rect 14356 1273 14841 1307
rect 14303 1267 14841 1273
rect 14303 1257 14372 1267
rect 14303 1255 14368 1257
rect 14187 917 14253 933
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14190 807 14250 867
rect 14308 807 14368 1255
rect 15372 1055 15432 1531
rect 14504 1010 15432 1055
rect 16072 1454 16132 1740
rect 16190 1714 16250 1740
rect 16308 1714 16368 1740
rect 16513 1714 16573 1740
rect 16072 1437 16208 1454
rect 16072 1382 16131 1437
rect 16189 1382 16208 1437
rect 16072 1367 16208 1382
rect 16072 1055 16132 1367
rect 16631 1322 16691 1740
rect 16749 1714 16809 1740
rect 16980 1714 17040 1740
rect 17098 1714 17158 1740
rect 17216 1714 17276 1740
rect 17334 1714 17394 1740
rect 17099 1554 17158 1714
rect 17099 1553 17162 1554
rect 17096 1537 17162 1553
rect 17096 1503 17112 1537
rect 17146 1503 17162 1537
rect 17096 1487 17162 1503
rect 17199 1438 17294 1453
rect 17199 1383 17218 1438
rect 17276 1415 17294 1438
rect 17452 1415 17512 1740
rect 17570 1714 17630 1740
rect 17807 1714 17867 1740
rect 17276 1383 17512 1415
rect 17199 1366 17512 1383
rect 16631 1265 17158 1322
rect 17098 1166 17158 1265
rect 17087 1153 17168 1166
rect 17087 1098 17100 1153
rect 17158 1098 17168 1153
rect 17087 1087 17168 1098
rect 16072 1010 16966 1055
rect 14504 807 14564 1010
rect 16906 807 16966 1010
rect 17098 807 17158 1087
rect 17216 807 17276 1366
rect 17925 1324 17985 1740
rect 18043 1714 18103 1740
rect 18280 1714 18340 1740
rect 18398 1714 18458 1740
rect 18406 1591 18472 1594
rect 18516 1591 18576 1740
rect 18406 1578 18576 1591
rect 18406 1544 18422 1578
rect 18456 1544 18576 1578
rect 18406 1531 18576 1544
rect 18406 1528 18472 1531
rect 17447 1307 17985 1324
rect 17447 1273 17466 1307
rect 17500 1273 17985 1307
rect 17447 1267 17985 1273
rect 17447 1257 17516 1267
rect 17447 1255 17512 1257
rect 17331 917 17397 933
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17334 807 17394 867
rect 17452 807 17512 1255
rect 18516 1055 18576 1531
rect 17648 1010 18576 1055
rect 19204 1458 19264 1744
rect 19322 1718 19382 1744
rect 19440 1718 19500 1744
rect 19645 1718 19705 1744
rect 19204 1441 19340 1458
rect 19204 1386 19263 1441
rect 19321 1386 19340 1441
rect 19204 1371 19340 1386
rect 19204 1059 19264 1371
rect 19763 1326 19823 1744
rect 19881 1718 19941 1744
rect 20112 1718 20172 1744
rect 20230 1718 20290 1744
rect 20348 1718 20408 1744
rect 20466 1718 20526 1744
rect 20231 1558 20290 1718
rect 20231 1557 20294 1558
rect 20228 1541 20294 1557
rect 20228 1507 20244 1541
rect 20278 1507 20294 1541
rect 20228 1491 20294 1507
rect 20331 1442 20426 1457
rect 20331 1387 20350 1442
rect 20408 1419 20426 1442
rect 20584 1419 20644 1744
rect 20702 1718 20762 1744
rect 20939 1718 20999 1744
rect 20408 1387 20644 1419
rect 20331 1370 20644 1387
rect 19763 1269 20290 1326
rect 20230 1170 20290 1269
rect 20219 1157 20300 1170
rect 20219 1102 20232 1157
rect 20290 1102 20300 1157
rect 20219 1091 20300 1102
rect 19204 1014 20098 1059
rect 17648 807 17708 1010
rect 20038 811 20098 1014
rect 20230 811 20290 1091
rect 20348 811 20408 1370
rect 21057 1328 21117 1744
rect 21175 1718 21235 1744
rect 21412 1718 21472 1744
rect 21530 1718 21590 1744
rect 21538 1595 21604 1598
rect 21648 1595 21708 1744
rect 21538 1582 21708 1595
rect 21538 1548 21554 1582
rect 21588 1548 21708 1582
rect 21538 1535 21708 1548
rect 21538 1532 21604 1535
rect 20579 1311 21117 1328
rect 20579 1277 20598 1311
rect 20632 1277 21117 1311
rect 20579 1271 21117 1277
rect 20579 1261 20648 1271
rect 20579 1259 20644 1261
rect 20463 921 20529 937
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20466 811 20526 871
rect 20584 811 20644 1259
rect 21648 1059 21708 1535
rect 20780 1014 21708 1059
rect 22348 1458 22408 1744
rect 22466 1718 22526 1744
rect 22584 1718 22644 1744
rect 22789 1718 22849 1744
rect 22348 1441 22484 1458
rect 22348 1386 22407 1441
rect 22465 1386 22484 1441
rect 22348 1371 22484 1386
rect 22348 1059 22408 1371
rect 22907 1326 22967 1744
rect 23025 1718 23085 1744
rect 23256 1718 23316 1744
rect 23374 1718 23434 1744
rect 23492 1718 23552 1744
rect 23610 1718 23670 1744
rect 23375 1558 23434 1718
rect 23375 1557 23438 1558
rect 23372 1541 23438 1557
rect 23372 1507 23388 1541
rect 23422 1507 23438 1541
rect 23372 1491 23438 1507
rect 23475 1442 23570 1457
rect 23475 1387 23494 1442
rect 23552 1419 23570 1442
rect 23728 1419 23788 1744
rect 23846 1718 23906 1744
rect 24083 1718 24143 1744
rect 23552 1387 23788 1419
rect 23475 1370 23788 1387
rect 22907 1269 23434 1326
rect 23374 1170 23434 1269
rect 23363 1157 23444 1170
rect 23363 1102 23376 1157
rect 23434 1102 23444 1157
rect 23363 1091 23444 1102
rect 22348 1014 23242 1059
rect 20780 811 20840 1014
rect 23182 811 23242 1014
rect 23374 811 23434 1091
rect 23492 811 23552 1370
rect 24201 1328 24261 1744
rect 24319 1718 24379 1744
rect 24556 1718 24616 1744
rect 24674 1718 24734 1744
rect 24682 1595 24748 1598
rect 24792 1595 24852 1744
rect 24682 1582 24852 1595
rect 24682 1548 24698 1582
rect 24732 1548 24852 1582
rect 24682 1535 24852 1548
rect 24682 1532 24748 1535
rect 23723 1311 24261 1328
rect 23723 1277 23742 1311
rect 23776 1277 24261 1311
rect 23723 1271 24261 1277
rect 23723 1261 23792 1271
rect 23723 1259 23788 1261
rect 23607 921 23673 937
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23610 811 23670 871
rect 23728 811 23788 1259
rect 24792 1059 24852 1535
rect 23924 1014 24852 1059
rect 23924 811 23984 1014
rect 10752 385 10812 411
rect 10870 385 10930 411
rect 10988 385 11048 411
rect 11106 385 11166 411
rect 7783 322 8218 330
rect 7783 288 7799 322
rect 7833 288 8218 322
rect 7783 279 8218 288
rect 10927 330 10993 338
rect 11302 330 11362 611
rect 13762 581 13822 607
rect 13954 381 14014 407
rect 14072 381 14132 407
rect 14190 381 14250 407
rect 14308 381 14368 407
rect 10927 322 11362 330
rect 10927 288 10943 322
rect 10977 288 11362 322
rect 10927 279 11362 288
rect 14129 326 14195 334
rect 14504 326 14564 607
rect 16906 581 16966 607
rect 17098 381 17158 407
rect 17216 381 17276 407
rect 17334 381 17394 407
rect 17452 381 17512 407
rect 14129 318 14564 326
rect 14129 284 14145 318
rect 14179 284 14564 318
rect 1507 268 1573 275
rect 4651 268 4717 275
rect 7783 272 7849 279
rect 10927 272 10993 279
rect 14129 275 14564 284
rect 17273 326 17339 334
rect 17648 326 17708 607
rect 20038 585 20098 611
rect 20230 385 20290 411
rect 20348 385 20408 411
rect 20466 385 20526 411
rect 20584 385 20644 411
rect 17273 318 17708 326
rect 17273 284 17289 318
rect 17323 284 17708 318
rect 17273 275 17708 284
rect 20405 330 20471 338
rect 20780 330 20840 611
rect 23182 585 23242 611
rect 23374 385 23434 411
rect 23492 385 23552 411
rect 23610 385 23670 411
rect 23728 385 23788 411
rect 20405 322 20840 330
rect 20405 288 20421 322
rect 20455 288 20840 322
rect 20405 279 20840 288
rect 23549 330 23615 338
rect 23924 330 23984 611
rect 23549 322 23984 330
rect 23549 288 23565 322
rect 23599 288 23984 322
rect 23549 279 23984 288
rect 14129 268 14195 275
rect 17273 268 17339 275
rect 20405 272 20471 279
rect 23549 272 23615 279
rect 747 -579 1043 -540
rect 747 -594 807 -579
rect 865 -594 925 -579
rect 983 -594 1043 -579
rect 1214 -579 1510 -540
rect 1214 -594 1274 -579
rect 1332 -594 1392 -579
rect 1450 -594 1510 -579
rect 1568 -579 1864 -540
rect 1568 -594 1628 -579
rect 1686 -594 1746 -579
rect 1804 -594 1864 -579
rect 2041 -579 2337 -540
rect 2041 -594 2101 -579
rect 2159 -594 2219 -579
rect 2277 -594 2337 -579
rect 3891 -579 4187 -540
rect 3891 -594 3951 -579
rect 4009 -594 4069 -579
rect 4127 -594 4187 -579
rect 4358 -579 4654 -540
rect 4358 -594 4418 -579
rect 4476 -594 4536 -579
rect 4594 -594 4654 -579
rect 4712 -579 5008 -540
rect 4712 -594 4772 -579
rect 4830 -594 4890 -579
rect 4948 -594 5008 -579
rect 5185 -579 5481 -540
rect 5185 -594 5245 -579
rect 5303 -594 5363 -579
rect 5421 -594 5481 -579
rect 7023 -575 7319 -536
rect 7023 -590 7083 -575
rect 7141 -590 7201 -575
rect 7259 -590 7319 -575
rect 7490 -575 7786 -536
rect 7490 -590 7550 -575
rect 7608 -590 7668 -575
rect 7726 -590 7786 -575
rect 7844 -575 8140 -536
rect 7844 -590 7904 -575
rect 7962 -590 8022 -575
rect 8080 -590 8140 -575
rect 8317 -575 8613 -536
rect 8317 -590 8377 -575
rect 8435 -590 8495 -575
rect 8553 -590 8613 -575
rect 10167 -575 10463 -536
rect 10167 -590 10227 -575
rect 10285 -590 10345 -575
rect 10403 -590 10463 -575
rect 10634 -575 10930 -536
rect 10634 -590 10694 -575
rect 10752 -590 10812 -575
rect 10870 -590 10930 -575
rect 10988 -575 11284 -536
rect 10988 -590 11048 -575
rect 11106 -590 11166 -575
rect 11224 -590 11284 -575
rect 11461 -575 11757 -536
rect 11461 -590 11521 -575
rect 11579 -590 11639 -575
rect 11697 -590 11757 -575
rect 13369 -579 13665 -540
rect 306 -778 602 -739
rect 306 -794 366 -778
rect 424 -794 484 -778
rect 542 -794 602 -778
rect 2514 -778 2810 -739
rect 2514 -794 2574 -778
rect 2632 -794 2692 -778
rect 2750 -794 2810 -778
rect 3450 -778 3746 -739
rect 3450 -794 3510 -778
rect 3568 -794 3628 -778
rect 3686 -794 3746 -778
rect 5658 -778 5954 -739
rect 5658 -794 5718 -778
rect 5776 -794 5836 -778
rect 5894 -794 5954 -778
rect 6582 -774 6878 -735
rect 6582 -790 6642 -774
rect 6700 -790 6760 -774
rect 6818 -790 6878 -774
rect 8790 -774 9086 -735
rect 8790 -790 8850 -774
rect 8908 -790 8968 -774
rect 9026 -790 9086 -774
rect 9726 -774 10022 -735
rect 9726 -790 9786 -774
rect 9844 -790 9904 -774
rect 9962 -790 10022 -774
rect 13369 -594 13429 -579
rect 13487 -594 13547 -579
rect 13605 -594 13665 -579
rect 13836 -579 14132 -540
rect 13836 -594 13896 -579
rect 13954 -594 14014 -579
rect 14072 -594 14132 -579
rect 14190 -579 14486 -540
rect 14190 -594 14250 -579
rect 14308 -594 14368 -579
rect 14426 -594 14486 -579
rect 14663 -579 14959 -540
rect 14663 -594 14723 -579
rect 14781 -594 14841 -579
rect 14899 -594 14959 -579
rect 16513 -579 16809 -540
rect 16513 -594 16573 -579
rect 16631 -594 16691 -579
rect 16749 -594 16809 -579
rect 16980 -579 17276 -540
rect 16980 -594 17040 -579
rect 17098 -594 17158 -579
rect 17216 -594 17276 -579
rect 17334 -579 17630 -540
rect 17334 -594 17394 -579
rect 17452 -594 17512 -579
rect 17570 -594 17630 -579
rect 17807 -579 18103 -540
rect 17807 -594 17867 -579
rect 17925 -594 17985 -579
rect 18043 -594 18103 -579
rect 19645 -575 19941 -536
rect 19645 -590 19705 -575
rect 19763 -590 19823 -575
rect 19881 -590 19941 -575
rect 20112 -575 20408 -536
rect 20112 -590 20172 -575
rect 20230 -590 20290 -575
rect 20348 -590 20408 -575
rect 20466 -575 20762 -536
rect 20466 -590 20526 -575
rect 20584 -590 20644 -575
rect 20702 -590 20762 -575
rect 20939 -575 21235 -536
rect 20939 -590 20999 -575
rect 21057 -590 21117 -575
rect 21175 -590 21235 -575
rect 22789 -575 23085 -536
rect 22789 -590 22849 -575
rect 22907 -590 22967 -575
rect 23025 -590 23085 -575
rect 23256 -575 23552 -536
rect 23256 -590 23316 -575
rect 23374 -590 23434 -575
rect 23492 -590 23552 -575
rect 23610 -575 23906 -536
rect 23610 -590 23670 -575
rect 23728 -590 23788 -575
rect 23846 -590 23906 -575
rect 24083 -575 24379 -536
rect 24083 -590 24143 -575
rect 24201 -590 24261 -575
rect 24319 -590 24379 -575
rect 11934 -774 12230 -735
rect 11934 -790 11994 -774
rect 12052 -790 12112 -774
rect 12170 -790 12230 -774
rect 12928 -778 13224 -739
rect 12928 -794 12988 -778
rect 13046 -794 13106 -778
rect 13164 -794 13224 -778
rect 306 -1280 366 -994
rect 424 -1020 484 -994
rect 542 -1020 602 -994
rect 747 -1020 807 -994
rect 306 -1297 442 -1280
rect 306 -1352 365 -1297
rect 423 -1352 442 -1297
rect 306 -1367 442 -1352
rect 306 -1679 366 -1367
rect 865 -1412 925 -994
rect 983 -1020 1043 -994
rect 1214 -1020 1274 -994
rect 1332 -1020 1392 -994
rect 1450 -1020 1510 -994
rect 1568 -1020 1628 -994
rect 1333 -1180 1392 -1020
rect 1333 -1181 1396 -1180
rect 1330 -1197 1396 -1181
rect 1330 -1231 1346 -1197
rect 1380 -1231 1396 -1197
rect 1330 -1247 1396 -1231
rect 1433 -1296 1528 -1281
rect 1433 -1351 1452 -1296
rect 1510 -1319 1528 -1296
rect 1686 -1319 1746 -994
rect 1804 -1020 1864 -994
rect 2041 -1020 2101 -994
rect 1510 -1351 1746 -1319
rect 1433 -1368 1746 -1351
rect 865 -1469 1392 -1412
rect 1332 -1568 1392 -1469
rect 1321 -1581 1402 -1568
rect 1321 -1636 1334 -1581
rect 1392 -1636 1402 -1581
rect 1321 -1647 1402 -1636
rect 306 -1724 1200 -1679
rect 1140 -1927 1200 -1724
rect 1332 -1927 1392 -1647
rect 1450 -1927 1510 -1368
rect 2159 -1410 2219 -994
rect 2277 -1020 2337 -994
rect 2514 -1020 2574 -994
rect 2632 -1020 2692 -994
rect 2640 -1143 2706 -1140
rect 2750 -1143 2810 -994
rect 2640 -1156 2810 -1143
rect 2640 -1190 2656 -1156
rect 2690 -1190 2810 -1156
rect 2640 -1203 2810 -1190
rect 2640 -1206 2706 -1203
rect 1681 -1427 2219 -1410
rect 1681 -1461 1700 -1427
rect 1734 -1461 2219 -1427
rect 1681 -1467 2219 -1461
rect 1681 -1477 1750 -1467
rect 1681 -1479 1746 -1477
rect 1565 -1817 1631 -1801
rect 1565 -1851 1581 -1817
rect 1615 -1851 1631 -1817
rect 1565 -1867 1631 -1851
rect 1568 -1927 1628 -1867
rect 1686 -1927 1746 -1479
rect 2750 -1679 2810 -1203
rect 1882 -1724 2810 -1679
rect 3450 -1280 3510 -994
rect 3568 -1020 3628 -994
rect 3686 -1020 3746 -994
rect 3891 -1020 3951 -994
rect 3450 -1297 3586 -1280
rect 3450 -1352 3509 -1297
rect 3567 -1352 3586 -1297
rect 3450 -1367 3586 -1352
rect 3450 -1679 3510 -1367
rect 4009 -1412 4069 -994
rect 4127 -1020 4187 -994
rect 4358 -1020 4418 -994
rect 4476 -1020 4536 -994
rect 4594 -1020 4654 -994
rect 4712 -1020 4772 -994
rect 4477 -1180 4536 -1020
rect 4477 -1181 4540 -1180
rect 4474 -1197 4540 -1181
rect 4474 -1231 4490 -1197
rect 4524 -1231 4540 -1197
rect 4474 -1247 4540 -1231
rect 4577 -1296 4672 -1281
rect 4577 -1351 4596 -1296
rect 4654 -1319 4672 -1296
rect 4830 -1319 4890 -994
rect 4948 -1020 5008 -994
rect 5185 -1020 5245 -994
rect 4654 -1351 4890 -1319
rect 4577 -1368 4890 -1351
rect 4009 -1469 4536 -1412
rect 4476 -1568 4536 -1469
rect 4465 -1581 4546 -1568
rect 4465 -1636 4478 -1581
rect 4536 -1636 4546 -1581
rect 4465 -1647 4546 -1636
rect 3450 -1724 4344 -1679
rect 1882 -1927 1942 -1724
rect 4284 -1927 4344 -1724
rect 4476 -1927 4536 -1647
rect 4594 -1927 4654 -1368
rect 5303 -1410 5363 -994
rect 5421 -1020 5481 -994
rect 5658 -1020 5718 -994
rect 5776 -1020 5836 -994
rect 5784 -1143 5850 -1140
rect 5894 -1143 5954 -994
rect 5784 -1156 5954 -1143
rect 5784 -1190 5800 -1156
rect 5834 -1190 5954 -1156
rect 5784 -1203 5954 -1190
rect 5784 -1206 5850 -1203
rect 4825 -1427 5363 -1410
rect 4825 -1461 4844 -1427
rect 4878 -1461 5363 -1427
rect 4825 -1467 5363 -1461
rect 4825 -1477 4894 -1467
rect 4825 -1479 4890 -1477
rect 4709 -1817 4775 -1801
rect 4709 -1851 4725 -1817
rect 4759 -1851 4775 -1817
rect 4709 -1867 4775 -1851
rect 4712 -1927 4772 -1867
rect 4830 -1927 4890 -1479
rect 5894 -1679 5954 -1203
rect 5026 -1724 5954 -1679
rect 6582 -1276 6642 -990
rect 6700 -1016 6760 -990
rect 6818 -1016 6878 -990
rect 7023 -1016 7083 -990
rect 6582 -1293 6718 -1276
rect 6582 -1348 6641 -1293
rect 6699 -1348 6718 -1293
rect 6582 -1363 6718 -1348
rect 6582 -1675 6642 -1363
rect 7141 -1408 7201 -990
rect 7259 -1016 7319 -990
rect 7490 -1016 7550 -990
rect 7608 -1016 7668 -990
rect 7726 -1016 7786 -990
rect 7844 -1016 7904 -990
rect 7609 -1176 7668 -1016
rect 7609 -1177 7672 -1176
rect 7606 -1193 7672 -1177
rect 7606 -1227 7622 -1193
rect 7656 -1227 7672 -1193
rect 7606 -1243 7672 -1227
rect 7709 -1292 7804 -1277
rect 7709 -1347 7728 -1292
rect 7786 -1315 7804 -1292
rect 7962 -1315 8022 -990
rect 8080 -1016 8140 -990
rect 8317 -1016 8377 -990
rect 7786 -1347 8022 -1315
rect 7709 -1364 8022 -1347
rect 7141 -1465 7668 -1408
rect 7608 -1564 7668 -1465
rect 7597 -1577 7678 -1564
rect 7597 -1632 7610 -1577
rect 7668 -1632 7678 -1577
rect 7597 -1643 7678 -1632
rect 6582 -1720 7476 -1675
rect 5026 -1927 5086 -1724
rect 7416 -1923 7476 -1720
rect 7608 -1923 7668 -1643
rect 7726 -1923 7786 -1364
rect 8435 -1406 8495 -990
rect 8553 -1016 8613 -990
rect 8790 -1016 8850 -990
rect 8908 -1016 8968 -990
rect 8916 -1139 8982 -1136
rect 9026 -1139 9086 -990
rect 8916 -1152 9086 -1139
rect 8916 -1186 8932 -1152
rect 8966 -1186 9086 -1152
rect 8916 -1199 9086 -1186
rect 8916 -1202 8982 -1199
rect 7957 -1423 8495 -1406
rect 7957 -1457 7976 -1423
rect 8010 -1457 8495 -1423
rect 7957 -1463 8495 -1457
rect 7957 -1473 8026 -1463
rect 7957 -1475 8022 -1473
rect 7841 -1813 7907 -1797
rect 7841 -1847 7857 -1813
rect 7891 -1847 7907 -1813
rect 7841 -1863 7907 -1847
rect 7844 -1923 7904 -1863
rect 7962 -1923 8022 -1475
rect 9026 -1675 9086 -1199
rect 8158 -1720 9086 -1675
rect 9726 -1276 9786 -990
rect 9844 -1016 9904 -990
rect 9962 -1016 10022 -990
rect 10167 -1016 10227 -990
rect 9726 -1293 9862 -1276
rect 9726 -1348 9785 -1293
rect 9843 -1348 9862 -1293
rect 9726 -1363 9862 -1348
rect 9726 -1675 9786 -1363
rect 10285 -1408 10345 -990
rect 10403 -1016 10463 -990
rect 10634 -1016 10694 -990
rect 10752 -1016 10812 -990
rect 10870 -1016 10930 -990
rect 10988 -1016 11048 -990
rect 10753 -1176 10812 -1016
rect 10753 -1177 10816 -1176
rect 10750 -1193 10816 -1177
rect 10750 -1227 10766 -1193
rect 10800 -1227 10816 -1193
rect 10750 -1243 10816 -1227
rect 10853 -1292 10948 -1277
rect 10853 -1347 10872 -1292
rect 10930 -1315 10948 -1292
rect 11106 -1315 11166 -990
rect 11224 -1016 11284 -990
rect 11461 -1016 11521 -990
rect 10930 -1347 11166 -1315
rect 10853 -1364 11166 -1347
rect 10285 -1465 10812 -1408
rect 10752 -1564 10812 -1465
rect 10741 -1577 10822 -1564
rect 10741 -1632 10754 -1577
rect 10812 -1632 10822 -1577
rect 10741 -1643 10822 -1632
rect 9726 -1720 10620 -1675
rect 8158 -1923 8218 -1720
rect 10560 -1923 10620 -1720
rect 10752 -1923 10812 -1643
rect 10870 -1923 10930 -1364
rect 11579 -1406 11639 -990
rect 11697 -1016 11757 -990
rect 11934 -1016 11994 -990
rect 12052 -1016 12112 -990
rect 12060 -1139 12126 -1136
rect 12170 -1139 12230 -990
rect 15136 -778 15432 -739
rect 15136 -794 15196 -778
rect 15254 -794 15314 -778
rect 15372 -794 15432 -778
rect 16072 -778 16368 -739
rect 16072 -794 16132 -778
rect 16190 -794 16250 -778
rect 16308 -794 16368 -778
rect 18280 -778 18576 -739
rect 18280 -794 18340 -778
rect 18398 -794 18458 -778
rect 18516 -794 18576 -778
rect 19204 -774 19500 -735
rect 19204 -790 19264 -774
rect 19322 -790 19382 -774
rect 19440 -790 19500 -774
rect 21412 -774 21708 -735
rect 21412 -790 21472 -774
rect 21530 -790 21590 -774
rect 21648 -790 21708 -774
rect 22348 -774 22644 -735
rect 22348 -790 22408 -774
rect 22466 -790 22526 -774
rect 22584 -790 22644 -774
rect 24556 -774 24852 -735
rect 24556 -790 24616 -774
rect 24674 -790 24734 -774
rect 24792 -790 24852 -774
rect 12060 -1152 12230 -1139
rect 12060 -1186 12076 -1152
rect 12110 -1186 12230 -1152
rect 12060 -1199 12230 -1186
rect 12060 -1202 12126 -1199
rect 11101 -1423 11639 -1406
rect 11101 -1457 11120 -1423
rect 11154 -1457 11639 -1423
rect 11101 -1463 11639 -1457
rect 11101 -1473 11170 -1463
rect 11101 -1475 11166 -1473
rect 10985 -1813 11051 -1797
rect 10985 -1847 11001 -1813
rect 11035 -1847 11051 -1813
rect 10985 -1863 11051 -1847
rect 10988 -1923 11048 -1863
rect 11106 -1923 11166 -1475
rect 12170 -1675 12230 -1199
rect 11302 -1720 12230 -1675
rect 12928 -1280 12988 -994
rect 13046 -1020 13106 -994
rect 13164 -1020 13224 -994
rect 13369 -1020 13429 -994
rect 12928 -1297 13064 -1280
rect 12928 -1352 12987 -1297
rect 13045 -1352 13064 -1297
rect 12928 -1367 13064 -1352
rect 12928 -1679 12988 -1367
rect 13487 -1412 13547 -994
rect 13605 -1020 13665 -994
rect 13836 -1020 13896 -994
rect 13954 -1020 14014 -994
rect 14072 -1020 14132 -994
rect 14190 -1020 14250 -994
rect 13955 -1180 14014 -1020
rect 13955 -1181 14018 -1180
rect 13952 -1197 14018 -1181
rect 13952 -1231 13968 -1197
rect 14002 -1231 14018 -1197
rect 13952 -1247 14018 -1231
rect 14055 -1296 14150 -1281
rect 14055 -1351 14074 -1296
rect 14132 -1319 14150 -1296
rect 14308 -1319 14368 -994
rect 14426 -1020 14486 -994
rect 14663 -1020 14723 -994
rect 14132 -1351 14368 -1319
rect 14055 -1368 14368 -1351
rect 13487 -1469 14014 -1412
rect 13954 -1568 14014 -1469
rect 13943 -1581 14024 -1568
rect 13943 -1636 13956 -1581
rect 14014 -1636 14024 -1581
rect 13943 -1647 14024 -1636
rect 11302 -1923 11362 -1720
rect 12928 -1724 13822 -1679
rect 1140 -2153 1200 -2127
rect 1332 -2353 1392 -2327
rect 1450 -2353 1510 -2327
rect 1568 -2353 1628 -2327
rect 1686 -2353 1746 -2327
rect 1507 -2408 1573 -2400
rect 1882 -2408 1942 -2127
rect 4284 -2153 4344 -2127
rect 4476 -2353 4536 -2327
rect 4594 -2353 4654 -2327
rect 4712 -2353 4772 -2327
rect 4830 -2353 4890 -2327
rect 1507 -2416 1942 -2408
rect 1507 -2450 1523 -2416
rect 1557 -2450 1942 -2416
rect 1507 -2459 1942 -2450
rect 4651 -2408 4717 -2400
rect 5026 -2408 5086 -2127
rect 7416 -2149 7476 -2123
rect 7608 -2349 7668 -2323
rect 7726 -2349 7786 -2323
rect 7844 -2349 7904 -2323
rect 7962 -2349 8022 -2323
rect 4651 -2416 5086 -2408
rect 4651 -2450 4667 -2416
rect 4701 -2450 5086 -2416
rect 4651 -2459 5086 -2450
rect 7783 -2404 7849 -2396
rect 8158 -2404 8218 -2123
rect 10560 -2149 10620 -2123
rect 13762 -1927 13822 -1724
rect 13954 -1927 14014 -1647
rect 14072 -1927 14132 -1368
rect 14781 -1410 14841 -994
rect 14899 -1020 14959 -994
rect 15136 -1020 15196 -994
rect 15254 -1020 15314 -994
rect 15262 -1143 15328 -1140
rect 15372 -1143 15432 -994
rect 15262 -1156 15432 -1143
rect 15262 -1190 15278 -1156
rect 15312 -1190 15432 -1156
rect 15262 -1203 15432 -1190
rect 15262 -1206 15328 -1203
rect 14303 -1427 14841 -1410
rect 14303 -1461 14322 -1427
rect 14356 -1461 14841 -1427
rect 14303 -1467 14841 -1461
rect 14303 -1477 14372 -1467
rect 14303 -1479 14368 -1477
rect 14187 -1817 14253 -1801
rect 14187 -1851 14203 -1817
rect 14237 -1851 14253 -1817
rect 14187 -1867 14253 -1851
rect 14190 -1927 14250 -1867
rect 14308 -1927 14368 -1479
rect 15372 -1679 15432 -1203
rect 14504 -1724 15432 -1679
rect 16072 -1280 16132 -994
rect 16190 -1020 16250 -994
rect 16308 -1020 16368 -994
rect 16513 -1020 16573 -994
rect 16072 -1297 16208 -1280
rect 16072 -1352 16131 -1297
rect 16189 -1352 16208 -1297
rect 16072 -1367 16208 -1352
rect 16072 -1679 16132 -1367
rect 16631 -1412 16691 -994
rect 16749 -1020 16809 -994
rect 16980 -1020 17040 -994
rect 17098 -1020 17158 -994
rect 17216 -1020 17276 -994
rect 17334 -1020 17394 -994
rect 17099 -1180 17158 -1020
rect 17099 -1181 17162 -1180
rect 17096 -1197 17162 -1181
rect 17096 -1231 17112 -1197
rect 17146 -1231 17162 -1197
rect 17096 -1247 17162 -1231
rect 17199 -1296 17294 -1281
rect 17199 -1351 17218 -1296
rect 17276 -1319 17294 -1296
rect 17452 -1319 17512 -994
rect 17570 -1020 17630 -994
rect 17807 -1020 17867 -994
rect 17276 -1351 17512 -1319
rect 17199 -1368 17512 -1351
rect 16631 -1469 17158 -1412
rect 17098 -1568 17158 -1469
rect 17087 -1581 17168 -1568
rect 17087 -1636 17100 -1581
rect 17158 -1636 17168 -1581
rect 17087 -1647 17168 -1636
rect 16072 -1724 16966 -1679
rect 14504 -1927 14564 -1724
rect 16906 -1927 16966 -1724
rect 17098 -1927 17158 -1647
rect 17216 -1927 17276 -1368
rect 17925 -1410 17985 -994
rect 18043 -1020 18103 -994
rect 18280 -1020 18340 -994
rect 18398 -1020 18458 -994
rect 18406 -1143 18472 -1140
rect 18516 -1143 18576 -994
rect 18406 -1156 18576 -1143
rect 18406 -1190 18422 -1156
rect 18456 -1190 18576 -1156
rect 18406 -1203 18576 -1190
rect 18406 -1206 18472 -1203
rect 17447 -1427 17985 -1410
rect 17447 -1461 17466 -1427
rect 17500 -1461 17985 -1427
rect 17447 -1467 17985 -1461
rect 17447 -1477 17516 -1467
rect 17447 -1479 17512 -1477
rect 17331 -1817 17397 -1801
rect 17331 -1851 17347 -1817
rect 17381 -1851 17397 -1817
rect 17331 -1867 17397 -1851
rect 17334 -1927 17394 -1867
rect 17452 -1927 17512 -1479
rect 18516 -1679 18576 -1203
rect 17648 -1724 18576 -1679
rect 19204 -1276 19264 -990
rect 19322 -1016 19382 -990
rect 19440 -1016 19500 -990
rect 19645 -1016 19705 -990
rect 19204 -1293 19340 -1276
rect 19204 -1348 19263 -1293
rect 19321 -1348 19340 -1293
rect 19204 -1363 19340 -1348
rect 19204 -1675 19264 -1363
rect 19763 -1408 19823 -990
rect 19881 -1016 19941 -990
rect 20112 -1016 20172 -990
rect 20230 -1016 20290 -990
rect 20348 -1016 20408 -990
rect 20466 -1016 20526 -990
rect 20231 -1176 20290 -1016
rect 20231 -1177 20294 -1176
rect 20228 -1193 20294 -1177
rect 20228 -1227 20244 -1193
rect 20278 -1227 20294 -1193
rect 20228 -1243 20294 -1227
rect 20331 -1292 20426 -1277
rect 20331 -1347 20350 -1292
rect 20408 -1315 20426 -1292
rect 20584 -1315 20644 -990
rect 20702 -1016 20762 -990
rect 20939 -1016 20999 -990
rect 20408 -1347 20644 -1315
rect 20331 -1364 20644 -1347
rect 19763 -1465 20290 -1408
rect 20230 -1564 20290 -1465
rect 20219 -1577 20300 -1564
rect 20219 -1632 20232 -1577
rect 20290 -1632 20300 -1577
rect 20219 -1643 20300 -1632
rect 19204 -1720 20098 -1675
rect 17648 -1927 17708 -1724
rect 20038 -1923 20098 -1720
rect 20230 -1923 20290 -1643
rect 20348 -1923 20408 -1364
rect 21057 -1406 21117 -990
rect 21175 -1016 21235 -990
rect 21412 -1016 21472 -990
rect 21530 -1016 21590 -990
rect 21538 -1139 21604 -1136
rect 21648 -1139 21708 -990
rect 21538 -1152 21708 -1139
rect 21538 -1186 21554 -1152
rect 21588 -1186 21708 -1152
rect 21538 -1199 21708 -1186
rect 21538 -1202 21604 -1199
rect 20579 -1423 21117 -1406
rect 20579 -1457 20598 -1423
rect 20632 -1457 21117 -1423
rect 20579 -1463 21117 -1457
rect 20579 -1473 20648 -1463
rect 20579 -1475 20644 -1473
rect 20463 -1813 20529 -1797
rect 20463 -1847 20479 -1813
rect 20513 -1847 20529 -1813
rect 20463 -1863 20529 -1847
rect 20466 -1923 20526 -1863
rect 20584 -1923 20644 -1475
rect 21648 -1675 21708 -1199
rect 20780 -1720 21708 -1675
rect 22348 -1276 22408 -990
rect 22466 -1016 22526 -990
rect 22584 -1016 22644 -990
rect 22789 -1016 22849 -990
rect 22348 -1293 22484 -1276
rect 22348 -1348 22407 -1293
rect 22465 -1348 22484 -1293
rect 22348 -1363 22484 -1348
rect 22348 -1675 22408 -1363
rect 22907 -1408 22967 -990
rect 23025 -1016 23085 -990
rect 23256 -1016 23316 -990
rect 23374 -1016 23434 -990
rect 23492 -1016 23552 -990
rect 23610 -1016 23670 -990
rect 23375 -1176 23434 -1016
rect 23375 -1177 23438 -1176
rect 23372 -1193 23438 -1177
rect 23372 -1227 23388 -1193
rect 23422 -1227 23438 -1193
rect 23372 -1243 23438 -1227
rect 23475 -1292 23570 -1277
rect 23475 -1347 23494 -1292
rect 23552 -1315 23570 -1292
rect 23728 -1315 23788 -990
rect 23846 -1016 23906 -990
rect 24083 -1016 24143 -990
rect 23552 -1347 23788 -1315
rect 23475 -1364 23788 -1347
rect 22907 -1465 23434 -1408
rect 23374 -1564 23434 -1465
rect 23363 -1577 23444 -1564
rect 23363 -1632 23376 -1577
rect 23434 -1632 23444 -1577
rect 23363 -1643 23444 -1632
rect 22348 -1720 23242 -1675
rect 20780 -1923 20840 -1720
rect 23182 -1923 23242 -1720
rect 23374 -1923 23434 -1643
rect 23492 -1923 23552 -1364
rect 24201 -1406 24261 -990
rect 24319 -1016 24379 -990
rect 24556 -1016 24616 -990
rect 24674 -1016 24734 -990
rect 24682 -1139 24748 -1136
rect 24792 -1139 24852 -990
rect 24682 -1152 24852 -1139
rect 24682 -1186 24698 -1152
rect 24732 -1186 24852 -1152
rect 24682 -1199 24852 -1186
rect 24682 -1202 24748 -1199
rect 23723 -1423 24261 -1406
rect 23723 -1457 23742 -1423
rect 23776 -1457 24261 -1423
rect 23723 -1463 24261 -1457
rect 23723 -1473 23792 -1463
rect 23723 -1475 23788 -1473
rect 23607 -1813 23673 -1797
rect 23607 -1847 23623 -1813
rect 23657 -1847 23673 -1813
rect 23607 -1863 23673 -1847
rect 23610 -1923 23670 -1863
rect 23728 -1923 23788 -1475
rect 24792 -1675 24852 -1199
rect 23924 -1720 24852 -1675
rect 23924 -1923 23984 -1720
rect 10752 -2349 10812 -2323
rect 10870 -2349 10930 -2323
rect 10988 -2349 11048 -2323
rect 11106 -2349 11166 -2323
rect 7783 -2412 8218 -2404
rect 7783 -2446 7799 -2412
rect 7833 -2446 8218 -2412
rect 7783 -2455 8218 -2446
rect 10927 -2404 10993 -2396
rect 11302 -2404 11362 -2123
rect 13762 -2153 13822 -2127
rect 13954 -2353 14014 -2327
rect 14072 -2353 14132 -2327
rect 14190 -2353 14250 -2327
rect 14308 -2353 14368 -2327
rect 10927 -2412 11362 -2404
rect 10927 -2446 10943 -2412
rect 10977 -2446 11362 -2412
rect 10927 -2455 11362 -2446
rect 14129 -2408 14195 -2400
rect 14504 -2408 14564 -2127
rect 16906 -2153 16966 -2127
rect 17098 -2353 17158 -2327
rect 17216 -2353 17276 -2327
rect 17334 -2353 17394 -2327
rect 17452 -2353 17512 -2327
rect 14129 -2416 14564 -2408
rect 14129 -2450 14145 -2416
rect 14179 -2450 14564 -2416
rect 1507 -2466 1573 -2459
rect 4651 -2466 4717 -2459
rect 7783 -2462 7849 -2455
rect 10927 -2462 10993 -2455
rect 14129 -2459 14564 -2450
rect 17273 -2408 17339 -2400
rect 17648 -2408 17708 -2127
rect 20038 -2149 20098 -2123
rect 20230 -2349 20290 -2323
rect 20348 -2349 20408 -2323
rect 20466 -2349 20526 -2323
rect 20584 -2349 20644 -2323
rect 17273 -2416 17708 -2408
rect 17273 -2450 17289 -2416
rect 17323 -2450 17708 -2416
rect 17273 -2459 17708 -2450
rect 20405 -2404 20471 -2396
rect 20780 -2404 20840 -2123
rect 23182 -2149 23242 -2123
rect 23374 -2349 23434 -2323
rect 23492 -2349 23552 -2323
rect 23610 -2349 23670 -2323
rect 23728 -2349 23788 -2323
rect 20405 -2412 20840 -2404
rect 20405 -2446 20421 -2412
rect 20455 -2446 20840 -2412
rect 20405 -2455 20840 -2446
rect 23549 -2404 23615 -2396
rect 23924 -2404 23984 -2123
rect 23549 -2412 23984 -2404
rect 23549 -2446 23565 -2412
rect 23599 -2446 23984 -2412
rect 23549 -2455 23984 -2446
rect 14129 -2466 14195 -2459
rect 17273 -2466 17339 -2459
rect 20405 -2462 20471 -2455
rect 23549 -2462 23615 -2455
rect 737 -3311 1033 -3272
rect 737 -3326 797 -3311
rect 855 -3326 915 -3311
rect 973 -3326 1033 -3311
rect 1204 -3311 1500 -3272
rect 1204 -3326 1264 -3311
rect 1322 -3326 1382 -3311
rect 1440 -3326 1500 -3311
rect 1558 -3311 1854 -3272
rect 1558 -3326 1618 -3311
rect 1676 -3326 1736 -3311
rect 1794 -3326 1854 -3311
rect 2031 -3311 2327 -3272
rect 2031 -3326 2091 -3311
rect 2149 -3326 2209 -3311
rect 2267 -3326 2327 -3311
rect 3881 -3311 4177 -3272
rect 3881 -3326 3941 -3311
rect 3999 -3326 4059 -3311
rect 4117 -3326 4177 -3311
rect 4348 -3311 4644 -3272
rect 4348 -3326 4408 -3311
rect 4466 -3326 4526 -3311
rect 4584 -3326 4644 -3311
rect 4702 -3311 4998 -3272
rect 4702 -3326 4762 -3311
rect 4820 -3326 4880 -3311
rect 4938 -3326 4998 -3311
rect 5175 -3311 5471 -3272
rect 5175 -3326 5235 -3311
rect 5293 -3326 5353 -3311
rect 5411 -3326 5471 -3311
rect 7013 -3307 7309 -3268
rect 7013 -3322 7073 -3307
rect 7131 -3322 7191 -3307
rect 7249 -3322 7309 -3307
rect 7480 -3307 7776 -3268
rect 7480 -3322 7540 -3307
rect 7598 -3322 7658 -3307
rect 7716 -3322 7776 -3307
rect 7834 -3307 8130 -3268
rect 7834 -3322 7894 -3307
rect 7952 -3322 8012 -3307
rect 8070 -3322 8130 -3307
rect 8307 -3307 8603 -3268
rect 8307 -3322 8367 -3307
rect 8425 -3322 8485 -3307
rect 8543 -3322 8603 -3307
rect 10157 -3307 10453 -3268
rect 10157 -3322 10217 -3307
rect 10275 -3322 10335 -3307
rect 10393 -3322 10453 -3307
rect 10624 -3307 10920 -3268
rect 10624 -3322 10684 -3307
rect 10742 -3322 10802 -3307
rect 10860 -3322 10920 -3307
rect 10978 -3307 11274 -3268
rect 10978 -3322 11038 -3307
rect 11096 -3322 11156 -3307
rect 11214 -3322 11274 -3307
rect 11451 -3307 11747 -3268
rect 11451 -3322 11511 -3307
rect 11569 -3322 11629 -3307
rect 11687 -3322 11747 -3307
rect 13359 -3311 13655 -3272
rect 296 -3510 592 -3471
rect 296 -3526 356 -3510
rect 414 -3526 474 -3510
rect 532 -3526 592 -3510
rect 2504 -3510 2800 -3471
rect 2504 -3526 2564 -3510
rect 2622 -3526 2682 -3510
rect 2740 -3526 2800 -3510
rect 3440 -3510 3736 -3471
rect 3440 -3526 3500 -3510
rect 3558 -3526 3618 -3510
rect 3676 -3526 3736 -3510
rect 5648 -3510 5944 -3471
rect 5648 -3526 5708 -3510
rect 5766 -3526 5826 -3510
rect 5884 -3526 5944 -3510
rect 6572 -3506 6868 -3467
rect 6572 -3522 6632 -3506
rect 6690 -3522 6750 -3506
rect 6808 -3522 6868 -3506
rect 8780 -3506 9076 -3467
rect 8780 -3522 8840 -3506
rect 8898 -3522 8958 -3506
rect 9016 -3522 9076 -3506
rect 9716 -3506 10012 -3467
rect 9716 -3522 9776 -3506
rect 9834 -3522 9894 -3506
rect 9952 -3522 10012 -3506
rect 13359 -3326 13419 -3311
rect 13477 -3326 13537 -3311
rect 13595 -3326 13655 -3311
rect 13826 -3311 14122 -3272
rect 13826 -3326 13886 -3311
rect 13944 -3326 14004 -3311
rect 14062 -3326 14122 -3311
rect 14180 -3311 14476 -3272
rect 14180 -3326 14240 -3311
rect 14298 -3326 14358 -3311
rect 14416 -3326 14476 -3311
rect 14653 -3311 14949 -3272
rect 14653 -3326 14713 -3311
rect 14771 -3326 14831 -3311
rect 14889 -3326 14949 -3311
rect 16503 -3311 16799 -3272
rect 16503 -3326 16563 -3311
rect 16621 -3326 16681 -3311
rect 16739 -3326 16799 -3311
rect 16970 -3311 17266 -3272
rect 16970 -3326 17030 -3311
rect 17088 -3326 17148 -3311
rect 17206 -3326 17266 -3311
rect 17324 -3311 17620 -3272
rect 17324 -3326 17384 -3311
rect 17442 -3326 17502 -3311
rect 17560 -3326 17620 -3311
rect 17797 -3311 18093 -3272
rect 17797 -3326 17857 -3311
rect 17915 -3326 17975 -3311
rect 18033 -3326 18093 -3311
rect 19635 -3307 19931 -3268
rect 19635 -3322 19695 -3307
rect 19753 -3322 19813 -3307
rect 19871 -3322 19931 -3307
rect 20102 -3307 20398 -3268
rect 20102 -3322 20162 -3307
rect 20220 -3322 20280 -3307
rect 20338 -3322 20398 -3307
rect 20456 -3307 20752 -3268
rect 20456 -3322 20516 -3307
rect 20574 -3322 20634 -3307
rect 20692 -3322 20752 -3307
rect 20929 -3307 21225 -3268
rect 20929 -3322 20989 -3307
rect 21047 -3322 21107 -3307
rect 21165 -3322 21225 -3307
rect 22779 -3307 23075 -3268
rect 22779 -3322 22839 -3307
rect 22897 -3322 22957 -3307
rect 23015 -3322 23075 -3307
rect 23246 -3307 23542 -3268
rect 23246 -3322 23306 -3307
rect 23364 -3322 23424 -3307
rect 23482 -3322 23542 -3307
rect 23600 -3307 23896 -3268
rect 23600 -3322 23660 -3307
rect 23718 -3322 23778 -3307
rect 23836 -3322 23896 -3307
rect 24073 -3307 24369 -3268
rect 24073 -3322 24133 -3307
rect 24191 -3322 24251 -3307
rect 24309 -3322 24369 -3307
rect 11924 -3506 12220 -3467
rect 11924 -3522 11984 -3506
rect 12042 -3522 12102 -3506
rect 12160 -3522 12220 -3506
rect 12918 -3510 13214 -3471
rect 12918 -3526 12978 -3510
rect 13036 -3526 13096 -3510
rect 13154 -3526 13214 -3510
rect 296 -4012 356 -3726
rect 414 -3752 474 -3726
rect 532 -3752 592 -3726
rect 737 -3752 797 -3726
rect 296 -4029 432 -4012
rect 296 -4084 355 -4029
rect 413 -4084 432 -4029
rect 296 -4099 432 -4084
rect 296 -4411 356 -4099
rect 855 -4144 915 -3726
rect 973 -3752 1033 -3726
rect 1204 -3752 1264 -3726
rect 1322 -3752 1382 -3726
rect 1440 -3752 1500 -3726
rect 1558 -3752 1618 -3726
rect 1323 -3912 1382 -3752
rect 1323 -3913 1386 -3912
rect 1320 -3929 1386 -3913
rect 1320 -3963 1336 -3929
rect 1370 -3963 1386 -3929
rect 1320 -3979 1386 -3963
rect 1423 -4028 1518 -4013
rect 1423 -4083 1442 -4028
rect 1500 -4051 1518 -4028
rect 1676 -4051 1736 -3726
rect 1794 -3752 1854 -3726
rect 2031 -3752 2091 -3726
rect 1500 -4083 1736 -4051
rect 1423 -4100 1736 -4083
rect 855 -4201 1382 -4144
rect 1322 -4300 1382 -4201
rect 1311 -4313 1392 -4300
rect 1311 -4368 1324 -4313
rect 1382 -4368 1392 -4313
rect 1311 -4379 1392 -4368
rect 296 -4456 1190 -4411
rect 1130 -4659 1190 -4456
rect 1322 -4659 1382 -4379
rect 1440 -4659 1500 -4100
rect 2149 -4142 2209 -3726
rect 2267 -3752 2327 -3726
rect 2504 -3752 2564 -3726
rect 2622 -3752 2682 -3726
rect 2630 -3875 2696 -3872
rect 2740 -3875 2800 -3726
rect 2630 -3888 2800 -3875
rect 2630 -3922 2646 -3888
rect 2680 -3922 2800 -3888
rect 2630 -3935 2800 -3922
rect 2630 -3938 2696 -3935
rect 1671 -4159 2209 -4142
rect 1671 -4193 1690 -4159
rect 1724 -4193 2209 -4159
rect 1671 -4199 2209 -4193
rect 1671 -4209 1740 -4199
rect 1671 -4211 1736 -4209
rect 1555 -4549 1621 -4533
rect 1555 -4583 1571 -4549
rect 1605 -4583 1621 -4549
rect 1555 -4599 1621 -4583
rect 1558 -4659 1618 -4599
rect 1676 -4659 1736 -4211
rect 2740 -4411 2800 -3935
rect 1872 -4456 2800 -4411
rect 3440 -4012 3500 -3726
rect 3558 -3752 3618 -3726
rect 3676 -3752 3736 -3726
rect 3881 -3752 3941 -3726
rect 3440 -4029 3576 -4012
rect 3440 -4084 3499 -4029
rect 3557 -4084 3576 -4029
rect 3440 -4099 3576 -4084
rect 3440 -4411 3500 -4099
rect 3999 -4144 4059 -3726
rect 4117 -3752 4177 -3726
rect 4348 -3752 4408 -3726
rect 4466 -3752 4526 -3726
rect 4584 -3752 4644 -3726
rect 4702 -3752 4762 -3726
rect 4467 -3912 4526 -3752
rect 4467 -3913 4530 -3912
rect 4464 -3929 4530 -3913
rect 4464 -3963 4480 -3929
rect 4514 -3963 4530 -3929
rect 4464 -3979 4530 -3963
rect 4567 -4028 4662 -4013
rect 4567 -4083 4586 -4028
rect 4644 -4051 4662 -4028
rect 4820 -4051 4880 -3726
rect 4938 -3752 4998 -3726
rect 5175 -3752 5235 -3726
rect 4644 -4083 4880 -4051
rect 4567 -4100 4880 -4083
rect 3999 -4201 4526 -4144
rect 4466 -4300 4526 -4201
rect 4455 -4313 4536 -4300
rect 4455 -4368 4468 -4313
rect 4526 -4368 4536 -4313
rect 4455 -4379 4536 -4368
rect 3440 -4456 4334 -4411
rect 1872 -4659 1932 -4456
rect 4274 -4659 4334 -4456
rect 4466 -4659 4526 -4379
rect 4584 -4659 4644 -4100
rect 5293 -4142 5353 -3726
rect 5411 -3752 5471 -3726
rect 5648 -3752 5708 -3726
rect 5766 -3752 5826 -3726
rect 5774 -3875 5840 -3872
rect 5884 -3875 5944 -3726
rect 5774 -3888 5944 -3875
rect 5774 -3922 5790 -3888
rect 5824 -3922 5944 -3888
rect 5774 -3935 5944 -3922
rect 5774 -3938 5840 -3935
rect 4815 -4159 5353 -4142
rect 4815 -4193 4834 -4159
rect 4868 -4193 5353 -4159
rect 4815 -4199 5353 -4193
rect 4815 -4209 4884 -4199
rect 4815 -4211 4880 -4209
rect 4699 -4549 4765 -4533
rect 4699 -4583 4715 -4549
rect 4749 -4583 4765 -4549
rect 4699 -4599 4765 -4583
rect 4702 -4659 4762 -4599
rect 4820 -4659 4880 -4211
rect 5884 -4411 5944 -3935
rect 5016 -4456 5944 -4411
rect 6572 -4008 6632 -3722
rect 6690 -3748 6750 -3722
rect 6808 -3748 6868 -3722
rect 7013 -3748 7073 -3722
rect 6572 -4025 6708 -4008
rect 6572 -4080 6631 -4025
rect 6689 -4080 6708 -4025
rect 6572 -4095 6708 -4080
rect 6572 -4407 6632 -4095
rect 7131 -4140 7191 -3722
rect 7249 -3748 7309 -3722
rect 7480 -3748 7540 -3722
rect 7598 -3748 7658 -3722
rect 7716 -3748 7776 -3722
rect 7834 -3748 7894 -3722
rect 7599 -3908 7658 -3748
rect 7599 -3909 7662 -3908
rect 7596 -3925 7662 -3909
rect 7596 -3959 7612 -3925
rect 7646 -3959 7662 -3925
rect 7596 -3975 7662 -3959
rect 7699 -4024 7794 -4009
rect 7699 -4079 7718 -4024
rect 7776 -4047 7794 -4024
rect 7952 -4047 8012 -3722
rect 8070 -3748 8130 -3722
rect 8307 -3748 8367 -3722
rect 7776 -4079 8012 -4047
rect 7699 -4096 8012 -4079
rect 7131 -4197 7658 -4140
rect 7598 -4296 7658 -4197
rect 7587 -4309 7668 -4296
rect 7587 -4364 7600 -4309
rect 7658 -4364 7668 -4309
rect 7587 -4375 7668 -4364
rect 6572 -4452 7466 -4407
rect 5016 -4659 5076 -4456
rect 7406 -4655 7466 -4452
rect 7598 -4655 7658 -4375
rect 7716 -4655 7776 -4096
rect 8425 -4138 8485 -3722
rect 8543 -3748 8603 -3722
rect 8780 -3748 8840 -3722
rect 8898 -3748 8958 -3722
rect 8906 -3871 8972 -3868
rect 9016 -3871 9076 -3722
rect 8906 -3884 9076 -3871
rect 8906 -3918 8922 -3884
rect 8956 -3918 9076 -3884
rect 8906 -3931 9076 -3918
rect 8906 -3934 8972 -3931
rect 7947 -4155 8485 -4138
rect 7947 -4189 7966 -4155
rect 8000 -4189 8485 -4155
rect 7947 -4195 8485 -4189
rect 7947 -4205 8016 -4195
rect 7947 -4207 8012 -4205
rect 7831 -4545 7897 -4529
rect 7831 -4579 7847 -4545
rect 7881 -4579 7897 -4545
rect 7831 -4595 7897 -4579
rect 7834 -4655 7894 -4595
rect 7952 -4655 8012 -4207
rect 9016 -4407 9076 -3931
rect 8148 -4452 9076 -4407
rect 9716 -4008 9776 -3722
rect 9834 -3748 9894 -3722
rect 9952 -3748 10012 -3722
rect 10157 -3748 10217 -3722
rect 9716 -4025 9852 -4008
rect 9716 -4080 9775 -4025
rect 9833 -4080 9852 -4025
rect 9716 -4095 9852 -4080
rect 9716 -4407 9776 -4095
rect 10275 -4140 10335 -3722
rect 10393 -3748 10453 -3722
rect 10624 -3748 10684 -3722
rect 10742 -3748 10802 -3722
rect 10860 -3748 10920 -3722
rect 10978 -3748 11038 -3722
rect 10743 -3908 10802 -3748
rect 10743 -3909 10806 -3908
rect 10740 -3925 10806 -3909
rect 10740 -3959 10756 -3925
rect 10790 -3959 10806 -3925
rect 10740 -3975 10806 -3959
rect 10843 -4024 10938 -4009
rect 10843 -4079 10862 -4024
rect 10920 -4047 10938 -4024
rect 11096 -4047 11156 -3722
rect 11214 -3748 11274 -3722
rect 11451 -3748 11511 -3722
rect 10920 -4079 11156 -4047
rect 10843 -4096 11156 -4079
rect 10275 -4197 10802 -4140
rect 10742 -4296 10802 -4197
rect 10731 -4309 10812 -4296
rect 10731 -4364 10744 -4309
rect 10802 -4364 10812 -4309
rect 10731 -4375 10812 -4364
rect 9716 -4452 10610 -4407
rect 8148 -4655 8208 -4452
rect 10550 -4655 10610 -4452
rect 10742 -4655 10802 -4375
rect 10860 -4655 10920 -4096
rect 11569 -4138 11629 -3722
rect 11687 -3748 11747 -3722
rect 11924 -3748 11984 -3722
rect 12042 -3748 12102 -3722
rect 12050 -3871 12116 -3868
rect 12160 -3871 12220 -3722
rect 15126 -3510 15422 -3471
rect 15126 -3526 15186 -3510
rect 15244 -3526 15304 -3510
rect 15362 -3526 15422 -3510
rect 16062 -3510 16358 -3471
rect 16062 -3526 16122 -3510
rect 16180 -3526 16240 -3510
rect 16298 -3526 16358 -3510
rect 18270 -3510 18566 -3471
rect 18270 -3526 18330 -3510
rect 18388 -3526 18448 -3510
rect 18506 -3526 18566 -3510
rect 19194 -3506 19490 -3467
rect 19194 -3522 19254 -3506
rect 19312 -3522 19372 -3506
rect 19430 -3522 19490 -3506
rect 21402 -3506 21698 -3467
rect 21402 -3522 21462 -3506
rect 21520 -3522 21580 -3506
rect 21638 -3522 21698 -3506
rect 22338 -3506 22634 -3467
rect 22338 -3522 22398 -3506
rect 22456 -3522 22516 -3506
rect 22574 -3522 22634 -3506
rect 24546 -3506 24842 -3467
rect 24546 -3522 24606 -3506
rect 24664 -3522 24724 -3506
rect 24782 -3522 24842 -3506
rect 12050 -3884 12220 -3871
rect 12050 -3918 12066 -3884
rect 12100 -3918 12220 -3884
rect 12050 -3931 12220 -3918
rect 12050 -3934 12116 -3931
rect 11091 -4155 11629 -4138
rect 11091 -4189 11110 -4155
rect 11144 -4189 11629 -4155
rect 11091 -4195 11629 -4189
rect 11091 -4205 11160 -4195
rect 11091 -4207 11156 -4205
rect 10975 -4545 11041 -4529
rect 10975 -4579 10991 -4545
rect 11025 -4579 11041 -4545
rect 10975 -4595 11041 -4579
rect 10978 -4655 11038 -4595
rect 11096 -4655 11156 -4207
rect 12160 -4407 12220 -3931
rect 11292 -4452 12220 -4407
rect 12918 -4012 12978 -3726
rect 13036 -3752 13096 -3726
rect 13154 -3752 13214 -3726
rect 13359 -3752 13419 -3726
rect 12918 -4029 13054 -4012
rect 12918 -4084 12977 -4029
rect 13035 -4084 13054 -4029
rect 12918 -4099 13054 -4084
rect 12918 -4411 12978 -4099
rect 13477 -4144 13537 -3726
rect 13595 -3752 13655 -3726
rect 13826 -3752 13886 -3726
rect 13944 -3752 14004 -3726
rect 14062 -3752 14122 -3726
rect 14180 -3752 14240 -3726
rect 13945 -3912 14004 -3752
rect 13945 -3913 14008 -3912
rect 13942 -3929 14008 -3913
rect 13942 -3963 13958 -3929
rect 13992 -3963 14008 -3929
rect 13942 -3979 14008 -3963
rect 14045 -4028 14140 -4013
rect 14045 -4083 14064 -4028
rect 14122 -4051 14140 -4028
rect 14298 -4051 14358 -3726
rect 14416 -3752 14476 -3726
rect 14653 -3752 14713 -3726
rect 14122 -4083 14358 -4051
rect 14045 -4100 14358 -4083
rect 13477 -4201 14004 -4144
rect 13944 -4300 14004 -4201
rect 13933 -4313 14014 -4300
rect 13933 -4368 13946 -4313
rect 14004 -4368 14014 -4313
rect 13933 -4379 14014 -4368
rect 11292 -4655 11352 -4452
rect 12918 -4456 13812 -4411
rect 1130 -4885 1190 -4859
rect 1322 -5085 1382 -5059
rect 1440 -5085 1500 -5059
rect 1558 -5085 1618 -5059
rect 1676 -5085 1736 -5059
rect 1497 -5140 1563 -5132
rect 1872 -5140 1932 -4859
rect 4274 -4885 4334 -4859
rect 4466 -5085 4526 -5059
rect 4584 -5085 4644 -5059
rect 4702 -5085 4762 -5059
rect 4820 -5085 4880 -5059
rect 1497 -5148 1932 -5140
rect 1497 -5182 1513 -5148
rect 1547 -5182 1932 -5148
rect 1497 -5191 1932 -5182
rect 4641 -5140 4707 -5132
rect 5016 -5140 5076 -4859
rect 7406 -4881 7466 -4855
rect 7598 -5081 7658 -5055
rect 7716 -5081 7776 -5055
rect 7834 -5081 7894 -5055
rect 7952 -5081 8012 -5055
rect 4641 -5148 5076 -5140
rect 4641 -5182 4657 -5148
rect 4691 -5182 5076 -5148
rect 4641 -5191 5076 -5182
rect 7773 -5136 7839 -5128
rect 8148 -5136 8208 -4855
rect 10550 -4881 10610 -4855
rect 13752 -4659 13812 -4456
rect 13944 -4659 14004 -4379
rect 14062 -4659 14122 -4100
rect 14771 -4142 14831 -3726
rect 14889 -3752 14949 -3726
rect 15126 -3752 15186 -3726
rect 15244 -3752 15304 -3726
rect 15252 -3875 15318 -3872
rect 15362 -3875 15422 -3726
rect 15252 -3888 15422 -3875
rect 15252 -3922 15268 -3888
rect 15302 -3922 15422 -3888
rect 15252 -3935 15422 -3922
rect 15252 -3938 15318 -3935
rect 14293 -4159 14831 -4142
rect 14293 -4193 14312 -4159
rect 14346 -4193 14831 -4159
rect 14293 -4199 14831 -4193
rect 14293 -4209 14362 -4199
rect 14293 -4211 14358 -4209
rect 14177 -4549 14243 -4533
rect 14177 -4583 14193 -4549
rect 14227 -4583 14243 -4549
rect 14177 -4599 14243 -4583
rect 14180 -4659 14240 -4599
rect 14298 -4659 14358 -4211
rect 15362 -4411 15422 -3935
rect 14494 -4456 15422 -4411
rect 16062 -4012 16122 -3726
rect 16180 -3752 16240 -3726
rect 16298 -3752 16358 -3726
rect 16503 -3752 16563 -3726
rect 16062 -4029 16198 -4012
rect 16062 -4084 16121 -4029
rect 16179 -4084 16198 -4029
rect 16062 -4099 16198 -4084
rect 16062 -4411 16122 -4099
rect 16621 -4144 16681 -3726
rect 16739 -3752 16799 -3726
rect 16970 -3752 17030 -3726
rect 17088 -3752 17148 -3726
rect 17206 -3752 17266 -3726
rect 17324 -3752 17384 -3726
rect 17089 -3912 17148 -3752
rect 17089 -3913 17152 -3912
rect 17086 -3929 17152 -3913
rect 17086 -3963 17102 -3929
rect 17136 -3963 17152 -3929
rect 17086 -3979 17152 -3963
rect 17189 -4028 17284 -4013
rect 17189 -4083 17208 -4028
rect 17266 -4051 17284 -4028
rect 17442 -4051 17502 -3726
rect 17560 -3752 17620 -3726
rect 17797 -3752 17857 -3726
rect 17266 -4083 17502 -4051
rect 17189 -4100 17502 -4083
rect 16621 -4201 17148 -4144
rect 17088 -4300 17148 -4201
rect 17077 -4313 17158 -4300
rect 17077 -4368 17090 -4313
rect 17148 -4368 17158 -4313
rect 17077 -4379 17158 -4368
rect 16062 -4456 16956 -4411
rect 14494 -4659 14554 -4456
rect 16896 -4659 16956 -4456
rect 17088 -4659 17148 -4379
rect 17206 -4659 17266 -4100
rect 17915 -4142 17975 -3726
rect 18033 -3752 18093 -3726
rect 18270 -3752 18330 -3726
rect 18388 -3752 18448 -3726
rect 18396 -3875 18462 -3872
rect 18506 -3875 18566 -3726
rect 18396 -3888 18566 -3875
rect 18396 -3922 18412 -3888
rect 18446 -3922 18566 -3888
rect 18396 -3935 18566 -3922
rect 18396 -3938 18462 -3935
rect 17437 -4159 17975 -4142
rect 17437 -4193 17456 -4159
rect 17490 -4193 17975 -4159
rect 17437 -4199 17975 -4193
rect 17437 -4209 17506 -4199
rect 17437 -4211 17502 -4209
rect 17321 -4549 17387 -4533
rect 17321 -4583 17337 -4549
rect 17371 -4583 17387 -4549
rect 17321 -4599 17387 -4583
rect 17324 -4659 17384 -4599
rect 17442 -4659 17502 -4211
rect 18506 -4411 18566 -3935
rect 17638 -4456 18566 -4411
rect 19194 -4008 19254 -3722
rect 19312 -3748 19372 -3722
rect 19430 -3748 19490 -3722
rect 19635 -3748 19695 -3722
rect 19194 -4025 19330 -4008
rect 19194 -4080 19253 -4025
rect 19311 -4080 19330 -4025
rect 19194 -4095 19330 -4080
rect 19194 -4407 19254 -4095
rect 19753 -4140 19813 -3722
rect 19871 -3748 19931 -3722
rect 20102 -3748 20162 -3722
rect 20220 -3748 20280 -3722
rect 20338 -3748 20398 -3722
rect 20456 -3748 20516 -3722
rect 20221 -3908 20280 -3748
rect 20221 -3909 20284 -3908
rect 20218 -3925 20284 -3909
rect 20218 -3959 20234 -3925
rect 20268 -3959 20284 -3925
rect 20218 -3975 20284 -3959
rect 20321 -4024 20416 -4009
rect 20321 -4079 20340 -4024
rect 20398 -4047 20416 -4024
rect 20574 -4047 20634 -3722
rect 20692 -3748 20752 -3722
rect 20929 -3748 20989 -3722
rect 20398 -4079 20634 -4047
rect 20321 -4096 20634 -4079
rect 19753 -4197 20280 -4140
rect 20220 -4296 20280 -4197
rect 20209 -4309 20290 -4296
rect 20209 -4364 20222 -4309
rect 20280 -4364 20290 -4309
rect 20209 -4375 20290 -4364
rect 19194 -4452 20088 -4407
rect 17638 -4659 17698 -4456
rect 20028 -4655 20088 -4452
rect 20220 -4655 20280 -4375
rect 20338 -4655 20398 -4096
rect 21047 -4138 21107 -3722
rect 21165 -3748 21225 -3722
rect 21402 -3748 21462 -3722
rect 21520 -3748 21580 -3722
rect 21528 -3871 21594 -3868
rect 21638 -3871 21698 -3722
rect 21528 -3884 21698 -3871
rect 21528 -3918 21544 -3884
rect 21578 -3918 21698 -3884
rect 21528 -3931 21698 -3918
rect 21528 -3934 21594 -3931
rect 20569 -4155 21107 -4138
rect 20569 -4189 20588 -4155
rect 20622 -4189 21107 -4155
rect 20569 -4195 21107 -4189
rect 20569 -4205 20638 -4195
rect 20569 -4207 20634 -4205
rect 20453 -4545 20519 -4529
rect 20453 -4579 20469 -4545
rect 20503 -4579 20519 -4545
rect 20453 -4595 20519 -4579
rect 20456 -4655 20516 -4595
rect 20574 -4655 20634 -4207
rect 21638 -4407 21698 -3931
rect 20770 -4452 21698 -4407
rect 22338 -4008 22398 -3722
rect 22456 -3748 22516 -3722
rect 22574 -3748 22634 -3722
rect 22779 -3748 22839 -3722
rect 22338 -4025 22474 -4008
rect 22338 -4080 22397 -4025
rect 22455 -4080 22474 -4025
rect 22338 -4095 22474 -4080
rect 22338 -4407 22398 -4095
rect 22897 -4140 22957 -3722
rect 23015 -3748 23075 -3722
rect 23246 -3748 23306 -3722
rect 23364 -3748 23424 -3722
rect 23482 -3748 23542 -3722
rect 23600 -3748 23660 -3722
rect 23365 -3908 23424 -3748
rect 23365 -3909 23428 -3908
rect 23362 -3925 23428 -3909
rect 23362 -3959 23378 -3925
rect 23412 -3959 23428 -3925
rect 23362 -3975 23428 -3959
rect 23465 -4024 23560 -4009
rect 23465 -4079 23484 -4024
rect 23542 -4047 23560 -4024
rect 23718 -4047 23778 -3722
rect 23836 -3748 23896 -3722
rect 24073 -3748 24133 -3722
rect 23542 -4079 23778 -4047
rect 23465 -4096 23778 -4079
rect 22897 -4197 23424 -4140
rect 23364 -4296 23424 -4197
rect 23353 -4309 23434 -4296
rect 23353 -4364 23366 -4309
rect 23424 -4364 23434 -4309
rect 23353 -4375 23434 -4364
rect 22338 -4452 23232 -4407
rect 20770 -4655 20830 -4452
rect 23172 -4655 23232 -4452
rect 23364 -4655 23424 -4375
rect 23482 -4655 23542 -4096
rect 24191 -4138 24251 -3722
rect 24309 -3748 24369 -3722
rect 24546 -3748 24606 -3722
rect 24664 -3748 24724 -3722
rect 24672 -3871 24738 -3868
rect 24782 -3871 24842 -3722
rect 24672 -3884 24842 -3871
rect 24672 -3918 24688 -3884
rect 24722 -3918 24842 -3884
rect 24672 -3931 24842 -3918
rect 24672 -3934 24738 -3931
rect 23713 -4155 24251 -4138
rect 23713 -4189 23732 -4155
rect 23766 -4189 24251 -4155
rect 23713 -4195 24251 -4189
rect 23713 -4205 23782 -4195
rect 23713 -4207 23778 -4205
rect 23597 -4545 23663 -4529
rect 23597 -4579 23613 -4545
rect 23647 -4579 23663 -4545
rect 23597 -4595 23663 -4579
rect 23600 -4655 23660 -4595
rect 23718 -4655 23778 -4207
rect 24782 -4407 24842 -3931
rect 23914 -4452 24842 -4407
rect 23914 -4655 23974 -4452
rect 10742 -5081 10802 -5055
rect 10860 -5081 10920 -5055
rect 10978 -5081 11038 -5055
rect 11096 -5081 11156 -5055
rect 7773 -5144 8208 -5136
rect 7773 -5178 7789 -5144
rect 7823 -5178 8208 -5144
rect 7773 -5187 8208 -5178
rect 10917 -5136 10983 -5128
rect 11292 -5136 11352 -4855
rect 13752 -4885 13812 -4859
rect 13944 -5085 14004 -5059
rect 14062 -5085 14122 -5059
rect 14180 -5085 14240 -5059
rect 14298 -5085 14358 -5059
rect 10917 -5144 11352 -5136
rect 10917 -5178 10933 -5144
rect 10967 -5178 11352 -5144
rect 10917 -5187 11352 -5178
rect 14119 -5140 14185 -5132
rect 14494 -5140 14554 -4859
rect 16896 -4885 16956 -4859
rect 17088 -5085 17148 -5059
rect 17206 -5085 17266 -5059
rect 17324 -5085 17384 -5059
rect 17442 -5085 17502 -5059
rect 14119 -5148 14554 -5140
rect 14119 -5182 14135 -5148
rect 14169 -5182 14554 -5148
rect 1497 -5198 1563 -5191
rect 4641 -5198 4707 -5191
rect 7773 -5194 7839 -5187
rect 10917 -5194 10983 -5187
rect 14119 -5191 14554 -5182
rect 17263 -5140 17329 -5132
rect 17638 -5140 17698 -4859
rect 20028 -4881 20088 -4855
rect 20220 -5081 20280 -5055
rect 20338 -5081 20398 -5055
rect 20456 -5081 20516 -5055
rect 20574 -5081 20634 -5055
rect 17263 -5148 17698 -5140
rect 17263 -5182 17279 -5148
rect 17313 -5182 17698 -5148
rect 17263 -5191 17698 -5182
rect 20395 -5136 20461 -5128
rect 20770 -5136 20830 -4855
rect 23172 -4881 23232 -4855
rect 23364 -5081 23424 -5055
rect 23482 -5081 23542 -5055
rect 23600 -5081 23660 -5055
rect 23718 -5081 23778 -5055
rect 20395 -5144 20830 -5136
rect 20395 -5178 20411 -5144
rect 20445 -5178 20830 -5144
rect 20395 -5187 20830 -5178
rect 23539 -5136 23605 -5128
rect 23914 -5136 23974 -4855
rect 23539 -5144 23974 -5136
rect 23539 -5178 23555 -5144
rect 23589 -5178 23974 -5144
rect 23539 -5187 23974 -5178
rect 14119 -5198 14185 -5191
rect 17263 -5198 17329 -5191
rect 20395 -5194 20461 -5187
rect 23539 -5194 23605 -5187
rect 16765 -6155 16825 -6129
rect 16883 -6155 16943 -6129
rect 17001 -6155 17061 -6129
rect 17503 -6151 17563 -6125
rect 17621 -6151 17681 -6125
rect 17739 -6151 17799 -6125
rect 517 -6256 813 -6205
rect 517 -6271 577 -6256
rect 635 -6271 695 -6256
rect 753 -6271 813 -6256
rect 871 -6271 931 -6245
rect 989 -6271 1049 -6245
rect 1107 -6271 1167 -6245
rect 2585 -6254 2881 -6203
rect 2585 -6269 2645 -6254
rect 2703 -6269 2763 -6254
rect 2821 -6269 2881 -6254
rect 2939 -6269 2999 -6243
rect 3057 -6269 3117 -6243
rect 3175 -6269 3235 -6243
rect 4654 -6256 4950 -6205
rect 33 -6471 93 -6445
rect 151 -6471 211 -6445
rect 269 -6471 329 -6445
rect 1354 -6454 1650 -6403
rect 1354 -6471 1414 -6454
rect 1472 -6471 1532 -6454
rect 1590 -6471 1650 -6454
rect 2101 -6469 2161 -6443
rect 2219 -6469 2279 -6443
rect 2337 -6469 2397 -6443
rect 4654 -6271 4714 -6256
rect 4772 -6271 4832 -6256
rect 4890 -6271 4950 -6256
rect 5008 -6271 5068 -6245
rect 5126 -6271 5186 -6245
rect 5244 -6271 5304 -6245
rect 6722 -6254 7018 -6203
rect 6722 -6269 6782 -6254
rect 6840 -6269 6900 -6254
rect 6958 -6269 7018 -6254
rect 7076 -6269 7136 -6243
rect 7194 -6269 7254 -6243
rect 7312 -6269 7372 -6243
rect 8791 -6254 9087 -6203
rect 8791 -6269 8851 -6254
rect 8909 -6269 8969 -6254
rect 9027 -6269 9087 -6254
rect 9145 -6269 9205 -6243
rect 9263 -6269 9323 -6243
rect 9381 -6269 9441 -6243
rect 10859 -6252 11155 -6201
rect 10859 -6267 10919 -6252
rect 10977 -6267 11037 -6252
rect 11095 -6267 11155 -6252
rect 11213 -6267 11273 -6241
rect 11331 -6267 11391 -6241
rect 11449 -6267 11509 -6241
rect 12928 -6254 13224 -6203
rect 3422 -6452 3718 -6401
rect 3422 -6469 3482 -6452
rect 3540 -6469 3600 -6452
rect 3658 -6469 3718 -6452
rect 4170 -6471 4230 -6445
rect 4288 -6471 4348 -6445
rect 4406 -6471 4466 -6445
rect 33 -6688 93 -6671
rect 151 -6688 211 -6671
rect 269 -6688 329 -6671
rect 517 -6688 577 -6671
rect 33 -6739 577 -6688
rect 635 -6697 695 -6671
rect 753 -6697 813 -6671
rect 871 -6690 931 -6671
rect 989 -6690 1049 -6671
rect 1107 -6690 1167 -6671
rect 1354 -6690 1414 -6671
rect 1472 -6690 1532 -6671
rect 158 -7018 218 -6739
rect 871 -6741 1414 -6690
rect 1456 -6697 1532 -6690
rect 1590 -6697 1650 -6671
rect 2101 -6686 2161 -6669
rect 2219 -6686 2279 -6669
rect 2337 -6686 2397 -6669
rect 2585 -6686 2645 -6669
rect 1456 -6741 1531 -6697
rect 2101 -6737 2645 -6686
rect 2703 -6695 2763 -6669
rect 2821 -6695 2881 -6669
rect 2939 -6688 2999 -6669
rect 3057 -6688 3117 -6669
rect 3175 -6688 3235 -6669
rect 3422 -6688 3482 -6669
rect 3540 -6688 3600 -6669
rect 1456 -6828 1516 -6741
rect 1388 -6838 1516 -6828
rect 1388 -6872 1404 -6838
rect 1438 -6872 1516 -6838
rect 460 -6941 756 -6881
rect 460 -6964 520 -6941
rect 578 -6964 638 -6941
rect 696 -6964 756 -6941
rect 814 -6940 1110 -6880
rect 1388 -6882 1516 -6872
rect 814 -6964 874 -6940
rect 932 -6964 992 -6940
rect 1050 -6964 1110 -6940
rect -6 -7032 218 -7018
rect -6 -7066 10 -7032
rect 44 -7066 218 -7032
rect -6 -7078 218 -7066
rect 158 -7591 218 -7078
rect 460 -7390 520 -7364
rect 428 -7531 495 -7524
rect 578 -7531 638 -7364
rect 696 -7390 756 -7364
rect 814 -7390 874 -7364
rect 428 -7540 638 -7531
rect 428 -7574 444 -7540
rect 478 -7574 638 -7540
rect 428 -7590 638 -7574
rect 158 -7607 309 -7591
rect 158 -7641 259 -7607
rect 293 -7641 309 -7607
rect 158 -7657 309 -7641
rect 158 -7696 218 -7657
rect 578 -7696 638 -7590
rect 932 -7531 992 -7364
rect 1050 -7390 1110 -7364
rect 1075 -7531 1142 -7524
rect 932 -7540 1142 -7531
rect 932 -7574 1092 -7540
rect 1126 -7574 1142 -7540
rect 932 -7590 1142 -7574
rect 694 -7624 760 -7608
rect 694 -7658 710 -7624
rect 744 -7658 760 -7624
rect 694 -7674 760 -7658
rect 812 -7623 878 -7608
rect 812 -7657 828 -7623
rect 862 -7657 878 -7623
rect 812 -7673 878 -7657
rect 696 -7696 756 -7674
rect 814 -7696 874 -7673
rect 932 -7696 992 -7590
rect 1456 -7592 1516 -6882
rect 2226 -7016 2286 -6737
rect 2939 -6739 3482 -6688
rect 3524 -6695 3600 -6688
rect 3658 -6695 3718 -6669
rect 5491 -6454 5787 -6403
rect 5491 -6471 5551 -6454
rect 5609 -6471 5669 -6454
rect 5727 -6471 5787 -6454
rect 6238 -6469 6298 -6443
rect 6356 -6469 6416 -6443
rect 6474 -6469 6534 -6443
rect 7559 -6452 7855 -6401
rect 7559 -6469 7619 -6452
rect 7677 -6469 7737 -6452
rect 7795 -6469 7855 -6452
rect 8307 -6469 8367 -6443
rect 8425 -6469 8485 -6443
rect 8543 -6469 8603 -6443
rect 9628 -6452 9924 -6401
rect 9628 -6469 9688 -6452
rect 9746 -6469 9806 -6452
rect 9864 -6469 9924 -6452
rect 10375 -6467 10435 -6441
rect 10493 -6467 10553 -6441
rect 10611 -6467 10671 -6441
rect 12928 -6269 12988 -6254
rect 13046 -6269 13106 -6254
rect 13164 -6269 13224 -6254
rect 13282 -6269 13342 -6243
rect 13400 -6269 13460 -6243
rect 13518 -6269 13578 -6243
rect 14996 -6252 15292 -6201
rect 14996 -6267 15056 -6252
rect 15114 -6267 15174 -6252
rect 15232 -6267 15292 -6252
rect 15350 -6267 15410 -6241
rect 15468 -6267 15528 -6241
rect 15586 -6267 15646 -6241
rect 11696 -6450 11992 -6399
rect 11696 -6467 11756 -6450
rect 11814 -6467 11874 -6450
rect 11932 -6467 11992 -6450
rect 12444 -6469 12504 -6443
rect 12562 -6469 12622 -6443
rect 12680 -6469 12740 -6443
rect 4170 -6688 4230 -6671
rect 4288 -6688 4348 -6671
rect 4406 -6688 4466 -6671
rect 4654 -6688 4714 -6671
rect 3524 -6739 3599 -6695
rect 4170 -6739 4714 -6688
rect 4772 -6697 4832 -6671
rect 4890 -6697 4950 -6671
rect 5008 -6690 5068 -6671
rect 5126 -6690 5186 -6671
rect 5244 -6690 5304 -6671
rect 5491 -6690 5551 -6671
rect 5609 -6690 5669 -6671
rect 3524 -6826 3584 -6739
rect 3456 -6836 3584 -6826
rect 3456 -6870 3472 -6836
rect 3506 -6870 3584 -6836
rect 2528 -6939 2824 -6879
rect 2528 -6962 2588 -6939
rect 2646 -6962 2706 -6939
rect 2764 -6962 2824 -6939
rect 2882 -6938 3178 -6878
rect 3456 -6880 3584 -6870
rect 2882 -6962 2942 -6938
rect 3000 -6962 3060 -6938
rect 3118 -6962 3178 -6938
rect 2062 -7030 2286 -7016
rect 2062 -7064 2078 -7030
rect 2112 -7064 2286 -7030
rect 2062 -7076 2286 -7064
rect 1366 -7608 1516 -7592
rect 1366 -7642 1382 -7608
rect 1416 -7642 1516 -7608
rect 1366 -7658 1516 -7642
rect 1456 -7696 1516 -7658
rect 2226 -7589 2286 -7076
rect 2528 -7388 2588 -7362
rect 2496 -7529 2563 -7522
rect 2646 -7529 2706 -7362
rect 2764 -7388 2824 -7362
rect 2882 -7388 2942 -7362
rect 2496 -7538 2706 -7529
rect 2496 -7572 2512 -7538
rect 2546 -7572 2706 -7538
rect 2496 -7588 2706 -7572
rect 2226 -7605 2377 -7589
rect 2226 -7639 2327 -7605
rect 2361 -7639 2377 -7605
rect 2226 -7655 2377 -7639
rect 2226 -7694 2286 -7655
rect 2646 -7694 2706 -7588
rect 3000 -7529 3060 -7362
rect 3118 -7388 3178 -7362
rect 3143 -7529 3210 -7522
rect 3000 -7538 3210 -7529
rect 3000 -7572 3160 -7538
rect 3194 -7572 3210 -7538
rect 3000 -7588 3210 -7572
rect 2762 -7622 2828 -7606
rect 2762 -7656 2778 -7622
rect 2812 -7656 2828 -7622
rect 2762 -7672 2828 -7656
rect 2880 -7621 2946 -7606
rect 2880 -7655 2896 -7621
rect 2930 -7655 2946 -7621
rect 2880 -7671 2946 -7655
rect 2764 -7694 2824 -7672
rect 2882 -7694 2942 -7671
rect 3000 -7694 3060 -7588
rect 3524 -7590 3584 -6880
rect 4295 -7018 4355 -6739
rect 5008 -6741 5551 -6690
rect 5593 -6697 5669 -6690
rect 5727 -6697 5787 -6671
rect 6238 -6686 6298 -6669
rect 6356 -6686 6416 -6669
rect 6474 -6686 6534 -6669
rect 6722 -6686 6782 -6669
rect 5593 -6741 5668 -6697
rect 6238 -6737 6782 -6686
rect 6840 -6695 6900 -6669
rect 6958 -6695 7018 -6669
rect 7076 -6688 7136 -6669
rect 7194 -6688 7254 -6669
rect 7312 -6688 7372 -6669
rect 7559 -6688 7619 -6669
rect 7677 -6688 7737 -6669
rect 5593 -6828 5653 -6741
rect 5525 -6838 5653 -6828
rect 5525 -6872 5541 -6838
rect 5575 -6872 5653 -6838
rect 4597 -6941 4893 -6881
rect 4597 -6964 4657 -6941
rect 4715 -6964 4775 -6941
rect 4833 -6964 4893 -6941
rect 4951 -6940 5247 -6880
rect 5525 -6882 5653 -6872
rect 4951 -6964 5011 -6940
rect 5069 -6964 5129 -6940
rect 5187 -6964 5247 -6940
rect 4131 -7032 4355 -7018
rect 4131 -7066 4147 -7032
rect 4181 -7066 4355 -7032
rect 4131 -7078 4355 -7066
rect 3434 -7606 3584 -7590
rect 3434 -7640 3450 -7606
rect 3484 -7640 3584 -7606
rect 3434 -7656 3584 -7640
rect 3524 -7694 3584 -7656
rect 4295 -7591 4355 -7078
rect 4597 -7390 4657 -7364
rect 4565 -7531 4632 -7524
rect 4715 -7531 4775 -7364
rect 4833 -7390 4893 -7364
rect 4951 -7390 5011 -7364
rect 4565 -7540 4775 -7531
rect 4565 -7574 4581 -7540
rect 4615 -7574 4775 -7540
rect 4565 -7590 4775 -7574
rect 4295 -7607 4446 -7591
rect 4295 -7641 4396 -7607
rect 4430 -7641 4446 -7607
rect 4295 -7657 4446 -7641
rect 158 -7922 218 -7896
rect 1456 -7922 1516 -7896
rect 2226 -7920 2286 -7894
rect 4295 -7696 4355 -7657
rect 4715 -7696 4775 -7590
rect 5069 -7531 5129 -7364
rect 5187 -7390 5247 -7364
rect 5212 -7531 5279 -7524
rect 5069 -7540 5279 -7531
rect 5069 -7574 5229 -7540
rect 5263 -7574 5279 -7540
rect 5069 -7590 5279 -7574
rect 4831 -7624 4897 -7608
rect 4831 -7658 4847 -7624
rect 4881 -7658 4897 -7624
rect 4831 -7674 4897 -7658
rect 4949 -7623 5015 -7608
rect 4949 -7657 4965 -7623
rect 4999 -7657 5015 -7623
rect 4949 -7673 5015 -7657
rect 4833 -7696 4893 -7674
rect 4951 -7696 5011 -7673
rect 5069 -7696 5129 -7590
rect 5593 -7592 5653 -6882
rect 6363 -7016 6423 -6737
rect 7076 -6739 7619 -6688
rect 7661 -6695 7737 -6688
rect 7795 -6695 7855 -6669
rect 8307 -6686 8367 -6669
rect 8425 -6686 8485 -6669
rect 8543 -6686 8603 -6669
rect 8791 -6686 8851 -6669
rect 7661 -6739 7736 -6695
rect 8307 -6737 8851 -6686
rect 8909 -6695 8969 -6669
rect 9027 -6695 9087 -6669
rect 9145 -6688 9205 -6669
rect 9263 -6688 9323 -6669
rect 9381 -6688 9441 -6669
rect 9628 -6688 9688 -6669
rect 9746 -6688 9806 -6669
rect 7661 -6826 7721 -6739
rect 7593 -6836 7721 -6826
rect 7593 -6870 7609 -6836
rect 7643 -6870 7721 -6836
rect 6665 -6939 6961 -6879
rect 6665 -6962 6725 -6939
rect 6783 -6962 6843 -6939
rect 6901 -6962 6961 -6939
rect 7019 -6938 7315 -6878
rect 7593 -6880 7721 -6870
rect 7019 -6962 7079 -6938
rect 7137 -6962 7197 -6938
rect 7255 -6962 7315 -6938
rect 6199 -7030 6423 -7016
rect 6199 -7064 6215 -7030
rect 6249 -7064 6423 -7030
rect 6199 -7076 6423 -7064
rect 5503 -7608 5653 -7592
rect 5503 -7642 5519 -7608
rect 5553 -7642 5653 -7608
rect 5503 -7658 5653 -7642
rect 5593 -7696 5653 -7658
rect 6363 -7589 6423 -7076
rect 6665 -7388 6725 -7362
rect 6633 -7529 6700 -7522
rect 6783 -7529 6843 -7362
rect 6901 -7388 6961 -7362
rect 7019 -7388 7079 -7362
rect 6633 -7538 6843 -7529
rect 6633 -7572 6649 -7538
rect 6683 -7572 6843 -7538
rect 6633 -7588 6843 -7572
rect 6363 -7605 6514 -7589
rect 6363 -7639 6464 -7605
rect 6498 -7639 6514 -7605
rect 6363 -7655 6514 -7639
rect 6363 -7694 6423 -7655
rect 6783 -7694 6843 -7588
rect 7137 -7529 7197 -7362
rect 7255 -7388 7315 -7362
rect 7280 -7529 7347 -7522
rect 7137 -7538 7347 -7529
rect 7137 -7572 7297 -7538
rect 7331 -7572 7347 -7538
rect 7137 -7588 7347 -7572
rect 6899 -7622 6965 -7606
rect 6899 -7656 6915 -7622
rect 6949 -7656 6965 -7622
rect 6899 -7672 6965 -7656
rect 7017 -7621 7083 -7606
rect 7017 -7655 7033 -7621
rect 7067 -7655 7083 -7621
rect 7017 -7671 7083 -7655
rect 6901 -7694 6961 -7672
rect 7019 -7694 7079 -7671
rect 7137 -7694 7197 -7588
rect 7661 -7590 7721 -6880
rect 8432 -7016 8492 -6737
rect 9145 -6739 9688 -6688
rect 9730 -6695 9806 -6688
rect 9864 -6695 9924 -6669
rect 10375 -6684 10435 -6667
rect 10493 -6684 10553 -6667
rect 10611 -6684 10671 -6667
rect 10859 -6684 10919 -6667
rect 9730 -6739 9805 -6695
rect 10375 -6735 10919 -6684
rect 10977 -6693 11037 -6667
rect 11095 -6693 11155 -6667
rect 11213 -6686 11273 -6667
rect 11331 -6686 11391 -6667
rect 11449 -6686 11509 -6667
rect 11696 -6686 11756 -6667
rect 11814 -6686 11874 -6667
rect 9730 -6826 9790 -6739
rect 9662 -6836 9790 -6826
rect 9662 -6870 9678 -6836
rect 9712 -6870 9790 -6836
rect 8734 -6939 9030 -6879
rect 8734 -6962 8794 -6939
rect 8852 -6962 8912 -6939
rect 8970 -6962 9030 -6939
rect 9088 -6938 9384 -6878
rect 9662 -6880 9790 -6870
rect 9088 -6962 9148 -6938
rect 9206 -6962 9266 -6938
rect 9324 -6962 9384 -6938
rect 8268 -7030 8492 -7016
rect 8268 -7064 8284 -7030
rect 8318 -7064 8492 -7030
rect 8268 -7076 8492 -7064
rect 7571 -7606 7721 -7590
rect 7571 -7640 7587 -7606
rect 7621 -7640 7721 -7606
rect 7571 -7656 7721 -7640
rect 7661 -7694 7721 -7656
rect 8432 -7589 8492 -7076
rect 8734 -7388 8794 -7362
rect 8702 -7529 8769 -7522
rect 8852 -7529 8912 -7362
rect 8970 -7388 9030 -7362
rect 9088 -7388 9148 -7362
rect 8702 -7538 8912 -7529
rect 8702 -7572 8718 -7538
rect 8752 -7572 8912 -7538
rect 8702 -7588 8912 -7572
rect 8432 -7605 8583 -7589
rect 8432 -7639 8533 -7605
rect 8567 -7639 8583 -7605
rect 8432 -7655 8583 -7639
rect 8432 -7694 8492 -7655
rect 8852 -7694 8912 -7588
rect 9206 -7529 9266 -7362
rect 9324 -7388 9384 -7362
rect 9349 -7529 9416 -7522
rect 9206 -7538 9416 -7529
rect 9206 -7572 9366 -7538
rect 9400 -7572 9416 -7538
rect 9206 -7588 9416 -7572
rect 8968 -7622 9034 -7606
rect 8968 -7656 8984 -7622
rect 9018 -7656 9034 -7622
rect 8968 -7672 9034 -7656
rect 9086 -7621 9152 -7606
rect 9086 -7655 9102 -7621
rect 9136 -7655 9152 -7621
rect 9086 -7671 9152 -7655
rect 8970 -7694 9030 -7672
rect 9088 -7694 9148 -7671
rect 9206 -7694 9266 -7588
rect 9730 -7590 9790 -6880
rect 10500 -7014 10560 -6735
rect 11213 -6737 11756 -6686
rect 11798 -6693 11874 -6686
rect 11932 -6693 11992 -6667
rect 13765 -6452 14061 -6401
rect 13765 -6469 13825 -6452
rect 13883 -6469 13943 -6452
rect 14001 -6469 14061 -6452
rect 14512 -6467 14572 -6441
rect 14630 -6467 14690 -6441
rect 14748 -6467 14808 -6441
rect 18241 -6155 18301 -6129
rect 18359 -6155 18419 -6129
rect 18477 -6155 18537 -6129
rect 16765 -6371 16825 -6355
rect 16883 -6371 16943 -6355
rect 17001 -6371 17061 -6355
rect 15833 -6450 16129 -6399
rect 16765 -6407 17061 -6371
rect 17503 -6373 17563 -6351
rect 17621 -6373 17681 -6351
rect 17739 -6373 17799 -6351
rect 18983 -6157 19043 -6131
rect 19101 -6157 19161 -6131
rect 19219 -6157 19279 -6131
rect 19723 -6157 19783 -6131
rect 19841 -6157 19901 -6131
rect 19959 -6157 20019 -6131
rect 20461 -6157 20521 -6131
rect 20579 -6157 20639 -6131
rect 20697 -6157 20757 -6131
rect 21199 -6157 21259 -6131
rect 21317 -6157 21377 -6131
rect 21435 -6157 21495 -6131
rect 21937 -6157 21997 -6131
rect 22055 -6157 22115 -6131
rect 22173 -6157 22233 -6131
rect 15833 -6467 15893 -6450
rect 15951 -6467 16011 -6450
rect 16069 -6467 16129 -6450
rect 16883 -6449 16943 -6407
rect 17503 -6409 17799 -6373
rect 18241 -6373 18301 -6355
rect 18359 -6373 18419 -6355
rect 18477 -6373 18537 -6355
rect 18241 -6409 18537 -6373
rect 18983 -6373 19043 -6357
rect 19101 -6373 19161 -6357
rect 19219 -6373 19279 -6357
rect 18983 -6409 19279 -6373
rect 19723 -6373 19783 -6357
rect 19841 -6373 19901 -6357
rect 19959 -6373 20019 -6357
rect 19723 -6409 20019 -6373
rect 20461 -6373 20521 -6357
rect 20579 -6373 20639 -6357
rect 20697 -6373 20757 -6357
rect 20461 -6409 20757 -6373
rect 21199 -6373 21259 -6357
rect 21317 -6373 21377 -6357
rect 21435 -6373 21495 -6357
rect 21199 -6409 21495 -6373
rect 21937 -6373 21997 -6357
rect 22055 -6373 22115 -6357
rect 22173 -6373 22233 -6357
rect 21937 -6409 22233 -6373
rect 16883 -6483 16895 -6449
rect 16929 -6483 16943 -6449
rect 16883 -6541 16943 -6483
rect 17621 -6451 17681 -6409
rect 17621 -6485 17633 -6451
rect 17667 -6485 17681 -6451
rect 17621 -6539 17681 -6485
rect 18359 -6451 18419 -6409
rect 18359 -6485 18371 -6451
rect 18405 -6485 18419 -6451
rect 12444 -6686 12504 -6669
rect 12562 -6686 12622 -6669
rect 12680 -6686 12740 -6669
rect 12928 -6686 12988 -6669
rect 11798 -6737 11873 -6693
rect 12444 -6737 12988 -6686
rect 13046 -6695 13106 -6669
rect 13164 -6695 13224 -6669
rect 13282 -6688 13342 -6669
rect 13400 -6688 13460 -6669
rect 13518 -6688 13578 -6669
rect 13765 -6688 13825 -6669
rect 13883 -6688 13943 -6669
rect 11798 -6824 11858 -6737
rect 11730 -6834 11858 -6824
rect 11730 -6868 11746 -6834
rect 11780 -6868 11858 -6834
rect 10802 -6937 11098 -6877
rect 10802 -6960 10862 -6937
rect 10920 -6960 10980 -6937
rect 11038 -6960 11098 -6937
rect 11156 -6936 11452 -6876
rect 11730 -6878 11858 -6868
rect 11156 -6960 11216 -6936
rect 11274 -6960 11334 -6936
rect 11392 -6960 11452 -6936
rect 10336 -7028 10560 -7014
rect 10336 -7062 10352 -7028
rect 10386 -7062 10560 -7028
rect 10336 -7074 10560 -7062
rect 9640 -7606 9790 -7590
rect 9640 -7640 9656 -7606
rect 9690 -7640 9790 -7606
rect 9640 -7656 9790 -7640
rect 9730 -7694 9790 -7656
rect 10500 -7587 10560 -7074
rect 10802 -7386 10862 -7360
rect 10770 -7527 10837 -7520
rect 10920 -7527 10980 -7360
rect 11038 -7386 11098 -7360
rect 11156 -7386 11216 -7360
rect 10770 -7536 10980 -7527
rect 10770 -7570 10786 -7536
rect 10820 -7570 10980 -7536
rect 10770 -7586 10980 -7570
rect 10500 -7603 10651 -7587
rect 10500 -7637 10601 -7603
rect 10635 -7637 10651 -7603
rect 10500 -7653 10651 -7637
rect 10500 -7692 10560 -7653
rect 10920 -7692 10980 -7586
rect 11274 -7527 11334 -7360
rect 11392 -7386 11452 -7360
rect 11417 -7527 11484 -7520
rect 11274 -7536 11484 -7527
rect 11274 -7570 11434 -7536
rect 11468 -7570 11484 -7536
rect 11274 -7586 11484 -7570
rect 11036 -7620 11102 -7604
rect 11036 -7654 11052 -7620
rect 11086 -7654 11102 -7620
rect 11036 -7670 11102 -7654
rect 11154 -7619 11220 -7604
rect 11154 -7653 11170 -7619
rect 11204 -7653 11220 -7619
rect 11154 -7669 11220 -7653
rect 11038 -7692 11098 -7670
rect 11156 -7692 11216 -7669
rect 11274 -7692 11334 -7586
rect 11798 -7588 11858 -6878
rect 12569 -7016 12629 -6737
rect 13282 -6739 13825 -6688
rect 13867 -6695 13943 -6688
rect 14001 -6695 14061 -6669
rect 14512 -6684 14572 -6667
rect 14630 -6684 14690 -6667
rect 14748 -6684 14808 -6667
rect 14996 -6684 15056 -6667
rect 13867 -6739 13942 -6695
rect 14512 -6735 15056 -6684
rect 15114 -6693 15174 -6667
rect 15232 -6693 15292 -6667
rect 15350 -6686 15410 -6667
rect 15468 -6686 15528 -6667
rect 15586 -6686 15646 -6667
rect 15833 -6686 15893 -6667
rect 15951 -6686 16011 -6667
rect 13867 -6826 13927 -6739
rect 13799 -6836 13927 -6826
rect 13799 -6870 13815 -6836
rect 13849 -6870 13927 -6836
rect 12871 -6939 13167 -6879
rect 12871 -6962 12931 -6939
rect 12989 -6962 13049 -6939
rect 13107 -6962 13167 -6939
rect 13225 -6938 13521 -6878
rect 13799 -6880 13927 -6870
rect 13225 -6962 13285 -6938
rect 13343 -6962 13403 -6938
rect 13461 -6962 13521 -6938
rect 12405 -7030 12629 -7016
rect 12405 -7064 12421 -7030
rect 12455 -7064 12629 -7030
rect 12405 -7076 12629 -7064
rect 11708 -7604 11858 -7588
rect 11708 -7638 11724 -7604
rect 11758 -7638 11858 -7604
rect 11708 -7654 11858 -7638
rect 11798 -7692 11858 -7654
rect 12569 -7589 12629 -7076
rect 12871 -7388 12931 -7362
rect 12839 -7529 12906 -7522
rect 12989 -7529 13049 -7362
rect 13107 -7388 13167 -7362
rect 13225 -7388 13285 -7362
rect 12839 -7538 13049 -7529
rect 12839 -7572 12855 -7538
rect 12889 -7572 13049 -7538
rect 12839 -7588 13049 -7572
rect 12569 -7605 12720 -7589
rect 12569 -7639 12670 -7605
rect 12704 -7639 12720 -7605
rect 12569 -7655 12720 -7639
rect 3524 -7920 3584 -7894
rect 4295 -7922 4355 -7896
rect 578 -8122 638 -8096
rect 696 -8122 756 -8096
rect 814 -8122 874 -8096
rect 932 -8122 992 -8096
rect 2646 -8120 2706 -8094
rect 2764 -8120 2824 -8094
rect 2882 -8120 2942 -8094
rect 3000 -8120 3060 -8094
rect 5593 -7922 5653 -7896
rect 6363 -7920 6423 -7894
rect 7661 -7920 7721 -7894
rect 8432 -7920 8492 -7894
rect 9730 -7920 9790 -7894
rect 10500 -7918 10560 -7892
rect 12569 -7694 12629 -7655
rect 12989 -7694 13049 -7588
rect 13343 -7529 13403 -7362
rect 13461 -7388 13521 -7362
rect 13486 -7529 13553 -7522
rect 13343 -7538 13553 -7529
rect 13343 -7572 13503 -7538
rect 13537 -7572 13553 -7538
rect 13343 -7588 13553 -7572
rect 13105 -7622 13171 -7606
rect 13105 -7656 13121 -7622
rect 13155 -7656 13171 -7622
rect 13105 -7672 13171 -7656
rect 13223 -7621 13289 -7606
rect 13223 -7655 13239 -7621
rect 13273 -7655 13289 -7621
rect 13223 -7671 13289 -7655
rect 13107 -7694 13167 -7672
rect 13225 -7694 13285 -7671
rect 13343 -7694 13403 -7588
rect 13867 -7590 13927 -6880
rect 14637 -7014 14697 -6735
rect 15350 -6737 15893 -6686
rect 15935 -6693 16011 -6686
rect 16069 -6693 16129 -6667
rect 15935 -6737 16010 -6693
rect 15935 -6824 15995 -6737
rect 18359 -6543 18419 -6485
rect 19101 -6451 19161 -6409
rect 19101 -6485 19113 -6451
rect 19147 -6485 19161 -6451
rect 19101 -6543 19161 -6485
rect 19841 -6451 19901 -6409
rect 19841 -6485 19853 -6451
rect 19887 -6485 19901 -6451
rect 19841 -6543 19901 -6485
rect 20579 -6451 20639 -6409
rect 20579 -6485 20591 -6451
rect 20625 -6485 20639 -6451
rect 20579 -6543 20639 -6485
rect 21317 -6451 21377 -6409
rect 21317 -6485 21329 -6451
rect 21363 -6485 21377 -6451
rect 21317 -6539 21377 -6485
rect 22055 -6451 22115 -6409
rect 22055 -6485 22067 -6451
rect 22101 -6485 22115 -6451
rect 22055 -6539 22115 -6485
rect 16883 -6767 16943 -6741
rect 17621 -6765 17681 -6739
rect 18359 -6769 18419 -6743
rect 19101 -6769 19161 -6743
rect 19841 -6769 19901 -6743
rect 20579 -6769 20639 -6743
rect 21317 -6765 21377 -6739
rect 22055 -6765 22115 -6739
rect 15867 -6834 15995 -6824
rect 15867 -6868 15883 -6834
rect 15917 -6868 15995 -6834
rect 14939 -6937 15235 -6877
rect 14939 -6960 14999 -6937
rect 15057 -6960 15117 -6937
rect 15175 -6960 15235 -6937
rect 15293 -6936 15589 -6876
rect 15867 -6878 15995 -6868
rect 15293 -6960 15353 -6936
rect 15411 -6960 15471 -6936
rect 15529 -6960 15589 -6936
rect 14473 -7028 14697 -7014
rect 14473 -7062 14489 -7028
rect 14523 -7062 14697 -7028
rect 14473 -7074 14697 -7062
rect 13777 -7606 13927 -7590
rect 13777 -7640 13793 -7606
rect 13827 -7640 13927 -7606
rect 13777 -7656 13927 -7640
rect 13867 -7694 13927 -7656
rect 14637 -7587 14697 -7074
rect 14939 -7386 14999 -7360
rect 14907 -7527 14974 -7520
rect 15057 -7527 15117 -7360
rect 15175 -7386 15235 -7360
rect 15293 -7386 15353 -7360
rect 14907 -7536 15117 -7527
rect 14907 -7570 14923 -7536
rect 14957 -7570 15117 -7536
rect 14907 -7586 15117 -7570
rect 14637 -7603 14788 -7587
rect 14637 -7637 14738 -7603
rect 14772 -7637 14788 -7603
rect 14637 -7653 14788 -7637
rect 14637 -7692 14697 -7653
rect 15057 -7692 15117 -7586
rect 15411 -7527 15471 -7360
rect 15529 -7386 15589 -7360
rect 15554 -7527 15621 -7520
rect 15411 -7536 15621 -7527
rect 15411 -7570 15571 -7536
rect 15605 -7570 15621 -7536
rect 15411 -7586 15621 -7570
rect 15173 -7620 15239 -7604
rect 15173 -7654 15189 -7620
rect 15223 -7654 15239 -7620
rect 15173 -7670 15239 -7654
rect 15291 -7619 15357 -7604
rect 15291 -7653 15307 -7619
rect 15341 -7653 15357 -7619
rect 15291 -7669 15357 -7653
rect 15175 -7692 15235 -7670
rect 15293 -7692 15353 -7669
rect 15411 -7692 15471 -7586
rect 15935 -7588 15995 -6878
rect 15845 -7604 15995 -7588
rect 15845 -7638 15861 -7604
rect 15895 -7638 15995 -7604
rect 15845 -7654 15995 -7638
rect 15935 -7692 15995 -7654
rect 11798 -7918 11858 -7892
rect 12569 -7920 12629 -7894
rect 4715 -8122 4775 -8096
rect 4833 -8122 4893 -8096
rect 4951 -8122 5011 -8096
rect 5069 -8122 5129 -8096
rect 6783 -8120 6843 -8094
rect 6901 -8120 6961 -8094
rect 7019 -8120 7079 -8094
rect 7137 -8120 7197 -8094
rect 8852 -8120 8912 -8094
rect 8970 -8120 9030 -8094
rect 9088 -8120 9148 -8094
rect 9206 -8120 9266 -8094
rect 10920 -8118 10980 -8092
rect 11038 -8118 11098 -8092
rect 11156 -8118 11216 -8092
rect 11274 -8118 11334 -8092
rect 13867 -7920 13927 -7894
rect 14637 -7918 14697 -7892
rect 15935 -7918 15995 -7892
rect 12989 -8120 13049 -8094
rect 13107 -8120 13167 -8094
rect 13225 -8120 13285 -8094
rect 13343 -8120 13403 -8094
rect 15057 -8118 15117 -8092
rect 15175 -8118 15235 -8092
rect 15293 -8118 15353 -8092
rect 15411 -8118 15471 -8092
<< polycont >>
rect 11874 4220 11908 4254
rect 13042 4220 13076 4254
rect 14210 4220 14244 4254
rect 15378 4220 15412 4254
rect 16552 4222 16586 4256
rect 17720 4222 17754 4256
rect 18888 4222 18922 4256
rect 20056 4222 20090 4256
rect 11874 4112 11908 4146
rect 13042 4112 13076 4146
rect 14210 4112 14244 4146
rect 968 3615 1002 3649
rect 850 3498 884 3532
rect 2416 3615 2450 3649
rect 2298 3498 2332 3532
rect 3914 3617 3948 3651
rect 3796 3500 3830 3534
rect 5362 3617 5396 3651
rect 5244 3500 5278 3534
rect 6882 3615 6916 3649
rect 6764 3498 6798 3532
rect 8330 3615 8364 3649
rect 8212 3498 8246 3532
rect 9828 3617 9862 3651
rect 9710 3500 9744 3534
rect 15378 4112 15412 4146
rect 16552 4114 16586 4148
rect 17720 4114 17754 4148
rect 11276 3617 11310 3651
rect 11158 3500 11192 3534
rect 12169 3349 12203 3383
rect 18888 4114 18922 4148
rect 20056 4114 20090 4148
rect 13337 3349 13371 3383
rect 14505 3349 14539 3383
rect 15673 3349 15707 3383
rect 16847 3351 16881 3385
rect 18015 3351 18049 3385
rect 497 2988 531 3022
rect 615 2988 649 3022
rect 1945 2988 1979 3022
rect 2063 2988 2097 3022
rect 3443 2990 3477 3024
rect 3561 2990 3595 3024
rect 4891 2990 4925 3024
rect 5009 2990 5043 3024
rect 6411 2988 6445 3022
rect 6529 2988 6563 3022
rect 7859 2988 7893 3022
rect 7977 2988 8011 3022
rect 9357 2990 9391 3024
rect 9475 2990 9509 3024
rect 10805 2990 10839 3024
rect 19183 3351 19217 3385
rect 20351 3351 20385 3385
rect 10923 2990 10957 3024
rect 365 1382 423 1437
rect 1346 1503 1380 1537
rect 1452 1383 1510 1438
rect 1334 1098 1392 1153
rect 2656 1544 2690 1578
rect 1700 1273 1734 1307
rect 1581 883 1615 917
rect 3509 1382 3567 1437
rect 4490 1503 4524 1537
rect 4596 1383 4654 1438
rect 4478 1098 4536 1153
rect 5800 1544 5834 1578
rect 4844 1273 4878 1307
rect 4725 883 4759 917
rect 6641 1386 6699 1441
rect 7622 1507 7656 1541
rect 7728 1387 7786 1442
rect 7610 1102 7668 1157
rect 8932 1548 8966 1582
rect 7976 1277 8010 1311
rect 7857 887 7891 921
rect 9785 1386 9843 1441
rect 10766 1507 10800 1541
rect 10872 1387 10930 1442
rect 10754 1102 10812 1157
rect 12076 1548 12110 1582
rect 11120 1277 11154 1311
rect 11001 887 11035 921
rect 12987 1382 13045 1437
rect 13968 1503 14002 1537
rect 14074 1383 14132 1438
rect 13956 1098 14014 1153
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 15278 1544 15312 1578
rect 14322 1273 14356 1307
rect 14203 883 14237 917
rect 16131 1382 16189 1437
rect 17112 1503 17146 1537
rect 17218 1383 17276 1438
rect 17100 1098 17158 1153
rect 18422 1544 18456 1578
rect 17466 1273 17500 1307
rect 17347 883 17381 917
rect 19263 1386 19321 1441
rect 20244 1507 20278 1541
rect 20350 1387 20408 1442
rect 20232 1102 20290 1157
rect 21554 1548 21588 1582
rect 20598 1277 20632 1311
rect 20479 887 20513 921
rect 22407 1386 22465 1441
rect 23388 1507 23422 1541
rect 23494 1387 23552 1442
rect 23376 1102 23434 1157
rect 24698 1548 24732 1582
rect 23742 1277 23776 1311
rect 23623 887 23657 921
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 23565 288 23599 322
rect 365 -1352 423 -1297
rect 1346 -1231 1380 -1197
rect 1452 -1351 1510 -1296
rect 1334 -1636 1392 -1581
rect 2656 -1190 2690 -1156
rect 1700 -1461 1734 -1427
rect 1581 -1851 1615 -1817
rect 3509 -1352 3567 -1297
rect 4490 -1231 4524 -1197
rect 4596 -1351 4654 -1296
rect 4478 -1636 4536 -1581
rect 5800 -1190 5834 -1156
rect 4844 -1461 4878 -1427
rect 4725 -1851 4759 -1817
rect 6641 -1348 6699 -1293
rect 7622 -1227 7656 -1193
rect 7728 -1347 7786 -1292
rect 7610 -1632 7668 -1577
rect 8932 -1186 8966 -1152
rect 7976 -1457 8010 -1423
rect 7857 -1847 7891 -1813
rect 9785 -1348 9843 -1293
rect 10766 -1227 10800 -1193
rect 10872 -1347 10930 -1292
rect 10754 -1632 10812 -1577
rect 12076 -1186 12110 -1152
rect 11120 -1457 11154 -1423
rect 11001 -1847 11035 -1813
rect 12987 -1352 13045 -1297
rect 13968 -1231 14002 -1197
rect 14074 -1351 14132 -1296
rect 13956 -1636 14014 -1581
rect 1523 -2450 1557 -2416
rect 4667 -2450 4701 -2416
rect 15278 -1190 15312 -1156
rect 14322 -1461 14356 -1427
rect 14203 -1851 14237 -1817
rect 16131 -1352 16189 -1297
rect 17112 -1231 17146 -1197
rect 17218 -1351 17276 -1296
rect 17100 -1636 17158 -1581
rect 18422 -1190 18456 -1156
rect 17466 -1461 17500 -1427
rect 17347 -1851 17381 -1817
rect 19263 -1348 19321 -1293
rect 20244 -1227 20278 -1193
rect 20350 -1347 20408 -1292
rect 20232 -1632 20290 -1577
rect 21554 -1186 21588 -1152
rect 20598 -1457 20632 -1423
rect 20479 -1847 20513 -1813
rect 22407 -1348 22465 -1293
rect 23388 -1227 23422 -1193
rect 23494 -1347 23552 -1292
rect 23376 -1632 23434 -1577
rect 24698 -1186 24732 -1152
rect 23742 -1457 23776 -1423
rect 23623 -1847 23657 -1813
rect 7799 -2446 7833 -2412
rect 10943 -2446 10977 -2412
rect 14145 -2450 14179 -2416
rect 17289 -2450 17323 -2416
rect 20421 -2446 20455 -2412
rect 23565 -2446 23599 -2412
rect 355 -4084 413 -4029
rect 1336 -3963 1370 -3929
rect 1442 -4083 1500 -4028
rect 1324 -4368 1382 -4313
rect 2646 -3922 2680 -3888
rect 1690 -4193 1724 -4159
rect 1571 -4583 1605 -4549
rect 3499 -4084 3557 -4029
rect 4480 -3963 4514 -3929
rect 4586 -4083 4644 -4028
rect 4468 -4368 4526 -4313
rect 5790 -3922 5824 -3888
rect 4834 -4193 4868 -4159
rect 4715 -4583 4749 -4549
rect 6631 -4080 6689 -4025
rect 7612 -3959 7646 -3925
rect 7718 -4079 7776 -4024
rect 7600 -4364 7658 -4309
rect 8922 -3918 8956 -3884
rect 7966 -4189 8000 -4155
rect 7847 -4579 7881 -4545
rect 9775 -4080 9833 -4025
rect 10756 -3959 10790 -3925
rect 10862 -4079 10920 -4024
rect 10744 -4364 10802 -4309
rect 12066 -3918 12100 -3884
rect 11110 -4189 11144 -4155
rect 10991 -4579 11025 -4545
rect 12977 -4084 13035 -4029
rect 13958 -3963 13992 -3929
rect 14064 -4083 14122 -4028
rect 13946 -4368 14004 -4313
rect 1513 -5182 1547 -5148
rect 4657 -5182 4691 -5148
rect 15268 -3922 15302 -3888
rect 14312 -4193 14346 -4159
rect 14193 -4583 14227 -4549
rect 16121 -4084 16179 -4029
rect 17102 -3963 17136 -3929
rect 17208 -4083 17266 -4028
rect 17090 -4368 17148 -4313
rect 18412 -3922 18446 -3888
rect 17456 -4193 17490 -4159
rect 17337 -4583 17371 -4549
rect 19253 -4080 19311 -4025
rect 20234 -3959 20268 -3925
rect 20340 -4079 20398 -4024
rect 20222 -4364 20280 -4309
rect 21544 -3918 21578 -3884
rect 20588 -4189 20622 -4155
rect 20469 -4579 20503 -4545
rect 22397 -4080 22455 -4025
rect 23378 -3959 23412 -3925
rect 23484 -4079 23542 -4024
rect 23366 -4364 23424 -4309
rect 24688 -3918 24722 -3884
rect 23732 -4189 23766 -4155
rect 23613 -4579 23647 -4545
rect 7789 -5178 7823 -5144
rect 10933 -5178 10967 -5144
rect 14135 -5182 14169 -5148
rect 17279 -5182 17313 -5148
rect 20411 -5178 20445 -5144
rect 23555 -5178 23589 -5144
rect 1404 -6872 1438 -6838
rect 10 -7066 44 -7032
rect 444 -7574 478 -7540
rect 259 -7641 293 -7607
rect 1092 -7574 1126 -7540
rect 710 -7658 744 -7624
rect 828 -7657 862 -7623
rect 3472 -6870 3506 -6836
rect 2078 -7064 2112 -7030
rect 1382 -7642 1416 -7608
rect 2512 -7572 2546 -7538
rect 2327 -7639 2361 -7605
rect 3160 -7572 3194 -7538
rect 2778 -7656 2812 -7622
rect 2896 -7655 2930 -7621
rect 5541 -6872 5575 -6838
rect 4147 -7066 4181 -7032
rect 3450 -7640 3484 -7606
rect 4581 -7574 4615 -7540
rect 4396 -7641 4430 -7607
rect 5229 -7574 5263 -7540
rect 4847 -7658 4881 -7624
rect 4965 -7657 4999 -7623
rect 7609 -6870 7643 -6836
rect 6215 -7064 6249 -7030
rect 5519 -7642 5553 -7608
rect 6649 -7572 6683 -7538
rect 6464 -7639 6498 -7605
rect 7297 -7572 7331 -7538
rect 6915 -7656 6949 -7622
rect 7033 -7655 7067 -7621
rect 9678 -6870 9712 -6836
rect 8284 -7064 8318 -7030
rect 7587 -7640 7621 -7606
rect 8718 -7572 8752 -7538
rect 8533 -7639 8567 -7605
rect 9366 -7572 9400 -7538
rect 8984 -7656 9018 -7622
rect 9102 -7655 9136 -7621
rect 16895 -6483 16929 -6449
rect 17633 -6485 17667 -6451
rect 18371 -6485 18405 -6451
rect 11746 -6868 11780 -6834
rect 10352 -7062 10386 -7028
rect 9656 -7640 9690 -7606
rect 10786 -7570 10820 -7536
rect 10601 -7637 10635 -7603
rect 11434 -7570 11468 -7536
rect 11052 -7654 11086 -7620
rect 11170 -7653 11204 -7619
rect 13815 -6870 13849 -6836
rect 12421 -7064 12455 -7030
rect 11724 -7638 11758 -7604
rect 12855 -7572 12889 -7538
rect 12670 -7639 12704 -7605
rect 13503 -7572 13537 -7538
rect 13121 -7656 13155 -7622
rect 13239 -7655 13273 -7621
rect 19113 -6485 19147 -6451
rect 19853 -6485 19887 -6451
rect 20591 -6485 20625 -6451
rect 21329 -6485 21363 -6451
rect 22067 -6485 22101 -6451
rect 15883 -6868 15917 -6834
rect 14489 -7062 14523 -7028
rect 13793 -7640 13827 -7606
rect 14923 -7570 14957 -7536
rect 14738 -7637 14772 -7603
rect 15571 -7570 15605 -7536
rect 15189 -7654 15223 -7620
rect 15307 -7653 15341 -7619
rect 15861 -7638 15895 -7604
<< locali >>
rect 12460 4332 12664 4344
rect 12460 4260 12492 4332
rect 12636 4260 12664 4332
rect 12460 4258 12522 4260
rect 12602 4258 12664 4260
rect 11858 4220 11874 4254
rect 11908 4220 11924 4254
rect 12460 4242 12664 4258
rect 13628 4332 13832 4344
rect 13628 4260 13660 4332
rect 13804 4260 13832 4332
rect 13628 4258 13690 4260
rect 13770 4258 13832 4260
rect 13026 4220 13042 4254
rect 13076 4220 13092 4254
rect 13628 4242 13832 4258
rect 14796 4332 15000 4344
rect 14796 4260 14828 4332
rect 14972 4260 15000 4332
rect 14796 4258 14858 4260
rect 14938 4258 15000 4260
rect 14194 4220 14210 4254
rect 14244 4220 14260 4254
rect 14796 4242 15000 4258
rect 15964 4332 16168 4344
rect 15964 4260 15996 4332
rect 16140 4260 16168 4332
rect 15964 4258 16026 4260
rect 16106 4258 16168 4260
rect 15362 4220 15378 4254
rect 15412 4220 15428 4254
rect 15964 4242 16168 4258
rect 17138 4334 17342 4346
rect 17138 4262 17170 4334
rect 17314 4262 17342 4334
rect 17138 4260 17200 4262
rect 17280 4260 17342 4262
rect 16536 4222 16552 4256
rect 16586 4222 16602 4256
rect 17138 4244 17342 4260
rect 18306 4334 18510 4346
rect 18306 4262 18338 4334
rect 18482 4262 18510 4334
rect 18306 4260 18368 4262
rect 18448 4260 18510 4262
rect 17704 4222 17720 4256
rect 17754 4222 17770 4256
rect 18306 4244 18510 4260
rect 19474 4334 19678 4346
rect 19474 4262 19506 4334
rect 19650 4262 19678 4334
rect 19474 4260 19536 4262
rect 19616 4260 19678 4262
rect 18872 4222 18888 4256
rect 18922 4222 18938 4256
rect 19474 4244 19678 4260
rect 20642 4334 20846 4346
rect 20642 4262 20674 4334
rect 20818 4262 20846 4334
rect 20642 4260 20704 4262
rect 20784 4260 20846 4262
rect 20040 4222 20056 4256
rect 20090 4222 20106 4256
rect 20642 4244 20846 4260
rect 490 4125 658 4141
rect 490 4055 506 4125
rect 642 4055 658 4125
rect 490 4039 658 4055
rect 1938 4125 2106 4141
rect 1938 4055 1954 4125
rect 2090 4055 2106 4125
rect 1938 4039 2106 4055
rect 3436 4127 3604 4143
rect 3436 4057 3452 4127
rect 3588 4057 3604 4127
rect 3436 4041 3604 4057
rect 4884 4127 5052 4143
rect 4884 4057 4900 4127
rect 5036 4057 5052 4127
rect 4884 4041 5052 4057
rect 6404 4125 6572 4141
rect 6404 4055 6420 4125
rect 6556 4055 6572 4125
rect 6404 4039 6572 4055
rect 7852 4125 8020 4141
rect 7852 4055 7868 4125
rect 8004 4055 8020 4125
rect 7852 4039 8020 4055
rect 9350 4127 9518 4143
rect 9350 4057 9366 4127
rect 9502 4057 9518 4127
rect 9350 4041 9518 4057
rect 10798 4127 10966 4143
rect 10798 4057 10814 4127
rect 10950 4057 10966 4127
rect 11858 4112 11874 4146
rect 11908 4112 11924 4146
rect 13026 4112 13042 4146
rect 13076 4112 13092 4146
rect 14194 4112 14210 4146
rect 14244 4112 14260 4146
rect 15362 4112 15378 4146
rect 15412 4112 15428 4146
rect 16536 4114 16552 4148
rect 16586 4114 16602 4148
rect 17704 4114 17720 4148
rect 17754 4114 17770 4148
rect 18872 4114 18888 4148
rect 18922 4114 18938 4148
rect 20040 4114 20056 4148
rect 20090 4114 20106 4148
rect 10798 4041 10966 4057
rect 11964 4082 11998 4098
rect 1027 3935 1297 3969
rect 201 3885 235 3901
rect 201 3693 235 3709
rect 319 3885 353 3901
rect 319 3693 353 3709
rect 437 3885 471 3901
rect 437 3693 471 3709
rect 555 3885 589 3901
rect 555 3693 589 3709
rect 673 3885 707 3901
rect 673 3693 707 3709
rect 791 3885 825 3901
rect 791 3693 825 3709
rect 909 3885 943 3901
rect 909 3693 943 3709
rect 1027 3885 1061 3935
rect 1027 3693 1061 3709
rect 1145 3885 1179 3901
rect 1145 3693 1179 3709
rect 1263 3885 1297 3935
rect 2475 3935 2745 3969
rect 1263 3693 1297 3709
rect 1649 3885 1683 3901
rect 1649 3693 1683 3709
rect 1767 3885 1801 3901
rect 1767 3693 1801 3709
rect 1885 3885 1919 3901
rect 1885 3693 1919 3709
rect 2003 3885 2037 3901
rect 2003 3693 2037 3709
rect 2121 3885 2155 3901
rect 2121 3693 2155 3709
rect 2239 3885 2273 3901
rect 2239 3693 2273 3709
rect 2357 3885 2391 3901
rect 2357 3693 2391 3709
rect 2475 3885 2509 3935
rect 2475 3693 2509 3709
rect 2593 3885 2627 3901
rect 2593 3693 2627 3709
rect 2711 3885 2745 3935
rect 3973 3937 4243 3971
rect 2711 3693 2745 3709
rect 3147 3887 3181 3903
rect 3147 3695 3181 3711
rect 3265 3887 3299 3903
rect 3265 3695 3299 3711
rect 3383 3887 3417 3903
rect 3383 3695 3417 3711
rect 3501 3887 3535 3903
rect 3501 3695 3535 3711
rect 3619 3887 3653 3903
rect 3619 3695 3653 3711
rect 3737 3887 3771 3903
rect 3737 3695 3771 3711
rect 3855 3887 3889 3903
rect 3855 3695 3889 3711
rect 3973 3887 4007 3937
rect 3973 3695 4007 3711
rect 4091 3887 4125 3903
rect 4091 3695 4125 3711
rect 4209 3887 4243 3937
rect 5421 3937 5691 3971
rect 4209 3695 4243 3711
rect 4595 3887 4629 3903
rect 4595 3695 4629 3711
rect 4713 3887 4747 3903
rect 4713 3695 4747 3711
rect 4831 3887 4865 3903
rect 4831 3695 4865 3711
rect 4949 3887 4983 3903
rect 4949 3695 4983 3711
rect 5067 3887 5101 3903
rect 5067 3695 5101 3711
rect 5185 3887 5219 3903
rect 5185 3695 5219 3711
rect 5303 3887 5337 3903
rect 5303 3695 5337 3711
rect 5421 3887 5455 3937
rect 5421 3695 5455 3711
rect 5539 3887 5573 3903
rect 5539 3695 5573 3711
rect 5657 3887 5691 3937
rect 6941 3935 7211 3969
rect 5657 3695 5691 3711
rect 6115 3885 6149 3901
rect 6115 3693 6149 3709
rect 6233 3885 6267 3901
rect 6233 3693 6267 3709
rect 6351 3885 6385 3901
rect 6351 3693 6385 3709
rect 6469 3885 6503 3901
rect 6469 3693 6503 3709
rect 6587 3885 6621 3901
rect 6587 3693 6621 3709
rect 6705 3885 6739 3901
rect 6705 3693 6739 3709
rect 6823 3885 6857 3901
rect 6823 3693 6857 3709
rect 6941 3885 6975 3935
rect 6941 3693 6975 3709
rect 7059 3885 7093 3901
rect 7059 3693 7093 3709
rect 7177 3885 7211 3935
rect 8389 3935 8659 3969
rect 7177 3693 7211 3709
rect 7563 3885 7597 3901
rect 7563 3693 7597 3709
rect 7681 3885 7715 3901
rect 7681 3693 7715 3709
rect 7799 3885 7833 3901
rect 7799 3693 7833 3709
rect 7917 3885 7951 3901
rect 7917 3693 7951 3709
rect 8035 3885 8069 3901
rect 8035 3693 8069 3709
rect 8153 3885 8187 3901
rect 8153 3693 8187 3709
rect 8271 3885 8305 3901
rect 8271 3693 8305 3709
rect 8389 3885 8423 3935
rect 8389 3693 8423 3709
rect 8507 3885 8541 3901
rect 8507 3693 8541 3709
rect 8625 3885 8659 3935
rect 9887 3937 10157 3971
rect 8625 3693 8659 3709
rect 9061 3887 9095 3903
rect 9061 3695 9095 3711
rect 9179 3887 9213 3903
rect 9179 3695 9213 3711
rect 9297 3887 9331 3903
rect 9297 3695 9331 3711
rect 9415 3887 9449 3903
rect 9415 3695 9449 3711
rect 9533 3887 9567 3903
rect 9533 3695 9567 3711
rect 9651 3887 9685 3903
rect 9651 3695 9685 3711
rect 9769 3887 9803 3903
rect 9769 3695 9803 3711
rect 9887 3887 9921 3937
rect 9887 3695 9921 3711
rect 10005 3887 10039 3903
rect 10005 3695 10039 3711
rect 10123 3887 10157 3937
rect 11335 3937 11605 3971
rect 10123 3695 10157 3711
rect 10509 3887 10543 3903
rect 10509 3695 10543 3711
rect 10627 3887 10661 3903
rect 10627 3695 10661 3711
rect 10745 3887 10779 3903
rect 10745 3695 10779 3711
rect 10863 3887 10897 3903
rect 10863 3695 10897 3711
rect 10981 3887 11015 3903
rect 10981 3695 11015 3711
rect 11099 3887 11133 3903
rect 11099 3695 11133 3711
rect 11217 3887 11251 3903
rect 11217 3695 11251 3711
rect 11335 3887 11369 3937
rect 11335 3695 11369 3711
rect 11453 3887 11487 3903
rect 11453 3695 11487 3711
rect 11571 3887 11605 3937
rect 11571 3695 11605 3711
rect 11964 3690 11998 3706
rect 12082 4082 12116 4098
rect 12082 3690 12116 3706
rect 12200 4082 12234 4098
rect 12200 3690 12234 3706
rect 12318 4082 12352 4098
rect 12318 3690 12352 3706
rect 12436 4082 12470 4098
rect 12436 3690 12470 3706
rect 12554 4082 12588 4098
rect 12554 3690 12588 3706
rect 12672 4082 12706 4098
rect 12672 3690 12706 3706
rect 13132 4082 13166 4098
rect 13132 3690 13166 3706
rect 13250 4082 13284 4098
rect 13250 3690 13284 3706
rect 13368 4082 13402 4098
rect 13368 3690 13402 3706
rect 13486 4082 13520 4098
rect 13486 3690 13520 3706
rect 13604 4082 13638 4098
rect 13604 3690 13638 3706
rect 13722 4082 13756 4098
rect 13722 3690 13756 3706
rect 13840 4082 13874 4098
rect 13840 3690 13874 3706
rect 14300 4080 14334 4096
rect 14300 3688 14334 3704
rect 14418 4080 14452 4096
rect 14418 3688 14452 3704
rect 14536 4080 14570 4096
rect 14536 3688 14570 3704
rect 14654 4080 14688 4096
rect 14654 3688 14688 3704
rect 14772 4080 14806 4096
rect 14772 3688 14806 3704
rect 14890 4080 14924 4096
rect 14890 3688 14924 3704
rect 15008 4080 15042 4096
rect 15008 3688 15042 3704
rect 15468 4082 15502 4098
rect 15468 3690 15502 3706
rect 15586 4082 15620 4098
rect 15586 3690 15620 3706
rect 15704 4082 15738 4098
rect 15704 3690 15738 3706
rect 15822 4082 15856 4098
rect 15822 3690 15856 3706
rect 15940 4082 15974 4098
rect 15940 3690 15974 3706
rect 16058 4082 16092 4098
rect 16058 3690 16092 3706
rect 16176 4082 16210 4098
rect 16176 3690 16210 3706
rect 16642 4084 16676 4100
rect 16642 3692 16676 3708
rect 16760 4084 16794 4100
rect 16760 3692 16794 3708
rect 16878 4084 16912 4100
rect 16878 3692 16912 3708
rect 16996 4084 17030 4100
rect 16996 3692 17030 3708
rect 17114 4084 17148 4100
rect 17114 3692 17148 3708
rect 17232 4084 17266 4100
rect 17232 3692 17266 3708
rect 17350 4084 17384 4100
rect 17350 3692 17384 3708
rect 17810 4082 17844 4098
rect 17810 3690 17844 3706
rect 17928 4082 17962 4098
rect 17928 3690 17962 3706
rect 18046 4082 18080 4098
rect 18046 3690 18080 3706
rect 18164 4082 18198 4098
rect 18164 3690 18198 3706
rect 18282 4082 18316 4098
rect 18282 3690 18316 3706
rect 18400 4082 18434 4098
rect 18400 3690 18434 3706
rect 18518 4082 18552 4098
rect 18518 3690 18552 3706
rect 18978 4084 19012 4100
rect 18978 3692 19012 3708
rect 19096 4084 19130 4100
rect 19096 3692 19130 3708
rect 19214 4084 19248 4100
rect 19214 3692 19248 3708
rect 19332 4084 19366 4100
rect 19332 3692 19366 3708
rect 19450 4084 19484 4100
rect 19450 3692 19484 3708
rect 19568 4084 19602 4100
rect 19568 3692 19602 3708
rect 19686 4084 19720 4100
rect 19686 3692 19720 3708
rect 20146 4082 20180 4098
rect 20146 3690 20180 3706
rect 20264 4082 20298 4098
rect 20264 3690 20298 3706
rect 20382 4082 20416 4098
rect 20382 3690 20416 3706
rect 20500 4082 20534 4098
rect 20500 3690 20534 3706
rect 20618 4082 20652 4098
rect 20618 3690 20652 3706
rect 20736 4082 20770 4098
rect 20736 3690 20770 3706
rect 20854 4082 20888 4098
rect 20854 3690 20888 3706
rect 952 3615 968 3649
rect 1002 3615 1018 3649
rect 2400 3615 2416 3649
rect 2450 3615 2466 3649
rect 3898 3617 3914 3651
rect 3948 3617 3964 3651
rect 5346 3617 5362 3651
rect 5396 3617 5412 3651
rect 6866 3615 6882 3649
rect 6916 3615 6932 3649
rect 8314 3615 8330 3649
rect 8364 3615 8380 3649
rect 9812 3617 9828 3651
rect 9862 3617 9878 3651
rect 11260 3617 11276 3651
rect 11310 3617 11326 3651
rect 834 3498 850 3532
rect 884 3498 900 3532
rect 2282 3498 2298 3532
rect 2332 3498 2348 3532
rect 3780 3500 3796 3534
rect 3830 3500 3846 3534
rect 5228 3500 5244 3534
rect 5278 3500 5294 3534
rect 6748 3498 6764 3532
rect 6798 3498 6814 3532
rect 8196 3498 8212 3532
rect 8246 3498 8262 3532
rect 9694 3500 9710 3534
rect 9744 3500 9760 3534
rect 11142 3500 11158 3534
rect 11192 3500 11208 3534
rect 438 3448 472 3464
rect 438 3056 472 3072
rect 556 3448 590 3464
rect 556 3056 590 3072
rect 674 3448 708 3464
rect 791 3448 825 3464
rect 791 3256 825 3272
rect 909 3448 943 3464
rect 909 3256 943 3272
rect 1886 3448 1920 3464
rect 674 3056 708 3072
rect 1886 3056 1920 3072
rect 2004 3448 2038 3464
rect 2004 3056 2038 3072
rect 2122 3448 2156 3464
rect 2239 3448 2273 3464
rect 2239 3256 2273 3272
rect 2357 3448 2391 3464
rect 2357 3256 2391 3272
rect 3384 3450 3418 3466
rect 2122 3056 2156 3072
rect 3384 3058 3418 3074
rect 3502 3450 3536 3466
rect 3502 3058 3536 3074
rect 3620 3450 3654 3466
rect 3737 3450 3771 3466
rect 3737 3258 3771 3274
rect 3855 3450 3889 3466
rect 3855 3258 3889 3274
rect 4832 3450 4866 3466
rect 3620 3058 3654 3074
rect 4832 3058 4866 3074
rect 4950 3450 4984 3466
rect 4950 3058 4984 3074
rect 5068 3450 5102 3466
rect 5185 3450 5219 3466
rect 5185 3258 5219 3274
rect 5303 3450 5337 3466
rect 5303 3258 5337 3274
rect 6352 3448 6386 3464
rect 5068 3058 5102 3074
rect 6352 3056 6386 3072
rect 6470 3448 6504 3464
rect 6470 3056 6504 3072
rect 6588 3448 6622 3464
rect 6705 3448 6739 3464
rect 6705 3256 6739 3272
rect 6823 3448 6857 3464
rect 6823 3256 6857 3272
rect 7800 3448 7834 3464
rect 6588 3056 6622 3072
rect 7800 3056 7834 3072
rect 7918 3448 7952 3464
rect 7918 3056 7952 3072
rect 8036 3448 8070 3464
rect 8153 3448 8187 3464
rect 8153 3256 8187 3272
rect 8271 3448 8305 3464
rect 8271 3256 8305 3272
rect 9298 3450 9332 3466
rect 8036 3056 8070 3072
rect 9298 3058 9332 3074
rect 9416 3450 9450 3466
rect 9416 3058 9450 3074
rect 9534 3450 9568 3466
rect 9651 3450 9685 3466
rect 9651 3258 9685 3274
rect 9769 3450 9803 3466
rect 9769 3258 9803 3274
rect 10746 3450 10780 3466
rect 9534 3058 9568 3074
rect 10746 3058 10780 3074
rect 10864 3450 10898 3466
rect 10864 3058 10898 3074
rect 10982 3450 11016 3466
rect 11099 3450 11133 3466
rect 11099 3258 11133 3274
rect 11217 3450 11251 3466
rect 15248 3420 16048 3454
rect 12153 3349 12169 3383
rect 12203 3349 12219 3383
rect 13321 3349 13337 3383
rect 13371 3349 13387 3383
rect 14489 3349 14505 3383
rect 14539 3349 14555 3383
rect 11217 3258 11251 3274
rect 11874 3296 11908 3312
rect 11874 3104 11908 3120
rect 11992 3296 12026 3312
rect 11992 3104 12026 3120
rect 12110 3296 12144 3312
rect 12110 3104 12144 3120
rect 12228 3296 12262 3312
rect 12228 3104 12262 3120
rect 12394 3292 12428 3308
rect 10982 3058 11016 3074
rect 481 2988 497 3022
rect 531 2988 547 3022
rect 599 2988 615 3022
rect 649 2988 665 3022
rect 1929 2988 1945 3022
rect 1979 2988 1995 3022
rect 2047 2988 2063 3022
rect 2097 2988 2113 3022
rect 3427 2990 3443 3024
rect 3477 2990 3493 3024
rect 3545 2990 3561 3024
rect 3595 2990 3611 3024
rect 4875 2990 4891 3024
rect 4925 2990 4941 3024
rect 4993 2990 5009 3024
rect 5043 2990 5059 3024
rect 6395 2988 6411 3022
rect 6445 2988 6461 3022
rect 6513 2988 6529 3022
rect 6563 2988 6579 3022
rect 7843 2988 7859 3022
rect 7893 2988 7909 3022
rect 7961 2988 7977 3022
rect 8011 2988 8027 3022
rect 9341 2990 9357 3024
rect 9391 2990 9407 3024
rect 9459 2990 9475 3024
rect 9509 2990 9525 3024
rect 10789 2990 10805 3024
rect 10839 2990 10855 3024
rect 10907 2990 10923 3024
rect 10957 2990 10973 3024
rect 12394 3016 12428 3116
rect 12512 3292 12546 3308
rect 12512 3100 12546 3116
rect 12630 3292 12664 3308
rect 12630 3016 12664 3116
rect 12748 3292 12782 3308
rect 12748 3100 12782 3116
rect 13042 3298 13076 3314
rect 13042 3106 13076 3122
rect 13160 3298 13194 3314
rect 13160 3106 13194 3122
rect 13278 3298 13312 3314
rect 13278 3106 13312 3122
rect 13396 3298 13430 3314
rect 13396 3106 13430 3122
rect 13561 3298 13595 3314
rect 12018 2992 12160 3004
rect 12018 2988 12058 2992
rect 12124 2988 12160 2992
rect 714 2917 882 2935
rect 714 2861 730 2917
rect 864 2861 882 2917
rect 714 2845 882 2861
rect 2162 2917 2330 2935
rect 2162 2861 2178 2917
rect 2312 2861 2330 2917
rect 2162 2845 2330 2861
rect 3660 2919 3828 2937
rect 3660 2863 3676 2919
rect 3810 2863 3828 2919
rect 3660 2847 3828 2863
rect 5108 2919 5276 2937
rect 5108 2863 5124 2919
rect 5258 2863 5276 2919
rect 5108 2847 5276 2863
rect 6628 2917 6796 2935
rect 6628 2861 6644 2917
rect 6778 2861 6796 2917
rect 6628 2845 6796 2861
rect 8076 2917 8244 2935
rect 8076 2861 8092 2917
rect 8226 2861 8244 2917
rect 8076 2845 8244 2861
rect 9574 2919 9742 2937
rect 9574 2863 9590 2919
rect 9724 2863 9742 2919
rect 9574 2847 9742 2863
rect 11022 2919 11190 2937
rect 11022 2863 11038 2919
rect 11172 2863 11190 2919
rect 12018 2922 12036 2988
rect 12154 2922 12160 2988
rect 12394 2982 12664 3016
rect 13561 3028 13595 3122
rect 13679 3298 13713 3314
rect 13679 3106 13713 3122
rect 13797 3298 13831 3314
rect 13797 3028 13831 3122
rect 13915 3298 13949 3314
rect 13915 3106 13949 3122
rect 14210 3298 14244 3314
rect 14210 3106 14244 3122
rect 14328 3298 14362 3314
rect 14328 3106 14362 3122
rect 14446 3298 14480 3314
rect 14446 3106 14480 3122
rect 14564 3298 14598 3314
rect 14564 3106 14598 3122
rect 14729 3298 14763 3314
rect 13186 2992 13328 3004
rect 13561 2994 13831 3028
rect 14729 3011 14763 3122
rect 14847 3298 14881 3314
rect 14847 3106 14881 3122
rect 14965 3298 14999 3314
rect 14965 3011 14999 3122
rect 15083 3298 15117 3314
rect 15083 3106 15117 3122
rect 13186 2988 13226 2992
rect 13292 2988 13328 2992
rect 12018 2896 12160 2922
rect 11022 2847 11190 2863
rect 12486 2809 12531 2982
rect 13186 2922 13204 2988
rect 13322 2922 13328 2988
rect 13186 2896 13328 2922
rect -134 2755 12531 2809
rect -134 1608 -42 2755
rect 13679 2721 13713 2994
rect 14354 2992 14496 3004
rect 14354 2988 14394 2992
rect 14460 2988 14496 2992
rect 14354 2922 14372 2988
rect 14490 2922 14496 2988
rect 14729 2975 14999 3011
rect 14354 2896 14496 2922
rect 3089 2667 13713 2721
rect 1430 2398 1658 2416
rect 1430 2322 1446 2398
rect 1642 2322 1658 2398
rect 1430 2306 1658 2322
rect 701 2181 971 2220
rect 701 2128 735 2181
rect 260 1979 530 2018
rect 260 1928 294 1979
rect 260 1736 294 1752
rect 378 1928 412 1944
rect 378 1701 412 1752
rect 496 1928 530 1979
rect 496 1736 530 1752
rect 614 1928 648 1944
rect 614 1701 648 1752
rect 701 1736 735 1752
rect 819 2128 853 2144
rect 378 1662 648 1701
rect 819 1701 853 1752
rect 937 2128 971 2181
rect 1168 2180 1438 2219
rect 937 1736 971 1752
rect 1055 2128 1089 2144
rect 1055 1701 1089 1752
rect 1168 2128 1202 2180
rect 1168 1736 1202 1752
rect 1286 2128 1320 2144
rect 1286 1701 1320 1752
rect 1404 2128 1438 2180
rect 1640 2180 1910 2219
rect 1404 1736 1438 1752
rect 1522 2128 1556 2144
rect 1522 1701 1556 1752
rect 1640 2128 1674 2180
rect 1640 1736 1674 1752
rect 1758 2128 1792 2144
rect 1758 1701 1792 1752
rect 1876 2128 1910 2180
rect 2113 2180 2383 2219
rect 1876 1736 1910 1752
rect 1995 2128 2029 2144
rect 1995 1701 2029 1752
rect 2113 2128 2147 2180
rect 2113 1736 2147 1752
rect 2231 2128 2265 2144
rect 2231 1701 2265 1752
rect 2349 2128 2383 2180
rect 2586 1978 2856 2015
rect 2349 1736 2383 1752
rect 2468 1928 2502 1944
rect 819 1662 2265 1701
rect 2468 1698 2502 1752
rect 2586 1928 2620 1978
rect 2586 1736 2620 1752
rect 2704 1928 2738 1944
rect 2704 1698 2738 1752
rect 2822 1928 2856 1978
rect 2822 1736 2856 1752
rect 2468 1659 2738 1698
rect -134 1167 -41 1608
rect 1346 1537 1380 1553
rect 2640 1544 2656 1578
rect 2690 1544 2706 1578
rect 1346 1487 1380 1503
rect 349 1437 441 1454
rect 349 1382 365 1437
rect 425 1382 441 1437
rect 349 1369 441 1382
rect 1434 1438 1526 1451
rect 1434 1383 1450 1438
rect 1510 1383 1526 1438
rect 1434 1366 1526 1383
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 1700 1307 1734 1323
rect 1700 1257 1734 1273
rect -134 1154 177 1167
rect -134 1094 121 1154
rect 170 1094 177 1154
rect -134 1081 177 1094
rect 1316 1153 1408 1166
rect 1316 1098 1332 1153
rect 1392 1098 1408 1153
rect 1316 1081 1408 1098
rect 3089 1158 3167 2667
rect 14815 2633 14864 2975
rect 6213 2585 14864 2633
rect 4574 2398 4802 2416
rect 4574 2322 4590 2398
rect 4786 2322 4802 2398
rect 4574 2306 4802 2322
rect 3845 2181 4115 2220
rect 3845 2128 3879 2181
rect 3404 1979 3674 2018
rect 3404 1928 3438 1979
rect 3404 1736 3438 1752
rect 3522 1928 3556 1944
rect 3522 1701 3556 1752
rect 3640 1928 3674 1979
rect 3640 1736 3674 1752
rect 3758 1928 3792 1944
rect 3758 1701 3792 1752
rect 3845 1736 3879 1752
rect 3963 2128 3997 2144
rect 3522 1662 3792 1701
rect 3963 1701 3997 1752
rect 4081 2128 4115 2181
rect 4312 2180 4582 2219
rect 4081 1736 4115 1752
rect 4199 2128 4233 2144
rect 4199 1701 4233 1752
rect 4312 2128 4346 2180
rect 4312 1736 4346 1752
rect 4430 2128 4464 2144
rect 4430 1701 4464 1752
rect 4548 2128 4582 2180
rect 4784 2180 5054 2219
rect 4548 1736 4582 1752
rect 4666 2128 4700 2144
rect 4666 1701 4700 1752
rect 4784 2128 4818 2180
rect 4784 1736 4818 1752
rect 4902 2128 4936 2144
rect 4902 1701 4936 1752
rect 5020 2128 5054 2180
rect 5257 2180 5527 2219
rect 5020 1736 5054 1752
rect 5139 2128 5173 2144
rect 5139 1701 5173 1752
rect 5257 2128 5291 2180
rect 5257 1736 5291 1752
rect 5375 2128 5409 2144
rect 5375 1701 5409 1752
rect 5493 2128 5527 2180
rect 5730 1978 6000 2015
rect 5493 1736 5527 1752
rect 5612 1928 5646 1944
rect 3963 1662 5409 1701
rect 5612 1698 5646 1752
rect 5730 1928 5764 1978
rect 5730 1736 5764 1752
rect 5848 1928 5882 1944
rect 5848 1698 5882 1752
rect 5966 1928 6000 1978
rect 5966 1736 6000 1752
rect 5612 1659 5882 1698
rect 4490 1537 4524 1553
rect 5784 1544 5800 1578
rect 5834 1544 5850 1578
rect 4490 1487 4524 1503
rect 3493 1437 3585 1454
rect 3493 1382 3509 1437
rect 3569 1382 3585 1437
rect 3493 1369 3585 1382
rect 4578 1438 4670 1451
rect 4578 1383 4594 1438
rect 4654 1383 4670 1438
rect 4578 1366 4670 1383
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 4844 1307 4878 1323
rect 4844 1257 4878 1273
rect 3089 1154 3318 1158
rect 3089 1094 3265 1154
rect 3314 1094 3318 1154
rect 3089 1090 3318 1094
rect 4460 1153 4552 1166
rect 4460 1098 4476 1153
rect 4536 1098 4552 1153
rect 4460 1081 4552 1098
rect 6213 1162 6281 2585
rect 15248 2551 15321 3420
rect 15657 3349 15673 3383
rect 15707 3349 15723 3383
rect 16014 3382 16048 3420
rect 15898 3348 16168 3382
rect 16831 3351 16847 3385
rect 16881 3351 16897 3385
rect 17999 3351 18015 3385
rect 18049 3351 18065 3385
rect 19167 3351 19183 3385
rect 19217 3351 19233 3385
rect 20335 3351 20351 3385
rect 20385 3351 20401 3385
rect 15378 3298 15412 3314
rect 15378 3106 15412 3122
rect 15496 3298 15530 3314
rect 15496 3106 15530 3122
rect 15614 3298 15648 3314
rect 15614 3106 15648 3122
rect 15732 3298 15766 3314
rect 15732 3106 15766 3122
rect 15898 3298 15932 3348
rect 15898 3106 15932 3122
rect 16016 3298 16050 3314
rect 16016 3106 16050 3122
rect 16134 3298 16168 3348
rect 16134 3106 16168 3122
rect 16252 3298 16286 3314
rect 16252 3106 16286 3122
rect 16552 3298 16586 3314
rect 16552 3106 16586 3122
rect 16670 3298 16704 3314
rect 16670 3106 16704 3122
rect 16788 3298 16822 3314
rect 16788 3106 16822 3122
rect 16906 3298 16940 3314
rect 16906 3106 16940 3122
rect 17070 3294 17104 3310
rect 17070 3018 17104 3118
rect 17188 3294 17222 3310
rect 17188 3102 17222 3118
rect 17306 3294 17340 3310
rect 17306 3018 17340 3118
rect 17424 3294 17458 3310
rect 17424 3102 17458 3118
rect 17720 3298 17754 3314
rect 17720 3106 17754 3122
rect 17838 3298 17872 3314
rect 17838 3106 17872 3122
rect 17956 3298 17990 3314
rect 17956 3106 17990 3122
rect 18074 3298 18108 3314
rect 18074 3106 18108 3122
rect 18239 3293 18273 3309
rect 15522 2992 15664 3004
rect 15522 2988 15562 2992
rect 15628 2988 15664 2992
rect 15522 2922 15540 2988
rect 15658 2922 15664 2988
rect 15522 2896 15664 2922
rect 16696 2994 16838 3006
rect 16696 2990 16736 2994
rect 16802 2990 16838 2994
rect 16696 2924 16714 2990
rect 16832 2924 16838 2990
rect 17070 2983 17340 3018
rect 18239 3032 18273 3117
rect 18357 3293 18391 3309
rect 18357 3101 18391 3117
rect 18475 3293 18509 3309
rect 18475 3032 18509 3117
rect 18593 3293 18627 3309
rect 18593 3101 18627 3117
rect 18888 3300 18922 3316
rect 18888 3108 18922 3124
rect 19006 3300 19040 3316
rect 19006 3108 19040 3124
rect 19124 3300 19158 3316
rect 19124 3108 19158 3124
rect 19242 3300 19276 3316
rect 19242 3108 19276 3124
rect 19407 3293 19441 3309
rect 17864 2994 18006 3006
rect 18239 2997 18509 3032
rect 19407 3032 19441 3117
rect 19525 3293 19559 3309
rect 19525 3101 19559 3117
rect 19643 3293 19677 3309
rect 19643 3032 19677 3117
rect 19761 3293 19795 3309
rect 19761 3101 19795 3117
rect 20056 3300 20090 3316
rect 20056 3108 20090 3124
rect 20174 3300 20208 3316
rect 20174 3108 20208 3124
rect 20292 3300 20326 3316
rect 20292 3108 20326 3124
rect 20410 3300 20444 3316
rect 20410 3108 20444 3124
rect 20575 3294 20609 3310
rect 17864 2990 17904 2994
rect 17970 2990 18006 2994
rect 16696 2898 16838 2924
rect 17192 2750 17250 2983
rect 17864 2924 17882 2990
rect 18000 2924 18006 2990
rect 17864 2898 18006 2924
rect 12329 2497 15321 2551
rect 15541 2691 17250 2750
rect 7706 2402 7934 2420
rect 7706 2326 7722 2402
rect 7918 2326 7934 2402
rect 7706 2310 7934 2326
rect 10850 2402 11078 2420
rect 10850 2326 10866 2402
rect 11062 2326 11078 2402
rect 10850 2310 11078 2326
rect 6977 2185 7247 2224
rect 6977 2132 7011 2185
rect 6536 1983 6806 2022
rect 6536 1932 6570 1983
rect 6536 1740 6570 1756
rect 6654 1932 6688 1948
rect 6654 1705 6688 1756
rect 6772 1932 6806 1983
rect 6772 1740 6806 1756
rect 6890 1932 6924 1948
rect 6890 1705 6924 1756
rect 6977 1740 7011 1756
rect 7095 2132 7129 2148
rect 6654 1666 6924 1705
rect 7095 1705 7129 1756
rect 7213 2132 7247 2185
rect 7444 2184 7714 2223
rect 7213 1740 7247 1756
rect 7331 2132 7365 2148
rect 7331 1705 7365 1756
rect 7444 2132 7478 2184
rect 7444 1740 7478 1756
rect 7562 2132 7596 2148
rect 7562 1705 7596 1756
rect 7680 2132 7714 2184
rect 7916 2184 8186 2223
rect 7680 1740 7714 1756
rect 7798 2132 7832 2148
rect 7798 1705 7832 1756
rect 7916 2132 7950 2184
rect 7916 1740 7950 1756
rect 8034 2132 8068 2148
rect 8034 1705 8068 1756
rect 8152 2132 8186 2184
rect 8389 2184 8659 2223
rect 8152 1740 8186 1756
rect 8271 2132 8305 2148
rect 8271 1705 8305 1756
rect 8389 2132 8423 2184
rect 8389 1740 8423 1756
rect 8507 2132 8541 2148
rect 8507 1705 8541 1756
rect 8625 2132 8659 2184
rect 10121 2185 10391 2224
rect 10121 2132 10155 2185
rect 8862 1982 9132 2019
rect 8625 1740 8659 1756
rect 8744 1932 8778 1948
rect 7095 1666 8541 1705
rect 8744 1702 8778 1756
rect 8862 1932 8896 1982
rect 8862 1740 8896 1756
rect 8980 1932 9014 1948
rect 8980 1702 9014 1756
rect 9098 1932 9132 1982
rect 9098 1740 9132 1756
rect 9680 1983 9950 2022
rect 9680 1932 9714 1983
rect 9680 1740 9714 1756
rect 9798 1932 9832 1948
rect 8744 1663 9014 1702
rect 9798 1705 9832 1756
rect 9916 1932 9950 1983
rect 9916 1740 9950 1756
rect 10034 1932 10068 1948
rect 10034 1705 10068 1756
rect 10121 1740 10155 1756
rect 10239 2132 10273 2148
rect 9798 1666 10068 1705
rect 10239 1705 10273 1756
rect 10357 2132 10391 2185
rect 10588 2184 10858 2223
rect 10357 1740 10391 1756
rect 10475 2132 10509 2148
rect 10475 1705 10509 1756
rect 10588 2132 10622 2184
rect 10588 1740 10622 1756
rect 10706 2132 10740 2148
rect 10706 1705 10740 1756
rect 10824 2132 10858 2184
rect 11060 2184 11330 2223
rect 10824 1740 10858 1756
rect 10942 2132 10976 2148
rect 10942 1705 10976 1756
rect 11060 2132 11094 2184
rect 11060 1740 11094 1756
rect 11178 2132 11212 2148
rect 11178 1705 11212 1756
rect 11296 2132 11330 2184
rect 11533 2184 11803 2223
rect 11296 1740 11330 1756
rect 11415 2132 11449 2148
rect 11415 1705 11449 1756
rect 11533 2132 11567 2184
rect 11533 1740 11567 1756
rect 11651 2132 11685 2148
rect 11651 1705 11685 1756
rect 11769 2132 11803 2184
rect 12006 1982 12276 2019
rect 11769 1740 11803 1756
rect 11888 1932 11922 1948
rect 10239 1666 11685 1705
rect 11888 1702 11922 1756
rect 12006 1932 12040 1982
rect 12006 1740 12040 1756
rect 12124 1932 12158 1948
rect 12124 1702 12158 1756
rect 12242 1932 12276 1982
rect 12242 1740 12276 1756
rect 11888 1663 12158 1702
rect 7622 1541 7656 1557
rect 8916 1548 8932 1582
rect 8966 1548 8982 1582
rect 7622 1491 7656 1507
rect 10766 1541 10800 1557
rect 12060 1548 12076 1582
rect 12110 1548 12126 1582
rect 10766 1491 10800 1507
rect 6625 1441 6717 1458
rect 6625 1386 6641 1441
rect 6701 1386 6717 1441
rect 6625 1373 6717 1386
rect 7710 1442 7802 1455
rect 7710 1387 7726 1442
rect 7786 1387 7802 1442
rect 7710 1370 7802 1387
rect 9769 1441 9861 1458
rect 9769 1386 9785 1441
rect 9845 1386 9861 1441
rect 9769 1373 9861 1386
rect 10854 1442 10946 1455
rect 10854 1387 10870 1442
rect 10930 1387 10946 1442
rect 10854 1370 10946 1387
rect 6393 1326 6450 1330
rect 6393 1266 6397 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 7976 1311 8010 1327
rect 7976 1261 8010 1277
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 11120 1311 11154 1327
rect 11120 1261 11154 1277
rect 6213 1158 6451 1162
rect 6213 1098 6397 1158
rect 6446 1098 6451 1158
rect 6213 1093 6451 1098
rect 7592 1157 7684 1170
rect 7592 1102 7608 1157
rect 7668 1102 7684 1157
rect 7592 1085 7684 1102
rect 10736 1163 10828 1170
rect 12329 1163 12401 2497
rect 14052 2398 14280 2416
rect 14052 2322 14068 2398
rect 14264 2322 14280 2398
rect 14052 2306 14280 2322
rect 13323 2181 13593 2220
rect 13323 2128 13357 2181
rect 12882 1979 13152 2018
rect 12882 1928 12916 1979
rect 12882 1736 12916 1752
rect 13000 1928 13034 1944
rect 13000 1701 13034 1752
rect 13118 1928 13152 1979
rect 13118 1736 13152 1752
rect 13236 1928 13270 1944
rect 13236 1701 13270 1752
rect 13323 1736 13357 1752
rect 13441 2128 13475 2144
rect 13000 1662 13270 1701
rect 13441 1701 13475 1752
rect 13559 2128 13593 2181
rect 13790 2180 14060 2219
rect 13559 1736 13593 1752
rect 13677 2128 13711 2144
rect 13677 1701 13711 1752
rect 13790 2128 13824 2180
rect 13790 1736 13824 1752
rect 13908 2128 13942 2144
rect 13908 1701 13942 1752
rect 14026 2128 14060 2180
rect 14262 2180 14532 2219
rect 14026 1736 14060 1752
rect 14144 2128 14178 2144
rect 14144 1701 14178 1752
rect 14262 2128 14296 2180
rect 14262 1736 14296 1752
rect 14380 2128 14414 2144
rect 14380 1701 14414 1752
rect 14498 2128 14532 2180
rect 14735 2180 15005 2219
rect 14498 1736 14532 1752
rect 14617 2128 14651 2144
rect 14617 1701 14651 1752
rect 14735 2128 14769 2180
rect 14735 1736 14769 1752
rect 14853 2128 14887 2144
rect 14853 1701 14887 1752
rect 14971 2128 15005 2180
rect 15208 1978 15478 2015
rect 14971 1736 15005 1752
rect 15090 1928 15124 1944
rect 13441 1662 14887 1701
rect 15090 1698 15124 1752
rect 15208 1928 15242 1978
rect 15208 1736 15242 1752
rect 15326 1928 15360 1944
rect 15326 1698 15360 1752
rect 15444 1928 15478 1978
rect 15444 1736 15478 1752
rect 15090 1659 15360 1698
rect 13968 1537 14002 1553
rect 15262 1544 15278 1578
rect 15312 1544 15328 1578
rect 13968 1487 14002 1503
rect 12971 1437 13063 1454
rect 12971 1382 12987 1437
rect 13047 1382 13063 1437
rect 12971 1369 13063 1382
rect 14056 1438 14148 1451
rect 14056 1383 14072 1438
rect 14132 1383 14148 1438
rect 14056 1366 14148 1383
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 14322 1307 14356 1323
rect 14322 1257 14356 1273
rect 10736 1157 12401 1163
rect 10736 1102 10754 1157
rect 10812 1102 12401 1157
rect 10736 1092 12401 1102
rect 13938 1158 14030 1166
rect 15541 1158 15620 2691
rect 18344 2655 18411 2997
rect 19032 2994 19174 3006
rect 19407 2997 19677 3032
rect 20575 3027 20609 3118
rect 20693 3294 20727 3310
rect 20693 3102 20727 3118
rect 20811 3294 20845 3310
rect 20811 3027 20845 3118
rect 20929 3294 20963 3310
rect 20929 3102 20963 3118
rect 19032 2990 19072 2994
rect 19138 2990 19174 2994
rect 19032 2924 19050 2990
rect 19168 2924 19174 2990
rect 19032 2898 19174 2924
rect 13938 1153 15620 1158
rect 13938 1098 13956 1153
rect 14014 1098 15620 1153
rect 10736 1085 10828 1092
rect 13938 1087 15620 1098
rect 15694 2591 18411 2655
rect 19521 2632 19564 2997
rect 20200 2994 20342 3006
rect 20200 2990 20240 2994
rect 20306 2990 20342 2994
rect 20575 2990 22009 3027
rect 20200 2924 20218 2990
rect 20336 2924 20342 2990
rect 20200 2898 20342 2924
rect 15694 1158 15762 2591
rect 18823 2573 19564 2632
rect 17196 2398 17424 2416
rect 17196 2322 17212 2398
rect 17408 2322 17424 2398
rect 17196 2306 17424 2322
rect 16467 2181 16737 2220
rect 16467 2128 16501 2181
rect 16026 1979 16296 2018
rect 16026 1928 16060 1979
rect 16026 1736 16060 1752
rect 16144 1928 16178 1944
rect 16144 1701 16178 1752
rect 16262 1928 16296 1979
rect 16262 1736 16296 1752
rect 16380 1928 16414 1944
rect 16380 1701 16414 1752
rect 16467 1736 16501 1752
rect 16585 2128 16619 2144
rect 16144 1662 16414 1701
rect 16585 1701 16619 1752
rect 16703 2128 16737 2181
rect 16934 2180 17204 2219
rect 16703 1736 16737 1752
rect 16821 2128 16855 2144
rect 16821 1701 16855 1752
rect 16934 2128 16968 2180
rect 16934 1736 16968 1752
rect 17052 2128 17086 2144
rect 17052 1701 17086 1752
rect 17170 2128 17204 2180
rect 17406 2180 17676 2219
rect 17170 1736 17204 1752
rect 17288 2128 17322 2144
rect 17288 1701 17322 1752
rect 17406 2128 17440 2180
rect 17406 1736 17440 1752
rect 17524 2128 17558 2144
rect 17524 1701 17558 1752
rect 17642 2128 17676 2180
rect 17879 2180 18149 2219
rect 17642 1736 17676 1752
rect 17761 2128 17795 2144
rect 17761 1701 17795 1752
rect 17879 2128 17913 2180
rect 17879 1736 17913 1752
rect 17997 2128 18031 2144
rect 17997 1701 18031 1752
rect 18115 2128 18149 2180
rect 18352 1978 18622 2015
rect 18115 1736 18149 1752
rect 18234 1928 18268 1944
rect 16585 1662 18031 1701
rect 18234 1698 18268 1752
rect 18352 1928 18386 1978
rect 18352 1736 18386 1752
rect 18470 1928 18504 1944
rect 18470 1698 18504 1752
rect 18588 1928 18622 1978
rect 18588 1736 18622 1752
rect 18234 1659 18504 1698
rect 17112 1537 17146 1553
rect 18406 1544 18422 1578
rect 18456 1544 18472 1578
rect 17112 1487 17146 1503
rect 18823 1520 18890 2573
rect 20328 2402 20556 2420
rect 20328 2326 20344 2402
rect 20540 2326 20556 2402
rect 20328 2310 20556 2326
rect 19599 2185 19869 2224
rect 19599 2132 19633 2185
rect 19158 1983 19428 2022
rect 19158 1932 19192 1983
rect 19158 1740 19192 1756
rect 19276 1932 19310 1948
rect 19276 1705 19310 1756
rect 19394 1932 19428 1983
rect 19394 1740 19428 1756
rect 19512 1932 19546 1948
rect 19512 1705 19546 1756
rect 19599 1740 19633 1756
rect 19717 2132 19751 2148
rect 19276 1666 19546 1705
rect 19717 1705 19751 1756
rect 19835 2132 19869 2185
rect 20066 2184 20336 2223
rect 19835 1740 19869 1756
rect 19953 2132 19987 2148
rect 19953 1705 19987 1756
rect 20066 2132 20100 2184
rect 20066 1740 20100 1756
rect 20184 2132 20218 2148
rect 20184 1705 20218 1756
rect 20302 2132 20336 2184
rect 20538 2184 20808 2223
rect 20302 1740 20336 1756
rect 20420 2132 20454 2148
rect 20420 1705 20454 1756
rect 20538 2132 20572 2184
rect 20538 1740 20572 1756
rect 20656 2132 20690 2148
rect 20656 1705 20690 1756
rect 20774 2132 20808 2184
rect 21011 2184 21281 2223
rect 20774 1740 20808 1756
rect 20893 2132 20927 2148
rect 20893 1705 20927 1756
rect 21011 2132 21045 2184
rect 21011 1740 21045 1756
rect 21129 2132 21163 2148
rect 21129 1705 21163 1756
rect 21247 2132 21281 2184
rect 21484 1982 21754 2019
rect 21247 1740 21281 1756
rect 21366 1932 21400 1948
rect 19717 1666 21163 1705
rect 21366 1702 21400 1756
rect 21484 1932 21518 1982
rect 21484 1740 21518 1756
rect 21602 1932 21636 1948
rect 21602 1702 21636 1756
rect 21720 1932 21754 1982
rect 21720 1740 21754 1756
rect 21366 1663 21636 1702
rect 20244 1541 20278 1557
rect 21538 1548 21554 1582
rect 21588 1548 21604 1582
rect 16115 1437 16207 1454
rect 16115 1382 16131 1437
rect 16191 1382 16207 1437
rect 16115 1369 16207 1382
rect 17200 1438 17292 1451
rect 17200 1383 17216 1438
rect 17276 1383 17292 1438
rect 17200 1366 17292 1383
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 17466 1307 17500 1323
rect 17466 1257 17500 1273
rect 15694 1154 15940 1158
rect 15694 1094 15887 1154
rect 15936 1094 15940 1154
rect 15694 1090 15940 1094
rect 17082 1153 17174 1166
rect 17082 1098 17098 1153
rect 17158 1098 17174 1153
rect 13938 1081 14030 1087
rect 17082 1081 17174 1098
rect 18823 1161 18891 1520
rect 20244 1491 20278 1507
rect 19247 1441 19339 1458
rect 19247 1386 19263 1441
rect 19323 1386 19339 1441
rect 19247 1373 19339 1386
rect 20332 1442 20424 1455
rect 20332 1387 20348 1442
rect 20408 1387 20424 1442
rect 20332 1370 20424 1387
rect 19015 1326 19072 1330
rect 19015 1266 19019 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 20598 1311 20632 1327
rect 20598 1261 20632 1277
rect 19015 1161 19072 1162
rect 18823 1158 19072 1161
rect 18823 1098 19019 1158
rect 19068 1098 19072 1158
rect 18823 1094 19072 1098
rect 20214 1157 20306 1170
rect 20214 1102 20230 1157
rect 20290 1102 20306 1157
rect 18823 1093 19069 1094
rect 20214 1085 20306 1102
rect 21971 1162 22009 2990
rect 23472 2402 23700 2420
rect 23472 2326 23488 2402
rect 23684 2326 23700 2402
rect 23472 2310 23700 2326
rect 22743 2185 23013 2224
rect 22743 2132 22777 2185
rect 22302 1983 22572 2022
rect 22302 1932 22336 1983
rect 22302 1740 22336 1756
rect 22420 1932 22454 1948
rect 22420 1705 22454 1756
rect 22538 1932 22572 1983
rect 22538 1740 22572 1756
rect 22656 1932 22690 1948
rect 22656 1705 22690 1756
rect 22743 1740 22777 1756
rect 22861 2132 22895 2148
rect 22420 1666 22690 1705
rect 22861 1705 22895 1756
rect 22979 2132 23013 2185
rect 23210 2184 23480 2223
rect 22979 1740 23013 1756
rect 23097 2132 23131 2148
rect 23097 1705 23131 1756
rect 23210 2132 23244 2184
rect 23210 1740 23244 1756
rect 23328 2132 23362 2148
rect 23328 1705 23362 1756
rect 23446 2132 23480 2184
rect 23682 2184 23952 2223
rect 23446 1740 23480 1756
rect 23564 2132 23598 2148
rect 23564 1705 23598 1756
rect 23682 2132 23716 2184
rect 23682 1740 23716 1756
rect 23800 2132 23834 2148
rect 23800 1705 23834 1756
rect 23918 2132 23952 2184
rect 24155 2184 24425 2223
rect 23918 1740 23952 1756
rect 24037 2132 24071 2148
rect 24037 1705 24071 1756
rect 24155 2132 24189 2184
rect 24155 1740 24189 1756
rect 24273 2132 24307 2148
rect 24273 1705 24307 1756
rect 24391 2132 24425 2184
rect 24628 1982 24898 2019
rect 24391 1740 24425 1756
rect 24510 1932 24544 1948
rect 22861 1666 24307 1705
rect 24510 1702 24544 1756
rect 24628 1932 24662 1982
rect 24628 1740 24662 1756
rect 24746 1932 24780 1948
rect 24746 1702 24780 1756
rect 24864 1932 24898 1982
rect 24864 1740 24898 1756
rect 24510 1663 24780 1702
rect 23388 1541 23422 1557
rect 24682 1548 24698 1582
rect 24732 1548 24748 1582
rect 23388 1491 23422 1507
rect 22391 1441 22483 1458
rect 22391 1386 22407 1441
rect 22467 1386 22483 1441
rect 22391 1373 22483 1386
rect 23476 1442 23568 1455
rect 23476 1387 23492 1442
rect 23552 1387 23568 1442
rect 23476 1370 23568 1387
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 23742 1311 23776 1327
rect 23742 1261 23776 1277
rect 21971 1158 22225 1162
rect 21971 1098 22163 1158
rect 22212 1098 22225 1158
rect 21971 1094 22225 1098
rect 23358 1157 23450 1170
rect 23358 1102 23374 1157
rect 23434 1102 23450 1157
rect 23358 1085 23450 1102
rect 1581 917 1615 933
rect 1581 867 1615 883
rect 4725 917 4759 933
rect 4725 867 4759 883
rect 7857 921 7891 937
rect 7857 871 7891 887
rect 11001 921 11035 937
rect 11001 871 11035 887
rect 14203 917 14237 933
rect 14203 867 14237 883
rect 17347 917 17381 933
rect 17347 867 17381 883
rect 20479 921 20513 937
rect 20479 871 20513 887
rect 23623 921 23657 937
rect 23623 871 23657 887
rect 1094 795 1128 811
rect 1094 603 1128 619
rect 1212 807 1246 811
rect 1286 807 1320 811
rect 1212 795 1320 807
rect 1246 619 1286 795
rect 1212 607 1286 619
rect 1212 603 1246 607
rect 1286 403 1320 419
rect 1404 795 1438 811
rect 1404 403 1438 419
rect 1522 795 1556 811
rect 1522 403 1556 419
rect 1640 795 1674 811
rect 1640 403 1674 419
rect 1758 807 1792 811
rect 1836 807 1870 811
rect 1758 795 1870 807
rect 1792 619 1836 795
rect 1792 607 1870 619
rect 1836 603 1870 607
rect 1954 795 1988 811
rect 1954 603 1988 619
rect 4238 795 4272 811
rect 4238 603 4272 619
rect 4356 807 4390 811
rect 4430 807 4464 811
rect 4356 795 4464 807
rect 4390 619 4430 795
rect 4356 607 4430 619
rect 4356 603 4390 607
rect 1758 403 1792 419
rect 4430 403 4464 419
rect 4548 795 4582 811
rect 4548 403 4582 419
rect 4666 795 4700 811
rect 4666 403 4700 419
rect 4784 795 4818 811
rect 4784 403 4818 419
rect 4902 807 4936 811
rect 4980 807 5014 811
rect 4902 795 5014 807
rect 4936 619 4980 795
rect 4936 607 5014 619
rect 4980 603 5014 607
rect 5098 795 5132 811
rect 5098 603 5132 619
rect 7370 799 7404 815
rect 7370 607 7404 623
rect 7488 811 7522 815
rect 7562 811 7596 815
rect 7488 799 7596 811
rect 7522 623 7562 799
rect 7488 611 7562 623
rect 7488 607 7522 611
rect 4902 403 4936 419
rect 7562 407 7596 423
rect 7680 799 7714 815
rect 7680 407 7714 423
rect 7798 799 7832 815
rect 7798 407 7832 423
rect 7916 799 7950 815
rect 7916 407 7950 423
rect 8034 811 8068 815
rect 8112 811 8146 815
rect 8034 799 8146 811
rect 8068 623 8112 799
rect 8068 611 8146 623
rect 8112 607 8146 611
rect 8230 799 8264 815
rect 8230 607 8264 623
rect 10514 799 10548 815
rect 10514 607 10548 623
rect 10632 811 10666 815
rect 10706 811 10740 815
rect 10632 799 10740 811
rect 10666 623 10706 799
rect 10632 611 10706 623
rect 10632 607 10666 611
rect 8034 407 8068 423
rect 10706 407 10740 423
rect 10824 799 10858 815
rect 10824 407 10858 423
rect 10942 799 10976 815
rect 10942 407 10976 423
rect 11060 799 11094 815
rect 11060 407 11094 423
rect 11178 811 11212 815
rect 11256 811 11290 815
rect 11178 799 11290 811
rect 11212 623 11256 799
rect 11212 611 11290 623
rect 11256 607 11290 611
rect 11374 799 11408 815
rect 11374 607 11408 623
rect 13716 795 13750 811
rect 13716 603 13750 619
rect 13834 807 13868 811
rect 13908 807 13942 811
rect 13834 795 13942 807
rect 13868 619 13908 795
rect 13834 607 13908 619
rect 13834 603 13868 607
rect 11178 407 11212 423
rect 13908 403 13942 419
rect 14026 795 14060 811
rect 14026 403 14060 419
rect 14144 795 14178 811
rect 14144 403 14178 419
rect 14262 795 14296 811
rect 14262 403 14296 419
rect 14380 807 14414 811
rect 14458 807 14492 811
rect 14380 795 14492 807
rect 14414 619 14458 795
rect 14414 607 14492 619
rect 14458 603 14492 607
rect 14576 795 14610 811
rect 14576 603 14610 619
rect 16860 795 16894 811
rect 16860 603 16894 619
rect 16978 807 17012 811
rect 17052 807 17086 811
rect 16978 795 17086 807
rect 17012 619 17052 795
rect 16978 607 17052 619
rect 16978 603 17012 607
rect 14380 403 14414 419
rect 17052 403 17086 419
rect 17170 795 17204 811
rect 17170 403 17204 419
rect 17288 795 17322 811
rect 17288 403 17322 419
rect 17406 795 17440 811
rect 17406 403 17440 419
rect 17524 807 17558 811
rect 17602 807 17636 811
rect 17524 795 17636 807
rect 17558 619 17602 795
rect 17558 607 17636 619
rect 17602 603 17636 607
rect 17720 795 17754 811
rect 17720 603 17754 619
rect 19992 799 20026 815
rect 19992 607 20026 623
rect 20110 811 20144 815
rect 20184 811 20218 815
rect 20110 799 20218 811
rect 20144 623 20184 799
rect 20110 611 20184 623
rect 20110 607 20144 611
rect 17524 403 17558 419
rect 20184 407 20218 423
rect 20302 799 20336 815
rect 20302 407 20336 423
rect 20420 799 20454 815
rect 20420 407 20454 423
rect 20538 799 20572 815
rect 20538 407 20572 423
rect 20656 811 20690 815
rect 20734 811 20768 815
rect 20656 799 20768 811
rect 20690 623 20734 799
rect 20690 611 20768 623
rect 20734 607 20768 611
rect 20852 799 20886 815
rect 20852 607 20886 623
rect 23136 799 23170 815
rect 23136 607 23170 623
rect 23254 811 23288 815
rect 23328 811 23362 815
rect 23254 799 23362 811
rect 23288 623 23328 799
rect 23254 611 23328 623
rect 23254 607 23288 611
rect 20656 407 20690 423
rect 23328 407 23362 423
rect 23446 799 23480 815
rect 23446 407 23480 423
rect 23564 799 23598 815
rect 23564 407 23598 423
rect 23682 799 23716 815
rect 23682 407 23716 423
rect 23800 811 23834 815
rect 23878 811 23912 815
rect 23800 799 23912 811
rect 23834 623 23878 799
rect 23834 611 23912 623
rect 23878 607 23912 611
rect 23996 799 24030 815
rect 23996 607 24030 623
rect 23800 407 23834 423
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 7764 170 7900 174
rect 1488 166 1624 170
rect 1488 152 1526 166
rect 1584 152 1624 166
rect 1488 106 1504 152
rect 1608 106 1624 152
rect 1488 84 1624 106
rect 4632 166 4768 170
rect 4632 152 4670 166
rect 4728 152 4768 166
rect 4632 106 4648 152
rect 4752 106 4768 152
rect 4632 84 4768 106
rect 7764 156 7802 170
rect 7860 156 7900 170
rect 7764 110 7780 156
rect 7884 110 7900 156
rect 7764 88 7900 110
rect 10908 170 11044 174
rect 20386 170 20522 174
rect 10908 156 10946 170
rect 11004 156 11044 170
rect 10908 110 10924 156
rect 11028 110 11044 156
rect 10908 88 11044 110
rect 14110 166 14246 170
rect 14110 152 14148 166
rect 14206 152 14246 166
rect 14110 106 14126 152
rect 14230 106 14246 152
rect 14110 84 14246 106
rect 17254 166 17390 170
rect 17254 152 17292 166
rect 17350 152 17390 166
rect 17254 106 17270 152
rect 17374 106 17390 152
rect 17254 84 17390 106
rect 20386 156 20424 170
rect 20482 156 20522 170
rect 20386 110 20402 156
rect 20506 110 20522 156
rect 20386 88 20522 110
rect 23530 170 23666 174
rect 23530 156 23568 170
rect 23626 156 23666 170
rect 23530 110 23546 156
rect 23650 110 23666 156
rect 23530 88 23666 110
rect 1430 -336 1658 -318
rect 1430 -412 1446 -336
rect 1642 -412 1658 -336
rect 1430 -428 1658 -412
rect 4574 -336 4802 -318
rect 4574 -412 4590 -336
rect 4786 -412 4802 -336
rect 4574 -428 4802 -412
rect 7706 -332 7934 -314
rect 7706 -408 7722 -332
rect 7918 -408 7934 -332
rect 7706 -424 7934 -408
rect 10850 -332 11078 -314
rect 10850 -408 10866 -332
rect 11062 -408 11078 -332
rect 10850 -424 11078 -408
rect 14052 -336 14280 -318
rect 14052 -412 14068 -336
rect 14264 -412 14280 -336
rect 14052 -428 14280 -412
rect 17196 -336 17424 -318
rect 17196 -412 17212 -336
rect 17408 -412 17424 -336
rect 17196 -428 17424 -412
rect 20328 -332 20556 -314
rect 20328 -408 20344 -332
rect 20540 -408 20556 -332
rect 20328 -424 20556 -408
rect 23472 -332 23700 -314
rect 23472 -408 23488 -332
rect 23684 -408 23700 -332
rect 23472 -424 23700 -408
rect 701 -553 971 -514
rect 701 -606 735 -553
rect 260 -755 530 -716
rect 260 -806 294 -755
rect 260 -998 294 -982
rect 378 -806 412 -790
rect 378 -1033 412 -982
rect 496 -806 530 -755
rect 496 -998 530 -982
rect 614 -806 648 -790
rect 614 -1033 648 -982
rect 701 -998 735 -982
rect 819 -606 853 -590
rect 378 -1072 648 -1033
rect 819 -1033 853 -982
rect 937 -606 971 -553
rect 1168 -554 1438 -515
rect 937 -998 971 -982
rect 1055 -606 1089 -590
rect 1055 -1033 1089 -982
rect 1168 -606 1202 -554
rect 1168 -998 1202 -982
rect 1286 -606 1320 -590
rect 1286 -1033 1320 -982
rect 1404 -606 1438 -554
rect 1640 -554 1910 -515
rect 1404 -998 1438 -982
rect 1522 -606 1556 -590
rect 1522 -1033 1556 -982
rect 1640 -606 1674 -554
rect 1640 -998 1674 -982
rect 1758 -606 1792 -590
rect 1758 -1033 1792 -982
rect 1876 -606 1910 -554
rect 2113 -554 2383 -515
rect 1876 -998 1910 -982
rect 1995 -606 2029 -590
rect 1995 -1033 2029 -982
rect 2113 -606 2147 -554
rect 2113 -998 2147 -982
rect 2231 -606 2265 -590
rect 2231 -1033 2265 -982
rect 2349 -606 2383 -554
rect 3845 -553 4115 -514
rect 3845 -606 3879 -553
rect 2586 -756 2856 -719
rect 2349 -998 2383 -982
rect 2468 -806 2502 -790
rect 819 -1072 2265 -1033
rect 2468 -1036 2502 -982
rect 2586 -806 2620 -756
rect 2586 -998 2620 -982
rect 2704 -806 2738 -790
rect 2704 -1036 2738 -982
rect 2822 -806 2856 -756
rect 2822 -998 2856 -982
rect 3404 -755 3674 -716
rect 3404 -806 3438 -755
rect 3404 -998 3438 -982
rect 3522 -806 3556 -790
rect 2468 -1075 2738 -1036
rect 3522 -1033 3556 -982
rect 3640 -806 3674 -755
rect 3640 -998 3674 -982
rect 3758 -806 3792 -790
rect 3758 -1033 3792 -982
rect 3845 -998 3879 -982
rect 3963 -606 3997 -590
rect 3522 -1072 3792 -1033
rect 3963 -1033 3997 -982
rect 4081 -606 4115 -553
rect 4312 -554 4582 -515
rect 4081 -998 4115 -982
rect 4199 -606 4233 -590
rect 4199 -1033 4233 -982
rect 4312 -606 4346 -554
rect 4312 -998 4346 -982
rect 4430 -606 4464 -590
rect 4430 -1033 4464 -982
rect 4548 -606 4582 -554
rect 4784 -554 5054 -515
rect 4548 -998 4582 -982
rect 4666 -606 4700 -590
rect 4666 -1033 4700 -982
rect 4784 -606 4818 -554
rect 4784 -998 4818 -982
rect 4902 -606 4936 -590
rect 4902 -1033 4936 -982
rect 5020 -606 5054 -554
rect 5257 -554 5527 -515
rect 5020 -998 5054 -982
rect 5139 -606 5173 -590
rect 5139 -1033 5173 -982
rect 5257 -606 5291 -554
rect 5257 -998 5291 -982
rect 5375 -606 5409 -590
rect 5375 -1033 5409 -982
rect 5493 -606 5527 -554
rect 6977 -549 7247 -510
rect 6977 -602 7011 -549
rect 5730 -756 6000 -719
rect 5493 -998 5527 -982
rect 5612 -806 5646 -790
rect 3963 -1072 5409 -1033
rect 5612 -1036 5646 -982
rect 5730 -806 5764 -756
rect 5730 -998 5764 -982
rect 5848 -806 5882 -790
rect 5848 -1036 5882 -982
rect 5966 -806 6000 -756
rect 5966 -998 6000 -982
rect 6536 -751 6806 -712
rect 6536 -802 6570 -751
rect 6536 -994 6570 -978
rect 6654 -802 6688 -786
rect 5612 -1075 5882 -1036
rect 6654 -1029 6688 -978
rect 6772 -802 6806 -751
rect 6772 -994 6806 -978
rect 6890 -802 6924 -786
rect 6890 -1029 6924 -978
rect 6977 -994 7011 -978
rect 7095 -602 7129 -586
rect 6654 -1068 6924 -1029
rect 7095 -1029 7129 -978
rect 7213 -602 7247 -549
rect 7444 -550 7714 -511
rect 7213 -994 7247 -978
rect 7331 -602 7365 -586
rect 7331 -1029 7365 -978
rect 7444 -602 7478 -550
rect 7444 -994 7478 -978
rect 7562 -602 7596 -586
rect 7562 -1029 7596 -978
rect 7680 -602 7714 -550
rect 7916 -550 8186 -511
rect 7680 -994 7714 -978
rect 7798 -602 7832 -586
rect 7798 -1029 7832 -978
rect 7916 -602 7950 -550
rect 7916 -994 7950 -978
rect 8034 -602 8068 -586
rect 8034 -1029 8068 -978
rect 8152 -602 8186 -550
rect 8389 -550 8659 -511
rect 8152 -994 8186 -978
rect 8271 -602 8305 -586
rect 8271 -1029 8305 -978
rect 8389 -602 8423 -550
rect 8389 -994 8423 -978
rect 8507 -602 8541 -586
rect 8507 -1029 8541 -978
rect 8625 -602 8659 -550
rect 10121 -549 10391 -510
rect 10121 -602 10155 -549
rect 8862 -752 9132 -715
rect 8625 -994 8659 -978
rect 8744 -802 8778 -786
rect 7095 -1068 8541 -1029
rect 8744 -1032 8778 -978
rect 8862 -802 8896 -752
rect 8862 -994 8896 -978
rect 8980 -802 9014 -786
rect 8980 -1032 9014 -978
rect 9098 -802 9132 -752
rect 9098 -994 9132 -978
rect 9680 -751 9950 -712
rect 9680 -802 9714 -751
rect 9680 -994 9714 -978
rect 9798 -802 9832 -786
rect 8744 -1071 9014 -1032
rect 9798 -1029 9832 -978
rect 9916 -802 9950 -751
rect 9916 -994 9950 -978
rect 10034 -802 10068 -786
rect 10034 -1029 10068 -978
rect 10121 -994 10155 -978
rect 10239 -602 10273 -586
rect 9798 -1068 10068 -1029
rect 10239 -1029 10273 -978
rect 10357 -602 10391 -549
rect 10588 -550 10858 -511
rect 10357 -994 10391 -978
rect 10475 -602 10509 -586
rect 10475 -1029 10509 -978
rect 10588 -602 10622 -550
rect 10588 -994 10622 -978
rect 10706 -602 10740 -586
rect 10706 -1029 10740 -978
rect 10824 -602 10858 -550
rect 11060 -550 11330 -511
rect 10824 -994 10858 -978
rect 10942 -602 10976 -586
rect 10942 -1029 10976 -978
rect 11060 -602 11094 -550
rect 11060 -994 11094 -978
rect 11178 -602 11212 -586
rect 11178 -1029 11212 -978
rect 11296 -602 11330 -550
rect 11533 -550 11803 -511
rect 11296 -994 11330 -978
rect 11415 -602 11449 -586
rect 11415 -1029 11449 -978
rect 11533 -602 11567 -550
rect 11533 -994 11567 -978
rect 11651 -602 11685 -586
rect 11651 -1029 11685 -978
rect 11769 -602 11803 -550
rect 13323 -553 13593 -514
rect 13323 -606 13357 -553
rect 12006 -752 12276 -715
rect 11769 -994 11803 -978
rect 11888 -802 11922 -786
rect 10239 -1068 11685 -1029
rect 11888 -1032 11922 -978
rect 12006 -802 12040 -752
rect 12006 -994 12040 -978
rect 12124 -802 12158 -786
rect 12124 -1032 12158 -978
rect 12242 -802 12276 -752
rect 12242 -994 12276 -978
rect 12882 -755 13152 -716
rect 12882 -806 12916 -755
rect 12882 -998 12916 -982
rect 13000 -806 13034 -790
rect 11888 -1071 12158 -1032
rect 13000 -1033 13034 -982
rect 13118 -806 13152 -755
rect 13118 -998 13152 -982
rect 13236 -806 13270 -790
rect 13236 -1033 13270 -982
rect 13323 -998 13357 -982
rect 13441 -606 13475 -590
rect 13000 -1072 13270 -1033
rect 13441 -1033 13475 -982
rect 13559 -606 13593 -553
rect 13790 -554 14060 -515
rect 13559 -998 13593 -982
rect 13677 -606 13711 -590
rect 13677 -1033 13711 -982
rect 13790 -606 13824 -554
rect 13790 -998 13824 -982
rect 13908 -606 13942 -590
rect 13908 -1033 13942 -982
rect 14026 -606 14060 -554
rect 14262 -554 14532 -515
rect 14026 -998 14060 -982
rect 14144 -606 14178 -590
rect 14144 -1033 14178 -982
rect 14262 -606 14296 -554
rect 14262 -998 14296 -982
rect 14380 -606 14414 -590
rect 14380 -1033 14414 -982
rect 14498 -606 14532 -554
rect 14735 -554 15005 -515
rect 14498 -998 14532 -982
rect 14617 -606 14651 -590
rect 14617 -1033 14651 -982
rect 14735 -606 14769 -554
rect 14735 -998 14769 -982
rect 14853 -606 14887 -590
rect 14853 -1033 14887 -982
rect 14971 -606 15005 -554
rect 16467 -553 16737 -514
rect 16467 -606 16501 -553
rect 15208 -756 15478 -719
rect 14971 -998 15005 -982
rect 15090 -806 15124 -790
rect 13441 -1072 14887 -1033
rect 15090 -1036 15124 -982
rect 15208 -806 15242 -756
rect 15208 -998 15242 -982
rect 15326 -806 15360 -790
rect 15326 -1036 15360 -982
rect 15444 -806 15478 -756
rect 15444 -998 15478 -982
rect 16026 -755 16296 -716
rect 16026 -806 16060 -755
rect 16026 -998 16060 -982
rect 16144 -806 16178 -790
rect 15090 -1075 15360 -1036
rect 16144 -1033 16178 -982
rect 16262 -806 16296 -755
rect 16262 -998 16296 -982
rect 16380 -806 16414 -790
rect 16380 -1033 16414 -982
rect 16467 -998 16501 -982
rect 16585 -606 16619 -590
rect 16144 -1072 16414 -1033
rect 16585 -1033 16619 -982
rect 16703 -606 16737 -553
rect 16934 -554 17204 -515
rect 16703 -998 16737 -982
rect 16821 -606 16855 -590
rect 16821 -1033 16855 -982
rect 16934 -606 16968 -554
rect 16934 -998 16968 -982
rect 17052 -606 17086 -590
rect 17052 -1033 17086 -982
rect 17170 -606 17204 -554
rect 17406 -554 17676 -515
rect 17170 -998 17204 -982
rect 17288 -606 17322 -590
rect 17288 -1033 17322 -982
rect 17406 -606 17440 -554
rect 17406 -998 17440 -982
rect 17524 -606 17558 -590
rect 17524 -1033 17558 -982
rect 17642 -606 17676 -554
rect 17879 -554 18149 -515
rect 17642 -998 17676 -982
rect 17761 -606 17795 -590
rect 17761 -1033 17795 -982
rect 17879 -606 17913 -554
rect 17879 -998 17913 -982
rect 17997 -606 18031 -590
rect 17997 -1033 18031 -982
rect 18115 -606 18149 -554
rect 19599 -549 19869 -510
rect 19599 -602 19633 -549
rect 18352 -756 18622 -719
rect 18115 -998 18149 -982
rect 18234 -806 18268 -790
rect 16585 -1072 18031 -1033
rect 18234 -1036 18268 -982
rect 18352 -806 18386 -756
rect 18352 -998 18386 -982
rect 18470 -806 18504 -790
rect 18470 -1036 18504 -982
rect 18588 -806 18622 -756
rect 18588 -998 18622 -982
rect 19158 -751 19428 -712
rect 19158 -802 19192 -751
rect 19158 -994 19192 -978
rect 19276 -802 19310 -786
rect 18234 -1075 18504 -1036
rect 19276 -1029 19310 -978
rect 19394 -802 19428 -751
rect 19394 -994 19428 -978
rect 19512 -802 19546 -786
rect 19512 -1029 19546 -978
rect 19599 -994 19633 -978
rect 19717 -602 19751 -586
rect 19276 -1068 19546 -1029
rect 19717 -1029 19751 -978
rect 19835 -602 19869 -549
rect 20066 -550 20336 -511
rect 19835 -994 19869 -978
rect 19953 -602 19987 -586
rect 19953 -1029 19987 -978
rect 20066 -602 20100 -550
rect 20066 -994 20100 -978
rect 20184 -602 20218 -586
rect 20184 -1029 20218 -978
rect 20302 -602 20336 -550
rect 20538 -550 20808 -511
rect 20302 -994 20336 -978
rect 20420 -602 20454 -586
rect 20420 -1029 20454 -978
rect 20538 -602 20572 -550
rect 20538 -994 20572 -978
rect 20656 -602 20690 -586
rect 20656 -1029 20690 -978
rect 20774 -602 20808 -550
rect 21011 -550 21281 -511
rect 20774 -994 20808 -978
rect 20893 -602 20927 -586
rect 20893 -1029 20927 -978
rect 21011 -602 21045 -550
rect 21011 -994 21045 -978
rect 21129 -602 21163 -586
rect 21129 -1029 21163 -978
rect 21247 -602 21281 -550
rect 22743 -549 23013 -510
rect 22743 -602 22777 -549
rect 21484 -752 21754 -715
rect 21247 -994 21281 -978
rect 21366 -802 21400 -786
rect 19717 -1068 21163 -1029
rect 21366 -1032 21400 -978
rect 21484 -802 21518 -752
rect 21484 -994 21518 -978
rect 21602 -802 21636 -786
rect 21602 -1032 21636 -978
rect 21720 -802 21754 -752
rect 21720 -994 21754 -978
rect 22302 -751 22572 -712
rect 22302 -802 22336 -751
rect 22302 -994 22336 -978
rect 22420 -802 22454 -786
rect 21366 -1071 21636 -1032
rect 22420 -1029 22454 -978
rect 22538 -802 22572 -751
rect 22538 -994 22572 -978
rect 22656 -802 22690 -786
rect 22656 -1029 22690 -978
rect 22743 -994 22777 -978
rect 22861 -602 22895 -586
rect 22420 -1068 22690 -1029
rect 22861 -1029 22895 -978
rect 22979 -602 23013 -549
rect 23210 -550 23480 -511
rect 22979 -994 23013 -978
rect 23097 -602 23131 -586
rect 23097 -1029 23131 -978
rect 23210 -602 23244 -550
rect 23210 -994 23244 -978
rect 23328 -602 23362 -586
rect 23328 -1029 23362 -978
rect 23446 -602 23480 -550
rect 23682 -550 23952 -511
rect 23446 -994 23480 -978
rect 23564 -602 23598 -586
rect 23564 -1029 23598 -978
rect 23682 -602 23716 -550
rect 23682 -994 23716 -978
rect 23800 -602 23834 -586
rect 23800 -1029 23834 -978
rect 23918 -602 23952 -550
rect 24155 -550 24425 -511
rect 23918 -994 23952 -978
rect 24037 -602 24071 -586
rect 24037 -1029 24071 -978
rect 24155 -602 24189 -550
rect 24155 -994 24189 -978
rect 24273 -602 24307 -586
rect 24273 -1029 24307 -978
rect 24391 -602 24425 -550
rect 24628 -752 24898 -715
rect 24391 -994 24425 -978
rect 24510 -802 24544 -786
rect 22861 -1068 24307 -1029
rect 24510 -1032 24544 -978
rect 24628 -802 24662 -752
rect 24628 -994 24662 -978
rect 24746 -802 24780 -786
rect 24746 -1032 24780 -978
rect 24864 -802 24898 -752
rect 24864 -994 24898 -978
rect 24510 -1071 24780 -1032
rect 1346 -1197 1380 -1181
rect 2640 -1190 2656 -1156
rect 2690 -1190 2706 -1156
rect 1346 -1247 1380 -1231
rect 4490 -1197 4524 -1181
rect 5784 -1190 5800 -1156
rect 5834 -1190 5850 -1156
rect 4490 -1247 4524 -1231
rect 7622 -1193 7656 -1177
rect 8916 -1186 8932 -1152
rect 8966 -1186 8982 -1152
rect 7622 -1243 7656 -1227
rect 10766 -1193 10800 -1177
rect 12060 -1186 12076 -1152
rect 12110 -1186 12126 -1152
rect 10766 -1243 10800 -1227
rect 13968 -1197 14002 -1181
rect 15262 -1190 15278 -1156
rect 15312 -1190 15328 -1156
rect 13968 -1247 14002 -1231
rect 17112 -1197 17146 -1181
rect 18406 -1190 18422 -1156
rect 18456 -1190 18472 -1156
rect 17112 -1247 17146 -1231
rect 20244 -1193 20278 -1177
rect 21538 -1186 21554 -1152
rect 21588 -1186 21604 -1152
rect 20244 -1243 20278 -1227
rect 23388 -1193 23422 -1177
rect 24682 -1186 24698 -1152
rect 24732 -1186 24748 -1152
rect 23388 -1243 23422 -1227
rect 349 -1297 441 -1280
rect 349 -1352 365 -1297
rect 425 -1352 441 -1297
rect 349 -1365 441 -1352
rect 1434 -1296 1526 -1283
rect 1434 -1351 1450 -1296
rect 1510 -1351 1526 -1296
rect 1434 -1368 1526 -1351
rect 3493 -1297 3585 -1280
rect 3493 -1352 3509 -1297
rect 3569 -1352 3585 -1297
rect 3493 -1365 3585 -1352
rect 4578 -1296 4670 -1283
rect 4578 -1351 4594 -1296
rect 4654 -1351 4670 -1296
rect 4578 -1368 4670 -1351
rect 6625 -1293 6717 -1276
rect 6625 -1348 6641 -1293
rect 6701 -1348 6717 -1293
rect 6625 -1361 6717 -1348
rect 7710 -1292 7802 -1279
rect 7710 -1347 7726 -1292
rect 7786 -1347 7802 -1292
rect 7710 -1364 7802 -1347
rect 9769 -1293 9861 -1276
rect 9769 -1348 9785 -1293
rect 9845 -1348 9861 -1293
rect 9769 -1361 9861 -1348
rect 10854 -1292 10946 -1279
rect 10854 -1347 10870 -1292
rect 10930 -1347 10946 -1292
rect 10854 -1364 10946 -1347
rect 12971 -1297 13063 -1280
rect 12971 -1352 12987 -1297
rect 13047 -1352 13063 -1297
rect 12971 -1365 13063 -1352
rect 14056 -1296 14148 -1283
rect 14056 -1351 14072 -1296
rect 14132 -1351 14148 -1296
rect 14056 -1368 14148 -1351
rect 15883 -1296 15940 -1292
rect 15883 -1356 15887 -1296
rect 15936 -1356 15940 -1296
rect 15883 -1360 15940 -1356
rect 16115 -1297 16207 -1280
rect 16115 -1352 16131 -1297
rect 16191 -1352 16207 -1297
rect 16115 -1365 16207 -1352
rect 17200 -1296 17292 -1283
rect 17200 -1351 17216 -1296
rect 17276 -1351 17292 -1296
rect 17200 -1368 17292 -1351
rect 19247 -1293 19339 -1276
rect 19247 -1348 19263 -1293
rect 19323 -1348 19339 -1293
rect 19247 -1361 19339 -1348
rect 20332 -1292 20424 -1279
rect 20332 -1347 20348 -1292
rect 20408 -1347 20424 -1292
rect 20332 -1364 20424 -1347
rect 22391 -1293 22483 -1276
rect 22391 -1348 22407 -1293
rect 22467 -1348 22483 -1293
rect 22391 -1361 22483 -1348
rect 23476 -1292 23568 -1279
rect 23476 -1347 23492 -1292
rect 23552 -1347 23568 -1292
rect 23476 -1364 23568 -1347
rect 6393 -1408 6450 -1404
rect 117 -1412 174 -1408
rect 117 -1472 121 -1412
rect 170 -1472 174 -1412
rect 117 -1476 174 -1472
rect 1700 -1427 1734 -1411
rect 1700 -1477 1734 -1461
rect 3261 -1412 3318 -1408
rect 3261 -1472 3265 -1412
rect 3314 -1472 3318 -1412
rect 3261 -1476 3318 -1472
rect 4844 -1427 4878 -1411
rect 4844 -1477 4878 -1461
rect 6393 -1468 6397 -1408
rect 6446 -1468 6450 -1408
rect 6393 -1472 6450 -1468
rect 7976 -1423 8010 -1407
rect 7976 -1473 8010 -1457
rect 9537 -1408 9594 -1404
rect 9537 -1468 9541 -1408
rect 9590 -1468 9594 -1408
rect 9537 -1472 9594 -1468
rect 11120 -1423 11154 -1407
rect 19015 -1408 19072 -1404
rect 11120 -1473 11154 -1457
rect 12739 -1412 12796 -1408
rect 12739 -1472 12743 -1412
rect 12792 -1472 12796 -1412
rect 12739 -1476 12796 -1472
rect 14322 -1427 14356 -1411
rect 14322 -1477 14356 -1461
rect 15883 -1412 15940 -1408
rect 15883 -1472 15887 -1412
rect 15936 -1472 15940 -1412
rect 15883 -1476 15940 -1472
rect 17466 -1427 17500 -1411
rect 17466 -1477 17500 -1461
rect 19015 -1468 19019 -1408
rect 19068 -1468 19072 -1408
rect 19015 -1472 19072 -1468
rect 20598 -1423 20632 -1407
rect 20598 -1473 20632 -1457
rect 22159 -1408 22216 -1404
rect 22159 -1468 22163 -1408
rect 22212 -1468 22216 -1408
rect 22159 -1472 22216 -1468
rect 23742 -1423 23776 -1407
rect 23742 -1473 23776 -1457
rect 117 -1580 174 -1576
rect 117 -1640 121 -1580
rect 170 -1640 174 -1580
rect 117 -1644 174 -1640
rect 1316 -1581 1408 -1568
rect 1316 -1636 1332 -1581
rect 1392 -1636 1408 -1581
rect 1316 -1653 1408 -1636
rect 3261 -1580 3318 -1576
rect 3261 -1640 3265 -1580
rect 3314 -1640 3318 -1580
rect 3261 -1644 3318 -1640
rect 4460 -1581 4552 -1568
rect 4460 -1636 4476 -1581
rect 4536 -1636 4552 -1581
rect 4460 -1653 4552 -1636
rect 6393 -1576 6450 -1572
rect 6393 -1636 6397 -1576
rect 6446 -1636 6450 -1576
rect 6393 -1640 6450 -1636
rect 7592 -1577 7684 -1564
rect 7592 -1632 7608 -1577
rect 7668 -1632 7684 -1577
rect 7592 -1649 7684 -1632
rect 9537 -1576 9594 -1572
rect 9537 -1636 9541 -1576
rect 9590 -1636 9594 -1576
rect 9537 -1640 9594 -1636
rect 10736 -1577 10828 -1564
rect 10736 -1632 10752 -1577
rect 10812 -1632 10828 -1577
rect 10736 -1649 10828 -1632
rect 12739 -1580 12796 -1576
rect 12739 -1640 12743 -1580
rect 12792 -1640 12796 -1580
rect 12739 -1644 12796 -1640
rect 13938 -1581 14030 -1568
rect 13938 -1636 13954 -1581
rect 14014 -1636 14030 -1581
rect 13938 -1653 14030 -1636
rect 15883 -1580 15940 -1576
rect 15883 -1640 15887 -1580
rect 15936 -1640 15940 -1580
rect 15883 -1644 15940 -1640
rect 17082 -1581 17174 -1568
rect 17082 -1636 17098 -1581
rect 17158 -1636 17174 -1581
rect 17082 -1653 17174 -1636
rect 19015 -1576 19072 -1572
rect 19015 -1636 19019 -1576
rect 19068 -1636 19072 -1576
rect 19015 -1640 19072 -1636
rect 20214 -1577 20306 -1564
rect 20214 -1632 20230 -1577
rect 20290 -1632 20306 -1577
rect 20214 -1649 20306 -1632
rect 22159 -1576 22216 -1572
rect 22159 -1636 22163 -1576
rect 22212 -1636 22216 -1576
rect 22159 -1640 22216 -1636
rect 23358 -1577 23450 -1564
rect 23358 -1632 23374 -1577
rect 23434 -1632 23450 -1577
rect 23358 -1649 23450 -1632
rect 1581 -1817 1615 -1801
rect 1581 -1867 1615 -1851
rect 4725 -1817 4759 -1801
rect 4725 -1867 4759 -1851
rect 7857 -1813 7891 -1797
rect 7857 -1863 7891 -1847
rect 11001 -1813 11035 -1797
rect 11001 -1863 11035 -1847
rect 14203 -1817 14237 -1801
rect 14203 -1867 14237 -1851
rect 17347 -1817 17381 -1801
rect 17347 -1867 17381 -1851
rect 20479 -1813 20513 -1797
rect 20479 -1863 20513 -1847
rect 23623 -1813 23657 -1797
rect 23623 -1863 23657 -1847
rect 1094 -1939 1128 -1923
rect 1094 -2131 1128 -2115
rect 1212 -1927 1246 -1923
rect 1286 -1927 1320 -1923
rect 1212 -1939 1320 -1927
rect 1246 -2115 1286 -1939
rect 1212 -2127 1286 -2115
rect 1212 -2131 1246 -2127
rect 1286 -2331 1320 -2315
rect 1404 -1939 1438 -1923
rect 1404 -2331 1438 -2315
rect 1522 -1939 1556 -1923
rect 1522 -2331 1556 -2315
rect 1640 -1939 1674 -1923
rect 1640 -2331 1674 -2315
rect 1758 -1927 1792 -1923
rect 1836 -1927 1870 -1923
rect 1758 -1939 1870 -1927
rect 1792 -2115 1836 -1939
rect 1792 -2127 1870 -2115
rect 1836 -2131 1870 -2127
rect 1954 -1939 1988 -1923
rect 1954 -2131 1988 -2115
rect 4238 -1939 4272 -1923
rect 4238 -2131 4272 -2115
rect 4356 -1927 4390 -1923
rect 4430 -1927 4464 -1923
rect 4356 -1939 4464 -1927
rect 4390 -2115 4430 -1939
rect 4356 -2127 4430 -2115
rect 4356 -2131 4390 -2127
rect 1758 -2331 1792 -2315
rect 4430 -2331 4464 -2315
rect 4548 -1939 4582 -1923
rect 4548 -2331 4582 -2315
rect 4666 -1939 4700 -1923
rect 4666 -2331 4700 -2315
rect 4784 -1939 4818 -1923
rect 4784 -2331 4818 -2315
rect 4902 -1927 4936 -1923
rect 4980 -1927 5014 -1923
rect 4902 -1939 5014 -1927
rect 4936 -2115 4980 -1939
rect 4936 -2127 5014 -2115
rect 4980 -2131 5014 -2127
rect 5098 -1939 5132 -1923
rect 5098 -2131 5132 -2115
rect 7370 -1935 7404 -1919
rect 7370 -2127 7404 -2111
rect 7488 -1923 7522 -1919
rect 7562 -1923 7596 -1919
rect 7488 -1935 7596 -1923
rect 7522 -2111 7562 -1935
rect 7488 -2123 7562 -2111
rect 7488 -2127 7522 -2123
rect 4902 -2331 4936 -2315
rect 7562 -2327 7596 -2311
rect 7680 -1935 7714 -1919
rect 7680 -2327 7714 -2311
rect 7798 -1935 7832 -1919
rect 7798 -2327 7832 -2311
rect 7916 -1935 7950 -1919
rect 7916 -2327 7950 -2311
rect 8034 -1923 8068 -1919
rect 8112 -1923 8146 -1919
rect 8034 -1935 8146 -1923
rect 8068 -2111 8112 -1935
rect 8068 -2123 8146 -2111
rect 8112 -2127 8146 -2123
rect 8230 -1935 8264 -1919
rect 8230 -2127 8264 -2111
rect 10514 -1935 10548 -1919
rect 10514 -2127 10548 -2111
rect 10632 -1923 10666 -1919
rect 10706 -1923 10740 -1919
rect 10632 -1935 10740 -1923
rect 10666 -2111 10706 -1935
rect 10632 -2123 10706 -2111
rect 10632 -2127 10666 -2123
rect 8034 -2327 8068 -2311
rect 10706 -2327 10740 -2311
rect 10824 -1935 10858 -1919
rect 10824 -2327 10858 -2311
rect 10942 -1935 10976 -1919
rect 10942 -2327 10976 -2311
rect 11060 -1935 11094 -1919
rect 11060 -2327 11094 -2311
rect 11178 -1923 11212 -1919
rect 11256 -1923 11290 -1919
rect 11178 -1935 11290 -1923
rect 11212 -2111 11256 -1935
rect 11212 -2123 11290 -2111
rect 11256 -2127 11290 -2123
rect 11374 -1935 11408 -1919
rect 11374 -2127 11408 -2111
rect 13716 -1939 13750 -1923
rect 13716 -2131 13750 -2115
rect 13834 -1927 13868 -1923
rect 13908 -1927 13942 -1923
rect 13834 -1939 13942 -1927
rect 13868 -2115 13908 -1939
rect 13834 -2127 13908 -2115
rect 13834 -2131 13868 -2127
rect 11178 -2327 11212 -2311
rect 13908 -2331 13942 -2315
rect 14026 -1939 14060 -1923
rect 14026 -2331 14060 -2315
rect 14144 -1939 14178 -1923
rect 14144 -2331 14178 -2315
rect 14262 -1939 14296 -1923
rect 14262 -2331 14296 -2315
rect 14380 -1927 14414 -1923
rect 14458 -1927 14492 -1923
rect 14380 -1939 14492 -1927
rect 14414 -2115 14458 -1939
rect 14414 -2127 14492 -2115
rect 14458 -2131 14492 -2127
rect 14576 -1939 14610 -1923
rect 14576 -2131 14610 -2115
rect 16860 -1939 16894 -1923
rect 16860 -2131 16894 -2115
rect 16978 -1927 17012 -1923
rect 17052 -1927 17086 -1923
rect 16978 -1939 17086 -1927
rect 17012 -2115 17052 -1939
rect 16978 -2127 17052 -2115
rect 16978 -2131 17012 -2127
rect 14380 -2331 14414 -2315
rect 17052 -2331 17086 -2315
rect 17170 -1939 17204 -1923
rect 17170 -2331 17204 -2315
rect 17288 -1939 17322 -1923
rect 17288 -2331 17322 -2315
rect 17406 -1939 17440 -1923
rect 17406 -2331 17440 -2315
rect 17524 -1927 17558 -1923
rect 17602 -1927 17636 -1923
rect 17524 -1939 17636 -1927
rect 17558 -2115 17602 -1939
rect 17558 -2127 17636 -2115
rect 17602 -2131 17636 -2127
rect 17720 -1939 17754 -1923
rect 17720 -2131 17754 -2115
rect 19992 -1935 20026 -1919
rect 19992 -2127 20026 -2111
rect 20110 -1923 20144 -1919
rect 20184 -1923 20218 -1919
rect 20110 -1935 20218 -1923
rect 20144 -2111 20184 -1935
rect 20110 -2123 20184 -2111
rect 20110 -2127 20144 -2123
rect 17524 -2331 17558 -2315
rect 20184 -2327 20218 -2311
rect 20302 -1935 20336 -1919
rect 20302 -2327 20336 -2311
rect 20420 -1935 20454 -1919
rect 20420 -2327 20454 -2311
rect 20538 -1935 20572 -1919
rect 20538 -2327 20572 -2311
rect 20656 -1923 20690 -1919
rect 20734 -1923 20768 -1919
rect 20656 -1935 20768 -1923
rect 20690 -2111 20734 -1935
rect 20690 -2123 20768 -2111
rect 20734 -2127 20768 -2123
rect 20852 -1935 20886 -1919
rect 20852 -2127 20886 -2111
rect 23136 -1935 23170 -1919
rect 23136 -2127 23170 -2111
rect 23254 -1923 23288 -1919
rect 23328 -1923 23362 -1919
rect 23254 -1935 23362 -1923
rect 23288 -2111 23328 -1935
rect 23254 -2123 23328 -2111
rect 23254 -2127 23288 -2123
rect 20656 -2327 20690 -2311
rect 23328 -2327 23362 -2311
rect 23446 -1935 23480 -1919
rect 23446 -2327 23480 -2311
rect 23564 -1935 23598 -1919
rect 23564 -2327 23598 -2311
rect 23682 -1935 23716 -1919
rect 23682 -2327 23716 -2311
rect 23800 -1923 23834 -1919
rect 23878 -1923 23912 -1919
rect 23800 -1935 23912 -1923
rect 23834 -2111 23878 -1935
rect 23834 -2123 23912 -2111
rect 23878 -2127 23912 -2123
rect 23996 -1935 24030 -1919
rect 23996 -2127 24030 -2111
rect 23800 -2327 23834 -2311
rect 1507 -2450 1523 -2416
rect 1557 -2450 1573 -2416
rect 4651 -2450 4667 -2416
rect 4701 -2450 4717 -2416
rect 7783 -2446 7799 -2412
rect 7833 -2446 7849 -2412
rect 10927 -2446 10943 -2412
rect 10977 -2446 10993 -2412
rect 14129 -2450 14145 -2416
rect 14179 -2450 14195 -2416
rect 17273 -2450 17289 -2416
rect 17323 -2450 17339 -2416
rect 20405 -2446 20421 -2412
rect 20455 -2446 20471 -2412
rect 23549 -2446 23565 -2412
rect 23599 -2446 23615 -2412
rect 7764 -2564 7900 -2560
rect 1488 -2568 1624 -2564
rect 1488 -2582 1526 -2568
rect 1584 -2582 1624 -2568
rect 1488 -2628 1504 -2582
rect 1608 -2628 1624 -2582
rect 1488 -2650 1624 -2628
rect 4632 -2568 4768 -2564
rect 4632 -2582 4670 -2568
rect 4728 -2582 4768 -2568
rect 4632 -2628 4648 -2582
rect 4752 -2628 4768 -2582
rect 4632 -2650 4768 -2628
rect 7764 -2578 7802 -2564
rect 7860 -2578 7900 -2564
rect 7764 -2624 7780 -2578
rect 7884 -2624 7900 -2578
rect 7764 -2646 7900 -2624
rect 10908 -2564 11044 -2560
rect 20386 -2564 20522 -2560
rect 10908 -2578 10946 -2564
rect 11004 -2578 11044 -2564
rect 10908 -2624 10924 -2578
rect 11028 -2624 11044 -2578
rect 10908 -2646 11044 -2624
rect 14110 -2568 14246 -2564
rect 14110 -2582 14148 -2568
rect 14206 -2582 14246 -2568
rect 14110 -2628 14126 -2582
rect 14230 -2628 14246 -2582
rect 14110 -2650 14246 -2628
rect 17254 -2568 17390 -2564
rect 17254 -2582 17292 -2568
rect 17350 -2582 17390 -2568
rect 17254 -2628 17270 -2582
rect 17374 -2628 17390 -2582
rect 17254 -2650 17390 -2628
rect 20386 -2578 20424 -2564
rect 20482 -2578 20522 -2564
rect 20386 -2624 20402 -2578
rect 20506 -2624 20522 -2578
rect 20386 -2646 20522 -2624
rect 23530 -2564 23666 -2560
rect 23530 -2578 23568 -2564
rect 23626 -2578 23666 -2564
rect 23530 -2624 23546 -2578
rect 23650 -2624 23666 -2578
rect 23530 -2646 23666 -2624
rect 1420 -3068 1648 -3050
rect 1420 -3144 1436 -3068
rect 1632 -3144 1648 -3068
rect 1420 -3160 1648 -3144
rect 4564 -3068 4792 -3050
rect 4564 -3144 4580 -3068
rect 4776 -3144 4792 -3068
rect 4564 -3160 4792 -3144
rect 7696 -3064 7924 -3046
rect 7696 -3140 7712 -3064
rect 7908 -3140 7924 -3064
rect 7696 -3156 7924 -3140
rect 10840 -3064 11068 -3046
rect 10840 -3140 10856 -3064
rect 11052 -3140 11068 -3064
rect 10840 -3156 11068 -3140
rect 14042 -3068 14270 -3050
rect 14042 -3144 14058 -3068
rect 14254 -3144 14270 -3068
rect 14042 -3160 14270 -3144
rect 17186 -3068 17414 -3050
rect 17186 -3144 17202 -3068
rect 17398 -3144 17414 -3068
rect 17186 -3160 17414 -3144
rect 20318 -3064 20546 -3046
rect 20318 -3140 20334 -3064
rect 20530 -3140 20546 -3064
rect 20318 -3156 20546 -3140
rect 23462 -3064 23690 -3046
rect 23462 -3140 23478 -3064
rect 23674 -3140 23690 -3064
rect 23462 -3156 23690 -3140
rect 691 -3285 961 -3246
rect 691 -3338 725 -3285
rect 250 -3487 520 -3448
rect 250 -3538 284 -3487
rect 250 -3730 284 -3714
rect 368 -3538 402 -3522
rect 368 -3765 402 -3714
rect 486 -3538 520 -3487
rect 486 -3730 520 -3714
rect 604 -3538 638 -3522
rect 604 -3765 638 -3714
rect 691 -3730 725 -3714
rect 809 -3338 843 -3322
rect 368 -3804 638 -3765
rect 809 -3765 843 -3714
rect 927 -3338 961 -3285
rect 1158 -3286 1428 -3247
rect 927 -3730 961 -3714
rect 1045 -3338 1079 -3322
rect 1045 -3765 1079 -3714
rect 1158 -3338 1192 -3286
rect 1158 -3730 1192 -3714
rect 1276 -3338 1310 -3322
rect 1276 -3765 1310 -3714
rect 1394 -3338 1428 -3286
rect 1630 -3286 1900 -3247
rect 1394 -3730 1428 -3714
rect 1512 -3338 1546 -3322
rect 1512 -3765 1546 -3714
rect 1630 -3338 1664 -3286
rect 1630 -3730 1664 -3714
rect 1748 -3338 1782 -3322
rect 1748 -3765 1782 -3714
rect 1866 -3338 1900 -3286
rect 2103 -3286 2373 -3247
rect 1866 -3730 1900 -3714
rect 1985 -3338 2019 -3322
rect 1985 -3765 2019 -3714
rect 2103 -3338 2137 -3286
rect 2103 -3730 2137 -3714
rect 2221 -3338 2255 -3322
rect 2221 -3765 2255 -3714
rect 2339 -3338 2373 -3286
rect 3835 -3285 4105 -3246
rect 3835 -3338 3869 -3285
rect 2576 -3488 2846 -3451
rect 2339 -3730 2373 -3714
rect 2458 -3538 2492 -3522
rect 809 -3804 2255 -3765
rect 2458 -3768 2492 -3714
rect 2576 -3538 2610 -3488
rect 2576 -3730 2610 -3714
rect 2694 -3538 2728 -3522
rect 2694 -3768 2728 -3714
rect 2812 -3538 2846 -3488
rect 2812 -3730 2846 -3714
rect 3394 -3487 3664 -3448
rect 3394 -3538 3428 -3487
rect 3394 -3730 3428 -3714
rect 3512 -3538 3546 -3522
rect 2458 -3807 2728 -3768
rect 3512 -3765 3546 -3714
rect 3630 -3538 3664 -3487
rect 3630 -3730 3664 -3714
rect 3748 -3538 3782 -3522
rect 3748 -3765 3782 -3714
rect 3835 -3730 3869 -3714
rect 3953 -3338 3987 -3322
rect 3512 -3804 3782 -3765
rect 3953 -3765 3987 -3714
rect 4071 -3338 4105 -3285
rect 4302 -3286 4572 -3247
rect 4071 -3730 4105 -3714
rect 4189 -3338 4223 -3322
rect 4189 -3765 4223 -3714
rect 4302 -3338 4336 -3286
rect 4302 -3730 4336 -3714
rect 4420 -3338 4454 -3322
rect 4420 -3765 4454 -3714
rect 4538 -3338 4572 -3286
rect 4774 -3286 5044 -3247
rect 4538 -3730 4572 -3714
rect 4656 -3338 4690 -3322
rect 4656 -3765 4690 -3714
rect 4774 -3338 4808 -3286
rect 4774 -3730 4808 -3714
rect 4892 -3338 4926 -3322
rect 4892 -3765 4926 -3714
rect 5010 -3338 5044 -3286
rect 5247 -3286 5517 -3247
rect 5010 -3730 5044 -3714
rect 5129 -3338 5163 -3322
rect 5129 -3765 5163 -3714
rect 5247 -3338 5281 -3286
rect 5247 -3730 5281 -3714
rect 5365 -3338 5399 -3322
rect 5365 -3765 5399 -3714
rect 5483 -3338 5517 -3286
rect 6967 -3281 7237 -3242
rect 6967 -3334 7001 -3281
rect 5720 -3488 5990 -3451
rect 5483 -3730 5517 -3714
rect 5602 -3538 5636 -3522
rect 3953 -3804 5399 -3765
rect 5602 -3768 5636 -3714
rect 5720 -3538 5754 -3488
rect 5720 -3730 5754 -3714
rect 5838 -3538 5872 -3522
rect 5838 -3768 5872 -3714
rect 5956 -3538 5990 -3488
rect 5956 -3730 5990 -3714
rect 6526 -3483 6796 -3444
rect 6526 -3534 6560 -3483
rect 6526 -3726 6560 -3710
rect 6644 -3534 6678 -3518
rect 5602 -3807 5872 -3768
rect 6644 -3761 6678 -3710
rect 6762 -3534 6796 -3483
rect 6762 -3726 6796 -3710
rect 6880 -3534 6914 -3518
rect 6880 -3761 6914 -3710
rect 6967 -3726 7001 -3710
rect 7085 -3334 7119 -3318
rect 6644 -3800 6914 -3761
rect 7085 -3761 7119 -3710
rect 7203 -3334 7237 -3281
rect 7434 -3282 7704 -3243
rect 7203 -3726 7237 -3710
rect 7321 -3334 7355 -3318
rect 7321 -3761 7355 -3710
rect 7434 -3334 7468 -3282
rect 7434 -3726 7468 -3710
rect 7552 -3334 7586 -3318
rect 7552 -3761 7586 -3710
rect 7670 -3334 7704 -3282
rect 7906 -3282 8176 -3243
rect 7670 -3726 7704 -3710
rect 7788 -3334 7822 -3318
rect 7788 -3761 7822 -3710
rect 7906 -3334 7940 -3282
rect 7906 -3726 7940 -3710
rect 8024 -3334 8058 -3318
rect 8024 -3761 8058 -3710
rect 8142 -3334 8176 -3282
rect 8379 -3282 8649 -3243
rect 8142 -3726 8176 -3710
rect 8261 -3334 8295 -3318
rect 8261 -3761 8295 -3710
rect 8379 -3334 8413 -3282
rect 8379 -3726 8413 -3710
rect 8497 -3334 8531 -3318
rect 8497 -3761 8531 -3710
rect 8615 -3334 8649 -3282
rect 10111 -3281 10381 -3242
rect 10111 -3334 10145 -3281
rect 8852 -3484 9122 -3447
rect 8615 -3726 8649 -3710
rect 8734 -3534 8768 -3518
rect 7085 -3800 8531 -3761
rect 8734 -3764 8768 -3710
rect 8852 -3534 8886 -3484
rect 8852 -3726 8886 -3710
rect 8970 -3534 9004 -3518
rect 8970 -3764 9004 -3710
rect 9088 -3534 9122 -3484
rect 9088 -3726 9122 -3710
rect 9670 -3483 9940 -3444
rect 9670 -3534 9704 -3483
rect 9670 -3726 9704 -3710
rect 9788 -3534 9822 -3518
rect 8734 -3803 9004 -3764
rect 9788 -3761 9822 -3710
rect 9906 -3534 9940 -3483
rect 9906 -3726 9940 -3710
rect 10024 -3534 10058 -3518
rect 10024 -3761 10058 -3710
rect 10111 -3726 10145 -3710
rect 10229 -3334 10263 -3318
rect 9788 -3800 10058 -3761
rect 10229 -3761 10263 -3710
rect 10347 -3334 10381 -3281
rect 10578 -3282 10848 -3243
rect 10347 -3726 10381 -3710
rect 10465 -3334 10499 -3318
rect 10465 -3761 10499 -3710
rect 10578 -3334 10612 -3282
rect 10578 -3726 10612 -3710
rect 10696 -3334 10730 -3318
rect 10696 -3761 10730 -3710
rect 10814 -3334 10848 -3282
rect 11050 -3282 11320 -3243
rect 10814 -3726 10848 -3710
rect 10932 -3334 10966 -3318
rect 10932 -3761 10966 -3710
rect 11050 -3334 11084 -3282
rect 11050 -3726 11084 -3710
rect 11168 -3334 11202 -3318
rect 11168 -3761 11202 -3710
rect 11286 -3334 11320 -3282
rect 11523 -3282 11793 -3243
rect 11286 -3726 11320 -3710
rect 11405 -3334 11439 -3318
rect 11405 -3761 11439 -3710
rect 11523 -3334 11557 -3282
rect 11523 -3726 11557 -3710
rect 11641 -3334 11675 -3318
rect 11641 -3761 11675 -3710
rect 11759 -3334 11793 -3282
rect 13313 -3285 13583 -3246
rect 13313 -3338 13347 -3285
rect 11996 -3484 12266 -3447
rect 11759 -3726 11793 -3710
rect 11878 -3534 11912 -3518
rect 10229 -3800 11675 -3761
rect 11878 -3764 11912 -3710
rect 11996 -3534 12030 -3484
rect 11996 -3726 12030 -3710
rect 12114 -3534 12148 -3518
rect 12114 -3764 12148 -3710
rect 12232 -3534 12266 -3484
rect 12232 -3726 12266 -3710
rect 12872 -3487 13142 -3448
rect 12872 -3538 12906 -3487
rect 12872 -3730 12906 -3714
rect 12990 -3538 13024 -3522
rect 11878 -3803 12148 -3764
rect 12990 -3765 13024 -3714
rect 13108 -3538 13142 -3487
rect 13108 -3730 13142 -3714
rect 13226 -3538 13260 -3522
rect 13226 -3765 13260 -3714
rect 13313 -3730 13347 -3714
rect 13431 -3338 13465 -3322
rect 12990 -3804 13260 -3765
rect 13431 -3765 13465 -3714
rect 13549 -3338 13583 -3285
rect 13780 -3286 14050 -3247
rect 13549 -3730 13583 -3714
rect 13667 -3338 13701 -3322
rect 13667 -3765 13701 -3714
rect 13780 -3338 13814 -3286
rect 13780 -3730 13814 -3714
rect 13898 -3338 13932 -3322
rect 13898 -3765 13932 -3714
rect 14016 -3338 14050 -3286
rect 14252 -3286 14522 -3247
rect 14016 -3730 14050 -3714
rect 14134 -3338 14168 -3322
rect 14134 -3765 14168 -3714
rect 14252 -3338 14286 -3286
rect 14252 -3730 14286 -3714
rect 14370 -3338 14404 -3322
rect 14370 -3765 14404 -3714
rect 14488 -3338 14522 -3286
rect 14725 -3286 14995 -3247
rect 14488 -3730 14522 -3714
rect 14607 -3338 14641 -3322
rect 14607 -3765 14641 -3714
rect 14725 -3338 14759 -3286
rect 14725 -3730 14759 -3714
rect 14843 -3338 14877 -3322
rect 14843 -3765 14877 -3714
rect 14961 -3338 14995 -3286
rect 16457 -3285 16727 -3246
rect 16457 -3338 16491 -3285
rect 15198 -3488 15468 -3451
rect 14961 -3730 14995 -3714
rect 15080 -3538 15114 -3522
rect 13431 -3804 14877 -3765
rect 15080 -3768 15114 -3714
rect 15198 -3538 15232 -3488
rect 15198 -3730 15232 -3714
rect 15316 -3538 15350 -3522
rect 15316 -3768 15350 -3714
rect 15434 -3538 15468 -3488
rect 15434 -3730 15468 -3714
rect 16016 -3487 16286 -3448
rect 16016 -3538 16050 -3487
rect 16016 -3730 16050 -3714
rect 16134 -3538 16168 -3522
rect 15080 -3807 15350 -3768
rect 16134 -3765 16168 -3714
rect 16252 -3538 16286 -3487
rect 16252 -3730 16286 -3714
rect 16370 -3538 16404 -3522
rect 16370 -3765 16404 -3714
rect 16457 -3730 16491 -3714
rect 16575 -3338 16609 -3322
rect 16134 -3804 16404 -3765
rect 16575 -3765 16609 -3714
rect 16693 -3338 16727 -3285
rect 16924 -3286 17194 -3247
rect 16693 -3730 16727 -3714
rect 16811 -3338 16845 -3322
rect 16811 -3765 16845 -3714
rect 16924 -3338 16958 -3286
rect 16924 -3730 16958 -3714
rect 17042 -3338 17076 -3322
rect 17042 -3765 17076 -3714
rect 17160 -3338 17194 -3286
rect 17396 -3286 17666 -3247
rect 17160 -3730 17194 -3714
rect 17278 -3338 17312 -3322
rect 17278 -3765 17312 -3714
rect 17396 -3338 17430 -3286
rect 17396 -3730 17430 -3714
rect 17514 -3338 17548 -3322
rect 17514 -3765 17548 -3714
rect 17632 -3338 17666 -3286
rect 17869 -3286 18139 -3247
rect 17632 -3730 17666 -3714
rect 17751 -3338 17785 -3322
rect 17751 -3765 17785 -3714
rect 17869 -3338 17903 -3286
rect 17869 -3730 17903 -3714
rect 17987 -3338 18021 -3322
rect 17987 -3765 18021 -3714
rect 18105 -3338 18139 -3286
rect 19589 -3281 19859 -3242
rect 19589 -3334 19623 -3281
rect 18342 -3488 18612 -3451
rect 18105 -3730 18139 -3714
rect 18224 -3538 18258 -3522
rect 16575 -3804 18021 -3765
rect 18224 -3768 18258 -3714
rect 18342 -3538 18376 -3488
rect 18342 -3730 18376 -3714
rect 18460 -3538 18494 -3522
rect 18460 -3768 18494 -3714
rect 18578 -3538 18612 -3488
rect 18578 -3730 18612 -3714
rect 19148 -3483 19418 -3444
rect 19148 -3534 19182 -3483
rect 19148 -3726 19182 -3710
rect 19266 -3534 19300 -3518
rect 18224 -3807 18494 -3768
rect 19266 -3761 19300 -3710
rect 19384 -3534 19418 -3483
rect 19384 -3726 19418 -3710
rect 19502 -3534 19536 -3518
rect 19502 -3761 19536 -3710
rect 19589 -3726 19623 -3710
rect 19707 -3334 19741 -3318
rect 19266 -3800 19536 -3761
rect 19707 -3761 19741 -3710
rect 19825 -3334 19859 -3281
rect 20056 -3282 20326 -3243
rect 19825 -3726 19859 -3710
rect 19943 -3334 19977 -3318
rect 19943 -3761 19977 -3710
rect 20056 -3334 20090 -3282
rect 20056 -3726 20090 -3710
rect 20174 -3334 20208 -3318
rect 20174 -3761 20208 -3710
rect 20292 -3334 20326 -3282
rect 20528 -3282 20798 -3243
rect 20292 -3726 20326 -3710
rect 20410 -3334 20444 -3318
rect 20410 -3761 20444 -3710
rect 20528 -3334 20562 -3282
rect 20528 -3726 20562 -3710
rect 20646 -3334 20680 -3318
rect 20646 -3761 20680 -3710
rect 20764 -3334 20798 -3282
rect 21001 -3282 21271 -3243
rect 20764 -3726 20798 -3710
rect 20883 -3334 20917 -3318
rect 20883 -3761 20917 -3710
rect 21001 -3334 21035 -3282
rect 21001 -3726 21035 -3710
rect 21119 -3334 21153 -3318
rect 21119 -3761 21153 -3710
rect 21237 -3334 21271 -3282
rect 22733 -3281 23003 -3242
rect 22733 -3334 22767 -3281
rect 21474 -3484 21744 -3447
rect 21237 -3726 21271 -3710
rect 21356 -3534 21390 -3518
rect 19707 -3800 21153 -3761
rect 21356 -3764 21390 -3710
rect 21474 -3534 21508 -3484
rect 21474 -3726 21508 -3710
rect 21592 -3534 21626 -3518
rect 21592 -3764 21626 -3710
rect 21710 -3534 21744 -3484
rect 21710 -3726 21744 -3710
rect 22292 -3483 22562 -3444
rect 22292 -3534 22326 -3483
rect 22292 -3726 22326 -3710
rect 22410 -3534 22444 -3518
rect 21356 -3803 21626 -3764
rect 22410 -3761 22444 -3710
rect 22528 -3534 22562 -3483
rect 22528 -3726 22562 -3710
rect 22646 -3534 22680 -3518
rect 22646 -3761 22680 -3710
rect 22733 -3726 22767 -3710
rect 22851 -3334 22885 -3318
rect 22410 -3800 22680 -3761
rect 22851 -3761 22885 -3710
rect 22969 -3334 23003 -3281
rect 23200 -3282 23470 -3243
rect 22969 -3726 23003 -3710
rect 23087 -3334 23121 -3318
rect 23087 -3761 23121 -3710
rect 23200 -3334 23234 -3282
rect 23200 -3726 23234 -3710
rect 23318 -3334 23352 -3318
rect 23318 -3761 23352 -3710
rect 23436 -3334 23470 -3282
rect 23672 -3282 23942 -3243
rect 23436 -3726 23470 -3710
rect 23554 -3334 23588 -3318
rect 23554 -3761 23588 -3710
rect 23672 -3334 23706 -3282
rect 23672 -3726 23706 -3710
rect 23790 -3334 23824 -3318
rect 23790 -3761 23824 -3710
rect 23908 -3334 23942 -3282
rect 24145 -3282 24415 -3243
rect 23908 -3726 23942 -3710
rect 24027 -3334 24061 -3318
rect 24027 -3761 24061 -3710
rect 24145 -3334 24179 -3282
rect 24145 -3726 24179 -3710
rect 24263 -3334 24297 -3318
rect 24263 -3761 24297 -3710
rect 24381 -3334 24415 -3282
rect 24618 -3484 24888 -3447
rect 24381 -3726 24415 -3710
rect 24500 -3534 24534 -3518
rect 22851 -3800 24297 -3761
rect 24500 -3764 24534 -3710
rect 24618 -3534 24652 -3484
rect 24618 -3726 24652 -3710
rect 24736 -3534 24770 -3518
rect 24736 -3764 24770 -3710
rect 24854 -3534 24888 -3484
rect 24854 -3726 24888 -3710
rect 24500 -3803 24770 -3764
rect 1336 -3929 1370 -3913
rect 2630 -3922 2646 -3888
rect 2680 -3922 2696 -3888
rect 1336 -3979 1370 -3963
rect 4480 -3929 4514 -3913
rect 5774 -3922 5790 -3888
rect 5824 -3922 5840 -3888
rect 4480 -3979 4514 -3963
rect 7612 -3925 7646 -3909
rect 8906 -3918 8922 -3884
rect 8956 -3918 8972 -3884
rect 7612 -3975 7646 -3959
rect 10756 -3925 10790 -3909
rect 12050 -3918 12066 -3884
rect 12100 -3918 12116 -3884
rect 10756 -3975 10790 -3959
rect 13958 -3929 13992 -3913
rect 15252 -3922 15268 -3888
rect 15302 -3922 15318 -3888
rect 13958 -3979 13992 -3963
rect 17102 -3929 17136 -3913
rect 18396 -3922 18412 -3888
rect 18446 -3922 18462 -3888
rect 17102 -3979 17136 -3963
rect 20234 -3925 20268 -3909
rect 21528 -3918 21544 -3884
rect 21578 -3918 21594 -3884
rect 20234 -3975 20268 -3959
rect 23378 -3925 23412 -3909
rect 24672 -3918 24688 -3884
rect 24722 -3918 24738 -3884
rect 23378 -3975 23412 -3959
rect 107 -4028 164 -4024
rect 107 -4088 111 -4028
rect 160 -4088 164 -4028
rect 107 -4092 164 -4088
rect 339 -4029 431 -4012
rect 339 -4084 355 -4029
rect 415 -4084 431 -4029
rect 339 -4097 431 -4084
rect 1424 -4028 1516 -4015
rect 1424 -4083 1440 -4028
rect 1500 -4083 1516 -4028
rect 1424 -4100 1516 -4083
rect 3251 -4028 3308 -4024
rect 3251 -4088 3255 -4028
rect 3304 -4088 3308 -4028
rect 3251 -4092 3308 -4088
rect 3483 -4029 3575 -4012
rect 3483 -4084 3499 -4029
rect 3559 -4084 3575 -4029
rect 3483 -4097 3575 -4084
rect 4568 -4028 4660 -4015
rect 4568 -4083 4584 -4028
rect 4644 -4083 4660 -4028
rect 4568 -4100 4660 -4083
rect 6383 -4024 6440 -4020
rect 6383 -4084 6387 -4024
rect 6436 -4084 6440 -4024
rect 6383 -4088 6440 -4084
rect 6615 -4025 6707 -4008
rect 6615 -4080 6631 -4025
rect 6691 -4080 6707 -4025
rect 6615 -4093 6707 -4080
rect 7700 -4024 7792 -4011
rect 7700 -4079 7716 -4024
rect 7776 -4079 7792 -4024
rect 7700 -4096 7792 -4079
rect 9527 -4024 9584 -4020
rect 9527 -4084 9531 -4024
rect 9580 -4084 9584 -4024
rect 9527 -4088 9584 -4084
rect 9759 -4025 9851 -4008
rect 9759 -4080 9775 -4025
rect 9835 -4080 9851 -4025
rect 9759 -4093 9851 -4080
rect 10844 -4024 10936 -4011
rect 10844 -4079 10860 -4024
rect 10920 -4079 10936 -4024
rect 10844 -4096 10936 -4079
rect 12729 -4028 12786 -4024
rect 12729 -4088 12733 -4028
rect 12782 -4088 12786 -4028
rect 12729 -4092 12786 -4088
rect 12961 -4029 13053 -4012
rect 12961 -4084 12977 -4029
rect 13037 -4084 13053 -4029
rect 12961 -4097 13053 -4084
rect 14046 -4028 14138 -4015
rect 14046 -4083 14062 -4028
rect 14122 -4083 14138 -4028
rect 14046 -4100 14138 -4083
rect 15873 -4028 15930 -4024
rect 15873 -4088 15877 -4028
rect 15926 -4088 15930 -4028
rect 15873 -4092 15930 -4088
rect 16105 -4029 16197 -4012
rect 16105 -4084 16121 -4029
rect 16181 -4084 16197 -4029
rect 16105 -4097 16197 -4084
rect 17190 -4028 17282 -4015
rect 17190 -4083 17206 -4028
rect 17266 -4083 17282 -4028
rect 17190 -4100 17282 -4083
rect 19005 -4024 19062 -4020
rect 19005 -4084 19009 -4024
rect 19058 -4084 19062 -4024
rect 19005 -4088 19062 -4084
rect 19237 -4025 19329 -4008
rect 19237 -4080 19253 -4025
rect 19313 -4080 19329 -4025
rect 19237 -4093 19329 -4080
rect 20322 -4024 20414 -4011
rect 20322 -4079 20338 -4024
rect 20398 -4079 20414 -4024
rect 20322 -4096 20414 -4079
rect 22149 -4024 22206 -4020
rect 22149 -4084 22153 -4024
rect 22202 -4084 22206 -4024
rect 22149 -4088 22206 -4084
rect 22381 -4025 22473 -4008
rect 22381 -4080 22397 -4025
rect 22457 -4080 22473 -4025
rect 22381 -4093 22473 -4080
rect 23466 -4024 23558 -4011
rect 23466 -4079 23482 -4024
rect 23542 -4079 23558 -4024
rect 23466 -4096 23558 -4079
rect 6383 -4138 6440 -4136
rect 6185 -4140 6440 -4138
rect 9527 -4139 9584 -4136
rect 19005 -4138 19062 -4136
rect -173 -4144 -57 -4143
rect 107 -4144 164 -4140
rect 3251 -4142 3308 -4140
rect -173 -4204 111 -4144
rect 160 -4204 164 -4144
rect -173 -4208 164 -4204
rect 1690 -4159 1724 -4143
rect -172 -5770 -108 -4208
rect 1690 -4209 1724 -4193
rect 3055 -4144 3308 -4142
rect 3055 -4204 3255 -4144
rect 3304 -4204 3308 -4144
rect 3055 -4206 3308 -4204
rect 107 -4312 164 -4308
rect 107 -4372 111 -4312
rect 160 -4372 164 -4312
rect 107 -4376 164 -4372
rect 1306 -4313 1398 -4300
rect 1306 -4368 1322 -4313
rect 1382 -4368 1398 -4313
rect 1306 -4385 1398 -4368
rect 1571 -4549 1605 -4533
rect 1571 -4599 1605 -4583
rect 1084 -4671 1118 -4655
rect 1084 -4863 1118 -4847
rect 1202 -4659 1236 -4655
rect 1276 -4659 1310 -4655
rect 1202 -4671 1310 -4659
rect 1236 -4847 1276 -4671
rect 1202 -4859 1276 -4847
rect 1202 -4863 1236 -4859
rect 1276 -5063 1310 -5047
rect 1394 -4671 1428 -4655
rect 1394 -5063 1428 -5047
rect 1512 -4671 1546 -4655
rect 1512 -5063 1546 -5047
rect 1630 -4671 1664 -4655
rect 1630 -5063 1664 -5047
rect 1748 -4659 1782 -4655
rect 1826 -4659 1860 -4655
rect 1748 -4671 1860 -4659
rect 1782 -4847 1826 -4671
rect 1782 -4859 1860 -4847
rect 1826 -4863 1860 -4859
rect 1944 -4671 1978 -4655
rect 1944 -4863 1978 -4847
rect 1748 -5063 1782 -5047
rect 1497 -5182 1513 -5148
rect 1547 -5182 1563 -5148
rect 1478 -5300 1614 -5296
rect 1478 -5314 1516 -5300
rect 1574 -5314 1614 -5300
rect 1478 -5360 1494 -5314
rect 1598 -5360 1614 -5314
rect 1478 -5382 1614 -5360
rect -172 -5834 1827 -5770
rect 738 -6012 940 -5992
rect 738 -6056 772 -6012
rect 894 -6056 940 -6012
rect 738 -6066 824 -6056
rect 862 -6066 940 -6056
rect 738 -6084 940 -6066
rect 825 -6230 1095 -6195
rect 471 -6283 505 -6267
rect -13 -6429 257 -6394
rect -13 -6483 21 -6429
rect -13 -6675 21 -6659
rect 105 -6483 139 -6467
rect 105 -6675 139 -6659
rect 223 -6483 257 -6429
rect 223 -6675 257 -6659
rect 341 -6483 375 -6467
rect 341 -6675 375 -6659
rect 471 -6675 505 -6659
rect 589 -6283 623 -6267
rect 589 -6675 623 -6659
rect 707 -6283 741 -6267
rect 707 -6675 741 -6659
rect 825 -6283 859 -6230
rect 825 -6675 859 -6659
rect 943 -6283 977 -6267
rect 943 -6675 977 -6659
rect 1061 -6283 1095 -6230
rect 1061 -6675 1095 -6659
rect 1179 -6283 1213 -6267
rect 1179 -6675 1213 -6659
rect 1308 -6483 1342 -6467
rect 1308 -6675 1342 -6659
rect 1426 -6483 1460 -6467
rect 1426 -6675 1460 -6659
rect 1544 -6483 1578 -6467
rect 1544 -6675 1578 -6659
rect 1662 -6483 1696 -6467
rect 1662 -6675 1696 -6659
rect 1388 -6872 1394 -6838
rect 1448 -6872 1454 -6838
rect 414 -6976 448 -6960
rect -43 -7078 -6 -7018
rect -43 -7134 22 -7078
rect -43 -8560 21 -7134
rect 532 -6976 566 -6960
rect 414 -7368 448 -7352
rect 531 -7352 532 -7305
rect 650 -6976 684 -6960
rect 566 -7352 567 -7305
rect 531 -7410 567 -7352
rect 768 -6976 802 -6960
rect 650 -7368 684 -7352
rect 766 -7352 768 -7305
rect 766 -7410 802 -7352
rect 886 -6976 920 -6960
rect 886 -7368 920 -7352
rect 1004 -6976 1038 -6960
rect 1122 -6976 1156 -6960
rect 1038 -7352 1040 -7306
rect 1004 -7410 1040 -7352
rect 1122 -7368 1156 -7352
rect 531 -7450 1626 -7410
rect 550 -7451 1626 -7450
rect 428 -7540 495 -7524
rect 428 -7574 444 -7540
rect 478 -7574 495 -7540
rect 428 -7590 495 -7574
rect 259 -7607 293 -7591
rect 259 -7657 293 -7641
rect 605 -7692 639 -7451
rect 1763 -7397 1827 -5834
rect 3055 -5786 3119 -4206
rect 3251 -4208 3308 -4206
rect 4834 -4159 4868 -4143
rect 4834 -4209 4868 -4193
rect 6185 -4200 6387 -4140
rect 6436 -4200 6440 -4140
rect 6185 -4202 6440 -4200
rect 3251 -4312 3308 -4308
rect 3251 -4372 3255 -4312
rect 3304 -4372 3308 -4312
rect 3251 -4376 3308 -4372
rect 4450 -4313 4542 -4300
rect 4450 -4368 4466 -4313
rect 4526 -4368 4542 -4313
rect 4450 -4385 4542 -4368
rect 4715 -4549 4749 -4533
rect 4715 -4599 4749 -4583
rect 6185 -4642 6249 -4202
rect 6383 -4204 6440 -4202
rect 7966 -4155 8000 -4139
rect 7966 -4205 8000 -4189
rect 9311 -4140 9584 -4139
rect 9311 -4200 9531 -4140
rect 9580 -4200 9584 -4140
rect 9311 -4203 9584 -4200
rect 6383 -4308 6440 -4304
rect 6383 -4368 6387 -4308
rect 6436 -4368 6440 -4308
rect 6383 -4372 6440 -4368
rect 7582 -4309 7674 -4296
rect 7582 -4364 7598 -4309
rect 7658 -4364 7674 -4309
rect 7582 -4381 7674 -4364
rect 7847 -4545 7881 -4529
rect 7847 -4595 7881 -4579
rect 4228 -4671 4262 -4655
rect 4228 -4863 4262 -4847
rect 4346 -4659 4380 -4655
rect 4420 -4659 4454 -4655
rect 4346 -4671 4454 -4659
rect 4380 -4847 4420 -4671
rect 4346 -4859 4420 -4847
rect 4346 -4863 4380 -4859
rect 4420 -5063 4454 -5047
rect 4538 -4671 4572 -4655
rect 4538 -5063 4572 -5047
rect 4656 -4671 4690 -4655
rect 4656 -5063 4690 -5047
rect 4774 -4671 4808 -4655
rect 4774 -5063 4808 -5047
rect 4892 -4659 4926 -4655
rect 4970 -4659 5004 -4655
rect 4892 -4671 5004 -4659
rect 4926 -4847 4970 -4671
rect 4926 -4859 5004 -4847
rect 4970 -4863 5004 -4859
rect 5088 -4671 5122 -4655
rect 5088 -4863 5122 -4847
rect 5924 -4706 6249 -4642
rect 7360 -4667 7394 -4651
rect 4892 -5063 4926 -5047
rect 4641 -5182 4657 -5148
rect 4691 -5182 4707 -5148
rect 4622 -5300 4758 -5296
rect 4622 -5314 4660 -5300
rect 4718 -5314 4758 -5300
rect 4622 -5360 4638 -5314
rect 4742 -5360 4758 -5314
rect 4622 -5382 4758 -5360
rect 3055 -5850 3893 -5786
rect 2806 -6010 3008 -5990
rect 2806 -6054 2840 -6010
rect 2962 -6054 3008 -6010
rect 2806 -6064 2892 -6054
rect 2930 -6064 3008 -6054
rect 2806 -6082 3008 -6064
rect 2893 -6228 3163 -6193
rect 2539 -6281 2573 -6265
rect 2055 -6427 2325 -6392
rect 2055 -6481 2089 -6427
rect 2055 -6673 2089 -6657
rect 2173 -6481 2207 -6465
rect 2173 -6673 2207 -6657
rect 2291 -6481 2325 -6427
rect 2291 -6673 2325 -6657
rect 2409 -6481 2443 -6465
rect 2409 -6673 2443 -6657
rect 2539 -6673 2573 -6657
rect 2657 -6281 2691 -6265
rect 2657 -6673 2691 -6657
rect 2775 -6281 2809 -6265
rect 2775 -6673 2809 -6657
rect 2893 -6281 2927 -6228
rect 2893 -6673 2927 -6657
rect 3011 -6281 3045 -6265
rect 3011 -6673 3045 -6657
rect 3129 -6281 3163 -6228
rect 3129 -6673 3163 -6657
rect 3247 -6281 3281 -6265
rect 3247 -6673 3281 -6657
rect 3376 -6481 3410 -6465
rect 3376 -6673 3410 -6657
rect 3494 -6481 3528 -6465
rect 3494 -6673 3528 -6657
rect 3612 -6481 3646 -6465
rect 3612 -6673 3646 -6657
rect 3730 -6481 3764 -6465
rect 3730 -6673 3764 -6657
rect 3456 -6870 3462 -6836
rect 3516 -6870 3522 -6836
rect 2482 -6974 2516 -6958
rect 2600 -6974 2634 -6958
rect 2482 -7366 2516 -7350
rect 2599 -7350 2600 -7303
rect 2718 -6974 2752 -6958
rect 2634 -7350 2635 -7303
rect 1728 -7461 1827 -7397
rect 2599 -7408 2635 -7350
rect 2836 -6974 2870 -6958
rect 2718 -7366 2752 -7350
rect 2834 -7350 2836 -7303
rect 2834 -7408 2870 -7350
rect 2954 -6974 2988 -6958
rect 2954 -7366 2988 -7350
rect 3072 -6974 3106 -6958
rect 3190 -6974 3224 -6958
rect 3106 -7350 3108 -7304
rect 3072 -7408 3108 -7350
rect 3190 -7366 3224 -7350
rect 2599 -7448 3694 -7408
rect 2618 -7449 3694 -7448
rect 1075 -7540 1142 -7524
rect 1075 -7574 1092 -7540
rect 1126 -7574 1142 -7540
rect 1075 -7590 1142 -7574
rect 2496 -7538 2563 -7522
rect 2496 -7572 2512 -7538
rect 2546 -7572 2563 -7538
rect 2496 -7588 2563 -7572
rect 1382 -7608 1416 -7592
rect 694 -7658 710 -7624
rect 744 -7658 760 -7624
rect 812 -7657 828 -7623
rect 862 -7657 878 -7623
rect 1382 -7658 1416 -7642
rect 2327 -7605 2361 -7589
rect 2327 -7655 2361 -7639
rect 2673 -7690 2707 -7449
rect 3836 -7408 3892 -5850
rect 4875 -6012 5077 -5992
rect 4875 -6056 4909 -6012
rect 5031 -6056 5077 -6012
rect 4875 -6066 4961 -6056
rect 4999 -6066 5077 -6056
rect 4875 -6084 5077 -6066
rect 4962 -6230 5232 -6195
rect 4608 -6283 4642 -6267
rect 4124 -6429 4394 -6394
rect 4124 -6483 4158 -6429
rect 4124 -6675 4158 -6659
rect 4242 -6483 4276 -6467
rect 4242 -6675 4276 -6659
rect 4360 -6483 4394 -6429
rect 4360 -6675 4394 -6659
rect 4478 -6483 4512 -6467
rect 4478 -6675 4512 -6659
rect 4608 -6675 4642 -6659
rect 4726 -6283 4760 -6267
rect 4726 -6675 4760 -6659
rect 4844 -6283 4878 -6267
rect 4844 -6675 4878 -6659
rect 4962 -6283 4996 -6230
rect 4962 -6675 4996 -6659
rect 5080 -6283 5114 -6267
rect 5080 -6675 5114 -6659
rect 5198 -6283 5232 -6230
rect 5198 -6675 5232 -6659
rect 5316 -6283 5350 -6267
rect 5316 -6675 5350 -6659
rect 5445 -6483 5479 -6467
rect 5445 -6675 5479 -6659
rect 5563 -6483 5597 -6467
rect 5563 -6675 5597 -6659
rect 5681 -6483 5715 -6467
rect 5681 -6675 5715 -6659
rect 5799 -6483 5833 -6467
rect 5799 -6675 5833 -6659
rect 5525 -6872 5531 -6838
rect 5585 -6872 5591 -6838
rect 4551 -6976 4585 -6960
rect 4669 -6976 4703 -6960
rect 4551 -7368 4585 -7352
rect 4668 -7352 4669 -7305
rect 4787 -6976 4821 -6960
rect 4703 -7352 4704 -7305
rect 3796 -7449 3892 -7408
rect 4668 -7410 4704 -7352
rect 4905 -6976 4939 -6960
rect 4787 -7368 4821 -7352
rect 4903 -7352 4905 -7305
rect 4903 -7410 4939 -7352
rect 5023 -6976 5057 -6960
rect 5023 -7368 5057 -7352
rect 5141 -6976 5175 -6960
rect 5259 -6976 5293 -6960
rect 5175 -7352 5177 -7306
rect 5141 -7410 5177 -7352
rect 5259 -7368 5293 -7352
rect 4668 -7450 5763 -7410
rect 4687 -7451 5763 -7450
rect 3143 -7538 3210 -7522
rect 3143 -7572 3160 -7538
rect 3194 -7572 3210 -7538
rect 3143 -7588 3210 -7572
rect 4565 -7540 4632 -7524
rect 4565 -7574 4581 -7540
rect 4615 -7574 4632 -7540
rect 4565 -7590 4632 -7574
rect 3450 -7606 3484 -7590
rect 2762 -7656 2778 -7622
rect 2812 -7656 2828 -7622
rect 2880 -7655 2896 -7621
rect 2930 -7655 2946 -7621
rect 3450 -7656 3484 -7640
rect 4396 -7607 4430 -7591
rect 4396 -7657 4430 -7641
rect 112 -7708 146 -7692
rect 112 -7900 146 -7884
rect 230 -7708 264 -7692
rect 230 -7900 264 -7884
rect 532 -7708 566 -7692
rect 605 -7708 684 -7692
rect 605 -7738 650 -7708
rect 532 -8151 567 -8084
rect 650 -8100 684 -8084
rect 768 -7708 802 -7692
rect 768 -8100 802 -8084
rect 886 -7708 920 -7692
rect 1004 -7708 1038 -7692
rect 1410 -7708 1444 -7692
rect 1410 -7900 1444 -7884
rect 1528 -7708 1562 -7692
rect 1528 -7900 1562 -7884
rect 2180 -7706 2214 -7690
rect 2180 -7898 2214 -7882
rect 2298 -7706 2332 -7690
rect 2298 -7898 2332 -7882
rect 2600 -7706 2634 -7690
rect 886 -8100 920 -8084
rect 1003 -8151 1038 -8084
rect 532 -8186 1038 -8151
rect 2673 -7706 2752 -7690
rect 2673 -7736 2718 -7706
rect 2600 -8149 2635 -8082
rect 2718 -8098 2752 -8082
rect 2836 -7706 2870 -7690
rect 2836 -8098 2870 -8082
rect 2954 -7706 2988 -7690
rect 3072 -7706 3106 -7690
rect 3478 -7706 3512 -7690
rect 3478 -7898 3512 -7882
rect 3596 -7706 3630 -7690
rect 4742 -7692 4776 -7451
rect 5924 -7399 5988 -4706
rect 7360 -4859 7394 -4843
rect 7478 -4655 7512 -4651
rect 7552 -4655 7586 -4651
rect 7478 -4667 7586 -4655
rect 7512 -4843 7552 -4667
rect 7478 -4855 7552 -4843
rect 7478 -4859 7512 -4855
rect 7552 -5059 7586 -5043
rect 7670 -4667 7704 -4651
rect 7670 -5059 7704 -5043
rect 7788 -4667 7822 -4651
rect 7788 -5059 7822 -5043
rect 7906 -4667 7940 -4651
rect 7906 -5059 7940 -5043
rect 8024 -4655 8058 -4651
rect 8102 -4655 8136 -4651
rect 8024 -4667 8136 -4655
rect 8058 -4843 8102 -4667
rect 8058 -4855 8136 -4843
rect 8102 -4859 8136 -4855
rect 8220 -4667 8254 -4651
rect 8220 -4859 8254 -4843
rect 8024 -5059 8058 -5043
rect 7773 -5178 7789 -5144
rect 7823 -5178 7839 -5144
rect 7754 -5296 7890 -5292
rect 7754 -5310 7792 -5296
rect 7850 -5310 7890 -5296
rect 7754 -5356 7770 -5310
rect 7874 -5356 7890 -5310
rect 7754 -5378 7890 -5356
rect 9311 -5468 9375 -4203
rect 9527 -4204 9584 -4203
rect 11110 -4155 11144 -4139
rect 18789 -4140 19062 -4138
rect 12729 -4142 12786 -4140
rect 15873 -4141 15930 -4140
rect 11110 -4205 11144 -4189
rect 12485 -4144 12787 -4142
rect 12485 -4204 12733 -4144
rect 12782 -4204 12787 -4144
rect 12485 -4206 12787 -4204
rect 14312 -4159 14346 -4143
rect 9527 -4308 9584 -4304
rect 9527 -4368 9531 -4308
rect 9580 -4368 9584 -4308
rect 9527 -4372 9584 -4368
rect 10726 -4309 10818 -4296
rect 10726 -4364 10742 -4309
rect 10802 -4364 10818 -4309
rect 10726 -4381 10818 -4364
rect 10991 -4545 11025 -4529
rect 10991 -4595 11025 -4579
rect 10504 -4667 10538 -4651
rect 10504 -4859 10538 -4843
rect 10622 -4655 10656 -4651
rect 10696 -4655 10730 -4651
rect 10622 -4667 10730 -4655
rect 10656 -4843 10696 -4667
rect 10622 -4855 10696 -4843
rect 10622 -4859 10656 -4855
rect 10696 -5059 10730 -5043
rect 10814 -4667 10848 -4651
rect 10814 -5059 10848 -5043
rect 10932 -4667 10966 -4651
rect 10932 -5059 10966 -5043
rect 11050 -4667 11084 -4651
rect 11050 -5059 11084 -5043
rect 11168 -4655 11202 -4651
rect 11246 -4655 11280 -4651
rect 11168 -4667 11280 -4655
rect 11202 -4843 11246 -4667
rect 11202 -4855 11280 -4843
rect 11246 -4859 11280 -4855
rect 11364 -4667 11398 -4651
rect 11364 -4859 11398 -4843
rect 11168 -5059 11202 -5043
rect 10917 -5178 10933 -5144
rect 10967 -5178 10983 -5144
rect 10898 -5296 11034 -5292
rect 10898 -5310 10936 -5296
rect 10994 -5310 11034 -5296
rect 10898 -5356 10914 -5310
rect 11018 -5356 11034 -5310
rect 10898 -5378 11034 -5356
rect 12485 -5441 12549 -4206
rect 12729 -4208 12786 -4206
rect 14312 -4209 14346 -4193
rect 15647 -4144 15930 -4141
rect 15647 -4204 15877 -4144
rect 15926 -4204 15930 -4144
rect 15647 -4205 15930 -4204
rect 12729 -4312 12786 -4308
rect 12729 -4372 12733 -4312
rect 12782 -4372 12786 -4312
rect 12729 -4376 12786 -4372
rect 13928 -4313 14020 -4300
rect 13928 -4368 13944 -4313
rect 14004 -4368 14020 -4313
rect 13928 -4385 14020 -4368
rect 14193 -4549 14227 -4533
rect 14193 -4599 14227 -4583
rect 13706 -4671 13740 -4655
rect 13706 -4863 13740 -4847
rect 13824 -4659 13858 -4655
rect 13898 -4659 13932 -4655
rect 13824 -4671 13932 -4659
rect 13858 -4847 13898 -4671
rect 13824 -4859 13898 -4847
rect 13824 -4863 13858 -4859
rect 13898 -5063 13932 -5047
rect 14016 -4671 14050 -4655
rect 14016 -5063 14050 -5047
rect 14134 -4671 14168 -4655
rect 14134 -5063 14168 -5047
rect 14252 -4671 14286 -4655
rect 14252 -5063 14286 -5047
rect 14370 -4659 14404 -4655
rect 14448 -4659 14482 -4655
rect 14370 -4671 14482 -4659
rect 14404 -4847 14448 -4671
rect 14404 -4859 14482 -4847
rect 14448 -4863 14482 -4859
rect 14566 -4671 14600 -4655
rect 14566 -4863 14600 -4847
rect 14370 -5063 14404 -5047
rect 14119 -5182 14135 -5148
rect 14169 -5182 14185 -5148
rect 14100 -5300 14236 -5296
rect 14100 -5314 14138 -5300
rect 14196 -5314 14236 -5300
rect 14100 -5360 14116 -5314
rect 14220 -5360 14236 -5314
rect 14100 -5382 14236 -5360
rect 8005 -5532 9375 -5468
rect 10071 -5505 12549 -5441
rect 6943 -6010 7145 -5990
rect 6943 -6054 6977 -6010
rect 7099 -6054 7145 -6010
rect 6943 -6064 7029 -6054
rect 7067 -6064 7145 -6054
rect 6943 -6082 7145 -6064
rect 7030 -6228 7300 -6193
rect 6676 -6281 6710 -6265
rect 6192 -6427 6462 -6392
rect 6192 -6481 6226 -6427
rect 6192 -6673 6226 -6657
rect 6310 -6481 6344 -6465
rect 6310 -6673 6344 -6657
rect 6428 -6481 6462 -6427
rect 6428 -6673 6462 -6657
rect 6546 -6481 6580 -6465
rect 6546 -6673 6580 -6657
rect 6676 -6673 6710 -6657
rect 6794 -6281 6828 -6265
rect 6794 -6673 6828 -6657
rect 6912 -6281 6946 -6265
rect 6912 -6673 6946 -6657
rect 7030 -6281 7064 -6228
rect 7030 -6673 7064 -6657
rect 7148 -6281 7182 -6265
rect 7148 -6673 7182 -6657
rect 7266 -6281 7300 -6228
rect 7266 -6673 7300 -6657
rect 7384 -6281 7418 -6265
rect 7384 -6673 7418 -6657
rect 7513 -6481 7547 -6465
rect 7513 -6673 7547 -6657
rect 7631 -6481 7665 -6465
rect 7631 -6673 7665 -6657
rect 7749 -6481 7783 -6465
rect 7749 -6673 7783 -6657
rect 7867 -6481 7901 -6465
rect 7867 -6673 7901 -6657
rect 7593 -6870 7599 -6836
rect 7653 -6870 7659 -6836
rect 6619 -6974 6653 -6958
rect 6737 -6974 6771 -6958
rect 6619 -7366 6653 -7350
rect 6736 -7350 6737 -7303
rect 6855 -6974 6889 -6958
rect 6771 -7350 6772 -7303
rect 5865 -7463 5988 -7399
rect 6736 -7408 6772 -7350
rect 6973 -6974 7007 -6958
rect 6855 -7366 6889 -7350
rect 6971 -7350 6973 -7303
rect 6971 -7408 7007 -7350
rect 7091 -6974 7125 -6958
rect 7091 -7366 7125 -7350
rect 7209 -6974 7243 -6958
rect 7327 -6974 7361 -6958
rect 7243 -7350 7245 -7304
rect 7209 -7408 7245 -7350
rect 7327 -7366 7361 -7350
rect 6736 -7448 7831 -7408
rect 6755 -7449 7831 -7448
rect 5212 -7540 5279 -7524
rect 5212 -7574 5229 -7540
rect 5263 -7574 5279 -7540
rect 5212 -7590 5279 -7574
rect 6633 -7538 6700 -7522
rect 6633 -7572 6649 -7538
rect 6683 -7572 6700 -7538
rect 6633 -7588 6700 -7572
rect 5519 -7608 5553 -7592
rect 4831 -7658 4847 -7624
rect 4881 -7658 4897 -7624
rect 4949 -7657 4965 -7623
rect 4999 -7657 5015 -7623
rect 5519 -7658 5553 -7642
rect 6464 -7605 6498 -7589
rect 6464 -7655 6498 -7639
rect 6810 -7690 6844 -7449
rect 8005 -7395 8070 -5532
rect 9012 -6010 9214 -5990
rect 9012 -6054 9046 -6010
rect 9168 -6054 9214 -6010
rect 9012 -6064 9098 -6054
rect 9136 -6064 9214 -6054
rect 9012 -6082 9214 -6064
rect 9099 -6228 9369 -6193
rect 8745 -6281 8779 -6265
rect 8261 -6427 8531 -6392
rect 8261 -6481 8295 -6427
rect 8261 -6673 8295 -6657
rect 8379 -6481 8413 -6465
rect 8379 -6673 8413 -6657
rect 8497 -6481 8531 -6427
rect 8497 -6673 8531 -6657
rect 8615 -6481 8649 -6465
rect 8615 -6673 8649 -6657
rect 8745 -6673 8779 -6657
rect 8863 -6281 8897 -6265
rect 8863 -6673 8897 -6657
rect 8981 -6281 9015 -6265
rect 8981 -6673 9015 -6657
rect 9099 -6281 9133 -6228
rect 9099 -6673 9133 -6657
rect 9217 -6281 9251 -6265
rect 9217 -6673 9251 -6657
rect 9335 -6281 9369 -6228
rect 9335 -6673 9369 -6657
rect 9453 -6281 9487 -6265
rect 9453 -6673 9487 -6657
rect 9582 -6481 9616 -6465
rect 9582 -6673 9616 -6657
rect 9700 -6481 9734 -6465
rect 9700 -6673 9734 -6657
rect 9818 -6481 9852 -6465
rect 9818 -6673 9852 -6657
rect 9936 -6481 9970 -6465
rect 9936 -6673 9970 -6657
rect 9662 -6870 9668 -6836
rect 9722 -6870 9728 -6836
rect 8688 -6974 8722 -6958
rect 8806 -6974 8840 -6958
rect 8688 -7366 8722 -7350
rect 8805 -7350 8806 -7303
rect 8924 -6974 8958 -6958
rect 8840 -7350 8841 -7303
rect 7933 -7459 8070 -7395
rect 8805 -7408 8841 -7350
rect 9042 -6974 9076 -6958
rect 8924 -7366 8958 -7350
rect 9040 -7350 9042 -7303
rect 9040 -7408 9076 -7350
rect 9160 -6974 9194 -6958
rect 9160 -7366 9194 -7350
rect 9278 -6974 9312 -6958
rect 9396 -6974 9430 -6958
rect 9312 -7350 9314 -7304
rect 9278 -7408 9314 -7350
rect 9396 -7366 9430 -7350
rect 8805 -7448 9900 -7408
rect 8824 -7449 9900 -7448
rect 7280 -7538 7347 -7522
rect 7280 -7572 7297 -7538
rect 7331 -7572 7347 -7538
rect 7280 -7588 7347 -7572
rect 8702 -7538 8769 -7522
rect 8702 -7572 8718 -7538
rect 8752 -7572 8769 -7538
rect 8702 -7588 8769 -7572
rect 7587 -7606 7621 -7590
rect 6899 -7656 6915 -7622
rect 6949 -7656 6965 -7622
rect 7017 -7655 7033 -7621
rect 7067 -7655 7083 -7621
rect 7587 -7656 7621 -7640
rect 8533 -7605 8567 -7589
rect 8533 -7655 8567 -7639
rect 8879 -7690 8913 -7449
rect 10071 -7408 10135 -5505
rect 15647 -5539 15711 -4205
rect 15873 -4208 15930 -4205
rect 17456 -4159 17490 -4143
rect 17456 -4209 17490 -4193
rect 18789 -4200 19009 -4140
rect 19058 -4200 19062 -4140
rect 18789 -4202 19062 -4200
rect 15873 -4312 15930 -4308
rect 15873 -4372 15877 -4312
rect 15926 -4372 15930 -4312
rect 15873 -4376 15930 -4372
rect 17072 -4313 17164 -4300
rect 17072 -4368 17088 -4313
rect 17148 -4368 17164 -4313
rect 17072 -4385 17164 -4368
rect 17337 -4549 17371 -4533
rect 17337 -4599 17371 -4583
rect 16850 -4671 16884 -4655
rect 16850 -4863 16884 -4847
rect 16968 -4659 17002 -4655
rect 17042 -4659 17076 -4655
rect 16968 -4671 17076 -4659
rect 17002 -4847 17042 -4671
rect 16968 -4859 17042 -4847
rect 16968 -4863 17002 -4859
rect 17042 -5063 17076 -5047
rect 17160 -4671 17194 -4655
rect 17160 -5063 17194 -5047
rect 17278 -4671 17312 -4655
rect 17278 -5063 17312 -5047
rect 17396 -4671 17430 -4655
rect 17396 -5063 17430 -5047
rect 17514 -4659 17548 -4655
rect 17592 -4659 17626 -4655
rect 17514 -4671 17626 -4659
rect 17548 -4847 17592 -4671
rect 17548 -4859 17626 -4847
rect 17592 -4863 17626 -4859
rect 17710 -4671 17744 -4655
rect 17710 -4863 17744 -4847
rect 17514 -5063 17548 -5047
rect 17263 -5182 17279 -5148
rect 17313 -5182 17329 -5148
rect 17244 -5300 17380 -5296
rect 17244 -5314 17282 -5300
rect 17340 -5314 17380 -5300
rect 17244 -5360 17260 -5314
rect 17364 -5360 17380 -5314
rect 17244 -5382 17380 -5360
rect 12148 -5603 15711 -5539
rect 11080 -6008 11282 -5988
rect 11080 -6052 11114 -6008
rect 11236 -6052 11282 -6008
rect 11080 -6062 11166 -6052
rect 11204 -6062 11282 -6052
rect 11080 -6080 11282 -6062
rect 11167 -6226 11437 -6191
rect 10813 -6279 10847 -6263
rect 10329 -6425 10599 -6390
rect 10329 -6479 10363 -6425
rect 10329 -6671 10363 -6655
rect 10447 -6479 10481 -6463
rect 10447 -6671 10481 -6655
rect 10565 -6479 10599 -6425
rect 10565 -6671 10599 -6655
rect 10683 -6479 10717 -6463
rect 10683 -6671 10717 -6655
rect 10813 -6671 10847 -6655
rect 10931 -6279 10965 -6263
rect 10931 -6671 10965 -6655
rect 11049 -6279 11083 -6263
rect 11049 -6671 11083 -6655
rect 11167 -6279 11201 -6226
rect 11167 -6671 11201 -6655
rect 11285 -6279 11319 -6263
rect 11285 -6671 11319 -6655
rect 11403 -6279 11437 -6226
rect 11403 -6671 11437 -6655
rect 11521 -6279 11555 -6263
rect 11521 -6671 11555 -6655
rect 11650 -6479 11684 -6463
rect 11650 -6671 11684 -6655
rect 11768 -6479 11802 -6463
rect 11768 -6671 11802 -6655
rect 11886 -6479 11920 -6463
rect 11886 -6671 11920 -6655
rect 12004 -6479 12038 -6463
rect 12004 -6671 12038 -6655
rect 11730 -6868 11736 -6834
rect 11790 -6868 11796 -6834
rect 10756 -6972 10790 -6956
rect 10874 -6972 10908 -6956
rect 10756 -7364 10790 -7348
rect 10873 -7348 10874 -7301
rect 10992 -6972 11026 -6956
rect 10908 -7348 10909 -7301
rect 10002 -7449 10135 -7408
rect 10873 -7406 10909 -7348
rect 11110 -6972 11144 -6956
rect 10992 -7364 11026 -7348
rect 11108 -7348 11110 -7301
rect 11108 -7406 11144 -7348
rect 11228 -6972 11262 -6956
rect 11228 -7364 11262 -7348
rect 11346 -6972 11380 -6956
rect 11464 -6972 11498 -6956
rect 11380 -7348 11382 -7302
rect 11346 -7406 11382 -7348
rect 11464 -7364 11498 -7348
rect 10873 -7446 11968 -7406
rect 10892 -7447 11968 -7446
rect 9349 -7538 9416 -7522
rect 9349 -7572 9366 -7538
rect 9400 -7572 9416 -7538
rect 9349 -7588 9416 -7572
rect 10770 -7536 10837 -7520
rect 10770 -7570 10786 -7536
rect 10820 -7570 10837 -7536
rect 10770 -7586 10837 -7570
rect 9656 -7606 9690 -7590
rect 8968 -7656 8984 -7622
rect 9018 -7656 9034 -7622
rect 9086 -7655 9102 -7621
rect 9136 -7655 9152 -7621
rect 9656 -7656 9690 -7640
rect 10601 -7603 10635 -7587
rect 10601 -7653 10635 -7637
rect 10947 -7688 10981 -7447
rect 12148 -7406 12212 -5603
rect 18789 -5662 18853 -4202
rect 19005 -4204 19062 -4202
rect 20588 -4155 20622 -4139
rect 22149 -4140 22206 -4136
rect 20588 -4205 20622 -4189
rect 21929 -4200 22153 -4140
rect 22202 -4200 22206 -4140
rect 21929 -4204 22206 -4200
rect 23732 -4155 23766 -4139
rect 19005 -4308 19062 -4304
rect 19005 -4368 19009 -4308
rect 19058 -4368 19062 -4308
rect 19005 -4372 19062 -4368
rect 20204 -4309 20296 -4296
rect 20204 -4364 20220 -4309
rect 20280 -4364 20296 -4309
rect 20204 -4381 20296 -4364
rect 20469 -4545 20503 -4529
rect 20469 -4595 20503 -4579
rect 19982 -4667 20016 -4651
rect 19982 -4859 20016 -4843
rect 20100 -4655 20134 -4651
rect 20174 -4655 20208 -4651
rect 20100 -4667 20208 -4655
rect 20134 -4843 20174 -4667
rect 20100 -4855 20174 -4843
rect 20100 -4859 20134 -4855
rect 20174 -5059 20208 -5043
rect 20292 -4667 20326 -4651
rect 20292 -5059 20326 -5043
rect 20410 -4667 20444 -4651
rect 20410 -5059 20444 -5043
rect 20528 -4667 20562 -4651
rect 20528 -5059 20562 -5043
rect 20646 -4655 20680 -4651
rect 20724 -4655 20758 -4651
rect 20646 -4667 20758 -4655
rect 20680 -4843 20724 -4667
rect 20680 -4855 20758 -4843
rect 20724 -4859 20758 -4855
rect 20842 -4667 20876 -4651
rect 20842 -4859 20876 -4843
rect 20646 -5059 20680 -5043
rect 20395 -5178 20411 -5144
rect 20445 -5178 20461 -5144
rect 20376 -5296 20512 -5292
rect 20376 -5310 20414 -5296
rect 20472 -5310 20512 -5296
rect 20376 -5356 20392 -5310
rect 20496 -5356 20512 -5310
rect 20376 -5378 20512 -5356
rect 14226 -5726 18853 -5662
rect 13149 -6010 13351 -5990
rect 13149 -6054 13183 -6010
rect 13305 -6054 13351 -6010
rect 13149 -6064 13235 -6054
rect 13273 -6064 13351 -6054
rect 13149 -6082 13351 -6064
rect 13236 -6228 13506 -6193
rect 12882 -6281 12916 -6265
rect 12398 -6427 12668 -6392
rect 12398 -6481 12432 -6427
rect 12398 -6673 12432 -6657
rect 12516 -6481 12550 -6465
rect 12516 -6673 12550 -6657
rect 12634 -6481 12668 -6427
rect 12634 -6673 12668 -6657
rect 12752 -6481 12786 -6465
rect 12752 -6673 12786 -6657
rect 12882 -6673 12916 -6657
rect 13000 -6281 13034 -6265
rect 13000 -6673 13034 -6657
rect 13118 -6281 13152 -6265
rect 13118 -6673 13152 -6657
rect 13236 -6281 13270 -6228
rect 13236 -6673 13270 -6657
rect 13354 -6281 13388 -6265
rect 13354 -6673 13388 -6657
rect 13472 -6281 13506 -6228
rect 13472 -6673 13506 -6657
rect 13590 -6281 13624 -6265
rect 13590 -6673 13624 -6657
rect 13719 -6481 13753 -6465
rect 13719 -6673 13753 -6657
rect 13837 -6481 13871 -6465
rect 13837 -6673 13871 -6657
rect 13955 -6481 13989 -6465
rect 13955 -6673 13989 -6657
rect 14073 -6481 14107 -6465
rect 14073 -6673 14107 -6657
rect 13799 -6870 13805 -6836
rect 13859 -6870 13865 -6836
rect 12825 -6974 12859 -6958
rect 12943 -6974 12977 -6958
rect 12825 -7366 12859 -7350
rect 12942 -7350 12943 -7303
rect 13061 -6974 13095 -6958
rect 12977 -7350 12978 -7303
rect 12070 -7447 12212 -7406
rect 12942 -7408 12978 -7350
rect 13179 -6974 13213 -6958
rect 13061 -7366 13095 -7350
rect 13177 -7350 13179 -7303
rect 13177 -7408 13213 -7350
rect 13297 -6974 13331 -6958
rect 13297 -7366 13331 -7350
rect 13415 -6974 13449 -6958
rect 13533 -6974 13567 -6958
rect 13449 -7350 13451 -7304
rect 13415 -7408 13451 -7350
rect 13533 -7366 13567 -7350
rect 12942 -7448 14037 -7408
rect 12961 -7449 14037 -7448
rect 11417 -7536 11484 -7520
rect 11417 -7570 11434 -7536
rect 11468 -7570 11484 -7536
rect 11417 -7586 11484 -7570
rect 12839 -7538 12906 -7522
rect 12839 -7572 12855 -7538
rect 12889 -7572 12906 -7538
rect 12839 -7588 12906 -7572
rect 11724 -7604 11758 -7588
rect 11036 -7654 11052 -7620
rect 11086 -7654 11102 -7620
rect 11154 -7653 11170 -7619
rect 11204 -7653 11220 -7619
rect 11724 -7654 11758 -7638
rect 12670 -7605 12704 -7589
rect 12670 -7655 12704 -7639
rect 3596 -7898 3630 -7882
rect 4249 -7708 4283 -7692
rect 4249 -7900 4283 -7884
rect 4367 -7708 4401 -7692
rect 4367 -7900 4401 -7884
rect 4669 -7708 4703 -7692
rect 2954 -8098 2988 -8082
rect 3071 -8149 3106 -8082
rect 2600 -8184 3106 -8149
rect 4742 -7708 4821 -7692
rect 4742 -7738 4787 -7708
rect 4669 -8151 4704 -8084
rect 4787 -8100 4821 -8084
rect 4905 -7708 4939 -7692
rect 4905 -8100 4939 -8084
rect 5023 -7708 5057 -7692
rect 5141 -7708 5175 -7692
rect 5547 -7708 5581 -7692
rect 5547 -7900 5581 -7884
rect 5665 -7708 5699 -7692
rect 5665 -7900 5699 -7884
rect 6317 -7706 6351 -7690
rect 6317 -7898 6351 -7882
rect 6435 -7706 6469 -7690
rect 6435 -7898 6469 -7882
rect 6737 -7706 6771 -7690
rect 5023 -8100 5057 -8084
rect 5140 -8151 5175 -8084
rect 4669 -8186 5175 -8151
rect 6810 -7706 6889 -7690
rect 6810 -7736 6855 -7706
rect 6737 -8149 6772 -8082
rect 6855 -8098 6889 -8082
rect 6973 -7706 7007 -7690
rect 6973 -8098 7007 -8082
rect 7091 -7706 7125 -7690
rect 7209 -7706 7243 -7690
rect 7615 -7706 7649 -7690
rect 7615 -7898 7649 -7882
rect 7733 -7706 7767 -7690
rect 7733 -7898 7767 -7882
rect 8386 -7706 8420 -7690
rect 8386 -7898 8420 -7882
rect 8504 -7706 8538 -7690
rect 8504 -7898 8538 -7882
rect 8806 -7706 8840 -7690
rect 7091 -8098 7125 -8082
rect 7208 -8149 7243 -8082
rect 6737 -8184 7243 -8149
rect 8879 -7706 8958 -7690
rect 8879 -7736 8924 -7706
rect 8806 -8149 8841 -8082
rect 8924 -8098 8958 -8082
rect 9042 -7706 9076 -7690
rect 9042 -8098 9076 -8082
rect 9160 -7706 9194 -7690
rect 9278 -7706 9312 -7690
rect 9684 -7706 9718 -7690
rect 9684 -7898 9718 -7882
rect 9802 -7706 9836 -7690
rect 9802 -7898 9836 -7882
rect 10454 -7704 10488 -7688
rect 10454 -7896 10488 -7880
rect 10572 -7704 10606 -7688
rect 10572 -7896 10606 -7880
rect 10874 -7704 10908 -7688
rect 9160 -8098 9194 -8082
rect 9277 -8149 9312 -8082
rect 8806 -8184 9312 -8149
rect 10947 -7704 11026 -7688
rect 10947 -7734 10992 -7704
rect 10874 -8147 10909 -8080
rect 10992 -8096 11026 -8080
rect 11110 -7704 11144 -7688
rect 11110 -8096 11144 -8080
rect 11228 -7704 11262 -7688
rect 11346 -7704 11380 -7688
rect 11752 -7704 11786 -7688
rect 11752 -7896 11786 -7880
rect 11870 -7704 11904 -7688
rect 13016 -7690 13050 -7449
rect 14226 -7408 14290 -5726
rect 21929 -5760 21993 -4204
rect 23732 -4205 23766 -4189
rect 22149 -4308 22206 -4304
rect 22149 -4368 22153 -4308
rect 22202 -4368 22206 -4308
rect 22149 -4372 22206 -4368
rect 23348 -4309 23440 -4296
rect 23348 -4364 23364 -4309
rect 23424 -4364 23440 -4309
rect 23348 -4381 23440 -4364
rect 23613 -4545 23647 -4529
rect 23613 -4595 23647 -4579
rect 23126 -4667 23160 -4651
rect 23126 -4859 23160 -4843
rect 23244 -4655 23278 -4651
rect 23318 -4655 23352 -4651
rect 23244 -4667 23352 -4655
rect 23278 -4843 23318 -4667
rect 23244 -4855 23318 -4843
rect 23244 -4859 23278 -4855
rect 23318 -5059 23352 -5043
rect 23436 -4667 23470 -4651
rect 23436 -5059 23470 -5043
rect 23554 -4667 23588 -4651
rect 23554 -5059 23588 -5043
rect 23672 -4667 23706 -4651
rect 23672 -5059 23706 -5043
rect 23790 -4655 23824 -4651
rect 23868 -4655 23902 -4651
rect 23790 -4667 23902 -4655
rect 23824 -4843 23868 -4667
rect 23824 -4855 23902 -4843
rect 23868 -4859 23902 -4855
rect 23986 -4667 24020 -4651
rect 23986 -4859 24020 -4843
rect 23790 -5059 23824 -5043
rect 23539 -5178 23555 -5144
rect 23589 -5178 23605 -5144
rect 23520 -5296 23656 -5292
rect 23520 -5310 23558 -5296
rect 23616 -5310 23656 -5296
rect 23520 -5356 23536 -5310
rect 23640 -5356 23656 -5310
rect 23520 -5378 23656 -5356
rect 16277 -5824 21993 -5760
rect 15217 -6008 15419 -5988
rect 15217 -6052 15251 -6008
rect 15373 -6052 15419 -6008
rect 15217 -6062 15303 -6052
rect 15341 -6062 15419 -6052
rect 15217 -6080 15419 -6062
rect 15304 -6226 15574 -6191
rect 14950 -6279 14984 -6263
rect 14466 -6425 14736 -6390
rect 14466 -6479 14500 -6425
rect 14466 -6671 14500 -6655
rect 14584 -6479 14618 -6463
rect 14584 -6671 14618 -6655
rect 14702 -6479 14736 -6425
rect 14702 -6671 14736 -6655
rect 14820 -6479 14854 -6463
rect 14820 -6671 14854 -6655
rect 14950 -6671 14984 -6655
rect 15068 -6279 15102 -6263
rect 15068 -6671 15102 -6655
rect 15186 -6279 15220 -6263
rect 15186 -6671 15220 -6655
rect 15304 -6279 15338 -6226
rect 15304 -6671 15338 -6655
rect 15422 -6279 15456 -6263
rect 15422 -6671 15456 -6655
rect 15540 -6279 15574 -6226
rect 15540 -6671 15574 -6655
rect 15658 -6279 15692 -6263
rect 15658 -6671 15692 -6655
rect 15787 -6479 15821 -6463
rect 15787 -6671 15821 -6655
rect 15905 -6479 15939 -6463
rect 15905 -6671 15939 -6655
rect 16023 -6479 16057 -6463
rect 16023 -6671 16057 -6655
rect 16141 -6479 16175 -6463
rect 16141 -6671 16175 -6655
rect 15867 -6868 15873 -6834
rect 15927 -6868 15933 -6834
rect 14893 -6972 14927 -6956
rect 14473 -7083 14539 -7074
rect 15011 -6972 15045 -6956
rect 14893 -7364 14927 -7348
rect 15010 -7348 15011 -7301
rect 15129 -6972 15163 -6956
rect 15045 -7348 15046 -7301
rect 14139 -7449 14290 -7408
rect 15010 -7406 15046 -7348
rect 15247 -6972 15281 -6956
rect 15129 -7364 15163 -7348
rect 15245 -7348 15247 -7301
rect 15245 -7406 15281 -7348
rect 15365 -6972 15399 -6956
rect 15365 -7364 15399 -7348
rect 15483 -6972 15517 -6956
rect 15601 -6972 15635 -6956
rect 15517 -7348 15519 -7302
rect 15483 -7406 15519 -7348
rect 15601 -7364 15635 -7348
rect 15010 -7446 16105 -7406
rect 15029 -7447 16105 -7446
rect 13486 -7538 13553 -7522
rect 13486 -7572 13503 -7538
rect 13537 -7572 13553 -7538
rect 13486 -7588 13553 -7572
rect 14907 -7536 14974 -7520
rect 14907 -7570 14923 -7536
rect 14957 -7570 14974 -7536
rect 14907 -7586 14974 -7570
rect 13793 -7606 13827 -7590
rect 13105 -7656 13121 -7622
rect 13155 -7656 13171 -7622
rect 13223 -7655 13239 -7621
rect 13273 -7655 13289 -7621
rect 13793 -7656 13827 -7640
rect 14738 -7603 14772 -7587
rect 14738 -7653 14772 -7637
rect 15084 -7688 15118 -7447
rect 16277 -7406 16341 -5824
rect 16809 -5961 17023 -5957
rect 16809 -6023 16843 -5961
rect 16983 -6023 17023 -5961
rect 16809 -6041 17023 -6023
rect 17547 -5963 17761 -5959
rect 17547 -6025 17581 -5963
rect 17721 -6025 17761 -5963
rect 17547 -6043 17761 -6025
rect 18285 -5963 18499 -5959
rect 18285 -6025 18319 -5963
rect 18459 -6025 18499 -5963
rect 18285 -6043 18499 -6025
rect 19027 -5963 19241 -5959
rect 19027 -6025 19061 -5963
rect 19201 -6025 19241 -5963
rect 19027 -6043 19241 -6025
rect 19767 -5963 19981 -5959
rect 19767 -6025 19801 -5963
rect 19941 -6025 19981 -5963
rect 19767 -6043 19981 -6025
rect 20505 -5963 20719 -5959
rect 20505 -6025 20539 -5963
rect 20679 -6025 20719 -5963
rect 20505 -6043 20719 -6025
rect 21243 -5963 21457 -5959
rect 21243 -6025 21277 -5963
rect 21417 -6025 21457 -5963
rect 21243 -6043 21457 -6025
rect 21981 -5963 22195 -5959
rect 21981 -6025 22015 -5963
rect 22155 -6025 22195 -5963
rect 21981 -6043 22195 -6025
rect 16837 -6111 17107 -6077
rect 16719 -6167 16753 -6151
rect 16719 -6359 16753 -6343
rect 16837 -6167 16871 -6111
rect 16837 -6359 16871 -6343
rect 16955 -6167 16989 -6151
rect 16955 -6359 16989 -6343
rect 17073 -6167 17107 -6111
rect 17575 -6113 17845 -6079
rect 17073 -6359 17107 -6343
rect 17457 -6163 17491 -6147
rect 17457 -6355 17491 -6339
rect 17575 -6163 17609 -6113
rect 17575 -6355 17609 -6339
rect 17693 -6163 17727 -6147
rect 17693 -6355 17727 -6339
rect 17811 -6163 17845 -6113
rect 18313 -6113 18583 -6079
rect 17811 -6355 17845 -6339
rect 18195 -6167 18229 -6151
rect 18195 -6359 18229 -6343
rect 18313 -6167 18347 -6113
rect 18313 -6359 18347 -6343
rect 18431 -6167 18465 -6151
rect 18431 -6359 18465 -6343
rect 18549 -6167 18583 -6113
rect 19055 -6113 19325 -6079
rect 18549 -6359 18583 -6343
rect 18937 -6169 18971 -6153
rect 18937 -6361 18971 -6345
rect 19055 -6169 19089 -6113
rect 19055 -6361 19089 -6345
rect 19173 -6169 19207 -6153
rect 19173 -6361 19207 -6345
rect 19291 -6169 19325 -6113
rect 19795 -6113 20065 -6079
rect 19291 -6361 19325 -6345
rect 19677 -6169 19711 -6153
rect 19677 -6361 19711 -6345
rect 19795 -6169 19829 -6113
rect 19795 -6361 19829 -6345
rect 19913 -6169 19947 -6153
rect 19913 -6361 19947 -6345
rect 20031 -6169 20065 -6113
rect 20533 -6113 20803 -6079
rect 20031 -6361 20065 -6345
rect 20415 -6169 20449 -6153
rect 20415 -6361 20449 -6345
rect 20533 -6169 20567 -6113
rect 20533 -6361 20567 -6345
rect 20651 -6169 20685 -6153
rect 20651 -6361 20685 -6345
rect 20769 -6169 20803 -6113
rect 21271 -6113 21541 -6079
rect 20769 -6361 20803 -6345
rect 21153 -6169 21187 -6153
rect 21153 -6361 21187 -6345
rect 21271 -6169 21305 -6113
rect 21271 -6361 21305 -6345
rect 21389 -6169 21423 -6153
rect 21389 -6361 21423 -6345
rect 21507 -6169 21541 -6113
rect 22009 -6113 22279 -6079
rect 21507 -6361 21541 -6345
rect 21891 -6169 21925 -6153
rect 21891 -6361 21925 -6345
rect 22009 -6169 22043 -6113
rect 22009 -6361 22043 -6345
rect 22127 -6169 22161 -6153
rect 22127 -6361 22161 -6345
rect 22245 -6169 22279 -6113
rect 22245 -6361 22279 -6345
rect 16207 -7447 16341 -7406
rect 16649 -6483 16895 -6449
rect 16929 -6483 16945 -6449
rect 15554 -7536 15621 -7520
rect 15554 -7570 15571 -7536
rect 15605 -7570 15621 -7536
rect 15554 -7586 15621 -7570
rect 15861 -7604 15895 -7588
rect 15173 -7654 15189 -7620
rect 15223 -7654 15239 -7620
rect 15291 -7653 15307 -7619
rect 15341 -7653 15357 -7619
rect 15861 -7654 15895 -7638
rect 11870 -7896 11904 -7880
rect 12523 -7706 12557 -7690
rect 12523 -7898 12557 -7882
rect 12641 -7706 12675 -7690
rect 12641 -7898 12675 -7882
rect 12943 -7706 12977 -7690
rect 11228 -8096 11262 -8080
rect 11345 -8147 11380 -8080
rect 10874 -8182 11380 -8147
rect 13016 -7706 13095 -7690
rect 13016 -7736 13061 -7706
rect 12943 -8149 12978 -8082
rect 13061 -8098 13095 -8082
rect 13179 -7706 13213 -7690
rect 13179 -8098 13213 -8082
rect 13297 -7706 13331 -7690
rect 13415 -7706 13449 -7690
rect 13821 -7706 13855 -7690
rect 13821 -7898 13855 -7882
rect 13939 -7706 13973 -7690
rect 13939 -7898 13973 -7882
rect 14591 -7704 14625 -7688
rect 14591 -7896 14625 -7880
rect 14709 -7704 14743 -7688
rect 14709 -7896 14743 -7880
rect 15011 -7704 15045 -7688
rect 13297 -8098 13331 -8082
rect 13414 -8149 13449 -8082
rect 12943 -8184 13449 -8149
rect 15084 -7704 15163 -7688
rect 15084 -7734 15129 -7704
rect 15011 -8147 15046 -8080
rect 15129 -8096 15163 -8080
rect 15247 -7704 15281 -7688
rect 15247 -8096 15281 -8080
rect 15365 -7704 15399 -7688
rect 15483 -7704 15517 -7688
rect 15889 -7704 15923 -7688
rect 15889 -7896 15923 -7880
rect 16007 -7704 16041 -7688
rect 16007 -7896 16041 -7880
rect 15365 -8096 15399 -8080
rect 15482 -8147 15517 -8080
rect 15011 -8182 15517 -8147
rect 706 -8272 762 -8256
rect 812 -8272 870 -8256
rect 706 -8328 722 -8272
rect 854 -8328 870 -8272
rect 706 -8344 870 -8328
rect 2774 -8270 2830 -8254
rect 2880 -8270 2938 -8254
rect 2774 -8326 2790 -8270
rect 2922 -8326 2938 -8270
rect 2774 -8342 2938 -8326
rect 4843 -8272 4899 -8256
rect 4949 -8272 5007 -8256
rect 4843 -8328 4859 -8272
rect 4991 -8328 5007 -8272
rect 4843 -8344 5007 -8328
rect 6911 -8270 6967 -8254
rect 7017 -8270 7075 -8254
rect 6911 -8326 6927 -8270
rect 7059 -8326 7075 -8270
rect 6911 -8342 7075 -8326
rect 8980 -8270 9036 -8254
rect 9086 -8270 9144 -8254
rect 8980 -8326 8996 -8270
rect 9128 -8326 9144 -8270
rect 8980 -8342 9144 -8326
rect 11048 -8268 11104 -8252
rect 11154 -8268 11212 -8252
rect 11048 -8324 11064 -8268
rect 11196 -8324 11212 -8268
rect 11048 -8340 11212 -8324
rect 13117 -8270 13173 -8254
rect 13223 -8270 13281 -8254
rect 13117 -8326 13133 -8270
rect 13265 -8326 13281 -8270
rect 13117 -8342 13281 -8326
rect 15185 -8268 15241 -8252
rect 15291 -8268 15349 -8252
rect 15185 -8324 15201 -8268
rect 15333 -8324 15349 -8268
rect 15185 -8340 15349 -8324
rect 16649 -8560 16713 -6483
rect 17249 -6485 17633 -6451
rect 17667 -6485 17683 -6451
rect 17969 -6485 18371 -6451
rect 18405 -6485 18421 -6451
rect 18698 -6485 19113 -6451
rect 19147 -6485 19163 -6451
rect 19521 -6485 19853 -6451
rect 19887 -6485 19903 -6451
rect 20219 -6485 20591 -6451
rect 20625 -6485 20641 -6451
rect 16837 -6553 16871 -6537
rect 16837 -6745 16871 -6729
rect 16955 -6553 16989 -6537
rect 16955 -6745 16989 -6729
rect 16757 -6841 16941 -6821
rect 16757 -6911 16777 -6841
rect 16921 -6911 16941 -6841
rect 16757 -6917 16941 -6911
rect -43 -8624 16713 -8560
rect 17249 -8658 17313 -6485
rect 17575 -6551 17609 -6535
rect 17575 -6743 17609 -6727
rect 17693 -6551 17727 -6535
rect 17693 -6743 17727 -6727
rect 17495 -6843 17679 -6823
rect 17495 -6913 17515 -6843
rect 17659 -6913 17679 -6843
rect 17495 -6919 17679 -6913
rect 2007 -8659 17313 -8658
rect 2058 -8710 17313 -8659
rect 2007 -8722 17313 -8710
rect 17969 -8767 18033 -6485
rect 18313 -6555 18347 -6539
rect 18313 -6747 18347 -6731
rect 18431 -6555 18465 -6539
rect 18431 -6747 18465 -6731
rect 18233 -6843 18417 -6823
rect 18233 -6913 18253 -6843
rect 18397 -6913 18417 -6843
rect 18233 -6919 18417 -6913
rect 4089 -8818 18033 -8767
rect 4042 -8831 18033 -8818
rect 4042 -8832 4105 -8831
rect 18698 -8865 18762 -6485
rect 19055 -6555 19089 -6539
rect 19055 -6747 19089 -6731
rect 19173 -6555 19207 -6539
rect 19173 -6747 19207 -6731
rect 18975 -6843 19159 -6823
rect 18975 -6913 18995 -6843
rect 19139 -6913 19159 -6843
rect 18975 -6919 19159 -6913
rect 6080 -8867 18762 -8865
rect 6080 -8921 6089 -8867
rect 6136 -8921 18762 -8867
rect 6080 -8929 18762 -8921
rect 19521 -8973 19585 -6485
rect 20219 -6486 20598 -6485
rect 19795 -6555 19829 -6539
rect 19795 -6747 19829 -6731
rect 19913 -6555 19947 -6539
rect 19913 -6747 19947 -6731
rect 19715 -6843 19899 -6823
rect 19715 -6913 19735 -6843
rect 19879 -6913 19899 -6843
rect 19715 -6919 19899 -6913
rect 8179 -8977 19585 -8973
rect 8229 -9028 19585 -8977
rect 8179 -9037 19585 -9028
rect 20219 -9071 20283 -6486
rect 21009 -6491 21146 -6445
rect 21313 -6485 21329 -6451
rect 21363 -6485 21379 -6451
rect 21767 -6491 21883 -6445
rect 22051 -6485 22067 -6451
rect 22101 -6485 22117 -6451
rect 20533 -6555 20567 -6539
rect 20533 -6747 20567 -6731
rect 20651 -6555 20685 -6539
rect 20651 -6747 20685 -6731
rect 20453 -6843 20637 -6823
rect 20453 -6913 20473 -6843
rect 20617 -6913 20637 -6843
rect 20453 -6919 20637 -6913
rect 10250 -9072 20283 -9071
rect 10301 -9125 20283 -9072
rect 10250 -9135 20283 -9125
rect 21010 -9212 21074 -6491
rect 21271 -6551 21305 -6535
rect 21271 -6743 21305 -6727
rect 21389 -6551 21423 -6535
rect 21389 -6743 21423 -6727
rect 21191 -6843 21375 -6823
rect 21191 -6913 21211 -6843
rect 21355 -6913 21375 -6843
rect 21191 -6919 21375 -6913
rect 21767 -8710 21831 -6491
rect 22009 -6551 22043 -6535
rect 22009 -6743 22043 -6727
rect 22127 -6551 22161 -6535
rect 22127 -6743 22161 -6727
rect 21929 -6843 22113 -6823
rect 21929 -6913 21949 -6843
rect 22093 -6913 22113 -6843
rect 21929 -6919 22113 -6913
rect 12343 -9216 21074 -9212
rect 12343 -9267 12353 -9216
rect 12397 -9267 21074 -9216
rect 12343 -9276 21074 -9267
rect 21766 -9310 21831 -8710
rect 14421 -9311 21831 -9310
rect 14474 -9365 21831 -9311
rect 14421 -9374 21831 -9365
rect 14421 -9375 14502 -9374
<< viali >>
rect 12522 4260 12602 4330
rect 12522 4258 12602 4260
rect 11874 4220 11908 4254
rect 13690 4260 13770 4330
rect 13690 4258 13770 4260
rect 13042 4220 13076 4254
rect 14858 4260 14938 4330
rect 14858 4258 14938 4260
rect 14210 4220 14244 4254
rect 16026 4260 16106 4330
rect 16026 4258 16106 4260
rect 15378 4220 15412 4254
rect 17200 4262 17280 4332
rect 17200 4260 17280 4262
rect 16552 4222 16586 4256
rect 18368 4262 18448 4332
rect 18368 4260 18448 4262
rect 17720 4222 17754 4256
rect 19536 4262 19616 4332
rect 19536 4260 19616 4262
rect 18888 4222 18922 4256
rect 20704 4262 20784 4332
rect 20704 4260 20784 4262
rect 20056 4222 20090 4256
rect 542 4061 602 4123
rect 1990 4061 2050 4123
rect 3488 4063 3548 4125
rect 4936 4063 4996 4125
rect 6456 4061 6516 4123
rect 7904 4061 7964 4123
rect 9402 4063 9462 4125
rect 10850 4063 10910 4125
rect 11874 4112 11908 4146
rect 13042 4112 13076 4146
rect 14210 4112 14244 4146
rect 15378 4112 15412 4146
rect 16552 4114 16586 4148
rect 17720 4114 17754 4148
rect 18888 4114 18922 4148
rect 20056 4114 20090 4148
rect 201 3709 235 3885
rect 319 3709 353 3885
rect 437 3709 471 3885
rect 555 3709 589 3885
rect 673 3709 707 3885
rect 791 3709 825 3885
rect 909 3709 943 3885
rect 1027 3709 1061 3885
rect 1145 3709 1179 3885
rect 1263 3709 1297 3885
rect 1649 3709 1683 3885
rect 1767 3709 1801 3885
rect 1885 3709 1919 3885
rect 2003 3709 2037 3885
rect 2121 3709 2155 3885
rect 2239 3709 2273 3885
rect 2357 3709 2391 3885
rect 2475 3709 2509 3885
rect 2593 3709 2627 3885
rect 2711 3709 2745 3885
rect 3147 3711 3181 3887
rect 3265 3711 3299 3887
rect 3383 3711 3417 3887
rect 3501 3711 3535 3887
rect 3619 3711 3653 3887
rect 3737 3711 3771 3887
rect 3855 3711 3889 3887
rect 3973 3711 4007 3887
rect 4091 3711 4125 3887
rect 4209 3711 4243 3887
rect 4595 3711 4629 3887
rect 4713 3711 4747 3887
rect 4831 3711 4865 3887
rect 4949 3711 4983 3887
rect 5067 3711 5101 3887
rect 5185 3711 5219 3887
rect 5303 3711 5337 3887
rect 5421 3711 5455 3887
rect 5539 3711 5573 3887
rect 5657 3711 5691 3887
rect 6115 3709 6149 3885
rect 6233 3709 6267 3885
rect 6351 3709 6385 3885
rect 6469 3709 6503 3885
rect 6587 3709 6621 3885
rect 6705 3709 6739 3885
rect 6823 3709 6857 3885
rect 6941 3709 6975 3885
rect 7059 3709 7093 3885
rect 7177 3709 7211 3885
rect 7563 3709 7597 3885
rect 7681 3709 7715 3885
rect 7799 3709 7833 3885
rect 7917 3709 7951 3885
rect 8035 3709 8069 3885
rect 8153 3709 8187 3885
rect 8271 3709 8305 3885
rect 8389 3709 8423 3885
rect 8507 3709 8541 3885
rect 8625 3709 8659 3885
rect 9061 3711 9095 3887
rect 9179 3711 9213 3887
rect 9297 3711 9331 3887
rect 9415 3711 9449 3887
rect 9533 3711 9567 3887
rect 9651 3711 9685 3887
rect 9769 3711 9803 3887
rect 9887 3711 9921 3887
rect 10005 3711 10039 3887
rect 10123 3711 10157 3887
rect 10509 3711 10543 3887
rect 10627 3711 10661 3887
rect 10745 3711 10779 3887
rect 10863 3711 10897 3887
rect 10981 3711 11015 3887
rect 11099 3711 11133 3887
rect 11217 3711 11251 3887
rect 11335 3711 11369 3887
rect 11453 3711 11487 3887
rect 11571 3711 11605 3887
rect 11964 3706 11998 4082
rect 12082 3706 12116 4082
rect 12200 3706 12234 4082
rect 12318 3706 12352 4082
rect 12436 3706 12470 4082
rect 12554 3706 12588 4082
rect 12672 3706 12706 4082
rect 13132 3706 13166 4082
rect 13250 3706 13284 4082
rect 13368 3706 13402 4082
rect 13486 3706 13520 4082
rect 13604 3706 13638 4082
rect 13722 3706 13756 4082
rect 13840 3706 13874 4082
rect 14300 3704 14334 4080
rect 14418 3704 14452 4080
rect 14536 3704 14570 4080
rect 14654 3704 14688 4080
rect 14772 3704 14806 4080
rect 14890 3704 14924 4080
rect 15008 3704 15042 4080
rect 15468 3706 15502 4082
rect 15586 3706 15620 4082
rect 15704 3706 15738 4082
rect 15822 3706 15856 4082
rect 15940 3706 15974 4082
rect 16058 3706 16092 4082
rect 16176 3706 16210 4082
rect 16642 3708 16676 4084
rect 16760 3708 16794 4084
rect 16878 3708 16912 4084
rect 16996 3708 17030 4084
rect 17114 3708 17148 4084
rect 17232 3708 17266 4084
rect 17350 3708 17384 4084
rect 17810 3706 17844 4082
rect 17928 3706 17962 4082
rect 18046 3706 18080 4082
rect 18164 3706 18198 4082
rect 18282 3706 18316 4082
rect 18400 3706 18434 4082
rect 18518 3706 18552 4082
rect 18978 3708 19012 4084
rect 19096 3708 19130 4084
rect 19214 3708 19248 4084
rect 19332 3708 19366 4084
rect 19450 3708 19484 4084
rect 19568 3708 19602 4084
rect 19686 3708 19720 4084
rect 20146 3706 20180 4082
rect 20264 3706 20298 4082
rect 20382 3706 20416 4082
rect 20500 3706 20534 4082
rect 20618 3706 20652 4082
rect 20736 3706 20770 4082
rect 20854 3706 20888 4082
rect 968 3615 1002 3649
rect 2416 3615 2450 3649
rect 3914 3617 3948 3651
rect 5362 3617 5396 3651
rect 6882 3615 6916 3649
rect 8330 3615 8364 3649
rect 9828 3617 9862 3651
rect 11276 3617 11310 3651
rect 850 3498 884 3532
rect 2298 3498 2332 3532
rect 3796 3500 3830 3534
rect 5244 3500 5278 3534
rect 6764 3498 6798 3532
rect 8212 3498 8246 3532
rect 9710 3500 9744 3534
rect 11158 3500 11192 3534
rect 438 3072 472 3448
rect 556 3072 590 3448
rect 674 3072 708 3448
rect 791 3272 825 3448
rect 909 3272 943 3448
rect 1886 3072 1920 3448
rect 2004 3072 2038 3448
rect 2122 3072 2156 3448
rect 2239 3272 2273 3448
rect 2357 3272 2391 3448
rect 3384 3074 3418 3450
rect 3502 3074 3536 3450
rect 3620 3074 3654 3450
rect 3737 3274 3771 3450
rect 3855 3274 3889 3450
rect 4832 3074 4866 3450
rect 4950 3074 4984 3450
rect 5068 3074 5102 3450
rect 5185 3274 5219 3450
rect 5303 3274 5337 3450
rect 6352 3072 6386 3448
rect 6470 3072 6504 3448
rect 6588 3072 6622 3448
rect 6705 3272 6739 3448
rect 6823 3272 6857 3448
rect 7800 3072 7834 3448
rect 7918 3072 7952 3448
rect 8036 3072 8070 3448
rect 8153 3272 8187 3448
rect 8271 3272 8305 3448
rect 9298 3074 9332 3450
rect 9416 3074 9450 3450
rect 9534 3074 9568 3450
rect 9651 3274 9685 3450
rect 9769 3274 9803 3450
rect 10746 3074 10780 3450
rect 10864 3074 10898 3450
rect 10982 3074 11016 3450
rect 11099 3274 11133 3450
rect 11217 3274 11251 3450
rect 12169 3349 12203 3383
rect 13337 3349 13371 3383
rect 14505 3349 14539 3383
rect 11874 3120 11908 3296
rect 11992 3120 12026 3296
rect 12110 3120 12144 3296
rect 12228 3120 12262 3296
rect 12394 3116 12428 3292
rect 497 2988 531 3022
rect 615 2988 649 3022
rect 1945 2988 1979 3022
rect 2063 2988 2097 3022
rect 3443 2990 3477 3024
rect 3561 2990 3595 3024
rect 4891 2990 4925 3024
rect 5009 2990 5043 3024
rect 6411 2988 6445 3022
rect 6529 2988 6563 3022
rect 7859 2988 7893 3022
rect 7977 2988 8011 3022
rect 9357 2990 9391 3024
rect 9475 2990 9509 3024
rect 10805 2990 10839 3024
rect 10923 2990 10957 3024
rect 12512 3116 12546 3292
rect 12630 3116 12664 3292
rect 12748 3116 12782 3292
rect 13042 3122 13076 3298
rect 13160 3122 13194 3298
rect 13278 3122 13312 3298
rect 13396 3122 13430 3298
rect 13561 3122 13595 3298
rect 12058 2988 12124 2992
rect 770 2865 822 2911
rect 2218 2865 2270 2911
rect 3716 2867 3768 2913
rect 5164 2867 5216 2913
rect 6684 2865 6736 2911
rect 8132 2865 8184 2911
rect 9630 2867 9682 2913
rect 11078 2867 11130 2913
rect 12058 2922 12124 2988
rect 13679 3122 13713 3298
rect 13797 3122 13831 3298
rect 13915 3122 13949 3298
rect 14210 3122 14244 3298
rect 14328 3122 14362 3298
rect 14446 3122 14480 3298
rect 14564 3122 14598 3298
rect 14729 3122 14763 3298
rect 14847 3122 14881 3298
rect 14965 3122 14999 3298
rect 15083 3122 15117 3298
rect 13226 2988 13292 2992
rect 13226 2922 13292 2988
rect 14394 2988 14460 2992
rect 14394 2922 14460 2988
rect 1512 2324 1584 2378
rect 260 1752 294 1928
rect 378 1752 412 1928
rect 496 1752 530 1928
rect 614 1752 648 1928
rect 701 1752 735 2128
rect 819 1752 853 2128
rect 937 1752 971 2128
rect 1055 1752 1089 2128
rect 1168 1752 1202 2128
rect 1286 1752 1320 2128
rect 1404 1752 1438 2128
rect 1522 1752 1556 2128
rect 1640 1752 1674 2128
rect 1758 1752 1792 2128
rect 1876 1752 1910 2128
rect 1995 1752 2029 2128
rect 2113 1752 2147 2128
rect 2231 1752 2265 2128
rect 2349 1752 2383 2128
rect 2468 1752 2502 1928
rect 2586 1752 2620 1928
rect 2704 1752 2738 1928
rect 2822 1752 2856 1928
rect 2656 1544 2690 1578
rect 1346 1503 1380 1537
rect 365 1382 423 1437
rect 423 1382 425 1437
rect 1450 1383 1452 1438
rect 1452 1383 1510 1438
rect 121 1262 170 1322
rect 1700 1273 1734 1307
rect 121 1094 170 1154
rect 1332 1098 1334 1153
rect 1334 1098 1392 1153
rect 4656 2324 4728 2378
rect 3404 1752 3438 1928
rect 3522 1752 3556 1928
rect 3640 1752 3674 1928
rect 3758 1752 3792 1928
rect 3845 1752 3879 2128
rect 3963 1752 3997 2128
rect 4081 1752 4115 2128
rect 4199 1752 4233 2128
rect 4312 1752 4346 2128
rect 4430 1752 4464 2128
rect 4548 1752 4582 2128
rect 4666 1752 4700 2128
rect 4784 1752 4818 2128
rect 4902 1752 4936 2128
rect 5020 1752 5054 2128
rect 5139 1752 5173 2128
rect 5257 1752 5291 2128
rect 5375 1752 5409 2128
rect 5493 1752 5527 2128
rect 5612 1752 5646 1928
rect 5730 1752 5764 1928
rect 5848 1752 5882 1928
rect 5966 1752 6000 1928
rect 5800 1544 5834 1578
rect 4490 1503 4524 1537
rect 3509 1382 3567 1437
rect 3567 1382 3569 1437
rect 4594 1383 4596 1438
rect 4596 1383 4654 1438
rect 3265 1262 3314 1322
rect 4844 1273 4878 1307
rect 3265 1094 3314 1154
rect 4476 1098 4478 1153
rect 4478 1098 4536 1153
rect 15673 3349 15707 3383
rect 16847 3351 16881 3385
rect 18015 3351 18049 3385
rect 19183 3351 19217 3385
rect 20351 3351 20385 3385
rect 15378 3122 15412 3298
rect 15496 3122 15530 3298
rect 15614 3122 15648 3298
rect 15732 3122 15766 3298
rect 15898 3122 15932 3298
rect 16016 3122 16050 3298
rect 16134 3122 16168 3298
rect 16252 3122 16286 3298
rect 16552 3122 16586 3298
rect 16670 3122 16704 3298
rect 16788 3122 16822 3298
rect 16906 3122 16940 3298
rect 17070 3118 17104 3294
rect 17188 3118 17222 3294
rect 17306 3118 17340 3294
rect 17424 3118 17458 3294
rect 17720 3122 17754 3298
rect 17838 3122 17872 3298
rect 17956 3122 17990 3298
rect 18074 3122 18108 3298
rect 18239 3117 18273 3293
rect 15562 2988 15628 2992
rect 15562 2922 15628 2988
rect 16736 2990 16802 2994
rect 16736 2924 16802 2990
rect 18357 3117 18391 3293
rect 18475 3117 18509 3293
rect 18593 3117 18627 3293
rect 18888 3124 18922 3300
rect 19006 3124 19040 3300
rect 19124 3124 19158 3300
rect 19242 3124 19276 3300
rect 19407 3117 19441 3293
rect 19525 3117 19559 3293
rect 19643 3117 19677 3293
rect 19761 3117 19795 3293
rect 20056 3124 20090 3300
rect 20174 3124 20208 3300
rect 20292 3124 20326 3300
rect 20410 3124 20444 3300
rect 20575 3118 20609 3294
rect 17904 2990 17970 2994
rect 17904 2924 17970 2990
rect 7788 2328 7860 2382
rect 10932 2328 11004 2382
rect 6536 1756 6570 1932
rect 6654 1756 6688 1932
rect 6772 1756 6806 1932
rect 6890 1756 6924 1932
rect 6977 1756 7011 2132
rect 7095 1756 7129 2132
rect 7213 1756 7247 2132
rect 7331 1756 7365 2132
rect 7444 1756 7478 2132
rect 7562 1756 7596 2132
rect 7680 1756 7714 2132
rect 7798 1756 7832 2132
rect 7916 1756 7950 2132
rect 8034 1756 8068 2132
rect 8152 1756 8186 2132
rect 8271 1756 8305 2132
rect 8389 1756 8423 2132
rect 8507 1756 8541 2132
rect 8625 1756 8659 2132
rect 8744 1756 8778 1932
rect 8862 1756 8896 1932
rect 8980 1756 9014 1932
rect 9098 1756 9132 1932
rect 9680 1756 9714 1932
rect 9798 1756 9832 1932
rect 9916 1756 9950 1932
rect 10034 1756 10068 1932
rect 10121 1756 10155 2132
rect 10239 1756 10273 2132
rect 10357 1756 10391 2132
rect 10475 1756 10509 2132
rect 10588 1756 10622 2132
rect 10706 1756 10740 2132
rect 10824 1756 10858 2132
rect 10942 1756 10976 2132
rect 11060 1756 11094 2132
rect 11178 1756 11212 2132
rect 11296 1756 11330 2132
rect 11415 1756 11449 2132
rect 11533 1756 11567 2132
rect 11651 1756 11685 2132
rect 11769 1756 11803 2132
rect 11888 1756 11922 1932
rect 12006 1756 12040 1932
rect 12124 1756 12158 1932
rect 12242 1756 12276 1932
rect 8932 1548 8966 1582
rect 7622 1507 7656 1541
rect 12076 1548 12110 1582
rect 10766 1507 10800 1541
rect 6641 1386 6699 1441
rect 6699 1386 6701 1441
rect 7726 1387 7728 1442
rect 7728 1387 7786 1442
rect 9785 1386 9843 1441
rect 9843 1386 9845 1441
rect 10870 1387 10872 1442
rect 10872 1387 10930 1442
rect 6397 1266 6446 1326
rect 7976 1277 8010 1311
rect 9541 1266 9590 1326
rect 11120 1277 11154 1311
rect 6397 1098 6446 1158
rect 7608 1102 7610 1157
rect 7610 1102 7668 1157
rect 14134 2324 14206 2378
rect 12882 1752 12916 1928
rect 13000 1752 13034 1928
rect 13118 1752 13152 1928
rect 13236 1752 13270 1928
rect 13323 1752 13357 2128
rect 13441 1752 13475 2128
rect 13559 1752 13593 2128
rect 13677 1752 13711 2128
rect 13790 1752 13824 2128
rect 13908 1752 13942 2128
rect 14026 1752 14060 2128
rect 14144 1752 14178 2128
rect 14262 1752 14296 2128
rect 14380 1752 14414 2128
rect 14498 1752 14532 2128
rect 14617 1752 14651 2128
rect 14735 1752 14769 2128
rect 14853 1752 14887 2128
rect 14971 1752 15005 2128
rect 15090 1752 15124 1928
rect 15208 1752 15242 1928
rect 15326 1752 15360 1928
rect 15444 1752 15478 1928
rect 15278 1544 15312 1578
rect 13968 1503 14002 1537
rect 12987 1382 13045 1437
rect 13045 1382 13047 1437
rect 14072 1383 14074 1438
rect 14074 1383 14132 1438
rect 12743 1262 12792 1322
rect 14322 1273 14356 1307
rect 20693 3118 20727 3294
rect 20811 3118 20845 3294
rect 20929 3118 20963 3294
rect 19072 2990 19138 2994
rect 19072 2924 19138 2990
rect 20240 2990 20306 2994
rect 20240 2924 20306 2990
rect 17278 2324 17350 2378
rect 16026 1752 16060 1928
rect 16144 1752 16178 1928
rect 16262 1752 16296 1928
rect 16380 1752 16414 1928
rect 16467 1752 16501 2128
rect 16585 1752 16619 2128
rect 16703 1752 16737 2128
rect 16821 1752 16855 2128
rect 16934 1752 16968 2128
rect 17052 1752 17086 2128
rect 17170 1752 17204 2128
rect 17288 1752 17322 2128
rect 17406 1752 17440 2128
rect 17524 1752 17558 2128
rect 17642 1752 17676 2128
rect 17761 1752 17795 2128
rect 17879 1752 17913 2128
rect 17997 1752 18031 2128
rect 18115 1752 18149 2128
rect 18234 1752 18268 1928
rect 18352 1752 18386 1928
rect 18470 1752 18504 1928
rect 18588 1752 18622 1928
rect 18422 1544 18456 1578
rect 17112 1503 17146 1537
rect 20410 2328 20482 2382
rect 19158 1756 19192 1932
rect 19276 1756 19310 1932
rect 19394 1756 19428 1932
rect 19512 1756 19546 1932
rect 19599 1756 19633 2132
rect 19717 1756 19751 2132
rect 19835 1756 19869 2132
rect 19953 1756 19987 2132
rect 20066 1756 20100 2132
rect 20184 1756 20218 2132
rect 20302 1756 20336 2132
rect 20420 1756 20454 2132
rect 20538 1756 20572 2132
rect 20656 1756 20690 2132
rect 20774 1756 20808 2132
rect 20893 1756 20927 2132
rect 21011 1756 21045 2132
rect 21129 1756 21163 2132
rect 21247 1756 21281 2132
rect 21366 1756 21400 1932
rect 21484 1756 21518 1932
rect 21602 1756 21636 1932
rect 21720 1756 21754 1932
rect 21554 1548 21588 1582
rect 16131 1382 16189 1437
rect 16189 1382 16191 1437
rect 17216 1383 17218 1438
rect 17218 1383 17276 1438
rect 15887 1262 15936 1322
rect 17466 1273 17500 1307
rect 15887 1094 15936 1154
rect 17098 1098 17100 1153
rect 17100 1098 17158 1153
rect 20244 1507 20278 1541
rect 19263 1386 19321 1441
rect 19321 1386 19323 1441
rect 20348 1387 20350 1442
rect 20350 1387 20408 1442
rect 19019 1266 19068 1326
rect 20598 1277 20632 1311
rect 19019 1098 19068 1158
rect 20230 1102 20232 1157
rect 20232 1102 20290 1157
rect 23554 2328 23626 2382
rect 22302 1756 22336 1932
rect 22420 1756 22454 1932
rect 22538 1756 22572 1932
rect 22656 1756 22690 1932
rect 22743 1756 22777 2132
rect 22861 1756 22895 2132
rect 22979 1756 23013 2132
rect 23097 1756 23131 2132
rect 23210 1756 23244 2132
rect 23328 1756 23362 2132
rect 23446 1756 23480 2132
rect 23564 1756 23598 2132
rect 23682 1756 23716 2132
rect 23800 1756 23834 2132
rect 23918 1756 23952 2132
rect 24037 1756 24071 2132
rect 24155 1756 24189 2132
rect 24273 1756 24307 2132
rect 24391 1756 24425 2132
rect 24510 1756 24544 1932
rect 24628 1756 24662 1932
rect 24746 1756 24780 1932
rect 24864 1756 24898 1932
rect 24698 1548 24732 1582
rect 23388 1507 23422 1541
rect 22407 1386 22465 1441
rect 22465 1386 22467 1441
rect 23492 1387 23494 1442
rect 23494 1387 23552 1442
rect 22163 1266 22212 1326
rect 23742 1277 23776 1311
rect 22163 1098 22212 1158
rect 23374 1102 23376 1157
rect 23376 1102 23434 1157
rect 1581 883 1615 917
rect 4725 883 4759 917
rect 7857 887 7891 921
rect 11001 887 11035 921
rect 14203 883 14237 917
rect 17347 883 17381 917
rect 20479 887 20513 921
rect 23623 887 23657 921
rect 1094 619 1128 795
rect 1212 619 1246 795
rect 1286 419 1320 795
rect 1404 419 1438 795
rect 1522 419 1556 795
rect 1640 419 1674 795
rect 1758 419 1792 795
rect 1836 619 1870 795
rect 1954 619 1988 795
rect 4238 619 4272 795
rect 4356 619 4390 795
rect 4430 419 4464 795
rect 4548 419 4582 795
rect 4666 419 4700 795
rect 4784 419 4818 795
rect 4902 419 4936 795
rect 4980 619 5014 795
rect 5098 619 5132 795
rect 7370 623 7404 799
rect 7488 623 7522 799
rect 7562 423 7596 799
rect 7680 423 7714 799
rect 7798 423 7832 799
rect 7916 423 7950 799
rect 8034 423 8068 799
rect 8112 623 8146 799
rect 8230 623 8264 799
rect 10514 623 10548 799
rect 10632 623 10666 799
rect 10706 423 10740 799
rect 10824 423 10858 799
rect 10942 423 10976 799
rect 11060 423 11094 799
rect 11178 423 11212 799
rect 11256 623 11290 799
rect 11374 623 11408 799
rect 13716 619 13750 795
rect 13834 619 13868 795
rect 13908 419 13942 795
rect 14026 419 14060 795
rect 14144 419 14178 795
rect 14262 419 14296 795
rect 14380 419 14414 795
rect 14458 619 14492 795
rect 14576 619 14610 795
rect 16860 619 16894 795
rect 16978 619 17012 795
rect 17052 419 17086 795
rect 17170 419 17204 795
rect 17288 419 17322 795
rect 17406 419 17440 795
rect 17524 419 17558 795
rect 17602 619 17636 795
rect 17720 619 17754 795
rect 19992 623 20026 799
rect 20110 623 20144 799
rect 20184 423 20218 799
rect 20302 423 20336 799
rect 20420 423 20454 799
rect 20538 423 20572 799
rect 20656 423 20690 799
rect 20734 623 20768 799
rect 20852 623 20886 799
rect 23136 623 23170 799
rect 23254 623 23288 799
rect 23328 423 23362 799
rect 23446 423 23480 799
rect 23564 423 23598 799
rect 23682 423 23716 799
rect 23800 423 23834 799
rect 23878 623 23912 799
rect 23996 623 24030 799
rect 1523 284 1557 318
rect 4667 284 4701 318
rect 7799 288 7833 322
rect 10943 288 10977 322
rect 14145 284 14179 318
rect 17289 284 17323 318
rect 20421 288 20455 322
rect 23565 288 23599 322
rect 1526 152 1584 166
rect 1526 120 1584 152
rect 4670 152 4728 166
rect 4670 120 4728 152
rect 7802 156 7860 170
rect 7802 124 7860 156
rect 10946 156 11004 170
rect 10946 124 11004 156
rect 14148 152 14206 166
rect 14148 120 14206 152
rect 17292 152 17350 166
rect 17292 120 17350 152
rect 20424 156 20482 170
rect 20424 124 20482 156
rect 23568 156 23626 170
rect 23568 124 23626 156
rect 1512 -410 1584 -356
rect 4656 -410 4728 -356
rect 7788 -406 7860 -352
rect 10932 -406 11004 -352
rect 14134 -410 14206 -356
rect 17278 -410 17350 -356
rect 20410 -406 20482 -352
rect 23554 -406 23626 -352
rect 260 -982 294 -806
rect 378 -982 412 -806
rect 496 -982 530 -806
rect 614 -982 648 -806
rect 701 -982 735 -606
rect 819 -982 853 -606
rect 937 -982 971 -606
rect 1055 -982 1089 -606
rect 1168 -982 1202 -606
rect 1286 -982 1320 -606
rect 1404 -982 1438 -606
rect 1522 -982 1556 -606
rect 1640 -982 1674 -606
rect 1758 -982 1792 -606
rect 1876 -982 1910 -606
rect 1995 -982 2029 -606
rect 2113 -982 2147 -606
rect 2231 -982 2265 -606
rect 2349 -982 2383 -606
rect 2468 -982 2502 -806
rect 2586 -982 2620 -806
rect 2704 -982 2738 -806
rect 2822 -982 2856 -806
rect 3404 -982 3438 -806
rect 3522 -982 3556 -806
rect 3640 -982 3674 -806
rect 3758 -982 3792 -806
rect 3845 -982 3879 -606
rect 3963 -982 3997 -606
rect 4081 -982 4115 -606
rect 4199 -982 4233 -606
rect 4312 -982 4346 -606
rect 4430 -982 4464 -606
rect 4548 -982 4582 -606
rect 4666 -982 4700 -606
rect 4784 -982 4818 -606
rect 4902 -982 4936 -606
rect 5020 -982 5054 -606
rect 5139 -982 5173 -606
rect 5257 -982 5291 -606
rect 5375 -982 5409 -606
rect 5493 -982 5527 -606
rect 5612 -982 5646 -806
rect 5730 -982 5764 -806
rect 5848 -982 5882 -806
rect 5966 -982 6000 -806
rect 6536 -978 6570 -802
rect 6654 -978 6688 -802
rect 6772 -978 6806 -802
rect 6890 -978 6924 -802
rect 6977 -978 7011 -602
rect 7095 -978 7129 -602
rect 7213 -978 7247 -602
rect 7331 -978 7365 -602
rect 7444 -978 7478 -602
rect 7562 -978 7596 -602
rect 7680 -978 7714 -602
rect 7798 -978 7832 -602
rect 7916 -978 7950 -602
rect 8034 -978 8068 -602
rect 8152 -978 8186 -602
rect 8271 -978 8305 -602
rect 8389 -978 8423 -602
rect 8507 -978 8541 -602
rect 8625 -978 8659 -602
rect 8744 -978 8778 -802
rect 8862 -978 8896 -802
rect 8980 -978 9014 -802
rect 9098 -978 9132 -802
rect 9680 -978 9714 -802
rect 9798 -978 9832 -802
rect 9916 -978 9950 -802
rect 10034 -978 10068 -802
rect 10121 -978 10155 -602
rect 10239 -978 10273 -602
rect 10357 -978 10391 -602
rect 10475 -978 10509 -602
rect 10588 -978 10622 -602
rect 10706 -978 10740 -602
rect 10824 -978 10858 -602
rect 10942 -978 10976 -602
rect 11060 -978 11094 -602
rect 11178 -978 11212 -602
rect 11296 -978 11330 -602
rect 11415 -978 11449 -602
rect 11533 -978 11567 -602
rect 11651 -978 11685 -602
rect 11769 -978 11803 -602
rect 11888 -978 11922 -802
rect 12006 -978 12040 -802
rect 12124 -978 12158 -802
rect 12242 -978 12276 -802
rect 12882 -982 12916 -806
rect 13000 -982 13034 -806
rect 13118 -982 13152 -806
rect 13236 -982 13270 -806
rect 13323 -982 13357 -606
rect 13441 -982 13475 -606
rect 13559 -982 13593 -606
rect 13677 -982 13711 -606
rect 13790 -982 13824 -606
rect 13908 -982 13942 -606
rect 14026 -982 14060 -606
rect 14144 -982 14178 -606
rect 14262 -982 14296 -606
rect 14380 -982 14414 -606
rect 14498 -982 14532 -606
rect 14617 -982 14651 -606
rect 14735 -982 14769 -606
rect 14853 -982 14887 -606
rect 14971 -982 15005 -606
rect 15090 -982 15124 -806
rect 15208 -982 15242 -806
rect 15326 -982 15360 -806
rect 15444 -982 15478 -806
rect 16026 -982 16060 -806
rect 16144 -982 16178 -806
rect 16262 -982 16296 -806
rect 16380 -982 16414 -806
rect 16467 -982 16501 -606
rect 16585 -982 16619 -606
rect 16703 -982 16737 -606
rect 16821 -982 16855 -606
rect 16934 -982 16968 -606
rect 17052 -982 17086 -606
rect 17170 -982 17204 -606
rect 17288 -982 17322 -606
rect 17406 -982 17440 -606
rect 17524 -982 17558 -606
rect 17642 -982 17676 -606
rect 17761 -982 17795 -606
rect 17879 -982 17913 -606
rect 17997 -982 18031 -606
rect 18115 -982 18149 -606
rect 18234 -982 18268 -806
rect 18352 -982 18386 -806
rect 18470 -982 18504 -806
rect 18588 -982 18622 -806
rect 19158 -978 19192 -802
rect 19276 -978 19310 -802
rect 19394 -978 19428 -802
rect 19512 -978 19546 -802
rect 19599 -978 19633 -602
rect 19717 -978 19751 -602
rect 19835 -978 19869 -602
rect 19953 -978 19987 -602
rect 20066 -978 20100 -602
rect 20184 -978 20218 -602
rect 20302 -978 20336 -602
rect 20420 -978 20454 -602
rect 20538 -978 20572 -602
rect 20656 -978 20690 -602
rect 20774 -978 20808 -602
rect 20893 -978 20927 -602
rect 21011 -978 21045 -602
rect 21129 -978 21163 -602
rect 21247 -978 21281 -602
rect 21366 -978 21400 -802
rect 21484 -978 21518 -802
rect 21602 -978 21636 -802
rect 21720 -978 21754 -802
rect 22302 -978 22336 -802
rect 22420 -978 22454 -802
rect 22538 -978 22572 -802
rect 22656 -978 22690 -802
rect 22743 -978 22777 -602
rect 22861 -978 22895 -602
rect 22979 -978 23013 -602
rect 23097 -978 23131 -602
rect 23210 -978 23244 -602
rect 23328 -978 23362 -602
rect 23446 -978 23480 -602
rect 23564 -978 23598 -602
rect 23682 -978 23716 -602
rect 23800 -978 23834 -602
rect 23918 -978 23952 -602
rect 24037 -978 24071 -602
rect 24155 -978 24189 -602
rect 24273 -978 24307 -602
rect 24391 -978 24425 -602
rect 24510 -978 24544 -802
rect 24628 -978 24662 -802
rect 24746 -978 24780 -802
rect 24864 -978 24898 -802
rect 2656 -1190 2690 -1156
rect 1346 -1231 1380 -1197
rect 5800 -1190 5834 -1156
rect 4490 -1231 4524 -1197
rect 8932 -1186 8966 -1152
rect 7622 -1227 7656 -1193
rect 12076 -1186 12110 -1152
rect 10766 -1227 10800 -1193
rect 15278 -1190 15312 -1156
rect 13968 -1231 14002 -1197
rect 18422 -1190 18456 -1156
rect 17112 -1231 17146 -1197
rect 21554 -1186 21588 -1152
rect 20244 -1227 20278 -1193
rect 24698 -1186 24732 -1152
rect 23388 -1227 23422 -1193
rect 365 -1352 423 -1297
rect 423 -1352 425 -1297
rect 1450 -1351 1452 -1296
rect 1452 -1351 1510 -1296
rect 3509 -1352 3567 -1297
rect 3567 -1352 3569 -1297
rect 4594 -1351 4596 -1296
rect 4596 -1351 4654 -1296
rect 6641 -1348 6699 -1293
rect 6699 -1348 6701 -1293
rect 7726 -1347 7728 -1292
rect 7728 -1347 7786 -1292
rect 9785 -1348 9843 -1293
rect 9843 -1348 9845 -1293
rect 10870 -1347 10872 -1292
rect 10872 -1347 10930 -1292
rect 12987 -1352 13045 -1297
rect 13045 -1352 13047 -1297
rect 14072 -1351 14074 -1296
rect 14074 -1351 14132 -1296
rect 15887 -1356 15936 -1296
rect 16131 -1352 16189 -1297
rect 16189 -1352 16191 -1297
rect 17216 -1351 17218 -1296
rect 17218 -1351 17276 -1296
rect 19263 -1348 19321 -1293
rect 19321 -1348 19323 -1293
rect 20348 -1347 20350 -1292
rect 20350 -1347 20408 -1292
rect 22407 -1348 22465 -1293
rect 22465 -1348 22467 -1293
rect 23492 -1347 23494 -1292
rect 23494 -1347 23552 -1292
rect 121 -1472 170 -1412
rect 1700 -1461 1734 -1427
rect 3265 -1472 3314 -1412
rect 4844 -1461 4878 -1427
rect 6397 -1468 6446 -1408
rect 7976 -1457 8010 -1423
rect 9541 -1468 9590 -1408
rect 11120 -1457 11154 -1423
rect 12743 -1472 12792 -1412
rect 14322 -1461 14356 -1427
rect 15887 -1472 15936 -1412
rect 17466 -1461 17500 -1427
rect 19019 -1468 19068 -1408
rect 20598 -1457 20632 -1423
rect 22163 -1468 22212 -1408
rect 23742 -1457 23776 -1423
rect 121 -1640 170 -1580
rect 1332 -1636 1334 -1581
rect 1334 -1636 1392 -1581
rect 3265 -1640 3314 -1580
rect 4476 -1636 4478 -1581
rect 4478 -1636 4536 -1581
rect 6397 -1636 6446 -1576
rect 7608 -1632 7610 -1577
rect 7610 -1632 7668 -1577
rect 9541 -1636 9590 -1576
rect 10752 -1632 10754 -1577
rect 10754 -1632 10812 -1577
rect 12743 -1640 12792 -1580
rect 13954 -1636 13956 -1581
rect 13956 -1636 14014 -1581
rect 15887 -1640 15936 -1580
rect 17098 -1636 17100 -1581
rect 17100 -1636 17158 -1581
rect 19019 -1636 19068 -1576
rect 20230 -1632 20232 -1577
rect 20232 -1632 20290 -1577
rect 22163 -1636 22212 -1576
rect 23374 -1632 23376 -1577
rect 23376 -1632 23434 -1577
rect 1581 -1851 1615 -1817
rect 4725 -1851 4759 -1817
rect 7857 -1847 7891 -1813
rect 11001 -1847 11035 -1813
rect 14203 -1851 14237 -1817
rect 17347 -1851 17381 -1817
rect 20479 -1847 20513 -1813
rect 23623 -1847 23657 -1813
rect 1094 -2115 1128 -1939
rect 1212 -2115 1246 -1939
rect 1286 -2315 1320 -1939
rect 1404 -2315 1438 -1939
rect 1522 -2315 1556 -1939
rect 1640 -2315 1674 -1939
rect 1758 -2315 1792 -1939
rect 1836 -2115 1870 -1939
rect 1954 -2115 1988 -1939
rect 4238 -2115 4272 -1939
rect 4356 -2115 4390 -1939
rect 4430 -2315 4464 -1939
rect 4548 -2315 4582 -1939
rect 4666 -2315 4700 -1939
rect 4784 -2315 4818 -1939
rect 4902 -2315 4936 -1939
rect 4980 -2115 5014 -1939
rect 5098 -2115 5132 -1939
rect 7370 -2111 7404 -1935
rect 7488 -2111 7522 -1935
rect 7562 -2311 7596 -1935
rect 7680 -2311 7714 -1935
rect 7798 -2311 7832 -1935
rect 7916 -2311 7950 -1935
rect 8034 -2311 8068 -1935
rect 8112 -2111 8146 -1935
rect 8230 -2111 8264 -1935
rect 10514 -2111 10548 -1935
rect 10632 -2111 10666 -1935
rect 10706 -2311 10740 -1935
rect 10824 -2311 10858 -1935
rect 10942 -2311 10976 -1935
rect 11060 -2311 11094 -1935
rect 11178 -2311 11212 -1935
rect 11256 -2111 11290 -1935
rect 11374 -2111 11408 -1935
rect 13716 -2115 13750 -1939
rect 13834 -2115 13868 -1939
rect 13908 -2315 13942 -1939
rect 14026 -2315 14060 -1939
rect 14144 -2315 14178 -1939
rect 14262 -2315 14296 -1939
rect 14380 -2315 14414 -1939
rect 14458 -2115 14492 -1939
rect 14576 -2115 14610 -1939
rect 16860 -2115 16894 -1939
rect 16978 -2115 17012 -1939
rect 17052 -2315 17086 -1939
rect 17170 -2315 17204 -1939
rect 17288 -2315 17322 -1939
rect 17406 -2315 17440 -1939
rect 17524 -2315 17558 -1939
rect 17602 -2115 17636 -1939
rect 17720 -2115 17754 -1939
rect 19992 -2111 20026 -1935
rect 20110 -2111 20144 -1935
rect 20184 -2311 20218 -1935
rect 20302 -2311 20336 -1935
rect 20420 -2311 20454 -1935
rect 20538 -2311 20572 -1935
rect 20656 -2311 20690 -1935
rect 20734 -2111 20768 -1935
rect 20852 -2111 20886 -1935
rect 23136 -2111 23170 -1935
rect 23254 -2111 23288 -1935
rect 23328 -2311 23362 -1935
rect 23446 -2311 23480 -1935
rect 23564 -2311 23598 -1935
rect 23682 -2311 23716 -1935
rect 23800 -2311 23834 -1935
rect 23878 -2111 23912 -1935
rect 23996 -2111 24030 -1935
rect 1523 -2450 1557 -2416
rect 4667 -2450 4701 -2416
rect 7799 -2446 7833 -2412
rect 10943 -2446 10977 -2412
rect 14145 -2450 14179 -2416
rect 17289 -2450 17323 -2416
rect 20421 -2446 20455 -2412
rect 23565 -2446 23599 -2412
rect 1526 -2582 1584 -2568
rect 1526 -2614 1584 -2582
rect 4670 -2582 4728 -2568
rect 4670 -2614 4728 -2582
rect 7802 -2578 7860 -2564
rect 7802 -2610 7860 -2578
rect 10946 -2578 11004 -2564
rect 10946 -2610 11004 -2578
rect 14148 -2582 14206 -2568
rect 14148 -2614 14206 -2582
rect 17292 -2582 17350 -2568
rect 17292 -2614 17350 -2582
rect 20424 -2578 20482 -2564
rect 20424 -2610 20482 -2578
rect 23568 -2578 23626 -2564
rect 23568 -2610 23626 -2578
rect 1502 -3142 1574 -3088
rect 4646 -3142 4718 -3088
rect 7778 -3138 7850 -3084
rect 10922 -3138 10994 -3084
rect 14124 -3142 14196 -3088
rect 17268 -3142 17340 -3088
rect 20400 -3138 20472 -3084
rect 23544 -3138 23616 -3084
rect 250 -3714 284 -3538
rect 368 -3714 402 -3538
rect 486 -3714 520 -3538
rect 604 -3714 638 -3538
rect 691 -3714 725 -3338
rect 809 -3714 843 -3338
rect 927 -3714 961 -3338
rect 1045 -3714 1079 -3338
rect 1158 -3714 1192 -3338
rect 1276 -3714 1310 -3338
rect 1394 -3714 1428 -3338
rect 1512 -3714 1546 -3338
rect 1630 -3714 1664 -3338
rect 1748 -3714 1782 -3338
rect 1866 -3714 1900 -3338
rect 1985 -3714 2019 -3338
rect 2103 -3714 2137 -3338
rect 2221 -3714 2255 -3338
rect 2339 -3714 2373 -3338
rect 2458 -3714 2492 -3538
rect 2576 -3714 2610 -3538
rect 2694 -3714 2728 -3538
rect 2812 -3714 2846 -3538
rect 3394 -3714 3428 -3538
rect 3512 -3714 3546 -3538
rect 3630 -3714 3664 -3538
rect 3748 -3714 3782 -3538
rect 3835 -3714 3869 -3338
rect 3953 -3714 3987 -3338
rect 4071 -3714 4105 -3338
rect 4189 -3714 4223 -3338
rect 4302 -3714 4336 -3338
rect 4420 -3714 4454 -3338
rect 4538 -3714 4572 -3338
rect 4656 -3714 4690 -3338
rect 4774 -3714 4808 -3338
rect 4892 -3714 4926 -3338
rect 5010 -3714 5044 -3338
rect 5129 -3714 5163 -3338
rect 5247 -3714 5281 -3338
rect 5365 -3714 5399 -3338
rect 5483 -3714 5517 -3338
rect 5602 -3714 5636 -3538
rect 5720 -3714 5754 -3538
rect 5838 -3714 5872 -3538
rect 5956 -3714 5990 -3538
rect 6526 -3710 6560 -3534
rect 6644 -3710 6678 -3534
rect 6762 -3710 6796 -3534
rect 6880 -3710 6914 -3534
rect 6967 -3710 7001 -3334
rect 7085 -3710 7119 -3334
rect 7203 -3710 7237 -3334
rect 7321 -3710 7355 -3334
rect 7434 -3710 7468 -3334
rect 7552 -3710 7586 -3334
rect 7670 -3710 7704 -3334
rect 7788 -3710 7822 -3334
rect 7906 -3710 7940 -3334
rect 8024 -3710 8058 -3334
rect 8142 -3710 8176 -3334
rect 8261 -3710 8295 -3334
rect 8379 -3710 8413 -3334
rect 8497 -3710 8531 -3334
rect 8615 -3710 8649 -3334
rect 8734 -3710 8768 -3534
rect 8852 -3710 8886 -3534
rect 8970 -3710 9004 -3534
rect 9088 -3710 9122 -3534
rect 9670 -3710 9704 -3534
rect 9788 -3710 9822 -3534
rect 9906 -3710 9940 -3534
rect 10024 -3710 10058 -3534
rect 10111 -3710 10145 -3334
rect 10229 -3710 10263 -3334
rect 10347 -3710 10381 -3334
rect 10465 -3710 10499 -3334
rect 10578 -3710 10612 -3334
rect 10696 -3710 10730 -3334
rect 10814 -3710 10848 -3334
rect 10932 -3710 10966 -3334
rect 11050 -3710 11084 -3334
rect 11168 -3710 11202 -3334
rect 11286 -3710 11320 -3334
rect 11405 -3710 11439 -3334
rect 11523 -3710 11557 -3334
rect 11641 -3710 11675 -3334
rect 11759 -3710 11793 -3334
rect 11878 -3710 11912 -3534
rect 11996 -3710 12030 -3534
rect 12114 -3710 12148 -3534
rect 12232 -3710 12266 -3534
rect 12872 -3714 12906 -3538
rect 12990 -3714 13024 -3538
rect 13108 -3714 13142 -3538
rect 13226 -3714 13260 -3538
rect 13313 -3714 13347 -3338
rect 13431 -3714 13465 -3338
rect 13549 -3714 13583 -3338
rect 13667 -3714 13701 -3338
rect 13780 -3714 13814 -3338
rect 13898 -3714 13932 -3338
rect 14016 -3714 14050 -3338
rect 14134 -3714 14168 -3338
rect 14252 -3714 14286 -3338
rect 14370 -3714 14404 -3338
rect 14488 -3714 14522 -3338
rect 14607 -3714 14641 -3338
rect 14725 -3714 14759 -3338
rect 14843 -3714 14877 -3338
rect 14961 -3714 14995 -3338
rect 15080 -3714 15114 -3538
rect 15198 -3714 15232 -3538
rect 15316 -3714 15350 -3538
rect 15434 -3714 15468 -3538
rect 16016 -3714 16050 -3538
rect 16134 -3714 16168 -3538
rect 16252 -3714 16286 -3538
rect 16370 -3714 16404 -3538
rect 16457 -3714 16491 -3338
rect 16575 -3714 16609 -3338
rect 16693 -3714 16727 -3338
rect 16811 -3714 16845 -3338
rect 16924 -3714 16958 -3338
rect 17042 -3714 17076 -3338
rect 17160 -3714 17194 -3338
rect 17278 -3714 17312 -3338
rect 17396 -3714 17430 -3338
rect 17514 -3714 17548 -3338
rect 17632 -3714 17666 -3338
rect 17751 -3714 17785 -3338
rect 17869 -3714 17903 -3338
rect 17987 -3714 18021 -3338
rect 18105 -3714 18139 -3338
rect 18224 -3714 18258 -3538
rect 18342 -3714 18376 -3538
rect 18460 -3714 18494 -3538
rect 18578 -3714 18612 -3538
rect 19148 -3710 19182 -3534
rect 19266 -3710 19300 -3534
rect 19384 -3710 19418 -3534
rect 19502 -3710 19536 -3534
rect 19589 -3710 19623 -3334
rect 19707 -3710 19741 -3334
rect 19825 -3710 19859 -3334
rect 19943 -3710 19977 -3334
rect 20056 -3710 20090 -3334
rect 20174 -3710 20208 -3334
rect 20292 -3710 20326 -3334
rect 20410 -3710 20444 -3334
rect 20528 -3710 20562 -3334
rect 20646 -3710 20680 -3334
rect 20764 -3710 20798 -3334
rect 20883 -3710 20917 -3334
rect 21001 -3710 21035 -3334
rect 21119 -3710 21153 -3334
rect 21237 -3710 21271 -3334
rect 21356 -3710 21390 -3534
rect 21474 -3710 21508 -3534
rect 21592 -3710 21626 -3534
rect 21710 -3710 21744 -3534
rect 22292 -3710 22326 -3534
rect 22410 -3710 22444 -3534
rect 22528 -3710 22562 -3534
rect 22646 -3710 22680 -3534
rect 22733 -3710 22767 -3334
rect 22851 -3710 22885 -3334
rect 22969 -3710 23003 -3334
rect 23087 -3710 23121 -3334
rect 23200 -3710 23234 -3334
rect 23318 -3710 23352 -3334
rect 23436 -3710 23470 -3334
rect 23554 -3710 23588 -3334
rect 23672 -3710 23706 -3334
rect 23790 -3710 23824 -3334
rect 23908 -3710 23942 -3334
rect 24027 -3710 24061 -3334
rect 24145 -3710 24179 -3334
rect 24263 -3710 24297 -3334
rect 24381 -3710 24415 -3334
rect 24500 -3710 24534 -3534
rect 24618 -3710 24652 -3534
rect 24736 -3710 24770 -3534
rect 24854 -3710 24888 -3534
rect 2646 -3922 2680 -3888
rect 1336 -3963 1370 -3929
rect 5790 -3922 5824 -3888
rect 4480 -3963 4514 -3929
rect 8922 -3918 8956 -3884
rect 7612 -3959 7646 -3925
rect 12066 -3918 12100 -3884
rect 10756 -3959 10790 -3925
rect 15268 -3922 15302 -3888
rect 13958 -3963 13992 -3929
rect 18412 -3922 18446 -3888
rect 17102 -3963 17136 -3929
rect 21544 -3918 21578 -3884
rect 20234 -3959 20268 -3925
rect 24688 -3918 24722 -3884
rect 23378 -3959 23412 -3925
rect 111 -4088 160 -4028
rect 355 -4084 413 -4029
rect 413 -4084 415 -4029
rect 1440 -4083 1442 -4028
rect 1442 -4083 1500 -4028
rect 3255 -4088 3304 -4028
rect 3499 -4084 3557 -4029
rect 3557 -4084 3559 -4029
rect 4584 -4083 4586 -4028
rect 4586 -4083 4644 -4028
rect 6387 -4084 6436 -4024
rect 6631 -4080 6689 -4025
rect 6689 -4080 6691 -4025
rect 7716 -4079 7718 -4024
rect 7718 -4079 7776 -4024
rect 9531 -4084 9580 -4024
rect 9775 -4080 9833 -4025
rect 9833 -4080 9835 -4025
rect 10860 -4079 10862 -4024
rect 10862 -4079 10920 -4024
rect 12733 -4088 12782 -4028
rect 12977 -4084 13035 -4029
rect 13035 -4084 13037 -4029
rect 14062 -4083 14064 -4028
rect 14064 -4083 14122 -4028
rect 15877 -4088 15926 -4028
rect 16121 -4084 16179 -4029
rect 16179 -4084 16181 -4029
rect 17206 -4083 17208 -4028
rect 17208 -4083 17266 -4028
rect 19009 -4084 19058 -4024
rect 19253 -4080 19311 -4025
rect 19311 -4080 19313 -4025
rect 20338 -4079 20340 -4024
rect 20340 -4079 20398 -4024
rect 22153 -4084 22202 -4024
rect 22397 -4080 22455 -4025
rect 22455 -4080 22457 -4025
rect 23482 -4079 23484 -4024
rect 23484 -4079 23542 -4024
rect 111 -4204 160 -4144
rect 1690 -4193 1724 -4159
rect 3255 -4204 3304 -4144
rect 111 -4372 160 -4312
rect 1322 -4368 1324 -4313
rect 1324 -4368 1382 -4313
rect 1571 -4583 1605 -4549
rect 1084 -4847 1118 -4671
rect 1202 -4847 1236 -4671
rect 1276 -5047 1310 -4671
rect 1394 -5047 1428 -4671
rect 1512 -5047 1546 -4671
rect 1630 -5047 1664 -4671
rect 1748 -5047 1782 -4671
rect 1826 -4847 1860 -4671
rect 1944 -4847 1978 -4671
rect 1513 -5182 1547 -5148
rect 1516 -5314 1574 -5300
rect 1516 -5346 1574 -5314
rect 824 -6056 862 -6028
rect 824 -6066 862 -6056
rect -13 -6659 21 -6483
rect 105 -6659 139 -6483
rect 223 -6659 257 -6483
rect 341 -6659 375 -6483
rect 471 -6659 505 -6283
rect 589 -6659 623 -6283
rect 707 -6659 741 -6283
rect 825 -6659 859 -6283
rect 943 -6659 977 -6283
rect 1061 -6659 1095 -6283
rect 1179 -6659 1213 -6283
rect 1308 -6659 1342 -6483
rect 1426 -6659 1460 -6483
rect 1544 -6659 1578 -6483
rect 1662 -6659 1696 -6483
rect 1394 -6838 1448 -6828
rect 1394 -6872 1404 -6838
rect 1404 -6872 1438 -6838
rect 1438 -6872 1448 -6838
rect 1394 -6882 1448 -6872
rect -6 -7032 60 -7018
rect -6 -7066 10 -7032
rect 10 -7066 44 -7032
rect 44 -7066 60 -7032
rect -6 -7078 60 -7066
rect 414 -7352 448 -6976
rect 532 -7352 566 -6976
rect 650 -7352 684 -6976
rect 768 -7352 802 -6976
rect 886 -7352 920 -6976
rect 1004 -7352 1038 -6976
rect 1122 -7352 1156 -6976
rect 444 -7574 478 -7540
rect 259 -7641 293 -7607
rect 1626 -7482 1728 -7380
rect 4834 -4193 4868 -4159
rect 6387 -4200 6436 -4140
rect 3255 -4372 3304 -4312
rect 4466 -4368 4468 -4313
rect 4468 -4368 4526 -4313
rect 4715 -4583 4749 -4549
rect 7966 -4189 8000 -4155
rect 9531 -4200 9580 -4140
rect 6387 -4368 6436 -4308
rect 7598 -4364 7600 -4309
rect 7600 -4364 7658 -4309
rect 7847 -4579 7881 -4545
rect 4228 -4847 4262 -4671
rect 4346 -4847 4380 -4671
rect 4420 -5047 4454 -4671
rect 4538 -5047 4572 -4671
rect 4656 -5047 4690 -4671
rect 4774 -5047 4808 -4671
rect 4892 -5047 4926 -4671
rect 4970 -4847 5004 -4671
rect 5088 -4847 5122 -4671
rect 4657 -5182 4691 -5148
rect 4660 -5314 4718 -5300
rect 4660 -5346 4718 -5314
rect 2892 -6054 2930 -6026
rect 2892 -6064 2930 -6054
rect 2055 -6657 2089 -6481
rect 2173 -6657 2207 -6481
rect 2291 -6657 2325 -6481
rect 2409 -6657 2443 -6481
rect 2539 -6657 2573 -6281
rect 2657 -6657 2691 -6281
rect 2775 -6657 2809 -6281
rect 2893 -6657 2927 -6281
rect 3011 -6657 3045 -6281
rect 3129 -6657 3163 -6281
rect 3247 -6657 3281 -6281
rect 3376 -6657 3410 -6481
rect 3494 -6657 3528 -6481
rect 3612 -6657 3646 -6481
rect 3730 -6657 3764 -6481
rect 3462 -6836 3516 -6826
rect 3462 -6870 3472 -6836
rect 3472 -6870 3506 -6836
rect 3506 -6870 3516 -6836
rect 3462 -6880 3516 -6870
rect 2062 -7030 2128 -7016
rect 2062 -7064 2078 -7030
rect 2078 -7064 2112 -7030
rect 2112 -7064 2128 -7030
rect 2062 -7076 2128 -7064
rect 2482 -7350 2516 -6974
rect 2600 -7350 2634 -6974
rect 2718 -7350 2752 -6974
rect 2836 -7350 2870 -6974
rect 2954 -7350 2988 -6974
rect 3072 -7350 3106 -6974
rect 3190 -7350 3224 -6974
rect 1092 -7574 1126 -7540
rect 2512 -7572 2546 -7538
rect 710 -7658 744 -7624
rect 828 -7657 862 -7623
rect 1382 -7642 1416 -7608
rect 2327 -7639 2361 -7605
rect 3694 -7480 3796 -7378
rect 4961 -6056 4999 -6028
rect 4961 -6066 4999 -6056
rect 4124 -6659 4158 -6483
rect 4242 -6659 4276 -6483
rect 4360 -6659 4394 -6483
rect 4478 -6659 4512 -6483
rect 4608 -6659 4642 -6283
rect 4726 -6659 4760 -6283
rect 4844 -6659 4878 -6283
rect 4962 -6659 4996 -6283
rect 5080 -6659 5114 -6283
rect 5198 -6659 5232 -6283
rect 5316 -6659 5350 -6283
rect 5445 -6659 5479 -6483
rect 5563 -6659 5597 -6483
rect 5681 -6659 5715 -6483
rect 5799 -6659 5833 -6483
rect 5531 -6838 5585 -6828
rect 5531 -6872 5541 -6838
rect 5541 -6872 5575 -6838
rect 5575 -6872 5585 -6838
rect 5531 -6882 5585 -6872
rect 4131 -7032 4197 -7018
rect 4131 -7066 4147 -7032
rect 4147 -7066 4181 -7032
rect 4181 -7066 4197 -7032
rect 4131 -7078 4197 -7066
rect 4551 -7352 4585 -6976
rect 4669 -7352 4703 -6976
rect 4787 -7352 4821 -6976
rect 4905 -7352 4939 -6976
rect 5023 -7352 5057 -6976
rect 5141 -7352 5175 -6976
rect 5259 -7352 5293 -6976
rect 3160 -7572 3194 -7538
rect 4581 -7574 4615 -7540
rect 2778 -7656 2812 -7622
rect 2896 -7655 2930 -7621
rect 3450 -7640 3484 -7606
rect 4396 -7641 4430 -7607
rect 112 -7884 146 -7708
rect 230 -7884 264 -7708
rect 532 -8084 566 -7708
rect 650 -8084 684 -7708
rect 768 -8084 802 -7708
rect 886 -8084 920 -7708
rect 1004 -8084 1038 -7708
rect 1410 -7884 1444 -7708
rect 1528 -7884 1562 -7708
rect 2180 -7882 2214 -7706
rect 2298 -7882 2332 -7706
rect 2600 -8082 2634 -7706
rect 2718 -8082 2752 -7706
rect 2836 -8082 2870 -7706
rect 2954 -8082 2988 -7706
rect 3072 -8082 3106 -7706
rect 3478 -7882 3512 -7706
rect 5763 -7482 5865 -7380
rect 7360 -4843 7394 -4667
rect 7478 -4843 7512 -4667
rect 7552 -5043 7586 -4667
rect 7670 -5043 7704 -4667
rect 7788 -5043 7822 -4667
rect 7906 -5043 7940 -4667
rect 8024 -5043 8058 -4667
rect 8102 -4843 8136 -4667
rect 8220 -4843 8254 -4667
rect 7789 -5178 7823 -5144
rect 7792 -5310 7850 -5296
rect 7792 -5342 7850 -5310
rect 11110 -4189 11144 -4155
rect 12733 -4204 12782 -4144
rect 14312 -4193 14346 -4159
rect 9531 -4368 9580 -4308
rect 10742 -4364 10744 -4309
rect 10744 -4364 10802 -4309
rect 10991 -4579 11025 -4545
rect 10504 -4843 10538 -4667
rect 10622 -4843 10656 -4667
rect 10696 -5043 10730 -4667
rect 10814 -5043 10848 -4667
rect 10932 -5043 10966 -4667
rect 11050 -5043 11084 -4667
rect 11168 -5043 11202 -4667
rect 11246 -4843 11280 -4667
rect 11364 -4843 11398 -4667
rect 10933 -5178 10967 -5144
rect 10936 -5310 10994 -5296
rect 10936 -5342 10994 -5310
rect 15877 -4204 15926 -4144
rect 12733 -4372 12782 -4312
rect 13944 -4368 13946 -4313
rect 13946 -4368 14004 -4313
rect 14193 -4583 14227 -4549
rect 13706 -4847 13740 -4671
rect 13824 -4847 13858 -4671
rect 13898 -5047 13932 -4671
rect 14016 -5047 14050 -4671
rect 14134 -5047 14168 -4671
rect 14252 -5047 14286 -4671
rect 14370 -5047 14404 -4671
rect 14448 -4847 14482 -4671
rect 14566 -4847 14600 -4671
rect 14135 -5182 14169 -5148
rect 14138 -5314 14196 -5300
rect 14138 -5346 14196 -5314
rect 7029 -6054 7067 -6026
rect 7029 -6064 7067 -6054
rect 6192 -6657 6226 -6481
rect 6310 -6657 6344 -6481
rect 6428 -6657 6462 -6481
rect 6546 -6657 6580 -6481
rect 6676 -6657 6710 -6281
rect 6794 -6657 6828 -6281
rect 6912 -6657 6946 -6281
rect 7030 -6657 7064 -6281
rect 7148 -6657 7182 -6281
rect 7266 -6657 7300 -6281
rect 7384 -6657 7418 -6281
rect 7513 -6657 7547 -6481
rect 7631 -6657 7665 -6481
rect 7749 -6657 7783 -6481
rect 7867 -6657 7901 -6481
rect 7599 -6836 7653 -6826
rect 7599 -6870 7609 -6836
rect 7609 -6870 7643 -6836
rect 7643 -6870 7653 -6836
rect 7599 -6880 7653 -6870
rect 6199 -7030 6265 -7016
rect 6199 -7064 6215 -7030
rect 6215 -7064 6249 -7030
rect 6249 -7064 6265 -7030
rect 6199 -7076 6265 -7064
rect 6619 -7350 6653 -6974
rect 6737 -7350 6771 -6974
rect 6855 -7350 6889 -6974
rect 6973 -7350 7007 -6974
rect 7091 -7350 7125 -6974
rect 7209 -7350 7243 -6974
rect 7327 -7350 7361 -6974
rect 5229 -7574 5263 -7540
rect 6649 -7572 6683 -7538
rect 4847 -7658 4881 -7624
rect 4965 -7657 4999 -7623
rect 5519 -7642 5553 -7608
rect 6464 -7639 6498 -7605
rect 7831 -7480 7933 -7378
rect 9098 -6054 9136 -6026
rect 9098 -6064 9136 -6054
rect 8261 -6657 8295 -6481
rect 8379 -6657 8413 -6481
rect 8497 -6657 8531 -6481
rect 8615 -6657 8649 -6481
rect 8745 -6657 8779 -6281
rect 8863 -6657 8897 -6281
rect 8981 -6657 9015 -6281
rect 9099 -6657 9133 -6281
rect 9217 -6657 9251 -6281
rect 9335 -6657 9369 -6281
rect 9453 -6657 9487 -6281
rect 9582 -6657 9616 -6481
rect 9700 -6657 9734 -6481
rect 9818 -6657 9852 -6481
rect 9936 -6657 9970 -6481
rect 9668 -6836 9722 -6826
rect 9668 -6870 9678 -6836
rect 9678 -6870 9712 -6836
rect 9712 -6870 9722 -6836
rect 9668 -6880 9722 -6870
rect 8268 -7030 8334 -7016
rect 8268 -7064 8284 -7030
rect 8284 -7064 8318 -7030
rect 8318 -7064 8334 -7030
rect 8268 -7076 8334 -7064
rect 8688 -7350 8722 -6974
rect 8806 -7350 8840 -6974
rect 8924 -7350 8958 -6974
rect 9042 -7350 9076 -6974
rect 9160 -7350 9194 -6974
rect 9278 -7350 9312 -6974
rect 9396 -7350 9430 -6974
rect 7297 -7572 7331 -7538
rect 8718 -7572 8752 -7538
rect 6915 -7656 6949 -7622
rect 7033 -7655 7067 -7621
rect 7587 -7640 7621 -7606
rect 8533 -7639 8567 -7605
rect 9900 -7480 10002 -7378
rect 17456 -4193 17490 -4159
rect 19009 -4200 19058 -4140
rect 15877 -4372 15926 -4312
rect 17088 -4368 17090 -4313
rect 17090 -4368 17148 -4313
rect 17337 -4583 17371 -4549
rect 16850 -4847 16884 -4671
rect 16968 -4847 17002 -4671
rect 17042 -5047 17076 -4671
rect 17160 -5047 17194 -4671
rect 17278 -5047 17312 -4671
rect 17396 -5047 17430 -4671
rect 17514 -5047 17548 -4671
rect 17592 -4847 17626 -4671
rect 17710 -4847 17744 -4671
rect 17279 -5182 17313 -5148
rect 17282 -5314 17340 -5300
rect 17282 -5346 17340 -5314
rect 11166 -6052 11204 -6024
rect 11166 -6062 11204 -6052
rect 10329 -6655 10363 -6479
rect 10447 -6655 10481 -6479
rect 10565 -6655 10599 -6479
rect 10683 -6655 10717 -6479
rect 10813 -6655 10847 -6279
rect 10931 -6655 10965 -6279
rect 11049 -6655 11083 -6279
rect 11167 -6655 11201 -6279
rect 11285 -6655 11319 -6279
rect 11403 -6655 11437 -6279
rect 11521 -6655 11555 -6279
rect 11650 -6655 11684 -6479
rect 11768 -6655 11802 -6479
rect 11886 -6655 11920 -6479
rect 12004 -6655 12038 -6479
rect 11736 -6834 11790 -6824
rect 11736 -6868 11746 -6834
rect 11746 -6868 11780 -6834
rect 11780 -6868 11790 -6834
rect 11736 -6878 11790 -6868
rect 10336 -7028 10402 -7014
rect 10336 -7062 10352 -7028
rect 10352 -7062 10386 -7028
rect 10386 -7062 10402 -7028
rect 10336 -7074 10402 -7062
rect 10756 -7348 10790 -6972
rect 10874 -7348 10908 -6972
rect 10992 -7348 11026 -6972
rect 11110 -7348 11144 -6972
rect 11228 -7348 11262 -6972
rect 11346 -7348 11380 -6972
rect 11464 -7348 11498 -6972
rect 9366 -7572 9400 -7538
rect 10786 -7570 10820 -7536
rect 8984 -7656 9018 -7622
rect 9102 -7655 9136 -7621
rect 9656 -7640 9690 -7606
rect 10601 -7637 10635 -7603
rect 11968 -7478 12070 -7376
rect 20588 -4189 20622 -4155
rect 22153 -4200 22202 -4140
rect 23732 -4189 23766 -4155
rect 19009 -4368 19058 -4308
rect 20220 -4364 20222 -4309
rect 20222 -4364 20280 -4309
rect 20469 -4579 20503 -4545
rect 19982 -4843 20016 -4667
rect 20100 -4843 20134 -4667
rect 20174 -5043 20208 -4667
rect 20292 -5043 20326 -4667
rect 20410 -5043 20444 -4667
rect 20528 -5043 20562 -4667
rect 20646 -5043 20680 -4667
rect 20724 -4843 20758 -4667
rect 20842 -4843 20876 -4667
rect 20411 -5178 20445 -5144
rect 20414 -5310 20472 -5296
rect 20414 -5342 20472 -5310
rect 13235 -6054 13273 -6026
rect 13235 -6064 13273 -6054
rect 12398 -6657 12432 -6481
rect 12516 -6657 12550 -6481
rect 12634 -6657 12668 -6481
rect 12752 -6657 12786 -6481
rect 12882 -6657 12916 -6281
rect 13000 -6657 13034 -6281
rect 13118 -6657 13152 -6281
rect 13236 -6657 13270 -6281
rect 13354 -6657 13388 -6281
rect 13472 -6657 13506 -6281
rect 13590 -6657 13624 -6281
rect 13719 -6657 13753 -6481
rect 13837 -6657 13871 -6481
rect 13955 -6657 13989 -6481
rect 14073 -6657 14107 -6481
rect 13805 -6836 13859 -6826
rect 13805 -6870 13815 -6836
rect 13815 -6870 13849 -6836
rect 13849 -6870 13859 -6836
rect 13805 -6880 13859 -6870
rect 12405 -7030 12471 -7016
rect 12405 -7064 12421 -7030
rect 12421 -7064 12455 -7030
rect 12455 -7064 12471 -7030
rect 12405 -7076 12471 -7064
rect 12825 -7350 12859 -6974
rect 12943 -7350 12977 -6974
rect 13061 -7350 13095 -6974
rect 13179 -7350 13213 -6974
rect 13297 -7350 13331 -6974
rect 13415 -7350 13449 -6974
rect 13533 -7350 13567 -6974
rect 11434 -7570 11468 -7536
rect 12855 -7572 12889 -7538
rect 11052 -7654 11086 -7620
rect 11170 -7653 11204 -7619
rect 11724 -7638 11758 -7604
rect 12670 -7639 12704 -7605
rect 3596 -7882 3630 -7706
rect 4249 -7884 4283 -7708
rect 4367 -7884 4401 -7708
rect 4669 -8084 4703 -7708
rect 4787 -8084 4821 -7708
rect 4905 -8084 4939 -7708
rect 5023 -8084 5057 -7708
rect 5141 -8084 5175 -7708
rect 5547 -7884 5581 -7708
rect 5665 -7884 5699 -7708
rect 6317 -7882 6351 -7706
rect 6435 -7882 6469 -7706
rect 6737 -8082 6771 -7706
rect 6855 -8082 6889 -7706
rect 6973 -8082 7007 -7706
rect 7091 -8082 7125 -7706
rect 7209 -8082 7243 -7706
rect 7615 -7882 7649 -7706
rect 7733 -7882 7767 -7706
rect 8386 -7882 8420 -7706
rect 8504 -7882 8538 -7706
rect 8806 -8082 8840 -7706
rect 8924 -8082 8958 -7706
rect 9042 -8082 9076 -7706
rect 9160 -8082 9194 -7706
rect 9278 -8082 9312 -7706
rect 9684 -7882 9718 -7706
rect 9802 -7882 9836 -7706
rect 10454 -7880 10488 -7704
rect 10572 -7880 10606 -7704
rect 10874 -8080 10908 -7704
rect 10992 -8080 11026 -7704
rect 11110 -8080 11144 -7704
rect 11228 -8080 11262 -7704
rect 11346 -8080 11380 -7704
rect 11752 -7880 11786 -7704
rect 14037 -7480 14139 -7378
rect 22153 -4368 22202 -4308
rect 23364 -4364 23366 -4309
rect 23366 -4364 23424 -4309
rect 23613 -4579 23647 -4545
rect 23126 -4843 23160 -4667
rect 23244 -4843 23278 -4667
rect 23318 -5043 23352 -4667
rect 23436 -5043 23470 -4667
rect 23554 -5043 23588 -4667
rect 23672 -5043 23706 -4667
rect 23790 -5043 23824 -4667
rect 23868 -4843 23902 -4667
rect 23986 -4843 24020 -4667
rect 23555 -5178 23589 -5144
rect 23558 -5310 23616 -5296
rect 23558 -5342 23616 -5310
rect 15303 -6052 15341 -6024
rect 15303 -6062 15341 -6052
rect 14466 -6655 14500 -6479
rect 14584 -6655 14618 -6479
rect 14702 -6655 14736 -6479
rect 14820 -6655 14854 -6479
rect 14950 -6655 14984 -6279
rect 15068 -6655 15102 -6279
rect 15186 -6655 15220 -6279
rect 15304 -6655 15338 -6279
rect 15422 -6655 15456 -6279
rect 15540 -6655 15574 -6279
rect 15658 -6655 15692 -6279
rect 15787 -6655 15821 -6479
rect 15905 -6655 15939 -6479
rect 16023 -6655 16057 -6479
rect 16141 -6655 16175 -6479
rect 15873 -6834 15927 -6824
rect 15873 -6868 15883 -6834
rect 15883 -6868 15917 -6834
rect 15917 -6868 15927 -6834
rect 15873 -6878 15927 -6868
rect 14473 -7028 14539 -7014
rect 14473 -7062 14489 -7028
rect 14489 -7062 14523 -7028
rect 14523 -7062 14539 -7028
rect 14473 -7074 14539 -7062
rect 14893 -7348 14927 -6972
rect 15011 -7348 15045 -6972
rect 15129 -7348 15163 -6972
rect 15247 -7348 15281 -6972
rect 15365 -7348 15399 -6972
rect 15483 -7348 15517 -6972
rect 15601 -7348 15635 -6972
rect 13503 -7572 13537 -7538
rect 14923 -7570 14957 -7536
rect 13121 -7656 13155 -7622
rect 13239 -7655 13273 -7621
rect 13793 -7640 13827 -7606
rect 14738 -7637 14772 -7603
rect 16105 -7478 16207 -7376
rect 16863 -6017 16959 -5981
rect 17601 -6019 17697 -5983
rect 18339 -6019 18435 -5983
rect 19081 -6019 19177 -5983
rect 19821 -6019 19917 -5983
rect 20559 -6019 20655 -5983
rect 21297 -6019 21393 -5983
rect 22035 -6019 22131 -5983
rect 16719 -6343 16753 -6167
rect 16837 -6343 16871 -6167
rect 16955 -6343 16989 -6167
rect 17073 -6343 17107 -6167
rect 17457 -6339 17491 -6163
rect 17575 -6339 17609 -6163
rect 17693 -6339 17727 -6163
rect 17811 -6339 17845 -6163
rect 18195 -6343 18229 -6167
rect 18313 -6343 18347 -6167
rect 18431 -6343 18465 -6167
rect 18549 -6343 18583 -6167
rect 18937 -6345 18971 -6169
rect 19055 -6345 19089 -6169
rect 19173 -6345 19207 -6169
rect 19291 -6345 19325 -6169
rect 19677 -6345 19711 -6169
rect 19795 -6345 19829 -6169
rect 19913 -6345 19947 -6169
rect 20031 -6345 20065 -6169
rect 20415 -6345 20449 -6169
rect 20533 -6345 20567 -6169
rect 20651 -6345 20685 -6169
rect 20769 -6345 20803 -6169
rect 21153 -6345 21187 -6169
rect 21271 -6345 21305 -6169
rect 21389 -6345 21423 -6169
rect 21507 -6345 21541 -6169
rect 21891 -6345 21925 -6169
rect 22009 -6345 22043 -6169
rect 22127 -6345 22161 -6169
rect 22245 -6345 22279 -6169
rect 16895 -6483 16929 -6449
rect 15571 -7570 15605 -7536
rect 15189 -7654 15223 -7620
rect 15307 -7653 15341 -7619
rect 15861 -7638 15895 -7604
rect 11870 -7880 11904 -7704
rect 12523 -7882 12557 -7706
rect 12641 -7882 12675 -7706
rect 12943 -8082 12977 -7706
rect 13061 -8082 13095 -7706
rect 13179 -8082 13213 -7706
rect 13297 -8082 13331 -7706
rect 13415 -8082 13449 -7706
rect 13821 -7882 13855 -7706
rect 13939 -7882 13973 -7706
rect 14591 -7880 14625 -7704
rect 14709 -7880 14743 -7704
rect 15011 -8080 15045 -7704
rect 15129 -8080 15163 -7704
rect 15247 -8080 15281 -7704
rect 15365 -8080 15399 -7704
rect 15483 -8080 15517 -7704
rect 15889 -7880 15923 -7704
rect 16007 -7880 16041 -7704
rect 762 -8272 812 -8250
rect 762 -8292 812 -8272
rect 2830 -8270 2880 -8248
rect 2830 -8290 2880 -8270
rect 4899 -8272 4949 -8250
rect 4899 -8292 4949 -8272
rect 6967 -8270 7017 -8248
rect 6967 -8290 7017 -8270
rect 9036 -8270 9086 -8248
rect 9036 -8290 9086 -8270
rect 11104 -8268 11154 -8246
rect 11104 -8288 11154 -8268
rect 13173 -8270 13223 -8248
rect 13173 -8290 13223 -8270
rect 15241 -8268 15291 -8246
rect 15241 -8288 15291 -8268
rect 17633 -6485 17667 -6451
rect 18371 -6485 18405 -6451
rect 19113 -6485 19147 -6451
rect 19853 -6485 19887 -6451
rect 20591 -6485 20625 -6451
rect 16837 -6729 16871 -6553
rect 16955 -6729 16989 -6553
rect 16813 -6903 16891 -6849
rect 17575 -6727 17609 -6551
rect 17693 -6727 17727 -6551
rect 17551 -6905 17629 -6851
rect 2007 -8710 2058 -8659
rect 4042 -8818 4089 -8764
rect 18313 -6731 18347 -6555
rect 18431 -6731 18465 -6555
rect 18289 -6905 18367 -6851
rect 19055 -6731 19089 -6555
rect 19173 -6731 19207 -6555
rect 19031 -6905 19109 -6851
rect 6089 -8921 6136 -8867
rect 19795 -6731 19829 -6555
rect 19913 -6731 19947 -6555
rect 19771 -6905 19849 -6851
rect 8179 -9028 8229 -8977
rect 21146 -6491 21182 -6445
rect 21329 -6485 21363 -6451
rect 21883 -6491 21921 -6445
rect 22067 -6485 22101 -6451
rect 20533 -6731 20567 -6555
rect 20651 -6731 20685 -6555
rect 20509 -6905 20587 -6851
rect 10250 -9125 10301 -9072
rect 21271 -6727 21305 -6551
rect 21389 -6727 21423 -6551
rect 21247 -6905 21325 -6851
rect 22009 -6727 22043 -6551
rect 22127 -6727 22161 -6551
rect 21985 -6905 22063 -6851
rect 12353 -9267 12397 -9216
rect 14421 -9365 14474 -9311
<< metal1 >>
rect -2585 5863 -2478 5922
rect -2418 5863 -2408 5922
rect 10294 5901 20106 5907
rect 10294 5847 10304 5901
rect 10358 5847 20106 5901
rect 10294 5843 20106 5847
rect -1987 5813 10479 5814
rect -1987 5808 19968 5813
rect -1987 5754 10398 5808
rect 10452 5754 19968 5808
rect -1987 5750 19968 5754
rect -2585 5722 -2448 5725
rect -2585 5660 -2481 5722
rect -2421 5660 -2411 5722
rect -2585 5532 -2458 5536
rect -2585 5470 -2488 5532
rect -2428 5470 -2418 5532
rect -2585 5281 -2488 5350
rect -2428 5281 -2418 5350
rect -2585 5100 -2501 5163
rect -2440 5100 -2430 5163
rect -2585 4900 -2514 4972
rect -2443 4900 -2433 4972
rect -2585 3166 -2501 3167
rect -2585 3111 -2497 3166
rect -2443 3111 -2433 3166
rect -2583 2737 -2526 2791
rect -2470 2737 -2460 2791
rect -2610 -1289 -2505 -1283
rect -2610 -1364 -2507 -1289
rect -2445 -1364 -2435 -1289
rect -2609 -1616 -2504 -1610
rect -2609 -1691 -2506 -1616
rect -2444 -1691 -2434 -1616
rect -1987 -5557 -1908 5750
rect 10388 5749 19968 5750
rect 8759 5716 18938 5721
rect 8759 5662 8766 5716
rect 8820 5662 18938 5716
rect 8759 5657 18938 5662
rect -1711 5628 -1592 5629
rect -1711 5627 -359 5628
rect -1734 5621 18805 5627
rect -1734 5567 8941 5621
rect 8995 5567 18805 5621
rect -1734 5564 18805 5567
rect -2303 -5618 -2237 -5557
rect -2182 -5618 -2172 -5557
rect -1991 -5615 -1981 -5557
rect -1913 -5615 -1903 -5557
rect -2303 -5910 -2237 -5849
rect -2182 -5910 -2172 -5849
rect -2303 -6215 -2237 -6154
rect -2182 -6215 -2172 -6154
rect -2303 -6376 -2237 -6315
rect -2182 -6376 -2172 -6315
rect -2303 -6527 -2237 -6466
rect -2181 -6527 -2171 -6466
rect -2303 -6687 -2237 -6626
rect -2182 -6687 -2172 -6626
rect -2303 -6874 -2237 -6813
rect -2182 -6874 -2172 -6813
rect -2303 -7080 -2237 -7019
rect -2182 -7080 -2172 -7019
rect -1987 -9310 -1908 -5615
rect -1734 -5851 -1654 5564
rect 8631 5563 18805 5564
rect 7295 5531 17770 5535
rect 7295 5477 7305 5531
rect 7359 5477 17770 5531
rect 7295 5471 17770 5477
rect -1734 -5908 -1722 -5851
rect -1666 -5908 -1654 -5851
rect -1734 -9211 -1654 -5908
rect -1505 5441 7516 5443
rect -1505 5437 17642 5441
rect -1505 5383 7443 5437
rect 7497 5383 17642 5437
rect -1505 5379 17642 5383
rect -1505 -6159 -1441 5379
rect 7433 5377 17642 5379
rect 5793 5343 16602 5349
rect 5793 5289 5803 5343
rect 5857 5289 16602 5343
rect 5793 5285 16602 5289
rect 5969 5253 16452 5255
rect -1333 5249 16452 5253
rect -1333 5195 5982 5249
rect 6036 5195 16452 5249
rect -1514 -6212 -1504 -6159
rect -1443 -6212 -1433 -6159
rect -1505 -9112 -1441 -6212
rect -1333 -6316 -1254 5195
rect 5969 5191 16452 5195
rect 4337 5159 15428 5163
rect 4337 5105 4347 5159
rect 4401 5105 15428 5159
rect 4337 5100 15428 5105
rect 10383 5099 15428 5100
rect -1130 5070 -1056 5071
rect -1130 5069 10017 5070
rect -1130 5064 15254 5069
rect -1130 5010 4475 5064
rect 4529 5010 15254 5064
rect -1130 5006 15254 5010
rect -1339 -6374 -1329 -6316
rect -1259 -6374 -1249 -6316
rect -1333 -8984 -1254 -6374
rect -1130 -6466 -1056 5006
rect 10290 5005 15254 5006
rect 2887 4977 10020 4978
rect 2887 4973 14260 4977
rect 2887 4919 2894 4973
rect 2948 4919 14260 4973
rect 2887 4914 14260 4919
rect 10466 4913 14260 4914
rect -933 4883 10020 4884
rect -933 4878 14083 4883
rect -933 4829 3025 4878
rect -1137 -6524 -1127 -6466
rect -1059 -6524 -1049 -6466
rect -1130 -8865 -1056 -6524
rect -933 -6629 -869 4829
rect 3016 4824 3025 4829
rect 3079 4824 14083 4878
rect 3016 4820 14083 4824
rect 10466 4819 14083 4820
rect 1449 4791 8888 4792
rect 1449 4787 13092 4791
rect 1439 4733 1449 4787
rect 1503 4733 13092 4787
rect 1449 4728 13092 4733
rect 10464 4727 13092 4728
rect -694 4698 -168 4699
rect -703 4697 8888 4698
rect -703 4694 12936 4697
rect -703 4640 1559 4694
rect 1613 4640 12936 4694
rect -703 4634 12936 4640
rect -941 -6683 -931 -6629
rect -873 -6683 -863 -6629
rect -933 -8756 -869 -6683
rect -703 -6813 -639 4634
rect 10464 4633 12936 4634
rect -161 4541 11924 4605
rect -161 3468 -98 4541
rect -303 3467 -98 3468
rect -303 3408 -293 3467
rect -222 3408 -98 3467
rect -161 3192 -98 3408
rect 78 4447 11779 4511
rect 78 4248 141 4447
rect 78 3393 142 4248
rect 506 4123 642 4143
rect 506 4061 542 4123
rect 602 4061 642 4123
rect 506 4033 642 4061
rect 1954 4123 2090 4143
rect 1954 4061 1990 4123
rect 2050 4061 2090 4123
rect 1954 4033 2090 4061
rect 3452 4125 3588 4145
rect 3452 4063 3488 4125
rect 3548 4063 3588 4125
rect 3452 4035 3588 4063
rect 4900 4125 5036 4145
rect 4900 4063 4936 4125
rect 4996 4063 5036 4125
rect 4900 4035 5036 4063
rect 6420 4123 6556 4143
rect 6420 4061 6456 4123
rect 6516 4061 6556 4123
rect 202 4003 1179 4033
rect 202 3897 234 4003
rect 438 3897 470 4003
rect 674 3897 706 4003
rect 910 3897 942 4003
rect 1145 3897 1179 4003
rect 1650 4003 2627 4033
rect 1650 3897 1682 4003
rect 1886 3897 1918 4003
rect 2122 3897 2154 4003
rect 2358 3897 2390 4003
rect 2593 3897 2627 4003
rect 3148 4005 4125 4035
rect 3148 3899 3180 4005
rect 3384 3899 3416 4005
rect 3620 3899 3652 4005
rect 3856 3899 3888 4005
rect 4091 3899 4125 4005
rect 4596 4005 5573 4035
rect 6420 4033 6556 4061
rect 7868 4123 8004 4143
rect 7868 4061 7904 4123
rect 7964 4061 8004 4123
rect 7868 4033 8004 4061
rect 9366 4125 9502 4145
rect 9366 4063 9402 4125
rect 9462 4063 9502 4125
rect 9366 4035 9502 4063
rect 10814 4125 10950 4145
rect 10814 4063 10850 4125
rect 10910 4063 10950 4125
rect 10814 4035 10950 4063
rect 11724 4083 11779 4447
rect 11860 4356 11924 4541
rect 11824 4254 11924 4356
rect 11824 4220 11874 4254
rect 11908 4220 11924 4254
rect 12510 4330 12614 4336
rect 12510 4258 12522 4330
rect 12602 4258 12614 4330
rect 12510 4252 12614 4258
rect 11824 4194 11924 4220
rect 12545 4196 12580 4252
rect 11824 4146 11924 4166
rect 11824 4112 11874 4146
rect 11908 4112 11924 4146
rect 11824 4083 11924 4112
rect 12082 4155 12352 4183
rect 12082 4094 12116 4155
rect 12318 4094 12352 4155
rect 12436 4155 12706 4196
rect 12436 4094 12470 4155
rect 12672 4094 12706 4155
rect 12872 4166 12936 4633
rect 13028 4356 13092 4727
rect 12992 4254 13092 4356
rect 12992 4220 13042 4254
rect 13076 4220 13092 4254
rect 13678 4330 13782 4336
rect 13678 4258 13690 4330
rect 13770 4258 13782 4330
rect 13678 4252 13782 4258
rect 12992 4194 13092 4220
rect 13713 4196 13748 4252
rect 12872 4146 13092 4166
rect 12872 4112 13042 4146
rect 13076 4112 13092 4146
rect 12872 4102 13092 4112
rect 4596 3899 4628 4005
rect 4832 3899 4864 4005
rect 5068 3899 5100 4005
rect 5304 3899 5336 4005
rect 5539 3899 5573 4005
rect 6116 4003 7093 4033
rect 195 3885 241 3897
rect 195 3709 201 3885
rect 235 3709 241 3885
rect 195 3697 241 3709
rect 313 3885 359 3897
rect 313 3709 319 3885
rect 353 3709 359 3885
rect 313 3697 359 3709
rect 431 3885 477 3897
rect 431 3709 437 3885
rect 471 3709 477 3885
rect 431 3697 477 3709
rect 549 3885 595 3897
rect 549 3709 555 3885
rect 589 3709 595 3885
rect 549 3697 595 3709
rect 667 3885 713 3897
rect 667 3709 673 3885
rect 707 3709 713 3885
rect 667 3697 713 3709
rect 785 3885 831 3897
rect 785 3709 791 3885
rect 825 3709 831 3885
rect 785 3697 831 3709
rect 903 3885 949 3897
rect 903 3709 909 3885
rect 943 3709 949 3885
rect 903 3697 949 3709
rect 1021 3885 1067 3897
rect 1021 3709 1027 3885
rect 1061 3709 1067 3885
rect 1021 3697 1067 3709
rect 1139 3885 1185 3897
rect 1139 3709 1145 3885
rect 1179 3709 1185 3885
rect 1139 3697 1185 3709
rect 1257 3885 1303 3897
rect 1257 3709 1263 3885
rect 1297 3709 1303 3885
rect 1257 3697 1303 3709
rect 1643 3885 1689 3897
rect 1643 3709 1649 3885
rect 1683 3709 1689 3885
rect 1643 3697 1689 3709
rect 1761 3885 1807 3897
rect 1761 3709 1767 3885
rect 1801 3709 1807 3885
rect 1761 3697 1807 3709
rect 1879 3885 1925 3897
rect 1879 3709 1885 3885
rect 1919 3709 1925 3885
rect 1879 3697 1925 3709
rect 1997 3885 2043 3897
rect 1997 3709 2003 3885
rect 2037 3709 2043 3885
rect 1997 3697 2043 3709
rect 2115 3885 2161 3897
rect 2115 3709 2121 3885
rect 2155 3709 2161 3885
rect 2115 3697 2161 3709
rect 2233 3885 2279 3897
rect 2233 3709 2239 3885
rect 2273 3709 2279 3885
rect 2233 3697 2279 3709
rect 2351 3885 2397 3897
rect 2351 3709 2357 3885
rect 2391 3709 2397 3885
rect 2351 3697 2397 3709
rect 2469 3885 2515 3897
rect 2469 3709 2475 3885
rect 2509 3709 2515 3885
rect 2469 3697 2515 3709
rect 2587 3885 2633 3897
rect 2587 3709 2593 3885
rect 2627 3709 2633 3885
rect 2587 3697 2633 3709
rect 2705 3885 2751 3897
rect 2705 3709 2711 3885
rect 2745 3709 2751 3885
rect 2705 3697 2751 3709
rect 3141 3887 3187 3899
rect 3141 3711 3147 3887
rect 3181 3711 3187 3887
rect 3141 3699 3187 3711
rect 3259 3887 3305 3899
rect 3259 3711 3265 3887
rect 3299 3711 3305 3887
rect 3259 3699 3305 3711
rect 3377 3887 3423 3899
rect 3377 3711 3383 3887
rect 3417 3711 3423 3887
rect 3377 3699 3423 3711
rect 3495 3887 3541 3899
rect 3495 3711 3501 3887
rect 3535 3711 3541 3887
rect 3495 3699 3541 3711
rect 3613 3887 3659 3899
rect 3613 3711 3619 3887
rect 3653 3711 3659 3887
rect 3613 3699 3659 3711
rect 3731 3887 3777 3899
rect 3731 3711 3737 3887
rect 3771 3711 3777 3887
rect 3731 3699 3777 3711
rect 3849 3887 3895 3899
rect 3849 3711 3855 3887
rect 3889 3711 3895 3887
rect 3849 3699 3895 3711
rect 3967 3887 4013 3899
rect 3967 3711 3973 3887
rect 4007 3711 4013 3887
rect 3967 3699 4013 3711
rect 4085 3887 4131 3899
rect 4085 3711 4091 3887
rect 4125 3711 4131 3887
rect 4085 3699 4131 3711
rect 4203 3887 4249 3899
rect 4203 3711 4209 3887
rect 4243 3711 4249 3887
rect 4203 3699 4249 3711
rect 4589 3887 4635 3899
rect 4589 3711 4595 3887
rect 4629 3711 4635 3887
rect 4589 3699 4635 3711
rect 4707 3887 4753 3899
rect 4707 3711 4713 3887
rect 4747 3711 4753 3887
rect 4707 3699 4753 3711
rect 4825 3887 4871 3899
rect 4825 3711 4831 3887
rect 4865 3711 4871 3887
rect 4825 3699 4871 3711
rect 4943 3887 4989 3899
rect 4943 3711 4949 3887
rect 4983 3711 4989 3887
rect 4943 3699 4989 3711
rect 5061 3887 5107 3899
rect 5061 3711 5067 3887
rect 5101 3711 5107 3887
rect 5061 3699 5107 3711
rect 5179 3887 5225 3899
rect 5179 3711 5185 3887
rect 5219 3711 5225 3887
rect 5179 3699 5225 3711
rect 5297 3887 5343 3899
rect 5297 3711 5303 3887
rect 5337 3711 5343 3887
rect 5297 3699 5343 3711
rect 5415 3887 5461 3899
rect 5415 3711 5421 3887
rect 5455 3711 5461 3887
rect 5415 3699 5461 3711
rect 5533 3887 5579 3899
rect 5533 3711 5539 3887
rect 5573 3711 5579 3887
rect 5533 3699 5579 3711
rect 5651 3887 5697 3899
rect 6116 3897 6148 4003
rect 6352 3897 6384 4003
rect 6588 3897 6620 4003
rect 6824 3897 6856 4003
rect 7059 3897 7093 4003
rect 7564 4003 8541 4033
rect 7564 3897 7596 4003
rect 7800 3897 7832 4003
rect 8036 3897 8068 4003
rect 8272 3897 8304 4003
rect 8507 3897 8541 4003
rect 9062 4005 10039 4035
rect 9062 3899 9094 4005
rect 9298 3899 9330 4005
rect 9534 3899 9566 4005
rect 9770 3899 9802 4005
rect 10005 3899 10039 4005
rect 10510 4005 11487 4035
rect 11724 4014 11924 4083
rect 11958 4082 12004 4094
rect 10510 3899 10542 4005
rect 10746 3899 10778 4005
rect 10982 3899 11014 4005
rect 11218 3899 11250 4005
rect 11453 3899 11487 4005
rect 5651 3711 5657 3887
rect 5691 3711 5697 3887
rect 5651 3699 5697 3711
rect 6109 3885 6155 3897
rect 6109 3709 6115 3885
rect 6149 3709 6155 3885
rect 318 3603 354 3697
rect 554 3603 590 3697
rect 790 3604 826 3697
rect 952 3649 1018 3656
rect 952 3615 968 3649
rect 1002 3615 1018 3649
rect 952 3604 1018 3615
rect 790 3603 1018 3604
rect 318 3574 1018 3603
rect 318 3573 900 3574
rect 438 3460 472 3573
rect 834 3532 900 3573
rect 834 3498 850 3532
rect 884 3498 900 3532
rect 834 3491 900 3498
rect 1262 3464 1297 3697
rect 1766 3603 1802 3697
rect 2002 3603 2038 3697
rect 2238 3604 2274 3697
rect 2400 3649 2466 3656
rect 2400 3615 2416 3649
rect 2450 3615 2466 3649
rect 2400 3604 2466 3615
rect 2238 3603 2466 3604
rect 1766 3574 2466 3603
rect 1766 3573 2348 3574
rect 908 3460 1297 3464
rect 1886 3460 1920 3573
rect 2282 3532 2348 3573
rect 2282 3498 2298 3532
rect 2332 3498 2348 3532
rect 2282 3491 2348 3498
rect 2710 3464 2745 3697
rect 3264 3605 3300 3699
rect 3500 3605 3536 3699
rect 3736 3606 3772 3699
rect 3898 3651 3964 3658
rect 3898 3617 3914 3651
rect 3948 3617 3964 3651
rect 3898 3606 3964 3617
rect 3736 3605 3964 3606
rect 3264 3576 3964 3605
rect 3264 3575 3846 3576
rect 2356 3460 2745 3464
rect 3384 3462 3418 3575
rect 3780 3534 3846 3575
rect 3780 3500 3796 3534
rect 3830 3500 3846 3534
rect 3780 3493 3846 3500
rect 4208 3466 4243 3699
rect 4712 3605 4748 3699
rect 4948 3605 4984 3699
rect 5184 3606 5220 3699
rect 5346 3651 5412 3658
rect 5346 3617 5362 3651
rect 5396 3617 5412 3651
rect 5346 3606 5412 3617
rect 5184 3605 5412 3606
rect 4712 3576 5412 3605
rect 4712 3575 5294 3576
rect 3854 3462 4243 3466
rect 4832 3462 4866 3575
rect 5228 3534 5294 3575
rect 5228 3500 5244 3534
rect 5278 3500 5294 3534
rect 5228 3493 5294 3500
rect 5656 3466 5691 3699
rect 6109 3697 6155 3709
rect 6227 3885 6273 3897
rect 6227 3709 6233 3885
rect 6267 3709 6273 3885
rect 6227 3697 6273 3709
rect 6345 3885 6391 3897
rect 6345 3709 6351 3885
rect 6385 3709 6391 3885
rect 6345 3697 6391 3709
rect 6463 3885 6509 3897
rect 6463 3709 6469 3885
rect 6503 3709 6509 3885
rect 6463 3697 6509 3709
rect 6581 3885 6627 3897
rect 6581 3709 6587 3885
rect 6621 3709 6627 3885
rect 6581 3697 6627 3709
rect 6699 3885 6745 3897
rect 6699 3709 6705 3885
rect 6739 3709 6745 3885
rect 6699 3697 6745 3709
rect 6817 3885 6863 3897
rect 6817 3709 6823 3885
rect 6857 3709 6863 3885
rect 6817 3697 6863 3709
rect 6935 3885 6981 3897
rect 6935 3709 6941 3885
rect 6975 3709 6981 3885
rect 6935 3697 6981 3709
rect 7053 3885 7099 3897
rect 7053 3709 7059 3885
rect 7093 3709 7099 3885
rect 7053 3697 7099 3709
rect 7171 3885 7217 3897
rect 7171 3709 7177 3885
rect 7211 3709 7217 3885
rect 7171 3697 7217 3709
rect 7557 3885 7603 3897
rect 7557 3709 7563 3885
rect 7597 3709 7603 3885
rect 7557 3697 7603 3709
rect 7675 3885 7721 3897
rect 7675 3709 7681 3885
rect 7715 3709 7721 3885
rect 7675 3697 7721 3709
rect 7793 3885 7839 3897
rect 7793 3709 7799 3885
rect 7833 3709 7839 3885
rect 7793 3697 7839 3709
rect 7911 3885 7957 3897
rect 7911 3709 7917 3885
rect 7951 3709 7957 3885
rect 7911 3697 7957 3709
rect 8029 3885 8075 3897
rect 8029 3709 8035 3885
rect 8069 3709 8075 3885
rect 8029 3697 8075 3709
rect 8147 3885 8193 3897
rect 8147 3709 8153 3885
rect 8187 3709 8193 3885
rect 8147 3697 8193 3709
rect 8265 3885 8311 3897
rect 8265 3709 8271 3885
rect 8305 3709 8311 3885
rect 8265 3697 8311 3709
rect 8383 3885 8429 3897
rect 8383 3709 8389 3885
rect 8423 3709 8429 3885
rect 8383 3697 8429 3709
rect 8501 3885 8547 3897
rect 8501 3709 8507 3885
rect 8541 3709 8547 3885
rect 8501 3697 8547 3709
rect 8619 3885 8665 3897
rect 8619 3709 8625 3885
rect 8659 3709 8665 3885
rect 8619 3697 8665 3709
rect 9055 3887 9101 3899
rect 9055 3711 9061 3887
rect 9095 3711 9101 3887
rect 9055 3699 9101 3711
rect 9173 3887 9219 3899
rect 9173 3711 9179 3887
rect 9213 3711 9219 3887
rect 9173 3699 9219 3711
rect 9291 3887 9337 3899
rect 9291 3711 9297 3887
rect 9331 3711 9337 3887
rect 9291 3699 9337 3711
rect 9409 3887 9455 3899
rect 9409 3711 9415 3887
rect 9449 3711 9455 3887
rect 9409 3699 9455 3711
rect 9527 3887 9573 3899
rect 9527 3711 9533 3887
rect 9567 3711 9573 3887
rect 9527 3699 9573 3711
rect 9645 3887 9691 3899
rect 9645 3711 9651 3887
rect 9685 3711 9691 3887
rect 9645 3699 9691 3711
rect 9763 3887 9809 3899
rect 9763 3711 9769 3887
rect 9803 3711 9809 3887
rect 9763 3699 9809 3711
rect 9881 3887 9927 3899
rect 9881 3711 9887 3887
rect 9921 3711 9927 3887
rect 9881 3699 9927 3711
rect 9999 3887 10045 3899
rect 9999 3711 10005 3887
rect 10039 3711 10045 3887
rect 9999 3699 10045 3711
rect 10117 3887 10163 3899
rect 10117 3711 10123 3887
rect 10157 3711 10163 3887
rect 10117 3699 10163 3711
rect 10503 3887 10549 3899
rect 10503 3711 10509 3887
rect 10543 3711 10549 3887
rect 10503 3699 10549 3711
rect 10621 3887 10667 3899
rect 10621 3711 10627 3887
rect 10661 3711 10667 3887
rect 10621 3699 10667 3711
rect 10739 3887 10785 3899
rect 10739 3711 10745 3887
rect 10779 3711 10785 3887
rect 10739 3699 10785 3711
rect 10857 3887 10903 3899
rect 10857 3711 10863 3887
rect 10897 3711 10903 3887
rect 10857 3699 10903 3711
rect 10975 3887 11021 3899
rect 10975 3711 10981 3887
rect 11015 3711 11021 3887
rect 10975 3699 11021 3711
rect 11093 3887 11139 3899
rect 11093 3711 11099 3887
rect 11133 3711 11139 3887
rect 11093 3699 11139 3711
rect 11211 3887 11257 3899
rect 11211 3711 11217 3887
rect 11251 3711 11257 3887
rect 11211 3699 11257 3711
rect 11329 3887 11375 3899
rect 11329 3711 11335 3887
rect 11369 3711 11375 3887
rect 11329 3699 11375 3711
rect 11447 3887 11493 3899
rect 11447 3711 11453 3887
rect 11487 3711 11493 3887
rect 11447 3699 11493 3711
rect 11565 3887 11611 3899
rect 11565 3711 11571 3887
rect 11605 3711 11611 3887
rect 11565 3699 11611 3711
rect 11958 3706 11964 4082
rect 11998 3706 12004 4082
rect 6232 3603 6268 3697
rect 6468 3603 6504 3697
rect 6704 3604 6740 3697
rect 6866 3649 6932 3656
rect 6866 3615 6882 3649
rect 6916 3615 6932 3649
rect 6866 3604 6932 3615
rect 6704 3603 6932 3604
rect 6232 3574 6932 3603
rect 6232 3573 6814 3574
rect 5302 3462 5691 3466
rect -17 3371 142 3393
rect -17 3307 -7 3371
rect 62 3320 142 3371
rect 432 3448 478 3460
rect 62 3307 392 3320
rect -17 3296 392 3307
rect 78 3220 392 3296
rect -161 3092 280 3192
rect 202 2943 256 3092
rect 316 3028 370 3220
rect 432 3072 438 3448
rect 472 3072 478 3448
rect 432 3060 478 3072
rect 550 3448 596 3460
rect 550 3072 556 3448
rect 590 3072 596 3448
rect 550 3060 596 3072
rect 668 3448 714 3460
rect 668 3072 674 3448
rect 708 3099 714 3448
rect 785 3448 831 3460
rect 785 3272 791 3448
rect 825 3272 831 3448
rect 785 3265 831 3272
rect 903 3448 1297 3460
rect 903 3272 909 3448
rect 943 3442 1297 3448
rect 1880 3448 1926 3460
rect 943 3435 1298 3442
rect 943 3272 949 3435
rect 1190 3302 1298 3435
rect 1190 3280 1299 3302
rect 785 3260 834 3265
rect 903 3260 949 3272
rect 791 3099 834 3260
rect 708 3072 834 3099
rect 668 3060 834 3072
rect 674 3056 834 3060
rect 316 3022 547 3028
rect 316 2988 497 3022
rect 531 2988 547 3022
rect 316 2972 547 2988
rect 599 3022 665 3028
rect 599 2988 615 3022
rect 649 2988 665 3022
rect 599 2943 665 2988
rect 202 2935 665 2943
rect 202 2903 666 2935
rect 758 2919 834 3056
rect 754 2859 764 2919
rect 826 2859 836 2919
rect 1191 2753 1299 3280
rect 1740 3298 1840 3320
rect 1740 3244 1766 3298
rect 1820 3244 1840 3298
rect 1740 3220 1840 3244
rect 1628 3167 1728 3192
rect 1628 3112 1651 3167
rect 1705 3112 1728 3167
rect 1628 3092 1728 3112
rect 1650 2943 1704 3092
rect 1764 3028 1818 3220
rect 1880 3072 1886 3448
rect 1920 3072 1926 3448
rect 1880 3060 1926 3072
rect 1998 3448 2044 3460
rect 1998 3072 2004 3448
rect 2038 3072 2044 3448
rect 1998 3060 2044 3072
rect 2116 3448 2162 3460
rect 2116 3072 2122 3448
rect 2156 3099 2162 3448
rect 2233 3448 2279 3460
rect 2233 3272 2239 3448
rect 2273 3272 2279 3448
rect 2233 3265 2279 3272
rect 2351 3448 2745 3460
rect 2351 3272 2357 3448
rect 2391 3435 2745 3448
rect 2391 3272 2397 3435
rect 2233 3260 2282 3265
rect 2351 3260 2397 3272
rect 2239 3099 2282 3260
rect 2156 3072 2282 3099
rect 2116 3060 2282 3072
rect 2122 3056 2282 3060
rect 1764 3022 1995 3028
rect 1764 2988 1945 3022
rect 1979 2988 1995 3022
rect 1764 2972 1995 2988
rect 2047 3022 2113 3028
rect 2047 2988 2063 3022
rect 2097 2988 2113 3022
rect 2047 2943 2113 2988
rect 1650 2935 2113 2943
rect 1650 2903 2114 2935
rect 2206 2919 2282 3056
rect 2202 2859 2212 2919
rect 2274 2859 2284 2919
rect 1191 2624 1297 2753
rect -1 2578 1297 2624
rect 2641 2624 2745 3435
rect 3378 3450 3424 3462
rect 3238 3297 3338 3322
rect 3238 3243 3260 3297
rect 3314 3243 3338 3297
rect 3238 3222 3338 3243
rect 3126 3165 3226 3194
rect 3126 3111 3149 3165
rect 3203 3111 3226 3165
rect 3126 3094 3226 3111
rect 3148 2945 3202 3094
rect 3262 3030 3316 3222
rect 3378 3074 3384 3450
rect 3418 3074 3424 3450
rect 3378 3062 3424 3074
rect 3496 3450 3542 3462
rect 3496 3074 3502 3450
rect 3536 3074 3542 3450
rect 3496 3062 3542 3074
rect 3614 3450 3660 3462
rect 3614 3074 3620 3450
rect 3654 3101 3660 3450
rect 3731 3450 3777 3462
rect 3731 3274 3737 3450
rect 3771 3274 3777 3450
rect 3731 3267 3777 3274
rect 3849 3450 4243 3462
rect 3849 3274 3855 3450
rect 3889 3437 4243 3450
rect 3889 3274 3895 3437
rect 3731 3262 3780 3267
rect 3849 3262 3895 3274
rect 3737 3101 3780 3262
rect 3654 3074 3780 3101
rect 3614 3062 3780 3074
rect 3620 3058 3780 3062
rect 3262 3024 3493 3030
rect 3262 2990 3443 3024
rect 3477 2990 3493 3024
rect 3262 2974 3493 2990
rect 3545 3024 3611 3030
rect 3545 2990 3561 3024
rect 3595 2990 3611 3024
rect 3545 2945 3611 2990
rect 3148 2937 3611 2945
rect 3148 2905 3612 2937
rect 3704 2921 3780 3058
rect 3700 2861 3710 2921
rect 3772 2861 3782 2921
rect -1 2531 1296 2578
rect 2641 2531 3231 2624
rect -519 1444 -409 1451
rect -519 1356 -503 1444
rect -420 1366 -409 1444
rect -420 1356 -410 1366
rect -519 -1467 -410 1356
rect -1 1334 86 2531
rect 1160 2530 1296 2531
rect 1498 2324 1508 2384
rect 1588 2324 1598 2384
rect 1498 2284 1598 2324
rect 701 2227 2504 2284
rect 701 2140 735 2227
rect 1876 2140 1910 2227
rect 695 2128 741 2140
rect 695 1940 701 2128
rect 254 1928 300 1940
rect 254 1752 260 1928
rect 294 1752 300 1928
rect 254 1740 300 1752
rect 372 1928 418 1940
rect 372 1752 378 1928
rect 412 1752 418 1928
rect 372 1740 418 1752
rect 490 1928 536 1940
rect 490 1752 496 1928
rect 530 1752 536 1928
rect 490 1740 536 1752
rect 608 1928 701 1940
rect 608 1752 614 1928
rect 648 1752 701 1928
rect 735 1752 741 2128
rect 608 1740 741 1752
rect 813 2128 859 2140
rect 813 1752 819 2128
rect 853 1752 859 2128
rect 813 1740 859 1752
rect 931 2128 977 2140
rect 931 1752 937 2128
rect 971 1752 977 2128
rect 931 1740 977 1752
rect 1049 2128 1095 2140
rect 1049 1752 1055 2128
rect 1089 1752 1095 2128
rect 1049 1740 1095 1752
rect 1162 2128 1208 2140
rect 1162 1752 1168 2128
rect 1202 1752 1208 2128
rect 1162 1740 1208 1752
rect 1280 2128 1326 2140
rect 1280 1752 1286 2128
rect 1320 1752 1326 2128
rect 1280 1740 1326 1752
rect 1398 2128 1444 2140
rect 1398 1752 1404 2128
rect 1438 1752 1444 2128
rect 1398 1740 1444 1752
rect 1516 2128 1562 2140
rect 1516 1752 1522 2128
rect 1556 1752 1562 2128
rect 1516 1740 1562 1752
rect 1634 2128 1680 2140
rect 1634 1752 1640 2128
rect 1674 1752 1680 2128
rect 1634 1740 1680 1752
rect 1752 2128 1798 2140
rect 1752 1752 1758 2128
rect 1792 1752 1798 2128
rect 1752 1740 1798 1752
rect 1870 2128 1916 2140
rect 1870 1752 1876 2128
rect 1910 1752 1916 2128
rect 1870 1740 1916 1752
rect 1989 2128 2035 2140
rect 1989 1752 1995 2128
rect 2029 1752 2035 2128
rect 1989 1740 2035 1752
rect 2107 2128 2153 2140
rect 2107 1752 2113 2128
rect 2147 1752 2153 2128
rect 2107 1740 2153 1752
rect 2225 2128 2271 2140
rect 2225 1752 2231 2128
rect 2265 1752 2271 2128
rect 2225 1740 2271 1752
rect 2343 2128 2389 2140
rect 2343 1752 2349 2128
rect 2383 1752 2389 2128
rect 2467 1940 2504 2227
rect 2343 1740 2389 1752
rect 2462 1928 2508 1940
rect 2462 1752 2468 1928
rect 2502 1752 2508 1928
rect 2462 1740 2508 1752
rect 2580 1928 2626 1940
rect 2580 1752 2586 1928
rect 2620 1752 2626 1928
rect 2580 1740 2626 1752
rect 2698 1928 2744 1940
rect 2698 1752 2704 1928
rect 2738 1752 2744 1928
rect 2698 1740 2744 1752
rect 2816 1928 2862 1940
rect 2816 1752 2822 1928
rect 2856 1752 2862 1928
rect 2816 1740 2862 1752
rect 259 1554 294 1740
rect 1168 1656 1202 1740
rect 2349 1656 2383 1740
rect 1168 1614 2383 1656
rect 2349 1594 2383 1614
rect 2349 1578 2706 1594
rect 259 1537 1396 1554
rect 259 1503 1346 1537
rect 1380 1503 1396 1537
rect 2349 1544 2656 1578
rect 2690 1544 2706 1578
rect 2349 1528 2706 1544
rect 259 1487 1396 1503
rect -1 1326 176 1334
rect -1 1258 117 1326
rect 174 1258 184 1326
rect -1 1250 176 1258
rect 103 1158 176 1166
rect 103 1090 117 1158
rect 174 1090 184 1158
rect 103 1082 176 1090
rect 259 977 294 1487
rect 349 1441 441 1454
rect 349 1378 361 1441
rect 432 1378 441 1441
rect 349 1369 441 1378
rect 1434 1441 1526 1451
rect 1434 1379 1446 1441
rect 1516 1379 1526 1441
rect 1434 1366 1526 1379
rect 2822 1386 2857 1740
rect 1681 1324 1746 1327
rect 1681 1321 1750 1324
rect 1681 1261 1687 1321
rect 1746 1261 1756 1321
rect 1681 1257 1750 1261
rect 1681 1255 1746 1257
rect 2822 1240 3003 1386
rect 3144 1334 3231 2531
rect 4139 2588 4243 3437
rect 4826 3450 4872 3462
rect 4686 3300 4786 3322
rect 4686 3246 4710 3300
rect 4764 3246 4786 3300
rect 4686 3222 4786 3246
rect 4574 3170 4674 3194
rect 4574 3116 4597 3170
rect 4651 3116 4674 3170
rect 4574 3094 4674 3116
rect 4596 2945 4650 3094
rect 4710 3030 4764 3222
rect 4826 3074 4832 3450
rect 4866 3074 4872 3450
rect 4826 3062 4872 3074
rect 4944 3450 4990 3462
rect 4944 3074 4950 3450
rect 4984 3074 4990 3450
rect 4944 3062 4990 3074
rect 5062 3450 5108 3462
rect 5062 3074 5068 3450
rect 5102 3101 5108 3450
rect 5179 3450 5225 3462
rect 5179 3274 5185 3450
rect 5219 3274 5225 3450
rect 5179 3267 5225 3274
rect 5297 3450 5691 3462
rect 6352 3460 6386 3573
rect 6748 3532 6814 3573
rect 6748 3498 6764 3532
rect 6798 3498 6814 3532
rect 6748 3491 6814 3498
rect 7176 3464 7211 3697
rect 7680 3603 7716 3697
rect 7916 3603 7952 3697
rect 8152 3604 8188 3697
rect 8314 3649 8380 3656
rect 8314 3615 8330 3649
rect 8364 3615 8380 3649
rect 8314 3604 8380 3615
rect 8152 3603 8380 3604
rect 7680 3574 8380 3603
rect 7680 3573 8262 3574
rect 6822 3460 7211 3464
rect 7800 3460 7834 3573
rect 8196 3532 8262 3573
rect 8196 3498 8212 3532
rect 8246 3498 8262 3532
rect 8196 3491 8262 3498
rect 8624 3464 8659 3697
rect 9178 3605 9214 3699
rect 9414 3605 9450 3699
rect 9650 3606 9686 3699
rect 9812 3651 9878 3658
rect 9812 3617 9828 3651
rect 9862 3617 9878 3651
rect 9812 3606 9878 3617
rect 9650 3605 9878 3606
rect 9178 3576 9878 3605
rect 9178 3575 9760 3576
rect 8270 3460 8659 3464
rect 9298 3462 9332 3575
rect 9694 3534 9760 3575
rect 9694 3500 9710 3534
rect 9744 3500 9760 3534
rect 9694 3493 9760 3500
rect 10122 3466 10157 3699
rect 10626 3605 10662 3699
rect 10862 3605 10898 3699
rect 11098 3606 11134 3699
rect 11260 3651 11326 3658
rect 11260 3617 11276 3651
rect 11310 3617 11326 3651
rect 11260 3606 11326 3617
rect 11098 3605 11326 3606
rect 10626 3576 11326 3605
rect 10626 3575 11208 3576
rect 9768 3462 10157 3466
rect 10746 3462 10780 3575
rect 11142 3534 11208 3575
rect 11142 3500 11158 3534
rect 11192 3500 11208 3534
rect 11142 3493 11208 3500
rect 11570 3466 11605 3699
rect 11958 3694 12004 3706
rect 12076 4082 12122 4094
rect 12076 3706 12082 4082
rect 12116 3706 12122 4082
rect 12076 3694 12122 3706
rect 12194 4082 12240 4094
rect 12194 3706 12200 4082
rect 12234 3706 12240 4082
rect 12194 3694 12240 3706
rect 12312 4082 12358 4094
rect 12312 3706 12318 4082
rect 12352 3706 12358 4082
rect 12312 3694 12358 3706
rect 12430 4082 12476 4094
rect 12430 3706 12436 4082
rect 12470 3706 12476 4082
rect 12430 3694 12476 3706
rect 12548 4082 12594 4094
rect 12548 3706 12554 4082
rect 12588 3706 12594 4082
rect 12548 3694 12594 3706
rect 12666 4082 12712 4094
rect 12666 3706 12672 4082
rect 12706 3706 12712 4082
rect 12992 4014 13092 4102
rect 13250 4155 13520 4183
rect 13250 4094 13284 4155
rect 13486 4094 13520 4155
rect 13604 4155 13874 4196
rect 13604 4094 13638 4155
rect 13840 4094 13874 4155
rect 14019 4166 14083 4819
rect 14196 4356 14260 4913
rect 14160 4254 14260 4356
rect 14160 4220 14210 4254
rect 14244 4220 14260 4254
rect 14846 4330 14950 4336
rect 14846 4258 14858 4330
rect 14938 4258 14950 4330
rect 14846 4252 14950 4258
rect 14160 4194 14260 4220
rect 14881 4196 14916 4252
rect 14019 4146 14260 4166
rect 14019 4112 14210 4146
rect 14244 4112 14260 4146
rect 14019 4102 14260 4112
rect 13126 4082 13172 4094
rect 12666 3694 12712 3706
rect 13126 3706 13132 4082
rect 13166 3706 13172 4082
rect 13126 3694 13172 3706
rect 13244 4082 13290 4094
rect 13244 3706 13250 4082
rect 13284 3706 13290 4082
rect 13244 3694 13290 3706
rect 13362 4082 13408 4094
rect 13362 3706 13368 4082
rect 13402 3706 13408 4082
rect 13362 3694 13408 3706
rect 13480 4082 13526 4094
rect 13480 3706 13486 4082
rect 13520 3706 13526 4082
rect 13480 3694 13526 3706
rect 13598 4082 13644 4094
rect 13598 3706 13604 4082
rect 13638 3706 13644 4082
rect 13598 3694 13644 3706
rect 13716 4082 13762 4094
rect 13716 3706 13722 4082
rect 13756 3706 13762 4082
rect 13716 3694 13762 3706
rect 13834 4082 13880 4094
rect 13834 3706 13840 4082
rect 13874 3706 13880 4082
rect 14160 4014 14260 4102
rect 14418 4155 14688 4183
rect 14418 4092 14452 4155
rect 14654 4092 14688 4155
rect 14772 4155 15042 4196
rect 14772 4092 14806 4155
rect 15008 4092 15042 4155
rect 15190 4166 15254 5005
rect 15364 4356 15428 5099
rect 15328 4254 15428 4356
rect 15328 4220 15378 4254
rect 15412 4220 15428 4254
rect 16014 4330 16118 4336
rect 16014 4258 16026 4330
rect 16106 4258 16118 4330
rect 16014 4252 16118 4258
rect 15328 4194 15428 4220
rect 16049 4196 16084 4252
rect 15190 4146 15428 4166
rect 15190 4112 15378 4146
rect 15412 4112 15428 4146
rect 15190 4102 15428 4112
rect 14294 4080 14340 4092
rect 13834 3694 13880 3706
rect 14294 3704 14300 4080
rect 14334 3704 14340 4080
rect 11964 3651 11998 3694
rect 12200 3651 12234 3694
rect 11964 3623 12234 3651
rect 12318 3652 12352 3694
rect 12554 3652 12588 3694
rect 12318 3623 12588 3652
rect 11964 3575 11998 3623
rect 11964 3545 12027 3575
rect 11216 3462 11605 3466
rect 5297 3274 5303 3450
rect 5337 3437 5691 3450
rect 5337 3274 5343 3437
rect 5179 3262 5228 3267
rect 5297 3262 5343 3274
rect 5185 3101 5228 3262
rect 5102 3074 5228 3101
rect 5062 3062 5228 3074
rect 5068 3058 5228 3062
rect 4710 3024 4941 3030
rect 4710 2990 4891 3024
rect 4925 2990 4941 3024
rect 4710 2974 4941 2990
rect 4993 3024 5059 3030
rect 4993 2990 5009 3024
rect 5043 2990 5059 3024
rect 4993 2945 5059 2990
rect 4596 2937 5059 2945
rect 4596 2905 5060 2937
rect 5152 2921 5228 3058
rect 5148 2861 5158 2921
rect 5220 2861 5230 2921
rect 5587 2688 5691 3437
rect 6346 3448 6392 3460
rect 6206 3295 6306 3320
rect 6206 3241 6229 3295
rect 6283 3241 6306 3295
rect 6206 3220 6306 3241
rect 6094 3170 6194 3192
rect 6094 3116 6113 3170
rect 6167 3116 6194 3170
rect 6094 3092 6194 3116
rect 6116 2943 6170 3092
rect 6230 3028 6284 3220
rect 6346 3072 6352 3448
rect 6386 3072 6392 3448
rect 6346 3060 6392 3072
rect 6464 3448 6510 3460
rect 6464 3072 6470 3448
rect 6504 3072 6510 3448
rect 6464 3060 6510 3072
rect 6582 3448 6628 3460
rect 6582 3072 6588 3448
rect 6622 3099 6628 3448
rect 6699 3448 6745 3460
rect 6699 3272 6705 3448
rect 6739 3272 6745 3448
rect 6699 3265 6745 3272
rect 6817 3448 7211 3460
rect 6817 3272 6823 3448
rect 6857 3435 7211 3448
rect 6857 3272 6863 3435
rect 6699 3260 6748 3265
rect 6817 3260 6863 3272
rect 6705 3099 6748 3260
rect 6622 3072 6748 3099
rect 6582 3060 6748 3072
rect 6588 3056 6748 3060
rect 6230 3022 6461 3028
rect 6230 2988 6411 3022
rect 6445 2988 6461 3022
rect 6230 2972 6461 2988
rect 6513 3022 6579 3028
rect 6513 2988 6529 3022
rect 6563 2988 6579 3022
rect 6513 2943 6579 2988
rect 6116 2935 6579 2943
rect 6116 2903 6580 2935
rect 6672 2919 6748 3056
rect 6668 2859 6678 2919
rect 6740 2859 6750 2919
rect 7107 2693 7211 3435
rect 7794 3448 7840 3460
rect 7654 3302 7754 3320
rect 7654 3248 7677 3302
rect 7731 3248 7754 3302
rect 7654 3220 7754 3248
rect 7542 3164 7642 3192
rect 7542 3110 7565 3164
rect 7619 3110 7642 3164
rect 7542 3092 7642 3110
rect 7564 2943 7618 3092
rect 7678 3028 7732 3220
rect 7794 3072 7800 3448
rect 7834 3072 7840 3448
rect 7794 3060 7840 3072
rect 7912 3448 7958 3460
rect 7912 3072 7918 3448
rect 7952 3072 7958 3448
rect 7912 3060 7958 3072
rect 8030 3448 8076 3460
rect 8030 3072 8036 3448
rect 8070 3099 8076 3448
rect 8147 3448 8193 3460
rect 8147 3272 8153 3448
rect 8187 3272 8193 3448
rect 8147 3265 8193 3272
rect 8265 3448 8659 3460
rect 8265 3272 8271 3448
rect 8305 3435 8659 3448
rect 8305 3272 8311 3435
rect 8147 3260 8196 3265
rect 8265 3260 8311 3272
rect 8153 3099 8196 3260
rect 8070 3072 8196 3099
rect 8030 3060 8196 3072
rect 8036 3056 8196 3060
rect 7678 3022 7909 3028
rect 7678 2988 7859 3022
rect 7893 2988 7909 3022
rect 7678 2972 7909 2988
rect 7961 3022 8027 3028
rect 7961 2988 7977 3022
rect 8011 2988 8027 3022
rect 7961 2943 8027 2988
rect 7564 2935 8027 2943
rect 7564 2903 8028 2935
rect 8120 2919 8196 3056
rect 8116 2859 8126 2919
rect 8188 2859 8198 2919
rect 8555 2782 8659 3435
rect 9292 3450 9338 3462
rect 9152 3300 9252 3322
rect 9152 3246 9174 3300
rect 9228 3246 9252 3300
rect 9152 3222 9252 3246
rect 9040 3170 9140 3194
rect 9040 3116 9062 3170
rect 9116 3116 9140 3170
rect 9040 3094 9140 3116
rect 9062 2945 9116 3094
rect 9176 3030 9230 3222
rect 9292 3074 9298 3450
rect 9332 3074 9338 3450
rect 9292 3062 9338 3074
rect 9410 3450 9456 3462
rect 9410 3074 9416 3450
rect 9450 3074 9456 3450
rect 9410 3062 9456 3074
rect 9528 3450 9574 3462
rect 9528 3074 9534 3450
rect 9568 3101 9574 3450
rect 9645 3450 9691 3462
rect 9645 3274 9651 3450
rect 9685 3274 9691 3450
rect 9645 3267 9691 3274
rect 9763 3450 10157 3462
rect 9763 3274 9769 3450
rect 9803 3437 10157 3450
rect 9803 3274 9809 3437
rect 9645 3262 9694 3267
rect 9763 3262 9809 3274
rect 9651 3101 9694 3262
rect 9568 3074 9694 3101
rect 9528 3062 9694 3074
rect 9534 3058 9694 3062
rect 9176 3024 9407 3030
rect 9176 2990 9357 3024
rect 9391 2990 9407 3024
rect 9176 2974 9407 2990
rect 9459 3024 9525 3030
rect 9459 2990 9475 3024
rect 9509 2990 9525 3024
rect 9459 2945 9525 2990
rect 9062 2937 9525 2945
rect 9062 2905 9526 2937
rect 9618 2921 9694 3058
rect 9614 2861 9624 2921
rect 9686 2861 9696 2921
rect 8555 2722 9722 2782
rect 10053 2772 10157 3437
rect 10740 3450 10786 3462
rect 10600 3316 10700 3322
rect 10596 3228 10606 3316
rect 10692 3228 10702 3316
rect 10600 3222 10700 3228
rect 10488 3187 10588 3194
rect 10482 3099 10492 3187
rect 10578 3099 10588 3187
rect 10488 3094 10588 3099
rect 10510 2945 10564 3094
rect 10624 3030 10678 3222
rect 10740 3074 10746 3450
rect 10780 3074 10786 3450
rect 10740 3062 10786 3074
rect 10858 3450 10904 3462
rect 10858 3074 10864 3450
rect 10898 3074 10904 3450
rect 10858 3062 10904 3074
rect 10976 3450 11022 3462
rect 10976 3074 10982 3450
rect 11016 3101 11022 3450
rect 11093 3450 11139 3462
rect 11093 3274 11099 3450
rect 11133 3274 11139 3450
rect 11093 3267 11139 3274
rect 11211 3450 11605 3462
rect 11211 3274 11217 3450
rect 11251 3437 11605 3450
rect 11251 3274 11257 3437
rect 11093 3262 11142 3267
rect 11211 3262 11257 3274
rect 11099 3101 11142 3262
rect 11016 3074 11142 3101
rect 10976 3062 11142 3074
rect 10982 3058 11142 3062
rect 10624 3024 10855 3030
rect 10624 2990 10805 3024
rect 10839 2990 10855 3024
rect 10624 2974 10855 2990
rect 10907 3024 10973 3030
rect 10907 2990 10923 3024
rect 10957 2990 10973 3024
rect 10907 2945 10973 2990
rect 10510 2937 10973 2945
rect 10510 2905 10974 2937
rect 11066 2921 11142 3058
rect 11062 2861 11072 2921
rect 11134 2861 11144 2921
rect 11501 2848 11605 3437
rect 11992 3453 12027 3545
rect 12672 3510 12706 3694
rect 13132 3651 13166 3694
rect 13368 3651 13402 3694
rect 13132 3623 13402 3651
rect 13486 3652 13520 3694
rect 13722 3652 13756 3694
rect 13486 3623 13756 3652
rect 13132 3575 13166 3623
rect 13132 3545 13195 3575
rect 12672 3456 12781 3510
rect 11992 3417 12219 3453
rect 11992 3308 12027 3417
rect 12153 3383 12219 3417
rect 12153 3349 12169 3383
rect 12203 3349 12219 3383
rect 12153 3343 12219 3349
rect 11868 3296 11914 3308
rect 11868 3120 11874 3296
rect 11908 3120 11914 3296
rect 11868 3108 11914 3120
rect 11986 3296 12032 3308
rect 11986 3120 11992 3296
rect 12026 3120 12032 3296
rect 11986 3108 12032 3120
rect 12104 3296 12150 3308
rect 12104 3120 12110 3296
rect 12144 3120 12150 3296
rect 12104 3108 12150 3120
rect 12222 3296 12268 3308
rect 12630 3304 12663 3335
rect 12747 3304 12781 3456
rect 13160 3453 13195 3545
rect 13840 3510 13874 3694
rect 14294 3692 14340 3704
rect 14412 4080 14458 4092
rect 14412 3704 14418 4080
rect 14452 3704 14458 4080
rect 14412 3692 14458 3704
rect 14530 4080 14576 4092
rect 14530 3704 14536 4080
rect 14570 3704 14576 4080
rect 14530 3692 14576 3704
rect 14648 4080 14694 4092
rect 14648 3704 14654 4080
rect 14688 3704 14694 4080
rect 14648 3692 14694 3704
rect 14766 4080 14812 4092
rect 14766 3704 14772 4080
rect 14806 3704 14812 4080
rect 14766 3692 14812 3704
rect 14884 4080 14930 4092
rect 14884 3704 14890 4080
rect 14924 3704 14930 4080
rect 14884 3692 14930 3704
rect 15002 4080 15048 4092
rect 15002 3704 15008 4080
rect 15042 3704 15048 4080
rect 15328 4014 15428 4102
rect 15586 4155 15856 4183
rect 15586 4094 15620 4155
rect 15822 4094 15856 4155
rect 15940 4155 16210 4196
rect 15940 4094 15974 4155
rect 16176 4094 16210 4155
rect 16388 4168 16452 5191
rect 16538 4358 16602 5285
rect 16502 4256 16602 4358
rect 16502 4222 16552 4256
rect 16586 4222 16602 4256
rect 17188 4332 17292 4338
rect 17188 4260 17200 4332
rect 17280 4260 17292 4332
rect 17188 4254 17292 4260
rect 16502 4196 16602 4222
rect 17223 4198 17258 4254
rect 16388 4148 16602 4168
rect 16388 4114 16552 4148
rect 16586 4114 16602 4148
rect 16388 4104 16602 4114
rect 15462 4082 15508 4094
rect 15002 3692 15048 3704
rect 15462 3706 15468 4082
rect 15502 3706 15508 4082
rect 15462 3694 15508 3706
rect 15580 4082 15626 4094
rect 15580 3706 15586 4082
rect 15620 3706 15626 4082
rect 15580 3694 15626 3706
rect 15698 4082 15744 4094
rect 15698 3706 15704 4082
rect 15738 3706 15744 4082
rect 15698 3694 15744 3706
rect 15816 4082 15862 4094
rect 15816 3706 15822 4082
rect 15856 3706 15862 4082
rect 15816 3694 15862 3706
rect 15934 4082 15980 4094
rect 15934 3706 15940 4082
rect 15974 3706 15980 4082
rect 15934 3694 15980 3706
rect 16052 4082 16098 4094
rect 16052 3706 16058 4082
rect 16092 3706 16098 4082
rect 16052 3694 16098 3706
rect 16170 4082 16216 4094
rect 16170 3706 16176 4082
rect 16210 3706 16216 4082
rect 16502 4016 16602 4104
rect 16760 4157 17030 4185
rect 16760 4096 16794 4157
rect 16996 4096 17030 4157
rect 17114 4157 17384 4198
rect 17114 4096 17148 4157
rect 17350 4096 17384 4157
rect 17578 4168 17642 5377
rect 17670 4256 17770 5471
rect 17670 4222 17720 4256
rect 17754 4222 17770 4256
rect 18356 4332 18460 4338
rect 18356 4260 18368 4332
rect 18448 4260 18460 4332
rect 18356 4254 18460 4260
rect 17670 4196 17770 4222
rect 18391 4198 18426 4254
rect 17578 4148 17770 4168
rect 17578 4114 17720 4148
rect 17754 4114 17770 4148
rect 17578 4104 17770 4114
rect 16636 4084 16682 4096
rect 16170 3694 16216 3706
rect 16636 3708 16642 4084
rect 16676 3708 16682 4084
rect 16636 3696 16682 3708
rect 16754 4084 16800 4096
rect 16754 3708 16760 4084
rect 16794 3708 16800 4084
rect 16754 3696 16800 3708
rect 16872 4084 16918 4096
rect 16872 3708 16878 4084
rect 16912 3708 16918 4084
rect 16872 3696 16918 3708
rect 16990 4084 17036 4096
rect 16990 3708 16996 4084
rect 17030 3708 17036 4084
rect 16990 3696 17036 3708
rect 17108 4084 17154 4096
rect 17108 3708 17114 4084
rect 17148 3708 17154 4084
rect 17108 3696 17154 3708
rect 17226 4084 17272 4096
rect 17226 3708 17232 4084
rect 17266 3708 17272 4084
rect 17226 3696 17272 3708
rect 17344 4084 17390 4096
rect 17344 3708 17350 4084
rect 17384 3708 17390 4084
rect 17670 4016 17770 4104
rect 17928 4157 18198 4185
rect 17928 4094 17962 4157
rect 18164 4094 18198 4157
rect 18282 4157 18552 4198
rect 18282 4094 18316 4157
rect 18518 4094 18552 4157
rect 18741 4168 18805 5563
rect 18838 4256 18938 5657
rect 18838 4222 18888 4256
rect 18922 4222 18938 4256
rect 19524 4332 19628 4338
rect 19524 4260 19536 4332
rect 19616 4260 19628 4332
rect 19524 4254 19628 4260
rect 18838 4196 18938 4222
rect 19559 4198 19594 4254
rect 18741 4148 18938 4168
rect 18741 4114 18888 4148
rect 18922 4114 18938 4148
rect 18741 4104 18938 4114
rect 17804 4082 17850 4094
rect 17344 3696 17390 3708
rect 17804 3706 17810 4082
rect 17844 3706 17850 4082
rect 14300 3651 14334 3692
rect 14536 3651 14570 3692
rect 14300 3623 14570 3651
rect 14654 3652 14688 3692
rect 14890 3652 14924 3692
rect 14654 3623 14924 3652
rect 14300 3575 14334 3623
rect 14300 3545 14363 3575
rect 13840 3456 13949 3510
rect 13160 3417 13387 3453
rect 13160 3310 13195 3417
rect 13321 3383 13387 3417
rect 13321 3349 13337 3383
rect 13371 3349 13387 3383
rect 13321 3343 13387 3349
rect 13562 3310 13595 3314
rect 13798 3310 13831 3314
rect 13915 3310 13949 3456
rect 14328 3453 14363 3545
rect 15008 3510 15042 3692
rect 15468 3651 15502 3694
rect 15704 3651 15738 3694
rect 15468 3623 15738 3651
rect 15822 3652 15856 3694
rect 16058 3652 16092 3694
rect 15822 3623 16092 3652
rect 15468 3575 15502 3623
rect 15468 3545 15531 3575
rect 15008 3456 15117 3510
rect 14328 3417 14555 3453
rect 14328 3310 14363 3417
rect 14489 3383 14555 3417
rect 14489 3349 14505 3383
rect 14539 3349 14555 3383
rect 14489 3343 14555 3349
rect 14730 3310 14763 3314
rect 14966 3310 14999 3314
rect 15083 3310 15117 3456
rect 15496 3453 15531 3545
rect 16176 3510 16210 3694
rect 16642 3653 16676 3696
rect 16878 3653 16912 3696
rect 16642 3625 16912 3653
rect 16996 3654 17030 3696
rect 17232 3654 17266 3696
rect 16996 3625 17266 3654
rect 16642 3577 16676 3625
rect 16642 3547 16705 3577
rect 16176 3456 16285 3510
rect 15496 3417 15723 3453
rect 15496 3310 15531 3417
rect 15657 3383 15723 3417
rect 15657 3349 15673 3383
rect 15707 3349 15723 3383
rect 15657 3343 15723 3349
rect 15898 3310 15931 3314
rect 16134 3310 16167 3314
rect 16251 3310 16285 3456
rect 16670 3455 16705 3547
rect 17350 3512 17384 3696
rect 17804 3694 17850 3706
rect 17922 4082 17968 4094
rect 17922 3706 17928 4082
rect 17962 3706 17968 4082
rect 17922 3694 17968 3706
rect 18040 4082 18086 4094
rect 18040 3706 18046 4082
rect 18080 3706 18086 4082
rect 18040 3694 18086 3706
rect 18158 4082 18204 4094
rect 18158 3706 18164 4082
rect 18198 3706 18204 4082
rect 18158 3694 18204 3706
rect 18276 4082 18322 4094
rect 18276 3706 18282 4082
rect 18316 3706 18322 4082
rect 18276 3694 18322 3706
rect 18394 4082 18440 4094
rect 18394 3706 18400 4082
rect 18434 3706 18440 4082
rect 18394 3694 18440 3706
rect 18512 4082 18558 4094
rect 18512 3706 18518 4082
rect 18552 3706 18558 4082
rect 18838 4016 18938 4104
rect 19096 4157 19366 4185
rect 19096 4096 19130 4157
rect 19332 4096 19366 4157
rect 19450 4157 19720 4198
rect 19450 4096 19484 4157
rect 19686 4096 19720 4157
rect 19904 4169 19968 5749
rect 20006 4256 20106 5843
rect 20006 4222 20056 4256
rect 20090 4222 20106 4256
rect 20692 4332 20796 4338
rect 20692 4260 20704 4332
rect 20784 4260 20796 4332
rect 20692 4254 20796 4260
rect 20006 4197 20106 4222
rect 20727 4198 20762 4254
rect 19904 4148 20106 4169
rect 19904 4114 20056 4148
rect 20090 4114 20106 4148
rect 19904 4097 20106 4114
rect 20264 4157 20534 4185
rect 18972 4084 19018 4096
rect 18512 3694 18558 3706
rect 18972 3708 18978 4084
rect 19012 3708 19018 4084
rect 18972 3696 19018 3708
rect 19090 4084 19136 4096
rect 19090 3708 19096 4084
rect 19130 3708 19136 4084
rect 19090 3696 19136 3708
rect 19208 4084 19254 4096
rect 19208 3708 19214 4084
rect 19248 3708 19254 4084
rect 19208 3696 19254 3708
rect 19326 4084 19372 4096
rect 19326 3708 19332 4084
rect 19366 3708 19372 4084
rect 19326 3696 19372 3708
rect 19444 4084 19490 4096
rect 19444 3708 19450 4084
rect 19484 3708 19490 4084
rect 19444 3696 19490 3708
rect 19562 4084 19608 4096
rect 19562 3708 19568 4084
rect 19602 3708 19608 4084
rect 19562 3696 19608 3708
rect 19680 4084 19726 4096
rect 20264 4094 20298 4157
rect 20500 4094 20534 4157
rect 20618 4157 20888 4198
rect 20618 4094 20652 4157
rect 20854 4094 20888 4157
rect 19680 3708 19686 4084
rect 19720 3708 19726 4084
rect 19680 3696 19726 3708
rect 20140 4082 20186 4094
rect 20140 3706 20146 4082
rect 20180 3706 20186 4082
rect 17810 3653 17844 3694
rect 18046 3653 18080 3694
rect 17810 3625 18080 3653
rect 18164 3654 18198 3694
rect 18400 3654 18434 3694
rect 18164 3625 18434 3654
rect 17810 3577 17844 3625
rect 17810 3547 17873 3577
rect 17350 3458 17459 3512
rect 16670 3419 16897 3455
rect 16670 3310 16705 3419
rect 16831 3385 16897 3419
rect 16831 3351 16847 3385
rect 16881 3351 16897 3385
rect 16831 3345 16897 3351
rect 12222 3120 12228 3296
rect 12262 3243 12268 3296
rect 12388 3292 12434 3304
rect 12388 3243 12394 3292
rect 12262 3155 12394 3243
rect 12262 3120 12268 3155
rect 12222 3108 12268 3120
rect 12388 3116 12394 3155
rect 12428 3116 12434 3292
rect 11874 3071 11908 3108
rect 12110 3071 12144 3108
rect 12388 3104 12434 3116
rect 12506 3292 12552 3304
rect 12506 3116 12512 3292
rect 12546 3116 12552 3292
rect 12506 3104 12552 3116
rect 12624 3292 12670 3304
rect 12624 3116 12630 3292
rect 12664 3116 12670 3292
rect 12624 3104 12670 3116
rect 12742 3292 12788 3304
rect 12742 3116 12748 3292
rect 12782 3116 12788 3292
rect 12742 3104 12788 3116
rect 13036 3298 13082 3310
rect 13036 3122 13042 3298
rect 13076 3122 13082 3298
rect 13036 3110 13082 3122
rect 13154 3298 13200 3310
rect 13154 3122 13160 3298
rect 13194 3122 13200 3298
rect 13154 3110 13200 3122
rect 13272 3298 13318 3310
rect 13272 3122 13278 3298
rect 13312 3122 13318 3298
rect 13272 3110 13318 3122
rect 13390 3298 13436 3310
rect 13390 3122 13396 3298
rect 13430 3243 13436 3298
rect 13555 3298 13601 3310
rect 13555 3243 13561 3298
rect 13430 3155 13561 3243
rect 13430 3122 13436 3155
rect 13390 3110 13436 3122
rect 13555 3122 13561 3155
rect 13595 3122 13601 3298
rect 13555 3110 13601 3122
rect 13673 3298 13719 3310
rect 13673 3122 13679 3298
rect 13713 3122 13719 3298
rect 13673 3110 13719 3122
rect 13791 3298 13837 3310
rect 13791 3122 13797 3298
rect 13831 3122 13837 3298
rect 13791 3110 13837 3122
rect 13909 3298 13955 3310
rect 13909 3122 13915 3298
rect 13949 3122 13955 3298
rect 13909 3110 13955 3122
rect 14204 3298 14250 3310
rect 14204 3122 14210 3298
rect 14244 3122 14250 3298
rect 14204 3110 14250 3122
rect 14322 3298 14368 3310
rect 14322 3122 14328 3298
rect 14362 3122 14368 3298
rect 14322 3110 14368 3122
rect 14440 3298 14486 3310
rect 14440 3122 14446 3298
rect 14480 3122 14486 3298
rect 14440 3110 14486 3122
rect 14558 3298 14604 3310
rect 14558 3122 14564 3298
rect 14598 3243 14604 3298
rect 14723 3298 14769 3310
rect 14723 3243 14729 3298
rect 14598 3155 14729 3243
rect 14598 3122 14604 3155
rect 14558 3110 14604 3122
rect 14723 3122 14729 3155
rect 14763 3122 14769 3298
rect 14723 3110 14769 3122
rect 14841 3298 14887 3310
rect 14841 3122 14847 3298
rect 14881 3122 14887 3298
rect 14841 3110 14887 3122
rect 14959 3298 15005 3310
rect 14959 3122 14965 3298
rect 14999 3122 15005 3298
rect 14959 3110 15005 3122
rect 15077 3298 15123 3310
rect 15077 3122 15083 3298
rect 15117 3122 15123 3298
rect 15077 3110 15123 3122
rect 15372 3298 15418 3310
rect 15372 3122 15378 3298
rect 15412 3122 15418 3298
rect 15372 3110 15418 3122
rect 15490 3298 15536 3310
rect 15490 3122 15496 3298
rect 15530 3122 15536 3298
rect 15490 3110 15536 3122
rect 15608 3298 15654 3310
rect 15608 3122 15614 3298
rect 15648 3122 15654 3298
rect 15608 3110 15654 3122
rect 15726 3298 15772 3310
rect 15726 3122 15732 3298
rect 15766 3243 15772 3298
rect 15892 3298 15938 3310
rect 15892 3243 15898 3298
rect 15766 3155 15898 3243
rect 15766 3122 15772 3155
rect 15726 3110 15772 3122
rect 15892 3122 15898 3155
rect 15932 3122 15938 3298
rect 15892 3110 15938 3122
rect 16010 3298 16056 3310
rect 16010 3122 16016 3298
rect 16050 3122 16056 3298
rect 16010 3110 16056 3122
rect 16128 3298 16174 3310
rect 16128 3122 16134 3298
rect 16168 3122 16174 3298
rect 16128 3110 16174 3122
rect 16246 3298 16292 3310
rect 16246 3122 16252 3298
rect 16286 3122 16292 3298
rect 16246 3110 16292 3122
rect 16546 3298 16592 3310
rect 16546 3122 16552 3298
rect 16586 3122 16592 3298
rect 16546 3110 16592 3122
rect 16664 3298 16710 3310
rect 16664 3122 16670 3298
rect 16704 3122 16710 3298
rect 16664 3110 16710 3122
rect 16782 3298 16828 3310
rect 16782 3122 16788 3298
rect 16822 3122 16828 3298
rect 16782 3110 16828 3122
rect 16900 3298 16946 3310
rect 17072 3306 17105 3310
rect 17308 3306 17341 3310
rect 17425 3306 17459 3458
rect 17838 3455 17873 3547
rect 18518 3512 18552 3694
rect 18978 3653 19012 3696
rect 19214 3653 19248 3696
rect 18978 3625 19248 3653
rect 19332 3654 19366 3696
rect 19568 3654 19602 3696
rect 19332 3625 19602 3654
rect 18978 3577 19012 3625
rect 18978 3547 19041 3577
rect 18518 3458 18627 3512
rect 17838 3419 18065 3455
rect 17838 3310 17873 3419
rect 17999 3385 18065 3419
rect 17999 3351 18015 3385
rect 18049 3351 18065 3385
rect 17999 3345 18065 3351
rect 16900 3122 16906 3298
rect 16940 3245 16946 3298
rect 17064 3294 17110 3306
rect 17064 3245 17070 3294
rect 16940 3157 17070 3245
rect 16940 3122 16946 3157
rect 16900 3110 16946 3122
rect 17064 3118 17070 3157
rect 17104 3118 17110 3294
rect 11874 3032 12144 3071
rect 12511 3072 12544 3104
rect 12747 3072 12780 3104
rect 12511 3036 12780 3072
rect 13042 3071 13076 3110
rect 13278 3071 13312 3110
rect 13042 3032 13312 3071
rect 13679 3072 13712 3110
rect 13915 3072 13948 3110
rect 13679 3036 13948 3072
rect 14210 3071 14244 3110
rect 14446 3071 14480 3110
rect 14210 3032 14480 3071
rect 14847 3072 14880 3110
rect 15083 3072 15116 3110
rect 14847 3036 15116 3072
rect 15378 3071 15412 3110
rect 15614 3071 15648 3110
rect 15378 3032 15648 3071
rect 16015 3072 16048 3110
rect 16251 3072 16284 3110
rect 16015 3036 16284 3072
rect 16552 3073 16586 3110
rect 16788 3073 16822 3110
rect 17064 3106 17110 3118
rect 17182 3294 17228 3306
rect 17182 3118 17188 3294
rect 17222 3118 17228 3294
rect 17182 3106 17228 3118
rect 17300 3294 17346 3306
rect 17300 3118 17306 3294
rect 17340 3118 17346 3294
rect 17300 3106 17346 3118
rect 17418 3294 17464 3306
rect 17418 3118 17424 3294
rect 17458 3118 17464 3294
rect 17418 3106 17464 3118
rect 17714 3298 17760 3310
rect 17714 3122 17720 3298
rect 17754 3122 17760 3298
rect 17714 3110 17760 3122
rect 17832 3298 17878 3310
rect 17832 3122 17838 3298
rect 17872 3122 17878 3298
rect 17832 3110 17878 3122
rect 17950 3298 17996 3310
rect 17950 3122 17956 3298
rect 17990 3122 17996 3298
rect 17950 3110 17996 3122
rect 18068 3298 18114 3310
rect 18240 3305 18273 3309
rect 18476 3305 18509 3310
rect 18593 3305 18627 3458
rect 19006 3455 19041 3547
rect 19686 3512 19720 3696
rect 20140 3694 20186 3706
rect 20258 4082 20304 4094
rect 20258 3706 20264 4082
rect 20298 3706 20304 4082
rect 20258 3694 20304 3706
rect 20376 4082 20422 4094
rect 20376 3706 20382 4082
rect 20416 3706 20422 4082
rect 20376 3694 20422 3706
rect 20494 4082 20540 4094
rect 20494 3706 20500 4082
rect 20534 3706 20540 4082
rect 20494 3694 20540 3706
rect 20612 4082 20658 4094
rect 20612 3706 20618 4082
rect 20652 3706 20658 4082
rect 20612 3694 20658 3706
rect 20730 4082 20776 4094
rect 20730 3706 20736 4082
rect 20770 3706 20776 4082
rect 20730 3694 20776 3706
rect 20848 4082 20894 4094
rect 20848 3706 20854 4082
rect 20888 3706 20894 4082
rect 20848 3694 20894 3706
rect 20146 3653 20180 3694
rect 20382 3653 20416 3694
rect 20146 3625 20416 3653
rect 20500 3654 20534 3694
rect 20736 3654 20770 3694
rect 20500 3625 20770 3654
rect 20146 3577 20180 3625
rect 20146 3547 20209 3577
rect 19686 3458 19795 3512
rect 19006 3419 19233 3455
rect 19006 3312 19041 3419
rect 19167 3385 19233 3419
rect 19167 3351 19183 3385
rect 19217 3351 19233 3385
rect 19167 3345 19233 3351
rect 18068 3122 18074 3298
rect 18108 3245 18114 3298
rect 18233 3293 18279 3305
rect 18233 3245 18239 3293
rect 18108 3157 18239 3245
rect 18108 3122 18114 3157
rect 18068 3110 18114 3122
rect 18233 3117 18239 3157
rect 18273 3117 18279 3293
rect 16552 3034 16822 3073
rect 17189 3074 17222 3106
rect 17425 3074 17458 3106
rect 17189 3038 17458 3074
rect 17720 3073 17754 3110
rect 17956 3073 17990 3110
rect 18233 3105 18279 3117
rect 18351 3293 18397 3305
rect 18351 3117 18357 3293
rect 18391 3117 18397 3293
rect 18351 3105 18397 3117
rect 18469 3293 18515 3305
rect 18469 3117 18475 3293
rect 18509 3117 18515 3293
rect 18469 3105 18515 3117
rect 18587 3293 18633 3305
rect 18587 3117 18593 3293
rect 18627 3117 18633 3293
rect 18587 3105 18633 3117
rect 18882 3300 18928 3312
rect 18882 3124 18888 3300
rect 18922 3124 18928 3300
rect 18882 3112 18928 3124
rect 19000 3300 19046 3312
rect 19000 3124 19006 3300
rect 19040 3124 19046 3300
rect 19000 3112 19046 3124
rect 19118 3300 19164 3312
rect 19118 3124 19124 3300
rect 19158 3124 19164 3300
rect 19118 3112 19164 3124
rect 19236 3300 19282 3312
rect 19408 3305 19441 3309
rect 19644 3305 19677 3309
rect 19761 3305 19795 3458
rect 20174 3455 20209 3547
rect 20854 3512 20888 3694
rect 20854 3501 20963 3512
rect 20855 3458 20963 3501
rect 20174 3419 20401 3455
rect 20174 3312 20209 3419
rect 20335 3385 20401 3419
rect 20335 3351 20351 3385
rect 20385 3351 20401 3385
rect 20335 3345 20401 3351
rect 19236 3124 19242 3300
rect 19276 3245 19282 3300
rect 19401 3293 19447 3305
rect 19401 3245 19407 3293
rect 19276 3157 19407 3245
rect 19276 3124 19282 3157
rect 19236 3112 19282 3124
rect 19401 3117 19407 3157
rect 19441 3117 19447 3293
rect 17720 3034 17990 3073
rect 18357 3074 18390 3105
rect 18593 3074 18626 3105
rect 18357 3038 18626 3074
rect 18888 3073 18922 3112
rect 19124 3073 19158 3112
rect 19401 3105 19447 3117
rect 19519 3293 19565 3305
rect 19519 3117 19525 3293
rect 19559 3117 19565 3293
rect 19519 3105 19565 3117
rect 19637 3293 19683 3305
rect 19637 3117 19643 3293
rect 19677 3117 19683 3293
rect 19637 3105 19683 3117
rect 19755 3293 19801 3305
rect 19755 3117 19761 3293
rect 19795 3117 19801 3293
rect 19755 3105 19801 3117
rect 20050 3300 20096 3312
rect 20050 3124 20056 3300
rect 20090 3124 20096 3300
rect 20050 3112 20096 3124
rect 20168 3300 20214 3312
rect 20168 3124 20174 3300
rect 20208 3124 20214 3300
rect 20168 3112 20214 3124
rect 20286 3300 20332 3312
rect 20286 3124 20292 3300
rect 20326 3124 20332 3300
rect 20286 3112 20332 3124
rect 20404 3300 20450 3312
rect 20576 3306 20609 3310
rect 20812 3306 20845 3311
rect 20929 3306 20963 3458
rect 20404 3124 20410 3300
rect 20444 3245 20450 3300
rect 20569 3294 20615 3306
rect 20569 3245 20575 3294
rect 20444 3157 20575 3245
rect 20444 3124 20450 3157
rect 20404 3112 20450 3124
rect 20569 3118 20575 3157
rect 20609 3118 20615 3294
rect 18888 3034 19158 3073
rect 19525 3074 19558 3105
rect 19761 3074 19794 3105
rect 19525 3038 19794 3074
rect 20056 3073 20090 3112
rect 20292 3073 20326 3112
rect 20569 3106 20615 3118
rect 20687 3294 20733 3306
rect 20687 3118 20693 3294
rect 20727 3118 20733 3294
rect 20687 3106 20733 3118
rect 20805 3294 20851 3306
rect 20805 3118 20811 3294
rect 20845 3118 20851 3294
rect 20805 3106 20851 3118
rect 20923 3294 20969 3306
rect 20923 3118 20929 3294
rect 20963 3118 20969 3294
rect 20923 3106 20969 3118
rect 20056 3034 20326 3073
rect 20693 3074 20726 3106
rect 20929 3074 20962 3106
rect 20693 3038 20962 3074
rect 12074 3004 12108 3032
rect 13242 3004 13276 3032
rect 14410 3004 14444 3032
rect 15578 3004 15612 3032
rect 16752 3006 16786 3034
rect 17920 3006 17954 3034
rect 19088 3006 19122 3034
rect 20256 3006 20290 3034
rect 12052 2992 12130 3004
rect 12052 2922 12058 2992
rect 12124 2922 12130 2992
rect 12052 2910 12130 2922
rect 13220 2992 13298 3004
rect 13220 2922 13226 2992
rect 13292 2922 13298 2992
rect 13220 2910 13298 2922
rect 14388 2992 14466 3004
rect 14388 2922 14394 2992
rect 14460 2922 14466 2992
rect 14388 2910 14466 2922
rect 15556 2992 15634 3004
rect 15556 2922 15562 2992
rect 15628 2922 15634 2992
rect 15556 2910 15634 2922
rect 16730 2994 16808 3006
rect 16730 2924 16736 2994
rect 16802 2924 16808 2994
rect 16730 2912 16808 2924
rect 17898 2994 17976 3006
rect 17898 2924 17904 2994
rect 17970 2924 17976 2994
rect 17898 2912 17976 2924
rect 19066 2994 19144 3006
rect 19066 2924 19072 2994
rect 19138 2924 19144 2994
rect 19066 2912 19144 2924
rect 20234 2994 20312 3006
rect 20234 2924 20240 2994
rect 20306 2924 20312 2994
rect 20234 2912 20312 2924
rect 11501 2800 13001 2848
rect 12963 2795 13001 2800
rect 10053 2724 12931 2772
rect 9663 2695 9722 2722
rect 12884 2695 12931 2724
rect 12963 2723 16121 2795
rect 5587 2616 6532 2688
rect 7107 2620 9631 2693
rect 9663 2622 12856 2695
rect 12884 2622 16011 2695
rect 6453 2592 6532 2616
rect 9557 2593 9631 2620
rect 12770 2593 12856 2622
rect 15932 2593 16011 2622
rect 16049 2693 16121 2723
rect 16049 2621 19102 2693
rect 19030 2593 19102 2621
rect 4139 2520 6380 2588
rect 6453 2520 9524 2592
rect 9557 2520 12724 2593
rect 12770 2520 15870 2593
rect 15932 2521 19001 2593
rect 19030 2521 22145 2593
rect 4642 2324 4652 2384
rect 4732 2324 4742 2384
rect 4642 2284 4742 2324
rect 3845 2227 5648 2284
rect 3845 2140 3879 2227
rect 5020 2140 5054 2227
rect 3839 2128 3885 2140
rect 3839 1940 3845 2128
rect 3398 1928 3444 1940
rect 3398 1752 3404 1928
rect 3438 1752 3444 1928
rect 3398 1740 3444 1752
rect 3516 1928 3562 1940
rect 3516 1752 3522 1928
rect 3556 1752 3562 1928
rect 3516 1740 3562 1752
rect 3634 1928 3680 1940
rect 3634 1752 3640 1928
rect 3674 1752 3680 1928
rect 3634 1740 3680 1752
rect 3752 1928 3845 1940
rect 3752 1752 3758 1928
rect 3792 1752 3845 1928
rect 3879 1752 3885 2128
rect 3752 1740 3885 1752
rect 3957 2128 4003 2140
rect 3957 1752 3963 2128
rect 3997 1752 4003 2128
rect 3957 1740 4003 1752
rect 4075 2128 4121 2140
rect 4075 1752 4081 2128
rect 4115 1752 4121 2128
rect 4075 1740 4121 1752
rect 4193 2128 4239 2140
rect 4193 1752 4199 2128
rect 4233 1752 4239 2128
rect 4193 1740 4239 1752
rect 4306 2128 4352 2140
rect 4306 1752 4312 2128
rect 4346 1752 4352 2128
rect 4306 1740 4352 1752
rect 4424 2128 4470 2140
rect 4424 1752 4430 2128
rect 4464 1752 4470 2128
rect 4424 1740 4470 1752
rect 4542 2128 4588 2140
rect 4542 1752 4548 2128
rect 4582 1752 4588 2128
rect 4542 1740 4588 1752
rect 4660 2128 4706 2140
rect 4660 1752 4666 2128
rect 4700 1752 4706 2128
rect 4660 1740 4706 1752
rect 4778 2128 4824 2140
rect 4778 1752 4784 2128
rect 4818 1752 4824 2128
rect 4778 1740 4824 1752
rect 4896 2128 4942 2140
rect 4896 1752 4902 2128
rect 4936 1752 4942 2128
rect 4896 1740 4942 1752
rect 5014 2128 5060 2140
rect 5014 1752 5020 2128
rect 5054 1752 5060 2128
rect 5014 1740 5060 1752
rect 5133 2128 5179 2140
rect 5133 1752 5139 2128
rect 5173 1752 5179 2128
rect 5133 1740 5179 1752
rect 5251 2128 5297 2140
rect 5251 1752 5257 2128
rect 5291 1752 5297 2128
rect 5251 1740 5297 1752
rect 5369 2128 5415 2140
rect 5369 1752 5375 2128
rect 5409 1752 5415 2128
rect 5369 1740 5415 1752
rect 5487 2128 5533 2140
rect 5487 1752 5493 2128
rect 5527 1752 5533 2128
rect 5611 1940 5648 2227
rect 5487 1740 5533 1752
rect 5606 1928 5652 1940
rect 5606 1752 5612 1928
rect 5646 1752 5652 1928
rect 5606 1740 5652 1752
rect 5724 1928 5770 1940
rect 5724 1752 5730 1928
rect 5764 1752 5770 1928
rect 5724 1740 5770 1752
rect 5842 1928 5888 1940
rect 5842 1752 5848 1928
rect 5882 1752 5888 1928
rect 5842 1740 5888 1752
rect 5960 1928 6006 1940
rect 5960 1752 5966 1928
rect 6000 1752 6006 1928
rect 5960 1740 6006 1752
rect 3403 1554 3438 1740
rect 4312 1656 4346 1740
rect 5493 1656 5527 1740
rect 4312 1614 5527 1656
rect 5493 1594 5527 1614
rect 5493 1578 5850 1594
rect 3403 1537 4540 1554
rect 3403 1503 4490 1537
rect 4524 1503 4540 1537
rect 5493 1544 5800 1578
rect 5834 1544 5850 1578
rect 5493 1528 5850 1544
rect 3403 1487 4540 1503
rect 3144 1326 3320 1334
rect 3144 1258 3261 1326
rect 3318 1258 3328 1326
rect 3144 1250 3320 1258
rect 1316 1158 1408 1166
rect 1316 1093 1328 1158
rect 1396 1093 1408 1158
rect 1316 1081 1408 1093
rect 2822 978 2857 1240
rect 259 930 1631 977
rect 1953 931 2857 978
rect 1093 807 1127 930
rect 1565 917 1631 930
rect 1565 883 1581 917
rect 1615 883 1631 917
rect 1565 867 1631 883
rect 1954 807 1988 931
rect 1088 795 1134 807
rect 1088 619 1094 795
rect 1128 619 1134 795
rect 1088 607 1134 619
rect 1206 795 1326 807
rect 1206 619 1212 795
rect 1246 619 1286 795
rect 1206 607 1286 619
rect 1212 240 1246 607
rect 1280 419 1286 607
rect 1320 419 1326 795
rect 1280 407 1326 419
rect 1398 795 1444 807
rect 1398 419 1404 795
rect 1438 419 1444 795
rect 1398 407 1444 419
rect 1516 795 1562 807
rect 1516 419 1522 795
rect 1556 419 1562 795
rect 1516 407 1562 419
rect 1634 795 1680 807
rect 1634 419 1640 795
rect 1674 419 1680 795
rect 1634 407 1680 419
rect 1752 795 1876 807
rect 1752 419 1758 795
rect 1792 619 1836 795
rect 1870 619 1876 795
rect 1792 607 1876 619
rect 1948 795 1994 807
rect 1948 619 1954 795
rect 1988 619 1994 795
rect 1948 607 1994 619
rect 1792 419 1798 607
rect 1752 407 1798 419
rect 1522 334 1556 407
rect 1507 318 1573 334
rect 1507 284 1523 318
rect 1557 284 1573 318
rect 1507 268 1573 284
rect 1836 240 1870 607
rect 1212 188 1870 240
rect 1510 166 1602 188
rect 1510 114 1522 166
rect 1588 114 1602 166
rect 1510 110 1602 114
rect 2930 -14 3002 1240
rect 3250 1158 3320 1166
rect 3250 1090 3261 1158
rect 3318 1090 3328 1158
rect 3250 1082 3320 1090
rect 3403 977 3438 1487
rect 3493 1441 3585 1454
rect 3493 1378 3505 1441
rect 3576 1378 3585 1441
rect 3493 1369 3585 1378
rect 4578 1441 4670 1451
rect 4578 1379 4590 1441
rect 4660 1379 4670 1441
rect 4578 1366 4670 1379
rect 5966 1386 6001 1740
rect 4825 1324 4890 1327
rect 4825 1321 4894 1324
rect 4825 1261 4831 1321
rect 4890 1261 4900 1321
rect 4825 1257 4894 1261
rect 4825 1255 4890 1257
rect 5966 1240 6147 1386
rect 6293 1338 6380 2520
rect 7774 2328 7784 2388
rect 7864 2328 7874 2388
rect 7774 2288 7874 2328
rect 6977 2231 8780 2288
rect 6977 2144 7011 2231
rect 8152 2144 8186 2231
rect 6971 2132 7017 2144
rect 6971 1944 6977 2132
rect 6530 1932 6576 1944
rect 6530 1756 6536 1932
rect 6570 1756 6576 1932
rect 6530 1744 6576 1756
rect 6648 1932 6694 1944
rect 6648 1756 6654 1932
rect 6688 1756 6694 1932
rect 6648 1744 6694 1756
rect 6766 1932 6812 1944
rect 6766 1756 6772 1932
rect 6806 1756 6812 1932
rect 6766 1744 6812 1756
rect 6884 1932 6977 1944
rect 6884 1756 6890 1932
rect 6924 1756 6977 1932
rect 7011 1756 7017 2132
rect 6884 1744 7017 1756
rect 7089 2132 7135 2144
rect 7089 1756 7095 2132
rect 7129 1756 7135 2132
rect 7089 1744 7135 1756
rect 7207 2132 7253 2144
rect 7207 1756 7213 2132
rect 7247 1756 7253 2132
rect 7207 1744 7253 1756
rect 7325 2132 7371 2144
rect 7325 1756 7331 2132
rect 7365 1756 7371 2132
rect 7325 1744 7371 1756
rect 7438 2132 7484 2144
rect 7438 1756 7444 2132
rect 7478 1756 7484 2132
rect 7438 1744 7484 1756
rect 7556 2132 7602 2144
rect 7556 1756 7562 2132
rect 7596 1756 7602 2132
rect 7556 1744 7602 1756
rect 7674 2132 7720 2144
rect 7674 1756 7680 2132
rect 7714 1756 7720 2132
rect 7674 1744 7720 1756
rect 7792 2132 7838 2144
rect 7792 1756 7798 2132
rect 7832 1756 7838 2132
rect 7792 1744 7838 1756
rect 7910 2132 7956 2144
rect 7910 1756 7916 2132
rect 7950 1756 7956 2132
rect 7910 1744 7956 1756
rect 8028 2132 8074 2144
rect 8028 1756 8034 2132
rect 8068 1756 8074 2132
rect 8028 1744 8074 1756
rect 8146 2132 8192 2144
rect 8146 1756 8152 2132
rect 8186 1756 8192 2132
rect 8146 1744 8192 1756
rect 8265 2132 8311 2144
rect 8265 1756 8271 2132
rect 8305 1756 8311 2132
rect 8265 1744 8311 1756
rect 8383 2132 8429 2144
rect 8383 1756 8389 2132
rect 8423 1756 8429 2132
rect 8383 1744 8429 1756
rect 8501 2132 8547 2144
rect 8501 1756 8507 2132
rect 8541 1756 8547 2132
rect 8501 1744 8547 1756
rect 8619 2132 8665 2144
rect 8619 1756 8625 2132
rect 8659 1756 8665 2132
rect 8743 1944 8780 2231
rect 8619 1744 8665 1756
rect 8738 1932 8784 1944
rect 8738 1756 8744 1932
rect 8778 1756 8784 1932
rect 8738 1744 8784 1756
rect 8856 1932 8902 1944
rect 8856 1756 8862 1932
rect 8896 1756 8902 1932
rect 8856 1744 8902 1756
rect 8974 1932 9020 1944
rect 8974 1756 8980 1932
rect 9014 1756 9020 1932
rect 8974 1744 9020 1756
rect 9092 1932 9138 1944
rect 9092 1756 9098 1932
rect 9132 1756 9138 1932
rect 9092 1744 9138 1756
rect 6535 1558 6570 1744
rect 7444 1660 7478 1744
rect 8625 1660 8659 1744
rect 7444 1618 8659 1660
rect 8625 1598 8659 1618
rect 8625 1582 8982 1598
rect 6535 1541 7672 1558
rect 6535 1507 7622 1541
rect 7656 1507 7672 1541
rect 8625 1548 8932 1582
rect 8966 1548 8982 1582
rect 8625 1532 8982 1548
rect 6535 1491 7672 1507
rect 6293 1330 6452 1338
rect 6293 1262 6393 1330
rect 6450 1262 6460 1330
rect 6293 1254 6452 1262
rect 4460 1158 4552 1166
rect 4460 1093 4472 1158
rect 4540 1093 4552 1158
rect 4460 1081 4552 1093
rect 5966 978 6001 1240
rect 3403 930 4775 977
rect 5097 931 6001 978
rect 4237 807 4271 930
rect 4709 917 4775 930
rect 4709 883 4725 917
rect 4759 883 4775 917
rect 4709 867 4775 883
rect 5098 807 5132 931
rect 4232 795 4278 807
rect 4232 619 4238 795
rect 4272 619 4278 795
rect 4232 607 4278 619
rect 4350 795 4470 807
rect 4350 619 4356 795
rect 4390 619 4430 795
rect 4350 607 4430 619
rect 4356 240 4390 607
rect 4424 419 4430 607
rect 4464 419 4470 795
rect 4424 407 4470 419
rect 4542 795 4588 807
rect 4542 419 4548 795
rect 4582 419 4588 795
rect 4542 407 4588 419
rect 4660 795 4706 807
rect 4660 419 4666 795
rect 4700 419 4706 795
rect 4660 407 4706 419
rect 4778 795 4824 807
rect 4778 419 4784 795
rect 4818 419 4824 795
rect 4778 407 4824 419
rect 4896 795 5020 807
rect 4896 419 4902 795
rect 4936 619 4980 795
rect 5014 619 5020 795
rect 4936 607 5020 619
rect 5092 795 5138 807
rect 5092 619 5098 795
rect 5132 619 5138 795
rect 5092 607 5138 619
rect 4936 419 4942 607
rect 4896 407 4942 419
rect 4666 334 4700 407
rect 4651 318 4717 334
rect 4651 284 4667 318
rect 4701 284 4717 318
rect 4651 268 4717 284
rect 4980 240 5014 607
rect 4356 188 5014 240
rect 4654 166 4746 188
rect 4654 114 4666 166
rect 4732 114 4746 166
rect 4654 110 4746 114
rect 6073 -13 6145 1240
rect 6380 1162 6452 1170
rect 6380 1094 6393 1162
rect 6450 1094 6460 1162
rect 6380 1086 6452 1094
rect 6535 981 6570 1491
rect 6625 1445 6717 1458
rect 6625 1382 6637 1445
rect 6708 1382 6717 1445
rect 6625 1373 6717 1382
rect 7710 1445 7802 1455
rect 7710 1383 7722 1445
rect 7792 1383 7802 1445
rect 7710 1370 7802 1383
rect 9098 1390 9133 1744
rect 7957 1328 8022 1331
rect 7957 1325 8026 1328
rect 7957 1265 7963 1325
rect 8022 1265 8032 1325
rect 7957 1261 8026 1265
rect 7957 1259 8022 1261
rect 9098 1244 9278 1390
rect 9437 1338 9524 2520
rect 10918 2328 10928 2388
rect 11008 2328 11018 2388
rect 10918 2288 11018 2328
rect 10121 2231 11924 2288
rect 10121 2144 10155 2231
rect 11296 2144 11330 2231
rect 10115 2132 10161 2144
rect 10115 1944 10121 2132
rect 9674 1932 9720 1944
rect 9674 1756 9680 1932
rect 9714 1756 9720 1932
rect 9674 1744 9720 1756
rect 9792 1932 9838 1944
rect 9792 1756 9798 1932
rect 9832 1756 9838 1932
rect 9792 1744 9838 1756
rect 9910 1932 9956 1944
rect 9910 1756 9916 1932
rect 9950 1756 9956 1932
rect 9910 1744 9956 1756
rect 10028 1932 10121 1944
rect 10028 1756 10034 1932
rect 10068 1756 10121 1932
rect 10155 1756 10161 2132
rect 10028 1744 10161 1756
rect 10233 2132 10279 2144
rect 10233 1756 10239 2132
rect 10273 1756 10279 2132
rect 10233 1744 10279 1756
rect 10351 2132 10397 2144
rect 10351 1756 10357 2132
rect 10391 1756 10397 2132
rect 10351 1744 10397 1756
rect 10469 2132 10515 2144
rect 10469 1756 10475 2132
rect 10509 1756 10515 2132
rect 10469 1744 10515 1756
rect 10582 2132 10628 2144
rect 10582 1756 10588 2132
rect 10622 1756 10628 2132
rect 10582 1744 10628 1756
rect 10700 2132 10746 2144
rect 10700 1756 10706 2132
rect 10740 1756 10746 2132
rect 10700 1744 10746 1756
rect 10818 2132 10864 2144
rect 10818 1756 10824 2132
rect 10858 1756 10864 2132
rect 10818 1744 10864 1756
rect 10936 2132 10982 2144
rect 10936 1756 10942 2132
rect 10976 1756 10982 2132
rect 10936 1744 10982 1756
rect 11054 2132 11100 2144
rect 11054 1756 11060 2132
rect 11094 1756 11100 2132
rect 11054 1744 11100 1756
rect 11172 2132 11218 2144
rect 11172 1756 11178 2132
rect 11212 1756 11218 2132
rect 11172 1744 11218 1756
rect 11290 2132 11336 2144
rect 11290 1756 11296 2132
rect 11330 1756 11336 2132
rect 11290 1744 11336 1756
rect 11409 2132 11455 2144
rect 11409 1756 11415 2132
rect 11449 1756 11455 2132
rect 11409 1744 11455 1756
rect 11527 2132 11573 2144
rect 11527 1756 11533 2132
rect 11567 1756 11573 2132
rect 11527 1744 11573 1756
rect 11645 2132 11691 2144
rect 11645 1756 11651 2132
rect 11685 1756 11691 2132
rect 11645 1744 11691 1756
rect 11763 2132 11809 2144
rect 11763 1756 11769 2132
rect 11803 1756 11809 2132
rect 11887 1944 11924 2231
rect 11763 1744 11809 1756
rect 11882 1932 11928 1944
rect 11882 1756 11888 1932
rect 11922 1756 11928 1932
rect 11882 1744 11928 1756
rect 12000 1932 12046 1944
rect 12000 1756 12006 1932
rect 12040 1756 12046 1932
rect 12000 1744 12046 1756
rect 12118 1932 12164 1944
rect 12118 1756 12124 1932
rect 12158 1756 12164 1932
rect 12118 1744 12164 1756
rect 12236 1932 12282 1944
rect 12236 1756 12242 1932
rect 12276 1756 12282 1932
rect 12236 1744 12282 1756
rect 9679 1558 9714 1744
rect 10588 1660 10622 1744
rect 11769 1660 11803 1744
rect 10588 1618 11803 1660
rect 11769 1598 11803 1618
rect 11769 1582 12126 1598
rect 9679 1541 10816 1558
rect 9679 1507 10766 1541
rect 10800 1507 10816 1541
rect 11769 1548 12076 1582
rect 12110 1548 12126 1582
rect 11769 1532 12126 1548
rect 9679 1491 10816 1507
rect 9437 1330 9596 1338
rect 9437 1262 9537 1330
rect 9594 1262 9604 1330
rect 9437 1254 9596 1262
rect 7592 1162 7684 1170
rect 7592 1097 7604 1162
rect 7672 1097 7684 1162
rect 7592 1085 7684 1097
rect 9098 982 9133 1244
rect 6535 934 7907 981
rect 8229 935 9133 982
rect 7369 811 7403 934
rect 7841 921 7907 934
rect 7841 887 7857 921
rect 7891 887 7907 921
rect 7841 871 7907 887
rect 8230 811 8264 935
rect 7364 799 7410 811
rect 7364 623 7370 799
rect 7404 623 7410 799
rect 7364 611 7410 623
rect 7482 799 7602 811
rect 7482 623 7488 799
rect 7522 623 7562 799
rect 7482 611 7562 623
rect 7488 244 7522 611
rect 7556 423 7562 611
rect 7596 423 7602 799
rect 7556 411 7602 423
rect 7674 799 7720 811
rect 7674 423 7680 799
rect 7714 423 7720 799
rect 7674 411 7720 423
rect 7792 799 7838 811
rect 7792 423 7798 799
rect 7832 423 7838 799
rect 7792 411 7838 423
rect 7910 799 7956 811
rect 7910 423 7916 799
rect 7950 423 7956 799
rect 7910 411 7956 423
rect 8028 799 8152 811
rect 8028 423 8034 799
rect 8068 623 8112 799
rect 8146 623 8152 799
rect 8068 611 8152 623
rect 8224 799 8270 811
rect 8224 623 8230 799
rect 8264 623 8270 799
rect 8224 611 8270 623
rect 8068 423 8074 611
rect 8028 411 8074 423
rect 7798 338 7832 411
rect 7783 322 7849 338
rect 7783 288 7799 322
rect 7833 288 7849 322
rect 7783 272 7849 288
rect 8112 244 8146 611
rect 7488 192 8146 244
rect 7786 170 7878 192
rect 7786 118 7798 170
rect 7864 118 7878 170
rect 7786 114 7878 118
rect 9206 -13 9278 1244
rect 9679 981 9714 1491
rect 9769 1445 9861 1458
rect 9769 1382 9781 1445
rect 9852 1382 9861 1445
rect 9769 1373 9861 1382
rect 10854 1445 10946 1455
rect 10854 1383 10866 1445
rect 10936 1383 10946 1445
rect 10854 1370 10946 1383
rect 12242 1390 12277 1744
rect 11101 1328 11166 1331
rect 11101 1325 11170 1328
rect 11101 1265 11107 1325
rect 11166 1265 11176 1325
rect 11101 1261 11170 1265
rect 11101 1259 11166 1261
rect 12242 1244 12418 1390
rect 12637 1334 12724 2520
rect 14120 2324 14130 2384
rect 14210 2324 14220 2384
rect 14120 2284 14220 2324
rect 13323 2227 15126 2284
rect 13323 2140 13357 2227
rect 14498 2140 14532 2227
rect 13317 2128 13363 2140
rect 13317 1940 13323 2128
rect 12876 1928 12922 1940
rect 12876 1752 12882 1928
rect 12916 1752 12922 1928
rect 12876 1740 12922 1752
rect 12994 1928 13040 1940
rect 12994 1752 13000 1928
rect 13034 1752 13040 1928
rect 12994 1740 13040 1752
rect 13112 1928 13158 1940
rect 13112 1752 13118 1928
rect 13152 1752 13158 1928
rect 13112 1740 13158 1752
rect 13230 1928 13323 1940
rect 13230 1752 13236 1928
rect 13270 1752 13323 1928
rect 13357 1752 13363 2128
rect 13230 1740 13363 1752
rect 13435 2128 13481 2140
rect 13435 1752 13441 2128
rect 13475 1752 13481 2128
rect 13435 1740 13481 1752
rect 13553 2128 13599 2140
rect 13553 1752 13559 2128
rect 13593 1752 13599 2128
rect 13553 1740 13599 1752
rect 13671 2128 13717 2140
rect 13671 1752 13677 2128
rect 13711 1752 13717 2128
rect 13671 1740 13717 1752
rect 13784 2128 13830 2140
rect 13784 1752 13790 2128
rect 13824 1752 13830 2128
rect 13784 1740 13830 1752
rect 13902 2128 13948 2140
rect 13902 1752 13908 2128
rect 13942 1752 13948 2128
rect 13902 1740 13948 1752
rect 14020 2128 14066 2140
rect 14020 1752 14026 2128
rect 14060 1752 14066 2128
rect 14020 1740 14066 1752
rect 14138 2128 14184 2140
rect 14138 1752 14144 2128
rect 14178 1752 14184 2128
rect 14138 1740 14184 1752
rect 14256 2128 14302 2140
rect 14256 1752 14262 2128
rect 14296 1752 14302 2128
rect 14256 1740 14302 1752
rect 14374 2128 14420 2140
rect 14374 1752 14380 2128
rect 14414 1752 14420 2128
rect 14374 1740 14420 1752
rect 14492 2128 14538 2140
rect 14492 1752 14498 2128
rect 14532 1752 14538 2128
rect 14492 1740 14538 1752
rect 14611 2128 14657 2140
rect 14611 1752 14617 2128
rect 14651 1752 14657 2128
rect 14611 1740 14657 1752
rect 14729 2128 14775 2140
rect 14729 1752 14735 2128
rect 14769 1752 14775 2128
rect 14729 1740 14775 1752
rect 14847 2128 14893 2140
rect 14847 1752 14853 2128
rect 14887 1752 14893 2128
rect 14847 1740 14893 1752
rect 14965 2128 15011 2140
rect 14965 1752 14971 2128
rect 15005 1752 15011 2128
rect 15089 1940 15126 2227
rect 14965 1740 15011 1752
rect 15084 1928 15130 1940
rect 15084 1752 15090 1928
rect 15124 1752 15130 1928
rect 15084 1740 15130 1752
rect 15202 1928 15248 1940
rect 15202 1752 15208 1928
rect 15242 1752 15248 1928
rect 15202 1740 15248 1752
rect 15320 1928 15366 1940
rect 15320 1752 15326 1928
rect 15360 1752 15366 1928
rect 15320 1740 15366 1752
rect 15438 1928 15484 1940
rect 15438 1752 15444 1928
rect 15478 1752 15484 1928
rect 15438 1740 15484 1752
rect 12881 1554 12916 1740
rect 13790 1656 13824 1740
rect 14971 1656 15005 1740
rect 13790 1614 15005 1656
rect 14971 1594 15005 1614
rect 14971 1578 15328 1594
rect 12881 1537 14018 1554
rect 12881 1503 13968 1537
rect 14002 1503 14018 1537
rect 14971 1544 15278 1578
rect 15312 1544 15328 1578
rect 14971 1528 15328 1544
rect 12881 1487 14018 1503
rect 12637 1326 12798 1334
rect 12637 1258 12739 1326
rect 12796 1258 12806 1326
rect 12637 1250 12798 1258
rect 12242 982 12277 1244
rect 9679 934 11051 981
rect 11373 935 12277 982
rect 10513 811 10547 934
rect 10985 921 11051 934
rect 10985 887 11001 921
rect 11035 887 11051 921
rect 10985 871 11051 887
rect 11374 811 11408 935
rect 10508 799 10554 811
rect 10508 623 10514 799
rect 10548 623 10554 799
rect 10508 611 10554 623
rect 10626 799 10746 811
rect 10626 623 10632 799
rect 10666 623 10706 799
rect 10626 611 10706 623
rect 10632 244 10666 611
rect 10700 423 10706 611
rect 10740 423 10746 799
rect 10700 411 10746 423
rect 10818 799 10864 811
rect 10818 423 10824 799
rect 10858 423 10864 799
rect 10818 411 10864 423
rect 10936 799 10982 811
rect 10936 423 10942 799
rect 10976 423 10982 799
rect 10936 411 10982 423
rect 11054 799 11100 811
rect 11054 423 11060 799
rect 11094 423 11100 799
rect 11054 411 11100 423
rect 11172 799 11296 811
rect 11172 423 11178 799
rect 11212 623 11256 799
rect 11290 623 11296 799
rect 11212 611 11296 623
rect 11368 799 11414 811
rect 11368 623 11374 799
rect 11408 623 11414 799
rect 11368 611 11414 623
rect 11212 423 11218 611
rect 11172 411 11218 423
rect 10942 338 10976 411
rect 10927 322 10993 338
rect 10927 288 10943 322
rect 10977 288 10993 322
rect 10927 272 10993 288
rect 11256 244 11290 611
rect 10632 192 11290 244
rect 10930 170 11022 192
rect 10930 118 10942 170
rect 11008 118 11022 170
rect 10930 114 11022 118
rect 12346 -10 12418 1244
rect 12881 977 12916 1487
rect 12971 1441 13063 1454
rect 12971 1378 12983 1441
rect 13054 1378 13063 1441
rect 12971 1369 13063 1378
rect 14056 1441 14148 1451
rect 14056 1379 14068 1441
rect 14138 1379 14148 1441
rect 14056 1366 14148 1379
rect 15444 1386 15479 1740
rect 14303 1324 14368 1327
rect 14303 1321 14372 1324
rect 14303 1261 14309 1321
rect 14368 1261 14378 1321
rect 14303 1257 14372 1261
rect 14303 1255 14368 1257
rect 15444 1240 15625 1386
rect 15783 1334 15870 2520
rect 17264 2324 17274 2384
rect 17354 2324 17364 2384
rect 17264 2284 17364 2324
rect 16467 2227 18270 2284
rect 16467 2140 16501 2227
rect 17642 2140 17676 2227
rect 16461 2128 16507 2140
rect 16461 1940 16467 2128
rect 16020 1928 16066 1940
rect 16020 1752 16026 1928
rect 16060 1752 16066 1928
rect 16020 1740 16066 1752
rect 16138 1928 16184 1940
rect 16138 1752 16144 1928
rect 16178 1752 16184 1928
rect 16138 1740 16184 1752
rect 16256 1928 16302 1940
rect 16256 1752 16262 1928
rect 16296 1752 16302 1928
rect 16256 1740 16302 1752
rect 16374 1928 16467 1940
rect 16374 1752 16380 1928
rect 16414 1752 16467 1928
rect 16501 1752 16507 2128
rect 16374 1740 16507 1752
rect 16579 2128 16625 2140
rect 16579 1752 16585 2128
rect 16619 1752 16625 2128
rect 16579 1740 16625 1752
rect 16697 2128 16743 2140
rect 16697 1752 16703 2128
rect 16737 1752 16743 2128
rect 16697 1740 16743 1752
rect 16815 2128 16861 2140
rect 16815 1752 16821 2128
rect 16855 1752 16861 2128
rect 16815 1740 16861 1752
rect 16928 2128 16974 2140
rect 16928 1752 16934 2128
rect 16968 1752 16974 2128
rect 16928 1740 16974 1752
rect 17046 2128 17092 2140
rect 17046 1752 17052 2128
rect 17086 1752 17092 2128
rect 17046 1740 17092 1752
rect 17164 2128 17210 2140
rect 17164 1752 17170 2128
rect 17204 1752 17210 2128
rect 17164 1740 17210 1752
rect 17282 2128 17328 2140
rect 17282 1752 17288 2128
rect 17322 1752 17328 2128
rect 17282 1740 17328 1752
rect 17400 2128 17446 2140
rect 17400 1752 17406 2128
rect 17440 1752 17446 2128
rect 17400 1740 17446 1752
rect 17518 2128 17564 2140
rect 17518 1752 17524 2128
rect 17558 1752 17564 2128
rect 17518 1740 17564 1752
rect 17636 2128 17682 2140
rect 17636 1752 17642 2128
rect 17676 1752 17682 2128
rect 17636 1740 17682 1752
rect 17755 2128 17801 2140
rect 17755 1752 17761 2128
rect 17795 1752 17801 2128
rect 17755 1740 17801 1752
rect 17873 2128 17919 2140
rect 17873 1752 17879 2128
rect 17913 1752 17919 2128
rect 17873 1740 17919 1752
rect 17991 2128 18037 2140
rect 17991 1752 17997 2128
rect 18031 1752 18037 2128
rect 17991 1740 18037 1752
rect 18109 2128 18155 2140
rect 18109 1752 18115 2128
rect 18149 1752 18155 2128
rect 18233 1940 18270 2227
rect 18109 1740 18155 1752
rect 18228 1928 18274 1940
rect 18228 1752 18234 1928
rect 18268 1752 18274 1928
rect 18228 1740 18274 1752
rect 18346 1928 18392 1940
rect 18346 1752 18352 1928
rect 18386 1752 18392 1928
rect 18346 1740 18392 1752
rect 18464 1928 18510 1940
rect 18464 1752 18470 1928
rect 18504 1752 18510 1928
rect 18464 1740 18510 1752
rect 18582 1928 18628 1940
rect 18582 1752 18588 1928
rect 18622 1752 18628 1928
rect 18582 1740 18628 1752
rect 16025 1554 16060 1740
rect 16934 1656 16968 1740
rect 18115 1656 18149 1740
rect 16934 1614 18149 1656
rect 18115 1594 18149 1614
rect 18115 1578 18472 1594
rect 16025 1537 17162 1554
rect 16025 1503 17112 1537
rect 17146 1503 17162 1537
rect 18115 1544 18422 1578
rect 18456 1544 18472 1578
rect 18115 1528 18472 1544
rect 16025 1487 17162 1503
rect 15783 1326 15942 1334
rect 15783 1258 15883 1326
rect 15940 1258 15950 1326
rect 15783 1250 15942 1258
rect 15444 978 15479 1240
rect 12881 930 14253 977
rect 14575 931 15479 978
rect 13715 807 13749 930
rect 14187 917 14253 930
rect 14187 883 14203 917
rect 14237 883 14253 917
rect 14187 867 14253 883
rect 14576 807 14610 931
rect 13710 795 13756 807
rect 13710 619 13716 795
rect 13750 619 13756 795
rect 13710 607 13756 619
rect 13828 795 13948 807
rect 13828 619 13834 795
rect 13868 619 13908 795
rect 13828 607 13908 619
rect 13834 240 13868 607
rect 13902 419 13908 607
rect 13942 419 13948 795
rect 13902 407 13948 419
rect 14020 795 14066 807
rect 14020 419 14026 795
rect 14060 419 14066 795
rect 14020 407 14066 419
rect 14138 795 14184 807
rect 14138 419 14144 795
rect 14178 419 14184 795
rect 14138 407 14184 419
rect 14256 795 14302 807
rect 14256 419 14262 795
rect 14296 419 14302 795
rect 14256 407 14302 419
rect 14374 795 14498 807
rect 14374 419 14380 795
rect 14414 619 14458 795
rect 14492 619 14498 795
rect 14414 607 14498 619
rect 14570 795 14616 807
rect 14570 619 14576 795
rect 14610 619 14616 795
rect 14570 607 14616 619
rect 14414 419 14420 607
rect 14374 407 14420 419
rect 14144 334 14178 407
rect 14129 318 14195 334
rect 14129 284 14145 318
rect 14179 284 14195 318
rect 14129 268 14195 284
rect 14458 240 14492 607
rect 13834 188 14492 240
rect 14132 166 14224 188
rect 14132 114 14144 166
rect 14210 114 14224 166
rect 14132 110 14224 114
rect 15538 -10 15625 1240
rect 15872 1158 15942 1166
rect 15872 1090 15883 1158
rect 15940 1090 15950 1158
rect 15872 1082 15942 1090
rect 16025 977 16060 1487
rect 16115 1441 16207 1454
rect 16115 1378 16127 1441
rect 16198 1378 16207 1441
rect 16115 1369 16207 1378
rect 17200 1441 17292 1451
rect 17200 1379 17212 1441
rect 17282 1379 17292 1441
rect 17200 1366 17292 1379
rect 18588 1386 18623 1740
rect 17447 1324 17512 1327
rect 17447 1321 17516 1324
rect 17447 1261 17453 1321
rect 17512 1261 17522 1321
rect 17447 1257 17516 1261
rect 17447 1255 17512 1257
rect 18588 1253 18769 1386
rect 18914 1338 19001 2521
rect 20396 2328 20406 2388
rect 20486 2328 20496 2388
rect 20396 2288 20496 2328
rect 19599 2231 21402 2288
rect 19599 2144 19633 2231
rect 20774 2144 20808 2231
rect 19593 2132 19639 2144
rect 19593 1944 19599 2132
rect 19152 1932 19198 1944
rect 19152 1756 19158 1932
rect 19192 1756 19198 1932
rect 19152 1744 19198 1756
rect 19270 1932 19316 1944
rect 19270 1756 19276 1932
rect 19310 1756 19316 1932
rect 19270 1744 19316 1756
rect 19388 1932 19434 1944
rect 19388 1756 19394 1932
rect 19428 1756 19434 1932
rect 19388 1744 19434 1756
rect 19506 1932 19599 1944
rect 19506 1756 19512 1932
rect 19546 1756 19599 1932
rect 19633 1756 19639 2132
rect 19506 1744 19639 1756
rect 19711 2132 19757 2144
rect 19711 1756 19717 2132
rect 19751 1756 19757 2132
rect 19711 1744 19757 1756
rect 19829 2132 19875 2144
rect 19829 1756 19835 2132
rect 19869 1756 19875 2132
rect 19829 1744 19875 1756
rect 19947 2132 19993 2144
rect 19947 1756 19953 2132
rect 19987 1756 19993 2132
rect 19947 1744 19993 1756
rect 20060 2132 20106 2144
rect 20060 1756 20066 2132
rect 20100 1756 20106 2132
rect 20060 1744 20106 1756
rect 20178 2132 20224 2144
rect 20178 1756 20184 2132
rect 20218 1756 20224 2132
rect 20178 1744 20224 1756
rect 20296 2132 20342 2144
rect 20296 1756 20302 2132
rect 20336 1756 20342 2132
rect 20296 1744 20342 1756
rect 20414 2132 20460 2144
rect 20414 1756 20420 2132
rect 20454 1756 20460 2132
rect 20414 1744 20460 1756
rect 20532 2132 20578 2144
rect 20532 1756 20538 2132
rect 20572 1756 20578 2132
rect 20532 1744 20578 1756
rect 20650 2132 20696 2144
rect 20650 1756 20656 2132
rect 20690 1756 20696 2132
rect 20650 1744 20696 1756
rect 20768 2132 20814 2144
rect 20768 1756 20774 2132
rect 20808 1756 20814 2132
rect 20768 1744 20814 1756
rect 20887 2132 20933 2144
rect 20887 1756 20893 2132
rect 20927 1756 20933 2132
rect 20887 1744 20933 1756
rect 21005 2132 21051 2144
rect 21005 1756 21011 2132
rect 21045 1756 21051 2132
rect 21005 1744 21051 1756
rect 21123 2132 21169 2144
rect 21123 1756 21129 2132
rect 21163 1756 21169 2132
rect 21123 1744 21169 1756
rect 21241 2132 21287 2144
rect 21241 1756 21247 2132
rect 21281 1756 21287 2132
rect 21365 1944 21402 2231
rect 21241 1744 21287 1756
rect 21360 1932 21406 1944
rect 21360 1756 21366 1932
rect 21400 1756 21406 1932
rect 21360 1744 21406 1756
rect 21478 1932 21524 1944
rect 21478 1756 21484 1932
rect 21518 1756 21524 1932
rect 21478 1744 21524 1756
rect 21596 1932 21642 1944
rect 21596 1756 21602 1932
rect 21636 1756 21642 1932
rect 21596 1744 21642 1756
rect 21714 1932 21760 1944
rect 21714 1756 21720 1932
rect 21754 1756 21760 1932
rect 21714 1744 21760 1756
rect 19157 1558 19192 1744
rect 20066 1660 20100 1744
rect 21247 1660 21281 1744
rect 20066 1618 21281 1660
rect 21247 1598 21281 1618
rect 21247 1582 21604 1598
rect 19157 1541 20294 1558
rect 19157 1507 20244 1541
rect 20278 1507 20294 1541
rect 21247 1548 21554 1582
rect 21588 1548 21604 1582
rect 21247 1532 21604 1548
rect 19157 1491 20294 1507
rect 18914 1330 19074 1338
rect 18914 1262 19015 1330
rect 19072 1262 19082 1330
rect 18914 1254 19074 1262
rect 18588 1240 18770 1253
rect 17082 1158 17174 1166
rect 17082 1093 17094 1158
rect 17162 1093 17174 1158
rect 17082 1081 17174 1093
rect 18588 978 18623 1240
rect 16025 930 17397 977
rect 17719 931 18623 978
rect 16859 807 16893 930
rect 17331 917 17397 930
rect 17331 883 17347 917
rect 17381 883 17397 917
rect 17331 867 17397 883
rect 17720 807 17754 931
rect 16854 795 16900 807
rect 16854 619 16860 795
rect 16894 619 16900 795
rect 16854 607 16900 619
rect 16972 795 17092 807
rect 16972 619 16978 795
rect 17012 619 17052 795
rect 16972 607 17052 619
rect 16978 240 17012 607
rect 17046 419 17052 607
rect 17086 419 17092 795
rect 17046 407 17092 419
rect 17164 795 17210 807
rect 17164 419 17170 795
rect 17204 419 17210 795
rect 17164 407 17210 419
rect 17282 795 17328 807
rect 17282 419 17288 795
rect 17322 419 17328 795
rect 17282 407 17328 419
rect 17400 795 17446 807
rect 17400 419 17406 795
rect 17440 419 17446 795
rect 17400 407 17446 419
rect 17518 795 17642 807
rect 17518 419 17524 795
rect 17558 619 17602 795
rect 17636 619 17642 795
rect 17558 607 17642 619
rect 17714 795 17760 807
rect 17714 619 17720 795
rect 17754 619 17760 795
rect 17714 607 17760 619
rect 17558 419 17564 607
rect 17518 407 17564 419
rect 17288 334 17322 407
rect 17273 318 17339 334
rect 17273 284 17289 318
rect 17323 284 17339 318
rect 17273 268 17339 284
rect 17602 240 17636 607
rect 16978 188 17636 240
rect 17276 166 17368 188
rect 17276 114 17288 166
rect 17354 114 17368 166
rect 17276 110 17368 114
rect 18667 -10 18770 1240
rect 19003 1162 19074 1170
rect 19003 1094 19015 1162
rect 19072 1094 19082 1162
rect 19003 1086 19074 1094
rect 19157 981 19192 1491
rect 19247 1445 19339 1458
rect 19247 1382 19259 1445
rect 19330 1382 19339 1445
rect 19247 1373 19339 1382
rect 20332 1445 20424 1455
rect 20332 1383 20344 1445
rect 20414 1383 20424 1445
rect 20332 1370 20424 1383
rect 21720 1390 21755 1744
rect 20579 1328 20644 1331
rect 20579 1325 20648 1328
rect 20579 1265 20585 1325
rect 20644 1265 20654 1325
rect 20579 1261 20648 1265
rect 20579 1259 20644 1261
rect 21720 1244 21899 1390
rect 22058 1338 22145 2521
rect 23540 2328 23550 2388
rect 23630 2328 23640 2388
rect 23540 2288 23640 2328
rect 22743 2231 24546 2288
rect 22743 2144 22777 2231
rect 23918 2144 23952 2231
rect 22737 2132 22783 2144
rect 22737 1944 22743 2132
rect 22296 1932 22342 1944
rect 22296 1756 22302 1932
rect 22336 1756 22342 1932
rect 22296 1744 22342 1756
rect 22414 1932 22460 1944
rect 22414 1756 22420 1932
rect 22454 1756 22460 1932
rect 22414 1744 22460 1756
rect 22532 1932 22578 1944
rect 22532 1756 22538 1932
rect 22572 1756 22578 1932
rect 22532 1744 22578 1756
rect 22650 1932 22743 1944
rect 22650 1756 22656 1932
rect 22690 1756 22743 1932
rect 22777 1756 22783 2132
rect 22650 1744 22783 1756
rect 22855 2132 22901 2144
rect 22855 1756 22861 2132
rect 22895 1756 22901 2132
rect 22855 1744 22901 1756
rect 22973 2132 23019 2144
rect 22973 1756 22979 2132
rect 23013 1756 23019 2132
rect 22973 1744 23019 1756
rect 23091 2132 23137 2144
rect 23091 1756 23097 2132
rect 23131 1756 23137 2132
rect 23091 1744 23137 1756
rect 23204 2132 23250 2144
rect 23204 1756 23210 2132
rect 23244 1756 23250 2132
rect 23204 1744 23250 1756
rect 23322 2132 23368 2144
rect 23322 1756 23328 2132
rect 23362 1756 23368 2132
rect 23322 1744 23368 1756
rect 23440 2132 23486 2144
rect 23440 1756 23446 2132
rect 23480 1756 23486 2132
rect 23440 1744 23486 1756
rect 23558 2132 23604 2144
rect 23558 1756 23564 2132
rect 23598 1756 23604 2132
rect 23558 1744 23604 1756
rect 23676 2132 23722 2144
rect 23676 1756 23682 2132
rect 23716 1756 23722 2132
rect 23676 1744 23722 1756
rect 23794 2132 23840 2144
rect 23794 1756 23800 2132
rect 23834 1756 23840 2132
rect 23794 1744 23840 1756
rect 23912 2132 23958 2144
rect 23912 1756 23918 2132
rect 23952 1756 23958 2132
rect 23912 1744 23958 1756
rect 24031 2132 24077 2144
rect 24031 1756 24037 2132
rect 24071 1756 24077 2132
rect 24031 1744 24077 1756
rect 24149 2132 24195 2144
rect 24149 1756 24155 2132
rect 24189 1756 24195 2132
rect 24149 1744 24195 1756
rect 24267 2132 24313 2144
rect 24267 1756 24273 2132
rect 24307 1756 24313 2132
rect 24267 1744 24313 1756
rect 24385 2132 24431 2144
rect 24385 1756 24391 2132
rect 24425 1756 24431 2132
rect 24509 1944 24546 2231
rect 24385 1744 24431 1756
rect 24504 1932 24550 1944
rect 24504 1756 24510 1932
rect 24544 1756 24550 1932
rect 24504 1744 24550 1756
rect 24622 1932 24668 1944
rect 24622 1756 24628 1932
rect 24662 1756 24668 1932
rect 24622 1744 24668 1756
rect 24740 1932 24786 1944
rect 24740 1756 24746 1932
rect 24780 1756 24786 1932
rect 24740 1744 24786 1756
rect 24858 1932 24904 1944
rect 24858 1756 24864 1932
rect 24898 1756 24904 1932
rect 24858 1744 24904 1756
rect 22301 1558 22336 1744
rect 23210 1660 23244 1744
rect 24391 1660 24425 1744
rect 23210 1618 24425 1660
rect 24391 1598 24425 1618
rect 24391 1582 24748 1598
rect 22301 1541 23438 1558
rect 22301 1507 23388 1541
rect 23422 1507 23438 1541
rect 24391 1548 24698 1582
rect 24732 1548 24748 1582
rect 24391 1532 24748 1548
rect 22301 1491 23438 1507
rect 22058 1330 22218 1338
rect 22058 1262 22159 1330
rect 22216 1262 22226 1330
rect 22058 1254 22218 1262
rect 20214 1162 20306 1170
rect 20214 1097 20226 1162
rect 20294 1097 20306 1162
rect 20214 1085 20306 1097
rect 21720 982 21755 1244
rect 19157 934 20529 981
rect 20851 935 21755 982
rect 19991 811 20025 934
rect 20463 921 20529 934
rect 20463 887 20479 921
rect 20513 887 20529 921
rect 20463 871 20529 887
rect 20852 811 20886 935
rect 19986 799 20032 811
rect 19986 623 19992 799
rect 20026 623 20032 799
rect 19986 611 20032 623
rect 20104 799 20224 811
rect 20104 623 20110 799
rect 20144 623 20184 799
rect 20104 611 20184 623
rect 20110 244 20144 611
rect 20178 423 20184 611
rect 20218 423 20224 799
rect 20178 411 20224 423
rect 20296 799 20342 811
rect 20296 423 20302 799
rect 20336 423 20342 799
rect 20296 411 20342 423
rect 20414 799 20460 811
rect 20414 423 20420 799
rect 20454 423 20460 799
rect 20414 411 20460 423
rect 20532 799 20578 811
rect 20532 423 20538 799
rect 20572 423 20578 799
rect 20532 411 20578 423
rect 20650 799 20774 811
rect 20650 423 20656 799
rect 20690 623 20734 799
rect 20768 623 20774 799
rect 20690 611 20774 623
rect 20846 799 20892 811
rect 20846 623 20852 799
rect 20886 623 20892 799
rect 20846 611 20892 623
rect 20690 423 20696 611
rect 20650 411 20696 423
rect 20420 338 20454 411
rect 20405 322 20471 338
rect 20405 288 20421 322
rect 20455 288 20471 322
rect 20405 272 20471 288
rect 20734 244 20768 611
rect 20110 192 20768 244
rect 20408 170 20500 192
rect 20408 118 20420 170
rect 20486 118 20500 170
rect 20408 114 20500 118
rect 21808 -10 21899 1244
rect 22148 1162 22218 1170
rect 22148 1094 22159 1162
rect 22216 1094 22226 1162
rect 22148 1086 22218 1094
rect 22301 981 22336 1491
rect 22391 1445 22483 1458
rect 22391 1382 22403 1445
rect 22474 1382 22483 1445
rect 22391 1373 22483 1382
rect 23476 1445 23568 1455
rect 23476 1383 23488 1445
rect 23558 1383 23568 1445
rect 23476 1370 23568 1383
rect 24864 1390 24899 1744
rect 23723 1328 23788 1331
rect 23723 1325 23792 1328
rect 23723 1265 23729 1325
rect 23788 1265 23798 1325
rect 23723 1261 23792 1265
rect 23723 1259 23788 1261
rect 24864 1244 25045 1390
rect 23358 1162 23450 1170
rect 23358 1097 23370 1162
rect 23438 1097 23450 1162
rect 23358 1085 23450 1097
rect 24864 982 24899 1244
rect 22301 934 23673 981
rect 23995 935 24899 982
rect 23135 811 23169 934
rect 23607 921 23673 934
rect 23607 887 23623 921
rect 23657 887 23673 921
rect 23607 871 23673 887
rect 23996 811 24030 935
rect 23130 799 23176 811
rect 23130 623 23136 799
rect 23170 623 23176 799
rect 23130 611 23176 623
rect 23248 799 23368 811
rect 23248 623 23254 799
rect 23288 623 23328 799
rect 23248 611 23328 623
rect 23254 244 23288 611
rect 23322 423 23328 611
rect 23362 423 23368 799
rect 23322 411 23368 423
rect 23440 799 23486 811
rect 23440 423 23446 799
rect 23480 423 23486 799
rect 23440 411 23486 423
rect 23558 799 23604 811
rect 23558 423 23564 799
rect 23598 423 23604 799
rect 23558 411 23604 423
rect 23676 799 23722 811
rect 23676 423 23682 799
rect 23716 423 23722 799
rect 23676 411 23722 423
rect 23794 799 23918 811
rect 23794 423 23800 799
rect 23834 623 23878 799
rect 23912 623 23918 799
rect 23834 611 23918 623
rect 23990 799 24036 811
rect 23990 623 23996 799
rect 24030 623 24036 799
rect 23990 611 24036 623
rect 23834 423 23840 611
rect 23794 411 23840 423
rect 23564 338 23598 411
rect 23549 322 23615 338
rect 23549 288 23565 322
rect 23599 288 23615 322
rect 23549 272 23615 288
rect 23878 244 23912 611
rect 23254 192 23912 244
rect 23552 170 23644 192
rect 23552 118 23564 170
rect 23630 118 23644 170
rect 23552 114 23644 118
rect 24965 -9 25045 1244
rect 0 -78 3002 -14
rect 3144 -78 6145 -13
rect 6276 -78 9278 -13
rect 9420 -78 12418 -10
rect 12622 -78 15625 -10
rect 15766 -78 18770 -10
rect 18898 -78 21899 -10
rect 22042 -77 25045 -9
rect 0 -1400 72 -78
rect 1498 -410 1508 -350
rect 1588 -410 1598 -350
rect 1498 -450 1598 -410
rect 701 -507 2504 -450
rect 701 -594 735 -507
rect 1876 -594 1910 -507
rect 695 -606 741 -594
rect 695 -794 701 -606
rect 254 -806 300 -794
rect 254 -982 260 -806
rect 294 -982 300 -806
rect 254 -994 300 -982
rect 372 -806 418 -794
rect 372 -982 378 -806
rect 412 -982 418 -806
rect 372 -994 418 -982
rect 490 -806 536 -794
rect 490 -982 496 -806
rect 530 -982 536 -806
rect 490 -994 536 -982
rect 608 -806 701 -794
rect 608 -982 614 -806
rect 648 -982 701 -806
rect 735 -982 741 -606
rect 608 -994 741 -982
rect 813 -606 859 -594
rect 813 -982 819 -606
rect 853 -982 859 -606
rect 813 -994 859 -982
rect 931 -606 977 -594
rect 931 -982 937 -606
rect 971 -982 977 -606
rect 931 -994 977 -982
rect 1049 -606 1095 -594
rect 1049 -982 1055 -606
rect 1089 -982 1095 -606
rect 1049 -994 1095 -982
rect 1162 -606 1208 -594
rect 1162 -982 1168 -606
rect 1202 -982 1208 -606
rect 1162 -994 1208 -982
rect 1280 -606 1326 -594
rect 1280 -982 1286 -606
rect 1320 -982 1326 -606
rect 1280 -994 1326 -982
rect 1398 -606 1444 -594
rect 1398 -982 1404 -606
rect 1438 -982 1444 -606
rect 1398 -994 1444 -982
rect 1516 -606 1562 -594
rect 1516 -982 1522 -606
rect 1556 -982 1562 -606
rect 1516 -994 1562 -982
rect 1634 -606 1680 -594
rect 1634 -982 1640 -606
rect 1674 -982 1680 -606
rect 1634 -994 1680 -982
rect 1752 -606 1798 -594
rect 1752 -982 1758 -606
rect 1792 -982 1798 -606
rect 1752 -994 1798 -982
rect 1870 -606 1916 -594
rect 1870 -982 1876 -606
rect 1910 -982 1916 -606
rect 1870 -994 1916 -982
rect 1989 -606 2035 -594
rect 1989 -982 1995 -606
rect 2029 -982 2035 -606
rect 1989 -994 2035 -982
rect 2107 -606 2153 -594
rect 2107 -982 2113 -606
rect 2147 -982 2153 -606
rect 2107 -994 2153 -982
rect 2225 -606 2271 -594
rect 2225 -982 2231 -606
rect 2265 -982 2271 -606
rect 2225 -994 2271 -982
rect 2343 -606 2389 -594
rect 2343 -982 2349 -606
rect 2383 -982 2389 -606
rect 2467 -794 2504 -507
rect 2343 -994 2389 -982
rect 2462 -806 2508 -794
rect 2462 -982 2468 -806
rect 2502 -982 2508 -806
rect 2462 -994 2508 -982
rect 2580 -806 2626 -794
rect 2580 -982 2586 -806
rect 2620 -982 2626 -806
rect 2580 -994 2626 -982
rect 2698 -806 2744 -794
rect 2698 -982 2704 -806
rect 2738 -982 2744 -806
rect 2698 -994 2744 -982
rect 2816 -806 2862 -794
rect 2816 -982 2822 -806
rect 2856 -982 2862 -806
rect 2816 -994 2862 -982
rect 259 -1180 294 -994
rect 1168 -1078 1202 -994
rect 2349 -1078 2383 -994
rect 1168 -1120 2383 -1078
rect 2349 -1140 2383 -1120
rect 2349 -1156 2706 -1140
rect 259 -1197 1396 -1180
rect 259 -1231 1346 -1197
rect 1380 -1231 1396 -1197
rect 2349 -1190 2656 -1156
rect 2690 -1190 2706 -1156
rect 2349 -1206 2706 -1190
rect 259 -1247 1396 -1231
rect 0 -1408 176 -1400
rect -519 -1615 -409 -1467
rect 0 -1476 117 -1408
rect 174 -1476 184 -1408
rect 0 -1484 176 -1476
rect -519 -1685 -496 -1615
rect -429 -1685 -409 -1615
rect -519 -4016 -409 -1685
rect 0 -1576 176 -1568
rect 0 -1644 117 -1576
rect 174 -1644 184 -1576
rect 0 -1652 176 -1644
rect 0 -2840 84 -1652
rect 259 -1757 294 -1247
rect 349 -1293 441 -1280
rect 349 -1356 361 -1293
rect 432 -1356 441 -1293
rect 349 -1365 441 -1356
rect 1434 -1293 1526 -1283
rect 1434 -1355 1446 -1293
rect 1516 -1355 1526 -1293
rect 1434 -1368 1526 -1355
rect 2822 -1348 2857 -994
rect 1681 -1410 1746 -1407
rect 1681 -1413 1750 -1410
rect 1681 -1473 1687 -1413
rect 1746 -1473 1756 -1413
rect 1681 -1477 1750 -1473
rect 1681 -1479 1746 -1477
rect 2822 -1494 3003 -1348
rect 3144 -1400 3215 -78
rect 4642 -410 4652 -350
rect 4732 -410 4742 -350
rect 4642 -450 4742 -410
rect 3845 -507 5648 -450
rect 3845 -594 3879 -507
rect 5020 -594 5054 -507
rect 3839 -606 3885 -594
rect 3839 -794 3845 -606
rect 3398 -806 3444 -794
rect 3398 -982 3404 -806
rect 3438 -982 3444 -806
rect 3398 -994 3444 -982
rect 3516 -806 3562 -794
rect 3516 -982 3522 -806
rect 3556 -982 3562 -806
rect 3516 -994 3562 -982
rect 3634 -806 3680 -794
rect 3634 -982 3640 -806
rect 3674 -982 3680 -806
rect 3634 -994 3680 -982
rect 3752 -806 3845 -794
rect 3752 -982 3758 -806
rect 3792 -982 3845 -806
rect 3879 -982 3885 -606
rect 3752 -994 3885 -982
rect 3957 -606 4003 -594
rect 3957 -982 3963 -606
rect 3997 -982 4003 -606
rect 3957 -994 4003 -982
rect 4075 -606 4121 -594
rect 4075 -982 4081 -606
rect 4115 -982 4121 -606
rect 4075 -994 4121 -982
rect 4193 -606 4239 -594
rect 4193 -982 4199 -606
rect 4233 -982 4239 -606
rect 4193 -994 4239 -982
rect 4306 -606 4352 -594
rect 4306 -982 4312 -606
rect 4346 -982 4352 -606
rect 4306 -994 4352 -982
rect 4424 -606 4470 -594
rect 4424 -982 4430 -606
rect 4464 -982 4470 -606
rect 4424 -994 4470 -982
rect 4542 -606 4588 -594
rect 4542 -982 4548 -606
rect 4582 -982 4588 -606
rect 4542 -994 4588 -982
rect 4660 -606 4706 -594
rect 4660 -982 4666 -606
rect 4700 -982 4706 -606
rect 4660 -994 4706 -982
rect 4778 -606 4824 -594
rect 4778 -982 4784 -606
rect 4818 -982 4824 -606
rect 4778 -994 4824 -982
rect 4896 -606 4942 -594
rect 4896 -982 4902 -606
rect 4936 -982 4942 -606
rect 4896 -994 4942 -982
rect 5014 -606 5060 -594
rect 5014 -982 5020 -606
rect 5054 -982 5060 -606
rect 5014 -994 5060 -982
rect 5133 -606 5179 -594
rect 5133 -982 5139 -606
rect 5173 -982 5179 -606
rect 5133 -994 5179 -982
rect 5251 -606 5297 -594
rect 5251 -982 5257 -606
rect 5291 -982 5297 -606
rect 5251 -994 5297 -982
rect 5369 -606 5415 -594
rect 5369 -982 5375 -606
rect 5409 -982 5415 -606
rect 5369 -994 5415 -982
rect 5487 -606 5533 -594
rect 5487 -982 5493 -606
rect 5527 -982 5533 -606
rect 5611 -794 5648 -507
rect 5487 -994 5533 -982
rect 5606 -806 5652 -794
rect 5606 -982 5612 -806
rect 5646 -982 5652 -806
rect 5606 -994 5652 -982
rect 5724 -806 5770 -794
rect 5724 -982 5730 -806
rect 5764 -982 5770 -806
rect 5724 -994 5770 -982
rect 5842 -806 5888 -794
rect 5842 -982 5848 -806
rect 5882 -982 5888 -806
rect 5842 -994 5888 -982
rect 5960 -806 6006 -794
rect 5960 -982 5966 -806
rect 6000 -982 6006 -806
rect 5960 -994 6006 -982
rect 3403 -1180 3438 -994
rect 4312 -1078 4346 -994
rect 5493 -1078 5527 -994
rect 4312 -1120 5527 -1078
rect 5493 -1140 5527 -1120
rect 5493 -1156 5850 -1140
rect 3403 -1197 4540 -1180
rect 3403 -1231 4490 -1197
rect 4524 -1231 4540 -1197
rect 5493 -1190 5800 -1156
rect 5834 -1190 5850 -1156
rect 5493 -1206 5850 -1190
rect 3403 -1247 4540 -1231
rect 3144 -1408 3320 -1400
rect 3144 -1476 3261 -1408
rect 3318 -1476 3328 -1408
rect 3144 -1484 3320 -1476
rect 1316 -1576 1408 -1568
rect 1316 -1641 1328 -1576
rect 1396 -1641 1408 -1576
rect 1316 -1653 1408 -1641
rect 2822 -1756 2857 -1494
rect 259 -1804 1631 -1757
rect 1953 -1803 2857 -1756
rect 1093 -1927 1127 -1804
rect 1565 -1817 1631 -1804
rect 1565 -1851 1581 -1817
rect 1615 -1851 1631 -1817
rect 1565 -1867 1631 -1851
rect 1954 -1927 1988 -1803
rect 1088 -1939 1134 -1927
rect 1088 -2115 1094 -1939
rect 1128 -2115 1134 -1939
rect 1088 -2127 1134 -2115
rect 1206 -1939 1326 -1927
rect 1206 -2115 1212 -1939
rect 1246 -2115 1286 -1939
rect 1206 -2127 1286 -2115
rect 1212 -2494 1246 -2127
rect 1280 -2315 1286 -2127
rect 1320 -2315 1326 -1939
rect 1280 -2327 1326 -2315
rect 1398 -1939 1444 -1927
rect 1398 -2315 1404 -1939
rect 1438 -2315 1444 -1939
rect 1398 -2327 1444 -2315
rect 1516 -1939 1562 -1927
rect 1516 -2315 1522 -1939
rect 1556 -2315 1562 -1939
rect 1516 -2327 1562 -2315
rect 1634 -1939 1680 -1927
rect 1634 -2315 1640 -1939
rect 1674 -2315 1680 -1939
rect 1634 -2327 1680 -2315
rect 1752 -1939 1876 -1927
rect 1752 -2315 1758 -1939
rect 1792 -2115 1836 -1939
rect 1870 -2115 1876 -1939
rect 1792 -2127 1876 -2115
rect 1948 -1939 1994 -1927
rect 1948 -2115 1954 -1939
rect 1988 -2115 1994 -1939
rect 1948 -2127 1994 -2115
rect 1792 -2315 1798 -2127
rect 1752 -2327 1798 -2315
rect 1522 -2400 1556 -2327
rect 1507 -2416 1573 -2400
rect 1507 -2450 1523 -2416
rect 1557 -2450 1573 -2416
rect 1507 -2466 1573 -2450
rect 1836 -2494 1870 -2127
rect 1212 -2546 1870 -2494
rect 2930 -2537 3003 -1494
rect 3144 -1576 3320 -1568
rect 3144 -1644 3261 -1576
rect 3318 -1644 3328 -1576
rect 3144 -1649 3320 -1644
rect 3143 -1652 3320 -1649
rect 1510 -2568 1602 -2546
rect 1510 -2620 1522 -2568
rect 1588 -2620 1602 -2568
rect 2926 -2614 2936 -2537
rect 3000 -2614 3010 -2537
rect 2930 -2615 3003 -2614
rect 1510 -2624 1602 -2620
rect 3143 -2839 3218 -1652
rect 3403 -1757 3438 -1247
rect 3493 -1293 3585 -1280
rect 3493 -1356 3505 -1293
rect 3576 -1356 3585 -1293
rect 3493 -1365 3585 -1356
rect 4578 -1293 4670 -1283
rect 4578 -1355 4590 -1293
rect 4660 -1355 4670 -1293
rect 4578 -1368 4670 -1355
rect 5966 -1348 6001 -994
rect 4825 -1410 4890 -1407
rect 4825 -1413 4894 -1410
rect 4825 -1473 4831 -1413
rect 4890 -1473 4900 -1413
rect 4825 -1477 4894 -1473
rect 5966 -1476 6147 -1348
rect 6276 -1396 6347 -78
rect 7774 -406 7784 -346
rect 7864 -406 7874 -346
rect 7774 -446 7874 -406
rect 6977 -503 8780 -446
rect 6977 -590 7011 -503
rect 8152 -590 8186 -503
rect 6971 -602 7017 -590
rect 6971 -790 6977 -602
rect 6530 -802 6576 -790
rect 6530 -978 6536 -802
rect 6570 -978 6576 -802
rect 6530 -990 6576 -978
rect 6648 -802 6694 -790
rect 6648 -978 6654 -802
rect 6688 -978 6694 -802
rect 6648 -990 6694 -978
rect 6766 -802 6812 -790
rect 6766 -978 6772 -802
rect 6806 -978 6812 -802
rect 6766 -990 6812 -978
rect 6884 -802 6977 -790
rect 6884 -978 6890 -802
rect 6924 -978 6977 -802
rect 7011 -978 7017 -602
rect 6884 -990 7017 -978
rect 7089 -602 7135 -590
rect 7089 -978 7095 -602
rect 7129 -978 7135 -602
rect 7089 -990 7135 -978
rect 7207 -602 7253 -590
rect 7207 -978 7213 -602
rect 7247 -978 7253 -602
rect 7207 -990 7253 -978
rect 7325 -602 7371 -590
rect 7325 -978 7331 -602
rect 7365 -978 7371 -602
rect 7325 -990 7371 -978
rect 7438 -602 7484 -590
rect 7438 -978 7444 -602
rect 7478 -978 7484 -602
rect 7438 -990 7484 -978
rect 7556 -602 7602 -590
rect 7556 -978 7562 -602
rect 7596 -978 7602 -602
rect 7556 -990 7602 -978
rect 7674 -602 7720 -590
rect 7674 -978 7680 -602
rect 7714 -978 7720 -602
rect 7674 -990 7720 -978
rect 7792 -602 7838 -590
rect 7792 -978 7798 -602
rect 7832 -978 7838 -602
rect 7792 -990 7838 -978
rect 7910 -602 7956 -590
rect 7910 -978 7916 -602
rect 7950 -978 7956 -602
rect 7910 -990 7956 -978
rect 8028 -602 8074 -590
rect 8028 -978 8034 -602
rect 8068 -978 8074 -602
rect 8028 -990 8074 -978
rect 8146 -602 8192 -590
rect 8146 -978 8152 -602
rect 8186 -978 8192 -602
rect 8146 -990 8192 -978
rect 8265 -602 8311 -590
rect 8265 -978 8271 -602
rect 8305 -978 8311 -602
rect 8265 -990 8311 -978
rect 8383 -602 8429 -590
rect 8383 -978 8389 -602
rect 8423 -978 8429 -602
rect 8383 -990 8429 -978
rect 8501 -602 8547 -590
rect 8501 -978 8507 -602
rect 8541 -978 8547 -602
rect 8501 -990 8547 -978
rect 8619 -602 8665 -590
rect 8619 -978 8625 -602
rect 8659 -978 8665 -602
rect 8743 -790 8780 -503
rect 8619 -990 8665 -978
rect 8738 -802 8784 -790
rect 8738 -978 8744 -802
rect 8778 -978 8784 -802
rect 8738 -990 8784 -978
rect 8856 -802 8902 -790
rect 8856 -978 8862 -802
rect 8896 -978 8902 -802
rect 8856 -990 8902 -978
rect 8974 -802 9020 -790
rect 8974 -978 8980 -802
rect 9014 -978 9020 -802
rect 8974 -990 9020 -978
rect 9092 -802 9138 -790
rect 9092 -978 9098 -802
rect 9132 -978 9138 -802
rect 9092 -990 9138 -978
rect 6535 -1176 6570 -990
rect 7444 -1074 7478 -990
rect 8625 -1074 8659 -990
rect 7444 -1116 8659 -1074
rect 8625 -1136 8659 -1116
rect 8625 -1152 8982 -1136
rect 6535 -1193 7672 -1176
rect 6535 -1227 7622 -1193
rect 7656 -1227 7672 -1193
rect 8625 -1186 8932 -1152
rect 8966 -1186 8982 -1152
rect 8625 -1202 8982 -1186
rect 6535 -1243 7672 -1227
rect 6276 -1404 6452 -1396
rect 6276 -1472 6393 -1404
rect 6450 -1472 6460 -1404
rect 4825 -1479 4890 -1477
rect 5966 -1494 6148 -1476
rect 6276 -1480 6452 -1472
rect 4460 -1576 4552 -1568
rect 4460 -1641 4472 -1576
rect 4540 -1641 4552 -1576
rect 4460 -1653 4552 -1641
rect 5966 -1756 6001 -1494
rect 3403 -1804 4775 -1757
rect 5097 -1803 6001 -1756
rect 4237 -1927 4271 -1804
rect 4709 -1817 4775 -1804
rect 4709 -1851 4725 -1817
rect 4759 -1851 4775 -1817
rect 4709 -1867 4775 -1851
rect 5098 -1927 5132 -1803
rect 4232 -1939 4278 -1927
rect 4232 -2115 4238 -1939
rect 4272 -2115 4278 -1939
rect 4232 -2127 4278 -2115
rect 4350 -1939 4470 -1927
rect 4350 -2115 4356 -1939
rect 4390 -2115 4430 -1939
rect 4350 -2127 4430 -2115
rect 4356 -2494 4390 -2127
rect 4424 -2315 4430 -2127
rect 4464 -2315 4470 -1939
rect 4424 -2327 4470 -2315
rect 4542 -1939 4588 -1927
rect 4542 -2315 4548 -1939
rect 4582 -2315 4588 -1939
rect 4542 -2327 4588 -2315
rect 4660 -1939 4706 -1927
rect 4660 -2315 4666 -1939
rect 4700 -2315 4706 -1939
rect 4660 -2327 4706 -2315
rect 4778 -1939 4824 -1927
rect 4778 -2315 4784 -1939
rect 4818 -2315 4824 -1939
rect 4778 -2327 4824 -2315
rect 4896 -1939 5020 -1927
rect 4896 -2315 4902 -1939
rect 4936 -2115 4980 -1939
rect 5014 -2115 5020 -1939
rect 4936 -2127 5020 -2115
rect 5092 -1939 5138 -1927
rect 5092 -2115 5098 -1939
rect 5132 -2115 5138 -1939
rect 5092 -2127 5138 -2115
rect 4936 -2315 4942 -2127
rect 4896 -2327 4942 -2315
rect 4666 -2400 4700 -2327
rect 4651 -2416 4717 -2400
rect 4651 -2450 4667 -2416
rect 4701 -2450 4717 -2416
rect 4651 -2466 4717 -2450
rect 4980 -2494 5014 -2127
rect 4356 -2546 5014 -2494
rect 4654 -2568 4746 -2546
rect 4654 -2620 4666 -2568
rect 4732 -2620 4746 -2568
rect 6050 -2596 6148 -1494
rect 4654 -2624 4746 -2620
rect 6036 -2668 6046 -2596
rect 6114 -2646 6148 -2596
rect 6293 -1572 6452 -1564
rect 6293 -1640 6393 -1572
rect 6450 -1640 6460 -1572
rect 6293 -1648 6452 -1640
rect 6114 -2668 6124 -2646
rect 6293 -2839 6342 -1648
rect 6535 -1753 6570 -1243
rect 6625 -1289 6717 -1276
rect 6625 -1352 6637 -1289
rect 6708 -1352 6717 -1289
rect 6625 -1361 6717 -1352
rect 7710 -1289 7802 -1279
rect 7710 -1351 7722 -1289
rect 7792 -1351 7802 -1289
rect 7710 -1364 7802 -1351
rect 9098 -1344 9133 -990
rect 7957 -1406 8022 -1403
rect 7957 -1409 8026 -1406
rect 7957 -1469 7963 -1409
rect 8022 -1469 8032 -1409
rect 7957 -1473 8026 -1469
rect 7957 -1475 8022 -1473
rect 9098 -1490 9279 -1344
rect 9420 -1396 9491 -78
rect 10918 -406 10928 -346
rect 11008 -406 11018 -346
rect 10918 -446 11018 -406
rect 10121 -503 11924 -446
rect 10121 -590 10155 -503
rect 11296 -590 11330 -503
rect 10115 -602 10161 -590
rect 10115 -790 10121 -602
rect 9674 -802 9720 -790
rect 9674 -978 9680 -802
rect 9714 -978 9720 -802
rect 9674 -990 9720 -978
rect 9792 -802 9838 -790
rect 9792 -978 9798 -802
rect 9832 -978 9838 -802
rect 9792 -990 9838 -978
rect 9910 -802 9956 -790
rect 9910 -978 9916 -802
rect 9950 -978 9956 -802
rect 9910 -990 9956 -978
rect 10028 -802 10121 -790
rect 10028 -978 10034 -802
rect 10068 -978 10121 -802
rect 10155 -978 10161 -602
rect 10028 -990 10161 -978
rect 10233 -602 10279 -590
rect 10233 -978 10239 -602
rect 10273 -978 10279 -602
rect 10233 -990 10279 -978
rect 10351 -602 10397 -590
rect 10351 -978 10357 -602
rect 10391 -978 10397 -602
rect 10351 -990 10397 -978
rect 10469 -602 10515 -590
rect 10469 -978 10475 -602
rect 10509 -978 10515 -602
rect 10469 -990 10515 -978
rect 10582 -602 10628 -590
rect 10582 -978 10588 -602
rect 10622 -978 10628 -602
rect 10582 -990 10628 -978
rect 10700 -602 10746 -590
rect 10700 -978 10706 -602
rect 10740 -978 10746 -602
rect 10700 -990 10746 -978
rect 10818 -602 10864 -590
rect 10818 -978 10824 -602
rect 10858 -978 10864 -602
rect 10818 -990 10864 -978
rect 10936 -602 10982 -590
rect 10936 -978 10942 -602
rect 10976 -978 10982 -602
rect 10936 -990 10982 -978
rect 11054 -602 11100 -590
rect 11054 -978 11060 -602
rect 11094 -978 11100 -602
rect 11054 -990 11100 -978
rect 11172 -602 11218 -590
rect 11172 -978 11178 -602
rect 11212 -978 11218 -602
rect 11172 -990 11218 -978
rect 11290 -602 11336 -590
rect 11290 -978 11296 -602
rect 11330 -978 11336 -602
rect 11290 -990 11336 -978
rect 11409 -602 11455 -590
rect 11409 -978 11415 -602
rect 11449 -978 11455 -602
rect 11409 -990 11455 -978
rect 11527 -602 11573 -590
rect 11527 -978 11533 -602
rect 11567 -978 11573 -602
rect 11527 -990 11573 -978
rect 11645 -602 11691 -590
rect 11645 -978 11651 -602
rect 11685 -978 11691 -602
rect 11645 -990 11691 -978
rect 11763 -602 11809 -590
rect 11763 -978 11769 -602
rect 11803 -978 11809 -602
rect 11887 -790 11924 -503
rect 11763 -990 11809 -978
rect 11882 -802 11928 -790
rect 11882 -978 11888 -802
rect 11922 -978 11928 -802
rect 11882 -990 11928 -978
rect 12000 -802 12046 -790
rect 12000 -978 12006 -802
rect 12040 -978 12046 -802
rect 12000 -990 12046 -978
rect 12118 -802 12164 -790
rect 12118 -978 12124 -802
rect 12158 -978 12164 -802
rect 12118 -990 12164 -978
rect 12236 -802 12282 -790
rect 12236 -978 12242 -802
rect 12276 -978 12282 -802
rect 12236 -990 12282 -978
rect 9679 -1176 9714 -990
rect 10588 -1074 10622 -990
rect 11769 -1074 11803 -990
rect 10588 -1116 11803 -1074
rect 11769 -1136 11803 -1116
rect 11769 -1152 12126 -1136
rect 9679 -1193 10816 -1176
rect 9679 -1227 10766 -1193
rect 10800 -1227 10816 -1193
rect 11769 -1186 12076 -1152
rect 12110 -1186 12126 -1152
rect 11769 -1202 12126 -1186
rect 9679 -1243 10816 -1227
rect 9420 -1404 9596 -1396
rect 9420 -1472 9537 -1404
rect 9594 -1472 9604 -1404
rect 9420 -1480 9596 -1472
rect 7592 -1572 7684 -1564
rect 7592 -1637 7604 -1572
rect 7672 -1637 7684 -1572
rect 7592 -1649 7684 -1637
rect 9098 -1752 9133 -1490
rect 6535 -1800 7907 -1753
rect 8229 -1799 9133 -1752
rect 7369 -1923 7403 -1800
rect 7841 -1813 7907 -1800
rect 7841 -1847 7857 -1813
rect 7891 -1847 7907 -1813
rect 7841 -1863 7907 -1847
rect 8230 -1923 8264 -1799
rect 7364 -1935 7410 -1923
rect 7364 -2111 7370 -1935
rect 7404 -2111 7410 -1935
rect 7364 -2123 7410 -2111
rect 7482 -1935 7602 -1923
rect 7482 -2111 7488 -1935
rect 7522 -2111 7562 -1935
rect 7482 -2123 7562 -2111
rect 7488 -2490 7522 -2123
rect 7556 -2311 7562 -2123
rect 7596 -2311 7602 -1935
rect 7556 -2323 7602 -2311
rect 7674 -1935 7720 -1923
rect 7674 -2311 7680 -1935
rect 7714 -2311 7720 -1935
rect 7674 -2323 7720 -2311
rect 7792 -1935 7838 -1923
rect 7792 -2311 7798 -1935
rect 7832 -2311 7838 -1935
rect 7792 -2323 7838 -2311
rect 7910 -1935 7956 -1923
rect 7910 -2311 7916 -1935
rect 7950 -2311 7956 -1935
rect 7910 -2323 7956 -2311
rect 8028 -1935 8152 -1923
rect 8028 -2311 8034 -1935
rect 8068 -2111 8112 -1935
rect 8146 -2111 8152 -1935
rect 8068 -2123 8152 -2111
rect 8224 -1935 8270 -1923
rect 8224 -2111 8230 -1935
rect 8264 -2111 8270 -1935
rect 8224 -2123 8270 -2111
rect 8068 -2311 8074 -2123
rect 8028 -2323 8074 -2311
rect 7798 -2396 7832 -2323
rect 7783 -2412 7849 -2396
rect 7783 -2446 7799 -2412
rect 7833 -2446 7849 -2412
rect 7783 -2462 7849 -2446
rect 8112 -2490 8146 -2123
rect 7488 -2542 8146 -2490
rect 7786 -2564 7878 -2542
rect 7786 -2616 7798 -2564
rect 7864 -2616 7878 -2564
rect 7786 -2620 7878 -2616
rect 9188 -2722 9279 -1490
rect 9172 -2790 9182 -2722
rect 9249 -2788 9279 -2722
rect 9444 -1572 9596 -1564
rect 9444 -1640 9537 -1572
rect 9594 -1640 9604 -1572
rect 9444 -1648 9596 -1640
rect 9249 -2790 9259 -2788
rect 9444 -2839 9505 -1648
rect 9679 -1753 9714 -1243
rect 9769 -1289 9861 -1276
rect 9769 -1352 9781 -1289
rect 9852 -1352 9861 -1289
rect 9769 -1361 9861 -1352
rect 10854 -1289 10946 -1279
rect 10854 -1351 10866 -1289
rect 10936 -1351 10946 -1289
rect 10854 -1364 10946 -1351
rect 12242 -1344 12277 -990
rect 11101 -1406 11166 -1403
rect 11101 -1409 11170 -1406
rect 11101 -1469 11107 -1409
rect 11166 -1469 11176 -1409
rect 11101 -1473 11170 -1469
rect 11101 -1475 11166 -1473
rect 12242 -1490 12423 -1344
rect 12622 -1400 12693 -78
rect 14120 -410 14130 -350
rect 14210 -410 14220 -350
rect 14120 -450 14220 -410
rect 13323 -507 15126 -450
rect 13323 -594 13357 -507
rect 14498 -594 14532 -507
rect 13317 -606 13363 -594
rect 13317 -794 13323 -606
rect 12876 -806 12922 -794
rect 12876 -982 12882 -806
rect 12916 -982 12922 -806
rect 12876 -994 12922 -982
rect 12994 -806 13040 -794
rect 12994 -982 13000 -806
rect 13034 -982 13040 -806
rect 12994 -994 13040 -982
rect 13112 -806 13158 -794
rect 13112 -982 13118 -806
rect 13152 -982 13158 -806
rect 13112 -994 13158 -982
rect 13230 -806 13323 -794
rect 13230 -982 13236 -806
rect 13270 -982 13323 -806
rect 13357 -982 13363 -606
rect 13230 -994 13363 -982
rect 13435 -606 13481 -594
rect 13435 -982 13441 -606
rect 13475 -982 13481 -606
rect 13435 -994 13481 -982
rect 13553 -606 13599 -594
rect 13553 -982 13559 -606
rect 13593 -982 13599 -606
rect 13553 -994 13599 -982
rect 13671 -606 13717 -594
rect 13671 -982 13677 -606
rect 13711 -982 13717 -606
rect 13671 -994 13717 -982
rect 13784 -606 13830 -594
rect 13784 -982 13790 -606
rect 13824 -982 13830 -606
rect 13784 -994 13830 -982
rect 13902 -606 13948 -594
rect 13902 -982 13908 -606
rect 13942 -982 13948 -606
rect 13902 -994 13948 -982
rect 14020 -606 14066 -594
rect 14020 -982 14026 -606
rect 14060 -982 14066 -606
rect 14020 -994 14066 -982
rect 14138 -606 14184 -594
rect 14138 -982 14144 -606
rect 14178 -982 14184 -606
rect 14138 -994 14184 -982
rect 14256 -606 14302 -594
rect 14256 -982 14262 -606
rect 14296 -982 14302 -606
rect 14256 -994 14302 -982
rect 14374 -606 14420 -594
rect 14374 -982 14380 -606
rect 14414 -982 14420 -606
rect 14374 -994 14420 -982
rect 14492 -606 14538 -594
rect 14492 -982 14498 -606
rect 14532 -982 14538 -606
rect 14492 -994 14538 -982
rect 14611 -606 14657 -594
rect 14611 -982 14617 -606
rect 14651 -982 14657 -606
rect 14611 -994 14657 -982
rect 14729 -606 14775 -594
rect 14729 -982 14735 -606
rect 14769 -982 14775 -606
rect 14729 -994 14775 -982
rect 14847 -606 14893 -594
rect 14847 -982 14853 -606
rect 14887 -982 14893 -606
rect 14847 -994 14893 -982
rect 14965 -606 15011 -594
rect 14965 -982 14971 -606
rect 15005 -982 15011 -606
rect 15089 -794 15126 -507
rect 14965 -994 15011 -982
rect 15084 -806 15130 -794
rect 15084 -982 15090 -806
rect 15124 -982 15130 -806
rect 15084 -994 15130 -982
rect 15202 -806 15248 -794
rect 15202 -982 15208 -806
rect 15242 -982 15248 -806
rect 15202 -994 15248 -982
rect 15320 -806 15366 -794
rect 15320 -982 15326 -806
rect 15360 -982 15366 -806
rect 15320 -994 15366 -982
rect 15438 -806 15484 -794
rect 15438 -982 15444 -806
rect 15478 -982 15484 -806
rect 15438 -994 15484 -982
rect 12881 -1180 12916 -994
rect 13790 -1078 13824 -994
rect 14971 -1078 15005 -994
rect 13790 -1120 15005 -1078
rect 14971 -1140 15005 -1120
rect 14971 -1156 15328 -1140
rect 12881 -1197 14018 -1180
rect 12881 -1231 13968 -1197
rect 14002 -1231 14018 -1197
rect 14971 -1190 15278 -1156
rect 15312 -1190 15328 -1156
rect 14971 -1206 15328 -1190
rect 12881 -1247 14018 -1231
rect 12622 -1408 12798 -1400
rect 12622 -1476 12739 -1408
rect 12796 -1476 12806 -1408
rect 12622 -1484 12798 -1476
rect 10736 -1572 10828 -1564
rect 10736 -1637 10748 -1572
rect 10816 -1637 10828 -1572
rect 10736 -1649 10828 -1637
rect 12242 -1752 12277 -1490
rect 9679 -1800 11051 -1753
rect 11373 -1799 12277 -1752
rect 10513 -1923 10547 -1800
rect 10985 -1813 11051 -1800
rect 10985 -1847 11001 -1813
rect 11035 -1847 11051 -1813
rect 10985 -1863 11051 -1847
rect 11374 -1923 11408 -1799
rect 10508 -1935 10554 -1923
rect 10508 -2111 10514 -1935
rect 10548 -2111 10554 -1935
rect 10508 -2123 10554 -2111
rect 10626 -1935 10746 -1923
rect 10626 -2111 10632 -1935
rect 10666 -2111 10706 -1935
rect 10626 -2123 10706 -2111
rect 10632 -2490 10666 -2123
rect 10700 -2311 10706 -2123
rect 10740 -2311 10746 -1935
rect 10700 -2323 10746 -2311
rect 10818 -1935 10864 -1923
rect 10818 -2311 10824 -1935
rect 10858 -2311 10864 -1935
rect 10818 -2323 10864 -2311
rect 10936 -1935 10982 -1923
rect 10936 -2311 10942 -1935
rect 10976 -2311 10982 -1935
rect 10936 -2323 10982 -2311
rect 11054 -1935 11100 -1923
rect 11054 -2311 11060 -1935
rect 11094 -2311 11100 -1935
rect 11054 -2323 11100 -2311
rect 11172 -1935 11296 -1923
rect 11172 -2311 11178 -1935
rect 11212 -2111 11256 -1935
rect 11290 -2111 11296 -1935
rect 11212 -2123 11296 -2111
rect 11368 -1935 11414 -1923
rect 11368 -2111 11374 -1935
rect 11408 -2111 11414 -1935
rect 11368 -2123 11414 -2111
rect 11212 -2311 11218 -2123
rect 11172 -2323 11218 -2311
rect 10942 -2396 10976 -2323
rect 10927 -2412 10993 -2396
rect 10927 -2446 10943 -2412
rect 10977 -2446 10993 -2412
rect 10927 -2462 10993 -2446
rect 11256 -2490 11290 -2123
rect 12329 -2378 12422 -1490
rect 12319 -2447 12329 -2378
rect 12407 -2447 12422 -2378
rect 12622 -1576 12798 -1568
rect 12622 -1644 12739 -1576
rect 12796 -1644 12806 -1576
rect 12622 -1652 12798 -1644
rect 10632 -2542 11290 -2490
rect 10930 -2564 11022 -2542
rect 10930 -2616 10942 -2564
rect 11008 -2616 11022 -2564
rect 10930 -2620 11022 -2616
rect 12622 -2838 12698 -1652
rect 12881 -1757 12916 -1247
rect 12971 -1293 13063 -1280
rect 12971 -1356 12983 -1293
rect 13054 -1356 13063 -1293
rect 12971 -1365 13063 -1356
rect 14056 -1293 14148 -1283
rect 14056 -1355 14068 -1293
rect 14138 -1355 14148 -1293
rect 14056 -1368 14148 -1355
rect 15444 -1348 15479 -994
rect 14303 -1410 14368 -1407
rect 14303 -1413 14372 -1410
rect 14303 -1473 14309 -1413
rect 14368 -1473 14378 -1413
rect 15444 -1445 15625 -1348
rect 15766 -1400 15837 -78
rect 17264 -410 17274 -350
rect 17354 -410 17364 -350
rect 17264 -450 17364 -410
rect 16467 -507 18270 -450
rect 16467 -594 16501 -507
rect 17642 -594 17676 -507
rect 16461 -606 16507 -594
rect 16461 -794 16467 -606
rect 16020 -806 16066 -794
rect 16020 -982 16026 -806
rect 16060 -982 16066 -806
rect 16020 -994 16066 -982
rect 16138 -806 16184 -794
rect 16138 -982 16144 -806
rect 16178 -982 16184 -806
rect 16138 -994 16184 -982
rect 16256 -806 16302 -794
rect 16256 -982 16262 -806
rect 16296 -982 16302 -806
rect 16256 -994 16302 -982
rect 16374 -806 16467 -794
rect 16374 -982 16380 -806
rect 16414 -982 16467 -806
rect 16501 -982 16507 -606
rect 16374 -994 16507 -982
rect 16579 -606 16625 -594
rect 16579 -982 16585 -606
rect 16619 -982 16625 -606
rect 16579 -994 16625 -982
rect 16697 -606 16743 -594
rect 16697 -982 16703 -606
rect 16737 -982 16743 -606
rect 16697 -994 16743 -982
rect 16815 -606 16861 -594
rect 16815 -982 16821 -606
rect 16855 -982 16861 -606
rect 16815 -994 16861 -982
rect 16928 -606 16974 -594
rect 16928 -982 16934 -606
rect 16968 -982 16974 -606
rect 16928 -994 16974 -982
rect 17046 -606 17092 -594
rect 17046 -982 17052 -606
rect 17086 -982 17092 -606
rect 17046 -994 17092 -982
rect 17164 -606 17210 -594
rect 17164 -982 17170 -606
rect 17204 -982 17210 -606
rect 17164 -994 17210 -982
rect 17282 -606 17328 -594
rect 17282 -982 17288 -606
rect 17322 -982 17328 -606
rect 17282 -994 17328 -982
rect 17400 -606 17446 -594
rect 17400 -982 17406 -606
rect 17440 -982 17446 -606
rect 17400 -994 17446 -982
rect 17518 -606 17564 -594
rect 17518 -982 17524 -606
rect 17558 -982 17564 -606
rect 17518 -994 17564 -982
rect 17636 -606 17682 -594
rect 17636 -982 17642 -606
rect 17676 -982 17682 -606
rect 17636 -994 17682 -982
rect 17755 -606 17801 -594
rect 17755 -982 17761 -606
rect 17795 -982 17801 -606
rect 17755 -994 17801 -982
rect 17873 -606 17919 -594
rect 17873 -982 17879 -606
rect 17913 -982 17919 -606
rect 17873 -994 17919 -982
rect 17991 -606 18037 -594
rect 17991 -982 17997 -606
rect 18031 -982 18037 -606
rect 17991 -994 18037 -982
rect 18109 -606 18155 -594
rect 18109 -982 18115 -606
rect 18149 -982 18155 -606
rect 18233 -794 18270 -507
rect 18109 -994 18155 -982
rect 18228 -806 18274 -794
rect 18228 -982 18234 -806
rect 18268 -982 18274 -806
rect 18228 -994 18274 -982
rect 18346 -806 18392 -794
rect 18346 -982 18352 -806
rect 18386 -982 18392 -806
rect 18346 -994 18392 -982
rect 18464 -806 18510 -794
rect 18464 -982 18470 -806
rect 18504 -982 18510 -806
rect 18464 -994 18510 -982
rect 18582 -806 18628 -794
rect 18582 -982 18588 -806
rect 18622 -982 18628 -806
rect 18582 -994 18628 -982
rect 16025 -1180 16060 -994
rect 16934 -1078 16968 -994
rect 18115 -1078 18149 -994
rect 16934 -1120 18149 -1078
rect 18115 -1140 18149 -1120
rect 18115 -1156 18472 -1140
rect 16025 -1197 17162 -1180
rect 16025 -1231 17112 -1197
rect 17146 -1231 17162 -1197
rect 18115 -1190 18422 -1156
rect 18456 -1190 18472 -1156
rect 18115 -1206 18472 -1190
rect 16025 -1247 17162 -1231
rect 15876 -1292 15942 -1284
rect 15876 -1360 15883 -1292
rect 15940 -1360 15950 -1292
rect 15876 -1368 15942 -1360
rect 15766 -1408 15942 -1400
rect 14303 -1477 14372 -1473
rect 14303 -1479 14368 -1477
rect 15444 -1494 15627 -1445
rect 15766 -1476 15883 -1408
rect 15940 -1476 15950 -1408
rect 15766 -1484 15942 -1476
rect 13938 -1576 14030 -1568
rect 13938 -1641 13950 -1576
rect 14018 -1641 14030 -1576
rect 13938 -1653 14030 -1641
rect 15444 -1756 15479 -1494
rect 12881 -1804 14253 -1757
rect 14575 -1803 15479 -1756
rect 13715 -1927 13749 -1804
rect 14187 -1817 14253 -1804
rect 14187 -1851 14203 -1817
rect 14237 -1851 14253 -1817
rect 14187 -1867 14253 -1851
rect 14576 -1927 14610 -1803
rect 13710 -1939 13756 -1927
rect 13710 -2115 13716 -1939
rect 13750 -2115 13756 -1939
rect 13710 -2127 13756 -2115
rect 13828 -1939 13948 -1927
rect 13828 -2115 13834 -1939
rect 13868 -2115 13908 -1939
rect 13828 -2127 13908 -2115
rect 13834 -2494 13868 -2127
rect 13902 -2315 13908 -2127
rect 13942 -2315 13948 -1939
rect 13902 -2327 13948 -2315
rect 14020 -1939 14066 -1927
rect 14020 -2315 14026 -1939
rect 14060 -2315 14066 -1939
rect 14020 -2327 14066 -2315
rect 14138 -1939 14184 -1927
rect 14138 -2315 14144 -1939
rect 14178 -2315 14184 -1939
rect 14138 -2327 14184 -2315
rect 14256 -1939 14302 -1927
rect 14256 -2315 14262 -1939
rect 14296 -2315 14302 -1939
rect 14256 -2327 14302 -2315
rect 14374 -1939 14498 -1927
rect 14374 -2315 14380 -1939
rect 14414 -2115 14458 -1939
rect 14492 -2115 14498 -1939
rect 14414 -2127 14498 -2115
rect 14570 -1939 14616 -1927
rect 14570 -2115 14576 -1939
rect 14610 -2115 14616 -1939
rect 14570 -2127 14616 -2115
rect 14414 -2315 14420 -2127
rect 14374 -2327 14420 -2315
rect 14144 -2400 14178 -2327
rect 14129 -2416 14195 -2400
rect 14129 -2450 14145 -2416
rect 14179 -2450 14195 -2416
rect 14129 -2466 14195 -2450
rect 14458 -2494 14492 -2127
rect 15529 -2174 15627 -1494
rect 15790 -1576 15942 -1568
rect 15790 -1644 15883 -1576
rect 15940 -1644 15950 -1576
rect 15790 -1652 15942 -1644
rect 15519 -2269 15529 -2174
rect 15625 -2269 15635 -2174
rect 13834 -2546 14492 -2494
rect 14132 -2568 14224 -2546
rect 14132 -2620 14144 -2568
rect 14210 -2620 14224 -2568
rect 14132 -2624 14224 -2620
rect 15790 -2838 15847 -1652
rect 16025 -1757 16060 -1247
rect 16115 -1293 16207 -1280
rect 16115 -1356 16127 -1293
rect 16198 -1356 16207 -1293
rect 16115 -1365 16207 -1356
rect 17200 -1293 17292 -1283
rect 17200 -1355 17212 -1293
rect 17282 -1355 17292 -1293
rect 17200 -1368 17292 -1355
rect 18588 -1348 18623 -994
rect 17447 -1410 17512 -1407
rect 17447 -1413 17516 -1410
rect 17447 -1473 17453 -1413
rect 17512 -1473 17522 -1413
rect 17447 -1477 17516 -1473
rect 17447 -1479 17512 -1477
rect 18588 -1494 18769 -1348
rect 18898 -1396 18969 -78
rect 20396 -406 20406 -346
rect 20486 -406 20496 -346
rect 20396 -446 20496 -406
rect 19599 -503 21402 -446
rect 19599 -590 19633 -503
rect 20774 -590 20808 -503
rect 19593 -602 19639 -590
rect 19593 -790 19599 -602
rect 19152 -802 19198 -790
rect 19152 -978 19158 -802
rect 19192 -978 19198 -802
rect 19152 -990 19198 -978
rect 19270 -802 19316 -790
rect 19270 -978 19276 -802
rect 19310 -978 19316 -802
rect 19270 -990 19316 -978
rect 19388 -802 19434 -790
rect 19388 -978 19394 -802
rect 19428 -978 19434 -802
rect 19388 -990 19434 -978
rect 19506 -802 19599 -790
rect 19506 -978 19512 -802
rect 19546 -978 19599 -802
rect 19633 -978 19639 -602
rect 19506 -990 19639 -978
rect 19711 -602 19757 -590
rect 19711 -978 19717 -602
rect 19751 -978 19757 -602
rect 19711 -990 19757 -978
rect 19829 -602 19875 -590
rect 19829 -978 19835 -602
rect 19869 -978 19875 -602
rect 19829 -990 19875 -978
rect 19947 -602 19993 -590
rect 19947 -978 19953 -602
rect 19987 -978 19993 -602
rect 19947 -990 19993 -978
rect 20060 -602 20106 -590
rect 20060 -978 20066 -602
rect 20100 -978 20106 -602
rect 20060 -990 20106 -978
rect 20178 -602 20224 -590
rect 20178 -978 20184 -602
rect 20218 -978 20224 -602
rect 20178 -990 20224 -978
rect 20296 -602 20342 -590
rect 20296 -978 20302 -602
rect 20336 -978 20342 -602
rect 20296 -990 20342 -978
rect 20414 -602 20460 -590
rect 20414 -978 20420 -602
rect 20454 -978 20460 -602
rect 20414 -990 20460 -978
rect 20532 -602 20578 -590
rect 20532 -978 20538 -602
rect 20572 -978 20578 -602
rect 20532 -990 20578 -978
rect 20650 -602 20696 -590
rect 20650 -978 20656 -602
rect 20690 -978 20696 -602
rect 20650 -990 20696 -978
rect 20768 -602 20814 -590
rect 20768 -978 20774 -602
rect 20808 -978 20814 -602
rect 20768 -990 20814 -978
rect 20887 -602 20933 -590
rect 20887 -978 20893 -602
rect 20927 -978 20933 -602
rect 20887 -990 20933 -978
rect 21005 -602 21051 -590
rect 21005 -978 21011 -602
rect 21045 -978 21051 -602
rect 21005 -990 21051 -978
rect 21123 -602 21169 -590
rect 21123 -978 21129 -602
rect 21163 -978 21169 -602
rect 21123 -990 21169 -978
rect 21241 -602 21287 -590
rect 21241 -978 21247 -602
rect 21281 -978 21287 -602
rect 21365 -790 21402 -503
rect 21241 -990 21287 -978
rect 21360 -802 21406 -790
rect 21360 -978 21366 -802
rect 21400 -978 21406 -802
rect 21360 -990 21406 -978
rect 21478 -802 21524 -790
rect 21478 -978 21484 -802
rect 21518 -978 21524 -802
rect 21478 -990 21524 -978
rect 21596 -802 21642 -790
rect 21596 -978 21602 -802
rect 21636 -978 21642 -802
rect 21596 -990 21642 -978
rect 21714 -802 21760 -790
rect 21714 -978 21720 -802
rect 21754 -978 21760 -802
rect 21714 -990 21760 -978
rect 19157 -1176 19192 -990
rect 20066 -1074 20100 -990
rect 21247 -1074 21281 -990
rect 20066 -1116 21281 -1074
rect 21247 -1136 21281 -1116
rect 21247 -1152 21604 -1136
rect 19157 -1193 20294 -1176
rect 19157 -1227 20244 -1193
rect 20278 -1227 20294 -1193
rect 21247 -1186 21554 -1152
rect 21588 -1186 21604 -1152
rect 21247 -1202 21604 -1186
rect 19157 -1243 20294 -1227
rect 18898 -1404 19074 -1396
rect 18898 -1472 19015 -1404
rect 19072 -1472 19082 -1404
rect 18898 -1480 19074 -1472
rect 17082 -1576 17174 -1568
rect 17082 -1641 17094 -1576
rect 17162 -1641 17174 -1576
rect 17082 -1653 17174 -1641
rect 18588 -1756 18623 -1494
rect 16025 -1804 17397 -1757
rect 17719 -1803 18623 -1756
rect 16859 -1927 16893 -1804
rect 17331 -1817 17397 -1804
rect 17331 -1851 17347 -1817
rect 17381 -1851 17397 -1817
rect 17331 -1867 17397 -1851
rect 17720 -1927 17754 -1803
rect 16854 -1939 16900 -1927
rect 16854 -2115 16860 -1939
rect 16894 -2115 16900 -1939
rect 16854 -2127 16900 -2115
rect 16972 -1939 17092 -1927
rect 16972 -2115 16978 -1939
rect 17012 -2115 17052 -1939
rect 16972 -2127 17052 -2115
rect 16978 -2494 17012 -2127
rect 17046 -2315 17052 -2127
rect 17086 -2315 17092 -1939
rect 17046 -2327 17092 -2315
rect 17164 -1939 17210 -1927
rect 17164 -2315 17170 -1939
rect 17204 -2315 17210 -1939
rect 17164 -2327 17210 -2315
rect 17282 -1939 17328 -1927
rect 17282 -2315 17288 -1939
rect 17322 -2315 17328 -1939
rect 17282 -2327 17328 -2315
rect 17400 -1939 17446 -1927
rect 17400 -2315 17406 -1939
rect 17440 -2315 17446 -1939
rect 17400 -2327 17446 -2315
rect 17518 -1939 17642 -1927
rect 17518 -2315 17524 -1939
rect 17558 -2115 17602 -1939
rect 17636 -2115 17642 -1939
rect 17558 -2127 17642 -2115
rect 17714 -1939 17760 -1927
rect 17714 -2115 17720 -1939
rect 17754 -2115 17760 -1939
rect 18679 -1943 18769 -1494
rect 18678 -2036 18688 -1943
rect 18758 -2036 18769 -1943
rect 18679 -2044 18769 -2036
rect 18906 -1572 19074 -1564
rect 18906 -1640 19015 -1572
rect 19072 -1640 19082 -1572
rect 18906 -1648 19074 -1640
rect 17714 -2127 17760 -2115
rect 17558 -2315 17564 -2127
rect 17518 -2327 17564 -2315
rect 17288 -2400 17322 -2327
rect 17273 -2416 17339 -2400
rect 17273 -2450 17289 -2416
rect 17323 -2450 17339 -2416
rect 17273 -2466 17339 -2450
rect 17602 -2494 17636 -2127
rect 16978 -2546 17636 -2494
rect 17276 -2568 17368 -2546
rect 17276 -2620 17288 -2568
rect 17354 -2620 17368 -2568
rect 17276 -2624 17368 -2620
rect 0 -2900 2994 -2840
rect 3143 -2900 6137 -2839
rect 1488 -3142 1498 -3082
rect 1578 -3142 1588 -3082
rect 1488 -3182 1588 -3142
rect 691 -3239 2494 -3182
rect 691 -3326 725 -3239
rect 1866 -3326 1900 -3239
rect 685 -3338 731 -3326
rect 685 -3526 691 -3338
rect 244 -3538 290 -3526
rect 244 -3714 250 -3538
rect 284 -3714 290 -3538
rect 244 -3726 290 -3714
rect 362 -3538 408 -3526
rect 362 -3714 368 -3538
rect 402 -3714 408 -3538
rect 362 -3726 408 -3714
rect 480 -3538 526 -3526
rect 480 -3714 486 -3538
rect 520 -3714 526 -3538
rect 480 -3726 526 -3714
rect 598 -3538 691 -3526
rect 598 -3714 604 -3538
rect 638 -3714 691 -3538
rect 725 -3714 731 -3338
rect 598 -3726 731 -3714
rect 803 -3338 849 -3326
rect 803 -3714 809 -3338
rect 843 -3714 849 -3338
rect 803 -3726 849 -3714
rect 921 -3338 967 -3326
rect 921 -3714 927 -3338
rect 961 -3714 967 -3338
rect 921 -3726 967 -3714
rect 1039 -3338 1085 -3326
rect 1039 -3714 1045 -3338
rect 1079 -3714 1085 -3338
rect 1039 -3726 1085 -3714
rect 1152 -3338 1198 -3326
rect 1152 -3714 1158 -3338
rect 1192 -3714 1198 -3338
rect 1152 -3726 1198 -3714
rect 1270 -3338 1316 -3326
rect 1270 -3714 1276 -3338
rect 1310 -3714 1316 -3338
rect 1270 -3726 1316 -3714
rect 1388 -3338 1434 -3326
rect 1388 -3714 1394 -3338
rect 1428 -3714 1434 -3338
rect 1388 -3726 1434 -3714
rect 1506 -3338 1552 -3326
rect 1506 -3714 1512 -3338
rect 1546 -3714 1552 -3338
rect 1506 -3726 1552 -3714
rect 1624 -3338 1670 -3326
rect 1624 -3714 1630 -3338
rect 1664 -3714 1670 -3338
rect 1624 -3726 1670 -3714
rect 1742 -3338 1788 -3326
rect 1742 -3714 1748 -3338
rect 1782 -3714 1788 -3338
rect 1742 -3726 1788 -3714
rect 1860 -3338 1906 -3326
rect 1860 -3714 1866 -3338
rect 1900 -3714 1906 -3338
rect 1860 -3726 1906 -3714
rect 1979 -3338 2025 -3326
rect 1979 -3714 1985 -3338
rect 2019 -3714 2025 -3338
rect 1979 -3726 2025 -3714
rect 2097 -3338 2143 -3326
rect 2097 -3714 2103 -3338
rect 2137 -3714 2143 -3338
rect 2097 -3726 2143 -3714
rect 2215 -3338 2261 -3326
rect 2215 -3714 2221 -3338
rect 2255 -3714 2261 -3338
rect 2215 -3726 2261 -3714
rect 2333 -3338 2379 -3326
rect 2333 -3714 2339 -3338
rect 2373 -3714 2379 -3338
rect 2457 -3526 2494 -3239
rect 2333 -3726 2379 -3714
rect 2452 -3538 2498 -3526
rect 2452 -3714 2458 -3538
rect 2492 -3714 2498 -3538
rect 2452 -3726 2498 -3714
rect 2570 -3538 2616 -3526
rect 2570 -3714 2576 -3538
rect 2610 -3714 2616 -3538
rect 2570 -3726 2616 -3714
rect 2688 -3538 2734 -3526
rect 2688 -3714 2694 -3538
rect 2728 -3714 2734 -3538
rect 2688 -3726 2734 -3714
rect 2806 -3538 2852 -3526
rect 2806 -3714 2812 -3538
rect 2846 -3714 2852 -3538
rect 2806 -3726 2852 -3714
rect 249 -3912 284 -3726
rect 1158 -3810 1192 -3726
rect 2339 -3810 2373 -3726
rect 1158 -3852 2373 -3810
rect 2339 -3872 2373 -3852
rect 2339 -3888 2696 -3872
rect 249 -3929 1386 -3912
rect 249 -3963 1336 -3929
rect 1370 -3963 1386 -3929
rect 2339 -3922 2646 -3888
rect 2680 -3922 2696 -3888
rect 2339 -3938 2696 -3922
rect 249 -3979 1386 -3963
rect -519 -4024 166 -4016
rect -519 -4092 107 -4024
rect 164 -4092 174 -4024
rect -519 -4100 166 -4092
rect 91 -4140 166 -4132
rect 91 -4208 107 -4140
rect 164 -4208 174 -4140
rect 91 -4216 166 -4208
rect 32 -4308 166 -4300
rect 32 -4376 107 -4308
rect 164 -4376 174 -4308
rect 32 -4384 166 -4376
rect 32 -5815 96 -4384
rect 249 -4489 284 -3979
rect 339 -4025 431 -4012
rect 339 -4088 351 -4025
rect 422 -4088 431 -4025
rect 339 -4097 431 -4088
rect 1424 -4025 1516 -4015
rect 1424 -4087 1436 -4025
rect 1506 -4087 1516 -4025
rect 1424 -4100 1516 -4087
rect 2812 -4080 2847 -3726
rect 2922 -4080 2994 -2900
rect 4632 -3142 4642 -3082
rect 4722 -3142 4732 -3082
rect 4632 -3182 4732 -3142
rect 3835 -3239 5638 -3182
rect 3835 -3326 3869 -3239
rect 5010 -3326 5044 -3239
rect 3829 -3338 3875 -3326
rect 3829 -3526 3835 -3338
rect 3388 -3538 3434 -3526
rect 3388 -3714 3394 -3538
rect 3428 -3714 3434 -3538
rect 3388 -3726 3434 -3714
rect 3506 -3538 3552 -3526
rect 3506 -3714 3512 -3538
rect 3546 -3714 3552 -3538
rect 3506 -3726 3552 -3714
rect 3624 -3538 3670 -3526
rect 3624 -3714 3630 -3538
rect 3664 -3714 3670 -3538
rect 3624 -3726 3670 -3714
rect 3742 -3538 3835 -3526
rect 3742 -3714 3748 -3538
rect 3782 -3714 3835 -3538
rect 3869 -3714 3875 -3338
rect 3742 -3726 3875 -3714
rect 3947 -3338 3993 -3326
rect 3947 -3714 3953 -3338
rect 3987 -3714 3993 -3338
rect 3947 -3726 3993 -3714
rect 4065 -3338 4111 -3326
rect 4065 -3714 4071 -3338
rect 4105 -3714 4111 -3338
rect 4065 -3726 4111 -3714
rect 4183 -3338 4229 -3326
rect 4183 -3714 4189 -3338
rect 4223 -3714 4229 -3338
rect 4183 -3726 4229 -3714
rect 4296 -3338 4342 -3326
rect 4296 -3714 4302 -3338
rect 4336 -3714 4342 -3338
rect 4296 -3726 4342 -3714
rect 4414 -3338 4460 -3326
rect 4414 -3714 4420 -3338
rect 4454 -3714 4460 -3338
rect 4414 -3726 4460 -3714
rect 4532 -3338 4578 -3326
rect 4532 -3714 4538 -3338
rect 4572 -3714 4578 -3338
rect 4532 -3726 4578 -3714
rect 4650 -3338 4696 -3326
rect 4650 -3714 4656 -3338
rect 4690 -3714 4696 -3338
rect 4650 -3726 4696 -3714
rect 4768 -3338 4814 -3326
rect 4768 -3714 4774 -3338
rect 4808 -3714 4814 -3338
rect 4768 -3726 4814 -3714
rect 4886 -3338 4932 -3326
rect 4886 -3714 4892 -3338
rect 4926 -3714 4932 -3338
rect 4886 -3726 4932 -3714
rect 5004 -3338 5050 -3326
rect 5004 -3714 5010 -3338
rect 5044 -3714 5050 -3338
rect 5004 -3726 5050 -3714
rect 5123 -3338 5169 -3326
rect 5123 -3714 5129 -3338
rect 5163 -3714 5169 -3338
rect 5123 -3726 5169 -3714
rect 5241 -3338 5287 -3326
rect 5241 -3714 5247 -3338
rect 5281 -3714 5287 -3338
rect 5241 -3726 5287 -3714
rect 5359 -3338 5405 -3326
rect 5359 -3714 5365 -3338
rect 5399 -3714 5405 -3338
rect 5359 -3726 5405 -3714
rect 5477 -3338 5523 -3326
rect 5477 -3714 5483 -3338
rect 5517 -3714 5523 -3338
rect 5601 -3526 5638 -3239
rect 5477 -3726 5523 -3714
rect 5596 -3538 5642 -3526
rect 5596 -3714 5602 -3538
rect 5636 -3714 5642 -3538
rect 5596 -3726 5642 -3714
rect 5714 -3538 5760 -3526
rect 5714 -3714 5720 -3538
rect 5754 -3714 5760 -3538
rect 5714 -3726 5760 -3714
rect 5832 -3538 5878 -3526
rect 5832 -3714 5838 -3538
rect 5872 -3714 5878 -3538
rect 5832 -3726 5878 -3714
rect 5950 -3538 5996 -3526
rect 5950 -3714 5956 -3538
rect 5990 -3714 5996 -3538
rect 5950 -3726 5996 -3714
rect 3393 -3912 3428 -3726
rect 4302 -3810 4336 -3726
rect 5483 -3810 5517 -3726
rect 4302 -3852 5517 -3810
rect 5483 -3872 5517 -3852
rect 5483 -3888 5840 -3872
rect 3393 -3929 4530 -3912
rect 3393 -3963 4480 -3929
rect 4514 -3963 4530 -3929
rect 5483 -3922 5790 -3888
rect 5824 -3922 5840 -3888
rect 5483 -3938 5840 -3922
rect 3393 -3979 4530 -3963
rect 2812 -4088 2994 -4080
rect 3134 -4024 3310 -4016
rect 1671 -4142 1736 -4139
rect 1671 -4145 1740 -4142
rect 1671 -4205 1677 -4145
rect 1736 -4205 1746 -4145
rect 1671 -4209 1740 -4205
rect 1671 -4211 1736 -4209
rect 2812 -4226 2993 -4088
rect 3134 -4092 3251 -4024
rect 3308 -4092 3318 -4024
rect 3134 -4100 3310 -4092
rect 3239 -4140 3310 -4132
rect 3239 -4208 3251 -4140
rect 3308 -4208 3318 -4140
rect 3239 -4216 3310 -4208
rect 1306 -4308 1398 -4300
rect 1306 -4373 1318 -4308
rect 1386 -4373 1398 -4308
rect 1306 -4385 1398 -4373
rect 2812 -4488 2847 -4226
rect 249 -4536 1621 -4489
rect 1943 -4535 2847 -4488
rect 3176 -4308 3310 -4300
rect 3176 -4376 3251 -4308
rect 3308 -4376 3318 -4308
rect 3176 -4384 3310 -4376
rect 1083 -4659 1117 -4536
rect 1555 -4549 1621 -4536
rect 1555 -4583 1571 -4549
rect 1605 -4583 1621 -4549
rect 1555 -4599 1621 -4583
rect 1944 -4659 1978 -4535
rect 1078 -4671 1124 -4659
rect 1078 -4847 1084 -4671
rect 1118 -4847 1124 -4671
rect 1078 -4859 1124 -4847
rect 1196 -4671 1316 -4659
rect 1196 -4847 1202 -4671
rect 1236 -4847 1276 -4671
rect 1196 -4859 1276 -4847
rect 1202 -5226 1236 -4859
rect 1270 -5047 1276 -4859
rect 1310 -5047 1316 -4671
rect 1270 -5059 1316 -5047
rect 1388 -4671 1434 -4659
rect 1388 -5047 1394 -4671
rect 1428 -5047 1434 -4671
rect 1388 -5059 1434 -5047
rect 1506 -4671 1552 -4659
rect 1506 -5047 1512 -4671
rect 1546 -5047 1552 -4671
rect 1506 -5059 1552 -5047
rect 1624 -4671 1670 -4659
rect 1624 -5047 1630 -4671
rect 1664 -5047 1670 -4671
rect 1624 -5059 1670 -5047
rect 1742 -4671 1866 -4659
rect 1742 -5047 1748 -4671
rect 1782 -4847 1826 -4671
rect 1860 -4847 1866 -4671
rect 1782 -4859 1866 -4847
rect 1938 -4671 1984 -4659
rect 1938 -4847 1944 -4671
rect 1978 -4847 1984 -4671
rect 1938 -4859 1984 -4847
rect 1782 -5047 1788 -4859
rect 1742 -5059 1788 -5047
rect 1512 -5132 1546 -5059
rect 1497 -5148 1563 -5132
rect 1497 -5182 1513 -5148
rect 1547 -5182 1563 -5148
rect 1497 -5198 1563 -5182
rect 1826 -5226 1860 -4859
rect 1202 -5278 1860 -5226
rect 1500 -5300 1592 -5278
rect 1500 -5352 1512 -5300
rect 1578 -5352 1592 -5300
rect 1500 -5356 1592 -5352
rect 3176 -5706 3240 -4384
rect 3393 -4489 3428 -3979
rect 3483 -4025 3575 -4012
rect 3483 -4088 3495 -4025
rect 3566 -4088 3575 -4025
rect 3483 -4097 3575 -4088
rect 4568 -4025 4660 -4015
rect 4568 -4087 4580 -4025
rect 4650 -4087 4660 -4025
rect 4568 -4100 4660 -4087
rect 5956 -4080 5991 -3726
rect 6066 -4080 6137 -2900
rect 6293 -2900 9269 -2839
rect 9444 -2900 12414 -2839
rect 12622 -2899 15474 -2838
rect 15790 -2899 18759 -2838
rect 6293 -2902 6342 -2900
rect 7764 -3138 7774 -3078
rect 7854 -3138 7864 -3078
rect 7764 -3178 7864 -3138
rect 6967 -3235 8770 -3178
rect 6967 -3322 7001 -3235
rect 8142 -3322 8176 -3235
rect 6961 -3334 7007 -3322
rect 6961 -3522 6967 -3334
rect 6520 -3534 6566 -3522
rect 6520 -3710 6526 -3534
rect 6560 -3710 6566 -3534
rect 6520 -3722 6566 -3710
rect 6638 -3534 6684 -3522
rect 6638 -3710 6644 -3534
rect 6678 -3710 6684 -3534
rect 6638 -3722 6684 -3710
rect 6756 -3534 6802 -3522
rect 6756 -3710 6762 -3534
rect 6796 -3710 6802 -3534
rect 6756 -3722 6802 -3710
rect 6874 -3534 6967 -3522
rect 6874 -3710 6880 -3534
rect 6914 -3710 6967 -3534
rect 7001 -3710 7007 -3334
rect 6874 -3722 7007 -3710
rect 7079 -3334 7125 -3322
rect 7079 -3710 7085 -3334
rect 7119 -3710 7125 -3334
rect 7079 -3722 7125 -3710
rect 7197 -3334 7243 -3322
rect 7197 -3710 7203 -3334
rect 7237 -3710 7243 -3334
rect 7197 -3722 7243 -3710
rect 7315 -3334 7361 -3322
rect 7315 -3710 7321 -3334
rect 7355 -3710 7361 -3334
rect 7315 -3722 7361 -3710
rect 7428 -3334 7474 -3322
rect 7428 -3710 7434 -3334
rect 7468 -3710 7474 -3334
rect 7428 -3722 7474 -3710
rect 7546 -3334 7592 -3322
rect 7546 -3710 7552 -3334
rect 7586 -3710 7592 -3334
rect 7546 -3722 7592 -3710
rect 7664 -3334 7710 -3322
rect 7664 -3710 7670 -3334
rect 7704 -3710 7710 -3334
rect 7664 -3722 7710 -3710
rect 7782 -3334 7828 -3322
rect 7782 -3710 7788 -3334
rect 7822 -3710 7828 -3334
rect 7782 -3722 7828 -3710
rect 7900 -3334 7946 -3322
rect 7900 -3710 7906 -3334
rect 7940 -3710 7946 -3334
rect 7900 -3722 7946 -3710
rect 8018 -3334 8064 -3322
rect 8018 -3710 8024 -3334
rect 8058 -3710 8064 -3334
rect 8018 -3722 8064 -3710
rect 8136 -3334 8182 -3322
rect 8136 -3710 8142 -3334
rect 8176 -3710 8182 -3334
rect 8136 -3722 8182 -3710
rect 8255 -3334 8301 -3322
rect 8255 -3710 8261 -3334
rect 8295 -3710 8301 -3334
rect 8255 -3722 8301 -3710
rect 8373 -3334 8419 -3322
rect 8373 -3710 8379 -3334
rect 8413 -3710 8419 -3334
rect 8373 -3722 8419 -3710
rect 8491 -3334 8537 -3322
rect 8491 -3710 8497 -3334
rect 8531 -3710 8537 -3334
rect 8491 -3722 8537 -3710
rect 8609 -3334 8655 -3322
rect 8609 -3710 8615 -3334
rect 8649 -3710 8655 -3334
rect 8733 -3522 8770 -3235
rect 8609 -3722 8655 -3710
rect 8728 -3534 8774 -3522
rect 8728 -3710 8734 -3534
rect 8768 -3710 8774 -3534
rect 8728 -3722 8774 -3710
rect 8846 -3534 8892 -3522
rect 8846 -3710 8852 -3534
rect 8886 -3710 8892 -3534
rect 8846 -3722 8892 -3710
rect 8964 -3534 9010 -3522
rect 8964 -3710 8970 -3534
rect 9004 -3710 9010 -3534
rect 8964 -3722 9010 -3710
rect 9082 -3534 9128 -3522
rect 9082 -3710 9088 -3534
rect 9122 -3710 9128 -3534
rect 9082 -3722 9128 -3710
rect 6525 -3908 6560 -3722
rect 7434 -3806 7468 -3722
rect 8615 -3806 8649 -3722
rect 7434 -3848 8649 -3806
rect 8615 -3868 8649 -3848
rect 8615 -3884 8972 -3868
rect 6525 -3925 7662 -3908
rect 6525 -3959 7612 -3925
rect 7646 -3959 7662 -3925
rect 8615 -3918 8922 -3884
rect 8956 -3918 8972 -3884
rect 8615 -3934 8972 -3918
rect 6525 -3975 7662 -3959
rect 4815 -4142 4880 -4139
rect 4815 -4145 4884 -4142
rect 4815 -4205 4821 -4145
rect 4880 -4205 4890 -4145
rect 4815 -4209 4884 -4205
rect 4815 -4211 4880 -4209
rect 5956 -4226 6137 -4080
rect 6266 -4020 6442 -4012
rect 6266 -4088 6383 -4020
rect 6440 -4088 6450 -4020
rect 6266 -4096 6442 -4088
rect 6371 -4136 6442 -4128
rect 6371 -4204 6383 -4136
rect 6440 -4204 6450 -4136
rect 6371 -4212 6442 -4204
rect 4450 -4308 4542 -4300
rect 4450 -4373 4462 -4308
rect 4530 -4373 4542 -4308
rect 4450 -4385 4542 -4373
rect 5956 -4488 5991 -4226
rect 6266 -4304 6442 -4296
rect 6266 -4372 6383 -4304
rect 6440 -4372 6450 -4304
rect 6266 -4380 6442 -4372
rect 3393 -4536 4765 -4489
rect 5087 -4535 5991 -4488
rect 4227 -4659 4261 -4536
rect 4699 -4549 4765 -4536
rect 4699 -4583 4715 -4549
rect 4749 -4583 4765 -4549
rect 4699 -4599 4765 -4583
rect 5088 -4659 5122 -4535
rect 4222 -4671 4268 -4659
rect 4222 -4847 4228 -4671
rect 4262 -4847 4268 -4671
rect 4222 -4859 4268 -4847
rect 4340 -4671 4460 -4659
rect 4340 -4847 4346 -4671
rect 4380 -4847 4420 -4671
rect 4340 -4859 4420 -4847
rect 4346 -5226 4380 -4859
rect 4414 -5047 4420 -4859
rect 4454 -5047 4460 -4671
rect 4414 -5059 4460 -5047
rect 4532 -4671 4578 -4659
rect 4532 -5047 4538 -4671
rect 4572 -5047 4578 -4671
rect 4532 -5059 4578 -5047
rect 4650 -4671 4696 -4659
rect 4650 -5047 4656 -4671
rect 4690 -5047 4696 -4671
rect 4650 -5059 4696 -5047
rect 4768 -4671 4814 -4659
rect 4768 -5047 4774 -4671
rect 4808 -5047 4814 -4671
rect 4768 -5059 4814 -5047
rect 4886 -4671 5010 -4659
rect 4886 -5047 4892 -4671
rect 4926 -4847 4970 -4671
rect 5004 -4847 5010 -4671
rect 4926 -4859 5010 -4847
rect 5082 -4671 5128 -4659
rect 5082 -4847 5088 -4671
rect 5122 -4847 5128 -4671
rect 5082 -4859 5128 -4847
rect 4926 -5047 4932 -4859
rect 4886 -5059 4932 -5047
rect 4656 -5132 4690 -5059
rect 4641 -5148 4707 -5132
rect 4641 -5182 4657 -5148
rect 4691 -5182 4707 -5148
rect 4641 -5198 4707 -5182
rect 4970 -5226 5004 -4859
rect 4346 -5278 5004 -5226
rect 4644 -5300 4736 -5278
rect 4644 -5352 4656 -5300
rect 4722 -5352 4736 -5300
rect 4644 -5356 4736 -5352
rect 6308 -5470 6371 -4380
rect 6525 -4485 6560 -3975
rect 6615 -4021 6707 -4008
rect 6615 -4084 6627 -4021
rect 6698 -4084 6707 -4021
rect 6615 -4093 6707 -4084
rect 7700 -4021 7792 -4011
rect 7700 -4083 7712 -4021
rect 7782 -4083 7792 -4021
rect 7700 -4096 7792 -4083
rect 9088 -4076 9123 -3722
rect 9198 -4076 9269 -2900
rect 10908 -3138 10918 -3078
rect 10998 -3138 11008 -3078
rect 10908 -3178 11008 -3138
rect 10111 -3235 11914 -3178
rect 10111 -3322 10145 -3235
rect 11286 -3322 11320 -3235
rect 10105 -3334 10151 -3322
rect 10105 -3522 10111 -3334
rect 9664 -3534 9710 -3522
rect 9664 -3710 9670 -3534
rect 9704 -3710 9710 -3534
rect 9664 -3722 9710 -3710
rect 9782 -3534 9828 -3522
rect 9782 -3710 9788 -3534
rect 9822 -3710 9828 -3534
rect 9782 -3722 9828 -3710
rect 9900 -3534 9946 -3522
rect 9900 -3710 9906 -3534
rect 9940 -3710 9946 -3534
rect 9900 -3722 9946 -3710
rect 10018 -3534 10111 -3522
rect 10018 -3710 10024 -3534
rect 10058 -3710 10111 -3534
rect 10145 -3710 10151 -3334
rect 10018 -3722 10151 -3710
rect 10223 -3334 10269 -3322
rect 10223 -3710 10229 -3334
rect 10263 -3710 10269 -3334
rect 10223 -3722 10269 -3710
rect 10341 -3334 10387 -3322
rect 10341 -3710 10347 -3334
rect 10381 -3710 10387 -3334
rect 10341 -3722 10387 -3710
rect 10459 -3334 10505 -3322
rect 10459 -3710 10465 -3334
rect 10499 -3710 10505 -3334
rect 10459 -3722 10505 -3710
rect 10572 -3334 10618 -3322
rect 10572 -3710 10578 -3334
rect 10612 -3710 10618 -3334
rect 10572 -3722 10618 -3710
rect 10690 -3334 10736 -3322
rect 10690 -3710 10696 -3334
rect 10730 -3710 10736 -3334
rect 10690 -3722 10736 -3710
rect 10808 -3334 10854 -3322
rect 10808 -3710 10814 -3334
rect 10848 -3710 10854 -3334
rect 10808 -3722 10854 -3710
rect 10926 -3334 10972 -3322
rect 10926 -3710 10932 -3334
rect 10966 -3710 10972 -3334
rect 10926 -3722 10972 -3710
rect 11044 -3334 11090 -3322
rect 11044 -3710 11050 -3334
rect 11084 -3710 11090 -3334
rect 11044 -3722 11090 -3710
rect 11162 -3334 11208 -3322
rect 11162 -3710 11168 -3334
rect 11202 -3710 11208 -3334
rect 11162 -3722 11208 -3710
rect 11280 -3334 11326 -3322
rect 11280 -3710 11286 -3334
rect 11320 -3710 11326 -3334
rect 11280 -3722 11326 -3710
rect 11399 -3334 11445 -3322
rect 11399 -3710 11405 -3334
rect 11439 -3710 11445 -3334
rect 11399 -3722 11445 -3710
rect 11517 -3334 11563 -3322
rect 11517 -3710 11523 -3334
rect 11557 -3710 11563 -3334
rect 11517 -3722 11563 -3710
rect 11635 -3334 11681 -3322
rect 11635 -3710 11641 -3334
rect 11675 -3710 11681 -3334
rect 11635 -3722 11681 -3710
rect 11753 -3334 11799 -3322
rect 11753 -3710 11759 -3334
rect 11793 -3710 11799 -3334
rect 11877 -3522 11914 -3235
rect 11753 -3722 11799 -3710
rect 11872 -3534 11918 -3522
rect 11872 -3710 11878 -3534
rect 11912 -3710 11918 -3534
rect 11872 -3722 11918 -3710
rect 11990 -3534 12036 -3522
rect 11990 -3710 11996 -3534
rect 12030 -3710 12036 -3534
rect 11990 -3722 12036 -3710
rect 12108 -3534 12154 -3522
rect 12108 -3710 12114 -3534
rect 12148 -3710 12154 -3534
rect 12108 -3722 12154 -3710
rect 12226 -3534 12272 -3522
rect 12226 -3710 12232 -3534
rect 12266 -3710 12272 -3534
rect 12226 -3722 12272 -3710
rect 9669 -3908 9704 -3722
rect 10578 -3806 10612 -3722
rect 11759 -3806 11793 -3722
rect 10578 -3848 11793 -3806
rect 11759 -3868 11793 -3848
rect 11759 -3884 12116 -3868
rect 9669 -3925 10806 -3908
rect 9669 -3959 10756 -3925
rect 10790 -3959 10806 -3925
rect 11759 -3918 12066 -3884
rect 12100 -3918 12116 -3884
rect 11759 -3934 12116 -3918
rect 9669 -3975 10806 -3959
rect 7947 -4138 8012 -4135
rect 7947 -4141 8016 -4138
rect 7947 -4201 7953 -4141
rect 8012 -4201 8022 -4141
rect 7947 -4205 8016 -4201
rect 7947 -4207 8012 -4205
rect 9088 -4214 9269 -4076
rect 9410 -4020 9586 -4012
rect 9410 -4088 9527 -4020
rect 9584 -4088 9594 -4020
rect 9410 -4096 9586 -4088
rect 9516 -4136 9586 -4128
rect 9516 -4204 9527 -4136
rect 9584 -4204 9594 -4136
rect 9516 -4212 9586 -4204
rect 7582 -4304 7674 -4296
rect 7582 -4369 7594 -4304
rect 7662 -4369 7674 -4304
rect 7582 -4381 7674 -4369
rect 9088 -4484 9123 -4214
rect 6525 -4532 7897 -4485
rect 8219 -4531 9123 -4484
rect 9468 -4304 9586 -4296
rect 9468 -4372 9527 -4304
rect 9584 -4372 9594 -4304
rect 9468 -4380 9586 -4372
rect 7359 -4655 7393 -4532
rect 7831 -4545 7897 -4532
rect 7831 -4579 7847 -4545
rect 7881 -4579 7897 -4545
rect 7831 -4595 7897 -4579
rect 8220 -4655 8254 -4531
rect 7354 -4667 7400 -4655
rect 7354 -4843 7360 -4667
rect 7394 -4843 7400 -4667
rect 7354 -4855 7400 -4843
rect 7472 -4667 7592 -4655
rect 7472 -4843 7478 -4667
rect 7512 -4843 7552 -4667
rect 7472 -4855 7552 -4843
rect 7478 -5222 7512 -4855
rect 7546 -5043 7552 -4855
rect 7586 -5043 7592 -4667
rect 7546 -5055 7592 -5043
rect 7664 -4667 7710 -4655
rect 7664 -5043 7670 -4667
rect 7704 -5043 7710 -4667
rect 7664 -5055 7710 -5043
rect 7782 -4667 7828 -4655
rect 7782 -5043 7788 -4667
rect 7822 -5043 7828 -4667
rect 7782 -5055 7828 -5043
rect 7900 -4667 7946 -4655
rect 7900 -5043 7906 -4667
rect 7940 -5043 7946 -4667
rect 7900 -5055 7946 -5043
rect 8018 -4667 8142 -4655
rect 8018 -5043 8024 -4667
rect 8058 -4843 8102 -4667
rect 8136 -4843 8142 -4667
rect 8058 -4855 8142 -4843
rect 8214 -4667 8260 -4655
rect 8214 -4843 8220 -4667
rect 8254 -4843 8260 -4667
rect 8214 -4855 8260 -4843
rect 8058 -5043 8064 -4855
rect 8018 -5055 8064 -5043
rect 7788 -5128 7822 -5055
rect 7773 -5144 7839 -5128
rect 7773 -5178 7789 -5144
rect 7823 -5178 7839 -5144
rect 7773 -5194 7839 -5178
rect 8102 -5222 8136 -4855
rect 7478 -5274 8136 -5222
rect 7776 -5296 7868 -5274
rect 7776 -5348 7788 -5296
rect 7854 -5348 7868 -5296
rect 7776 -5352 7868 -5348
rect 9468 -5394 9516 -4380
rect 9669 -4485 9704 -3975
rect 9759 -4021 9851 -4008
rect 9759 -4084 9771 -4021
rect 9842 -4084 9851 -4021
rect 9759 -4093 9851 -4084
rect 10844 -4021 10936 -4011
rect 10844 -4083 10856 -4021
rect 10926 -4083 10936 -4021
rect 10844 -4096 10936 -4083
rect 12232 -4076 12267 -3722
rect 12343 -4076 12414 -2900
rect 14110 -3142 14120 -3082
rect 14200 -3142 14210 -3082
rect 14110 -3182 14210 -3142
rect 13313 -3239 15116 -3182
rect 13313 -3326 13347 -3239
rect 14488 -3326 14522 -3239
rect 13307 -3338 13353 -3326
rect 13307 -3526 13313 -3338
rect 12866 -3538 12912 -3526
rect 12866 -3714 12872 -3538
rect 12906 -3714 12912 -3538
rect 12866 -3726 12912 -3714
rect 12984 -3538 13030 -3526
rect 12984 -3714 12990 -3538
rect 13024 -3714 13030 -3538
rect 12984 -3726 13030 -3714
rect 13102 -3538 13148 -3526
rect 13102 -3714 13108 -3538
rect 13142 -3714 13148 -3538
rect 13102 -3726 13148 -3714
rect 13220 -3538 13313 -3526
rect 13220 -3714 13226 -3538
rect 13260 -3714 13313 -3538
rect 13347 -3714 13353 -3338
rect 13220 -3726 13353 -3714
rect 13425 -3338 13471 -3326
rect 13425 -3714 13431 -3338
rect 13465 -3714 13471 -3338
rect 13425 -3726 13471 -3714
rect 13543 -3338 13589 -3326
rect 13543 -3714 13549 -3338
rect 13583 -3714 13589 -3338
rect 13543 -3726 13589 -3714
rect 13661 -3338 13707 -3326
rect 13661 -3714 13667 -3338
rect 13701 -3714 13707 -3338
rect 13661 -3726 13707 -3714
rect 13774 -3338 13820 -3326
rect 13774 -3714 13780 -3338
rect 13814 -3714 13820 -3338
rect 13774 -3726 13820 -3714
rect 13892 -3338 13938 -3326
rect 13892 -3714 13898 -3338
rect 13932 -3714 13938 -3338
rect 13892 -3726 13938 -3714
rect 14010 -3338 14056 -3326
rect 14010 -3714 14016 -3338
rect 14050 -3714 14056 -3338
rect 14010 -3726 14056 -3714
rect 14128 -3338 14174 -3326
rect 14128 -3714 14134 -3338
rect 14168 -3714 14174 -3338
rect 14128 -3726 14174 -3714
rect 14246 -3338 14292 -3326
rect 14246 -3714 14252 -3338
rect 14286 -3714 14292 -3338
rect 14246 -3726 14292 -3714
rect 14364 -3338 14410 -3326
rect 14364 -3714 14370 -3338
rect 14404 -3714 14410 -3338
rect 14364 -3726 14410 -3714
rect 14482 -3338 14528 -3326
rect 14482 -3714 14488 -3338
rect 14522 -3714 14528 -3338
rect 14482 -3726 14528 -3714
rect 14601 -3338 14647 -3326
rect 14601 -3714 14607 -3338
rect 14641 -3714 14647 -3338
rect 14601 -3726 14647 -3714
rect 14719 -3338 14765 -3326
rect 14719 -3714 14725 -3338
rect 14759 -3714 14765 -3338
rect 14719 -3726 14765 -3714
rect 14837 -3338 14883 -3326
rect 14837 -3714 14843 -3338
rect 14877 -3714 14883 -3338
rect 14837 -3726 14883 -3714
rect 14955 -3338 15001 -3326
rect 14955 -3714 14961 -3338
rect 14995 -3714 15001 -3338
rect 15079 -3526 15116 -3239
rect 14955 -3726 15001 -3714
rect 15074 -3538 15120 -3526
rect 15074 -3714 15080 -3538
rect 15114 -3714 15120 -3538
rect 15074 -3726 15120 -3714
rect 15192 -3538 15238 -3526
rect 15192 -3714 15198 -3538
rect 15232 -3714 15238 -3538
rect 15192 -3726 15238 -3714
rect 15310 -3538 15356 -3526
rect 15310 -3714 15316 -3538
rect 15350 -3714 15356 -3538
rect 15310 -3726 15356 -3714
rect 15428 -3538 15474 -2899
rect 17254 -3142 17264 -3082
rect 17344 -3142 17354 -3082
rect 17254 -3182 17354 -3142
rect 16457 -3239 18260 -3182
rect 16457 -3326 16491 -3239
rect 17632 -3326 17666 -3239
rect 16451 -3338 16497 -3326
rect 16451 -3526 16457 -3338
rect 15428 -3714 15434 -3538
rect 15468 -3714 15474 -3538
rect 15428 -3726 15474 -3714
rect 16010 -3538 16056 -3526
rect 16010 -3714 16016 -3538
rect 16050 -3714 16056 -3538
rect 16010 -3726 16056 -3714
rect 16128 -3538 16174 -3526
rect 16128 -3714 16134 -3538
rect 16168 -3714 16174 -3538
rect 16128 -3726 16174 -3714
rect 16246 -3538 16292 -3526
rect 16246 -3714 16252 -3538
rect 16286 -3714 16292 -3538
rect 16246 -3726 16292 -3714
rect 16364 -3538 16457 -3526
rect 16364 -3714 16370 -3538
rect 16404 -3714 16457 -3538
rect 16491 -3714 16497 -3338
rect 16364 -3726 16497 -3714
rect 16569 -3338 16615 -3326
rect 16569 -3714 16575 -3338
rect 16609 -3714 16615 -3338
rect 16569 -3726 16615 -3714
rect 16687 -3338 16733 -3326
rect 16687 -3714 16693 -3338
rect 16727 -3714 16733 -3338
rect 16687 -3726 16733 -3714
rect 16805 -3338 16851 -3326
rect 16805 -3714 16811 -3338
rect 16845 -3714 16851 -3338
rect 16805 -3726 16851 -3714
rect 16918 -3338 16964 -3326
rect 16918 -3714 16924 -3338
rect 16958 -3714 16964 -3338
rect 16918 -3726 16964 -3714
rect 17036 -3338 17082 -3326
rect 17036 -3714 17042 -3338
rect 17076 -3714 17082 -3338
rect 17036 -3726 17082 -3714
rect 17154 -3338 17200 -3326
rect 17154 -3714 17160 -3338
rect 17194 -3714 17200 -3338
rect 17154 -3726 17200 -3714
rect 17272 -3338 17318 -3326
rect 17272 -3714 17278 -3338
rect 17312 -3714 17318 -3338
rect 17272 -3726 17318 -3714
rect 17390 -3338 17436 -3326
rect 17390 -3714 17396 -3338
rect 17430 -3714 17436 -3338
rect 17390 -3726 17436 -3714
rect 17508 -3338 17554 -3326
rect 17508 -3714 17514 -3338
rect 17548 -3714 17554 -3338
rect 17508 -3726 17554 -3714
rect 17626 -3338 17672 -3326
rect 17626 -3714 17632 -3338
rect 17666 -3714 17672 -3338
rect 17626 -3726 17672 -3714
rect 17745 -3338 17791 -3326
rect 17745 -3714 17751 -3338
rect 17785 -3714 17791 -3338
rect 17745 -3726 17791 -3714
rect 17863 -3338 17909 -3326
rect 17863 -3714 17869 -3338
rect 17903 -3714 17909 -3338
rect 17863 -3726 17909 -3714
rect 17981 -3338 18027 -3326
rect 17981 -3714 17987 -3338
rect 18021 -3714 18027 -3338
rect 17981 -3726 18027 -3714
rect 18099 -3338 18145 -3326
rect 18099 -3714 18105 -3338
rect 18139 -3714 18145 -3338
rect 18223 -3526 18260 -3239
rect 18099 -3726 18145 -3714
rect 18218 -3538 18264 -3526
rect 18218 -3714 18224 -3538
rect 18258 -3714 18264 -3538
rect 18218 -3726 18264 -3714
rect 18336 -3538 18382 -3526
rect 18336 -3714 18342 -3538
rect 18376 -3714 18382 -3538
rect 18336 -3726 18382 -3714
rect 18454 -3538 18500 -3526
rect 18454 -3714 18460 -3538
rect 18494 -3714 18500 -3538
rect 18454 -3726 18500 -3714
rect 18572 -3538 18618 -3526
rect 18572 -3714 18578 -3538
rect 18612 -3714 18618 -3538
rect 18572 -3726 18618 -3714
rect 12871 -3912 12906 -3726
rect 13780 -3810 13814 -3726
rect 14961 -3810 14995 -3726
rect 13780 -3852 14995 -3810
rect 14961 -3872 14995 -3852
rect 14961 -3888 15318 -3872
rect 12871 -3929 14008 -3912
rect 12871 -3963 13958 -3929
rect 13992 -3963 14008 -3929
rect 14961 -3922 15268 -3888
rect 15302 -3922 15318 -3888
rect 14961 -3938 15318 -3922
rect 12871 -3979 14008 -3963
rect 12612 -4024 12788 -4016
rect 11091 -4138 11156 -4135
rect 11091 -4141 11160 -4138
rect 11091 -4201 11097 -4141
rect 11156 -4201 11166 -4141
rect 11091 -4205 11160 -4201
rect 11091 -4207 11156 -4205
rect 12232 -4222 12413 -4076
rect 12612 -4092 12729 -4024
rect 12786 -4092 12796 -4024
rect 12612 -4100 12788 -4092
rect 12718 -4140 12788 -4132
rect 12718 -4208 12729 -4140
rect 12786 -4208 12796 -4140
rect 12718 -4216 12788 -4208
rect 10726 -4304 10818 -4296
rect 10726 -4369 10738 -4304
rect 10806 -4369 10818 -4304
rect 10726 -4381 10818 -4369
rect 12232 -4484 12267 -4222
rect 9669 -4532 11041 -4485
rect 11363 -4531 12267 -4484
rect 12672 -4308 12788 -4300
rect 12672 -4376 12729 -4308
rect 12786 -4376 12796 -4308
rect 12672 -4384 12788 -4376
rect 10503 -4655 10537 -4532
rect 10975 -4545 11041 -4532
rect 10975 -4579 10991 -4545
rect 11025 -4579 11041 -4545
rect 10975 -4595 11041 -4579
rect 11364 -4655 11398 -4531
rect 10498 -4667 10544 -4655
rect 10498 -4843 10504 -4667
rect 10538 -4843 10544 -4667
rect 10498 -4855 10544 -4843
rect 10616 -4667 10736 -4655
rect 10616 -4843 10622 -4667
rect 10656 -4843 10696 -4667
rect 10616 -4855 10696 -4843
rect 10622 -5222 10656 -4855
rect 10690 -5043 10696 -4855
rect 10730 -5043 10736 -4667
rect 10690 -5055 10736 -5043
rect 10808 -4667 10854 -4655
rect 10808 -5043 10814 -4667
rect 10848 -5043 10854 -4667
rect 10808 -5055 10854 -5043
rect 10926 -4667 10972 -4655
rect 10926 -5043 10932 -4667
rect 10966 -5043 10972 -4667
rect 10926 -5055 10972 -5043
rect 11044 -4667 11090 -4655
rect 11044 -5043 11050 -4667
rect 11084 -5043 11090 -4667
rect 11044 -5055 11090 -5043
rect 11162 -4667 11286 -4655
rect 11162 -5043 11168 -4667
rect 11202 -4843 11246 -4667
rect 11280 -4843 11286 -4667
rect 11202 -4855 11286 -4843
rect 11358 -4667 11404 -4655
rect 11358 -4843 11364 -4667
rect 11398 -4843 11404 -4667
rect 11358 -4855 11404 -4843
rect 11202 -5043 11208 -4855
rect 11162 -5055 11208 -5043
rect 10932 -5128 10966 -5055
rect 10917 -5144 10983 -5128
rect 10917 -5178 10933 -5144
rect 10967 -5178 10983 -5144
rect 10917 -5194 10983 -5178
rect 11246 -5222 11280 -4855
rect 10622 -5274 11280 -5222
rect 10920 -5296 11012 -5274
rect 10920 -5348 10932 -5296
rect 10998 -5348 11012 -5296
rect 10920 -5352 11012 -5348
rect 12672 -5391 12720 -4384
rect 12871 -4489 12906 -3979
rect 12961 -4025 13053 -4012
rect 12961 -4088 12973 -4025
rect 13044 -4088 13053 -4025
rect 12961 -4097 13053 -4088
rect 14046 -4025 14138 -4015
rect 14046 -4087 14058 -4025
rect 14128 -4087 14138 -4025
rect 14046 -4100 14138 -4087
rect 14293 -4142 14358 -4139
rect 14293 -4145 14362 -4142
rect 14293 -4205 14299 -4145
rect 14358 -4205 14368 -4145
rect 14293 -4209 14362 -4205
rect 14293 -4211 14358 -4209
rect 13928 -4308 14020 -4300
rect 13928 -4373 13940 -4308
rect 14008 -4373 14020 -4308
rect 13928 -4385 14020 -4373
rect 15434 -4488 15469 -3726
rect 16015 -3912 16050 -3726
rect 16924 -3810 16958 -3726
rect 18105 -3810 18139 -3726
rect 16924 -3852 18139 -3810
rect 18105 -3872 18139 -3852
rect 18105 -3888 18462 -3872
rect 16015 -3929 17152 -3912
rect 16015 -3963 17102 -3929
rect 17136 -3963 17152 -3929
rect 18105 -3922 18412 -3888
rect 18446 -3922 18462 -3888
rect 18105 -3938 18462 -3922
rect 16015 -3979 17152 -3963
rect 15756 -4024 15932 -4016
rect 15756 -4092 15873 -4024
rect 15930 -4092 15940 -4024
rect 15756 -4100 15932 -4092
rect 15861 -4140 15932 -4132
rect 15861 -4208 15873 -4140
rect 15930 -4208 15940 -4140
rect 15861 -4216 15932 -4208
rect 15814 -4300 15862 -4299
rect 15813 -4308 15932 -4300
rect 15813 -4376 15873 -4308
rect 15930 -4376 15940 -4308
rect 15813 -4384 15932 -4376
rect 12871 -4536 14243 -4489
rect 14565 -4535 15469 -4488
rect 13705 -4659 13739 -4536
rect 14177 -4549 14243 -4536
rect 14177 -4583 14193 -4549
rect 14227 -4583 14243 -4549
rect 14177 -4599 14243 -4583
rect 14566 -4659 14600 -4535
rect 13700 -4671 13746 -4659
rect 13700 -4847 13706 -4671
rect 13740 -4847 13746 -4671
rect 13700 -4859 13746 -4847
rect 13818 -4671 13938 -4659
rect 13818 -4847 13824 -4671
rect 13858 -4847 13898 -4671
rect 13818 -4859 13898 -4847
rect 13824 -5226 13858 -4859
rect 13892 -5047 13898 -4859
rect 13932 -5047 13938 -4671
rect 13892 -5059 13938 -5047
rect 14010 -4671 14056 -4659
rect 14010 -5047 14016 -4671
rect 14050 -5047 14056 -4671
rect 14010 -5059 14056 -5047
rect 14128 -4671 14174 -4659
rect 14128 -5047 14134 -4671
rect 14168 -5047 14174 -4671
rect 14128 -5059 14174 -5047
rect 14246 -4671 14292 -4659
rect 14246 -5047 14252 -4671
rect 14286 -5047 14292 -4671
rect 14246 -5059 14292 -5047
rect 14364 -4671 14488 -4659
rect 14364 -5047 14370 -4671
rect 14404 -4847 14448 -4671
rect 14482 -4847 14488 -4671
rect 14404 -4859 14488 -4847
rect 14560 -4671 14606 -4659
rect 14560 -4847 14566 -4671
rect 14600 -4847 14606 -4671
rect 14560 -4859 14606 -4847
rect 14404 -5047 14410 -4859
rect 14364 -5059 14410 -5047
rect 14134 -5132 14168 -5059
rect 14119 -5148 14185 -5132
rect 14119 -5182 14135 -5148
rect 14169 -5182 14185 -5148
rect 14119 -5198 14185 -5182
rect 14448 -5226 14482 -4859
rect 13824 -5278 14482 -5226
rect 14122 -5300 14214 -5278
rect 14122 -5352 14134 -5300
rect 14200 -5352 14214 -5300
rect 14122 -5356 14214 -5352
rect 15814 -5391 15862 -4384
rect 16015 -4489 16050 -3979
rect 16105 -4025 16197 -4012
rect 16105 -4088 16117 -4025
rect 16188 -4088 16197 -4025
rect 16105 -4097 16197 -4088
rect 17190 -4025 17282 -4015
rect 17190 -4087 17202 -4025
rect 17272 -4087 17282 -4025
rect 17190 -4100 17282 -4087
rect 18578 -4080 18613 -3726
rect 18688 -4080 18759 -2899
rect 18906 -2839 18986 -1648
rect 19157 -1753 19192 -1243
rect 19247 -1289 19339 -1276
rect 19247 -1352 19259 -1289
rect 19330 -1352 19339 -1289
rect 19247 -1361 19339 -1352
rect 20332 -1289 20424 -1279
rect 20332 -1351 20344 -1289
rect 20414 -1351 20424 -1289
rect 20332 -1364 20424 -1351
rect 21720 -1344 21755 -990
rect 20579 -1406 20644 -1403
rect 20579 -1409 20648 -1406
rect 20579 -1469 20585 -1409
rect 20644 -1469 20654 -1409
rect 20579 -1473 20648 -1469
rect 20579 -1475 20644 -1473
rect 21720 -1490 21901 -1344
rect 22042 -1396 22113 -77
rect 23540 -406 23550 -346
rect 23630 -406 23640 -346
rect 23540 -446 23640 -406
rect 22743 -503 24546 -446
rect 22743 -590 22777 -503
rect 23918 -590 23952 -503
rect 22737 -602 22783 -590
rect 22737 -790 22743 -602
rect 22296 -802 22342 -790
rect 22296 -978 22302 -802
rect 22336 -978 22342 -802
rect 22296 -990 22342 -978
rect 22414 -802 22460 -790
rect 22414 -978 22420 -802
rect 22454 -978 22460 -802
rect 22414 -990 22460 -978
rect 22532 -802 22578 -790
rect 22532 -978 22538 -802
rect 22572 -978 22578 -802
rect 22532 -990 22578 -978
rect 22650 -802 22743 -790
rect 22650 -978 22656 -802
rect 22690 -978 22743 -802
rect 22777 -978 22783 -602
rect 22650 -990 22783 -978
rect 22855 -602 22901 -590
rect 22855 -978 22861 -602
rect 22895 -978 22901 -602
rect 22855 -990 22901 -978
rect 22973 -602 23019 -590
rect 22973 -978 22979 -602
rect 23013 -978 23019 -602
rect 22973 -990 23019 -978
rect 23091 -602 23137 -590
rect 23091 -978 23097 -602
rect 23131 -978 23137 -602
rect 23091 -990 23137 -978
rect 23204 -602 23250 -590
rect 23204 -978 23210 -602
rect 23244 -978 23250 -602
rect 23204 -990 23250 -978
rect 23322 -602 23368 -590
rect 23322 -978 23328 -602
rect 23362 -978 23368 -602
rect 23322 -990 23368 -978
rect 23440 -602 23486 -590
rect 23440 -978 23446 -602
rect 23480 -978 23486 -602
rect 23440 -990 23486 -978
rect 23558 -602 23604 -590
rect 23558 -978 23564 -602
rect 23598 -978 23604 -602
rect 23558 -990 23604 -978
rect 23676 -602 23722 -590
rect 23676 -978 23682 -602
rect 23716 -978 23722 -602
rect 23676 -990 23722 -978
rect 23794 -602 23840 -590
rect 23794 -978 23800 -602
rect 23834 -978 23840 -602
rect 23794 -990 23840 -978
rect 23912 -602 23958 -590
rect 23912 -978 23918 -602
rect 23952 -978 23958 -602
rect 23912 -990 23958 -978
rect 24031 -602 24077 -590
rect 24031 -978 24037 -602
rect 24071 -978 24077 -602
rect 24031 -990 24077 -978
rect 24149 -602 24195 -590
rect 24149 -978 24155 -602
rect 24189 -978 24195 -602
rect 24149 -990 24195 -978
rect 24267 -602 24313 -590
rect 24267 -978 24273 -602
rect 24307 -978 24313 -602
rect 24267 -990 24313 -978
rect 24385 -602 24431 -590
rect 24385 -978 24391 -602
rect 24425 -978 24431 -602
rect 24509 -790 24546 -503
rect 24385 -990 24431 -978
rect 24504 -802 24550 -790
rect 24504 -978 24510 -802
rect 24544 -978 24550 -802
rect 24504 -990 24550 -978
rect 24622 -802 24668 -790
rect 24622 -978 24628 -802
rect 24662 -978 24668 -802
rect 24622 -990 24668 -978
rect 24740 -802 24786 -790
rect 24740 -978 24746 -802
rect 24780 -978 24786 -802
rect 24740 -990 24786 -978
rect 24858 -802 24904 -790
rect 24858 -978 24864 -802
rect 24898 -978 24904 -802
rect 24858 -990 24904 -978
rect 22301 -1176 22336 -990
rect 23210 -1074 23244 -990
rect 24391 -1074 24425 -990
rect 23210 -1116 24425 -1074
rect 24391 -1136 24425 -1116
rect 24391 -1152 24748 -1136
rect 22301 -1193 23438 -1176
rect 22301 -1227 23388 -1193
rect 23422 -1227 23438 -1193
rect 24391 -1186 24698 -1152
rect 24732 -1186 24748 -1152
rect 24391 -1202 24748 -1186
rect 22301 -1243 23438 -1227
rect 22042 -1404 22218 -1396
rect 22042 -1472 22159 -1404
rect 22216 -1472 22226 -1404
rect 22042 -1480 22218 -1472
rect 20214 -1572 20306 -1564
rect 20214 -1637 20226 -1572
rect 20294 -1637 20306 -1572
rect 20214 -1649 20306 -1637
rect 21720 -1752 21755 -1490
rect 19157 -1800 20529 -1753
rect 20851 -1799 21755 -1752
rect 21805 -1784 21901 -1490
rect 19991 -1923 20025 -1800
rect 20463 -1813 20529 -1800
rect 20463 -1847 20479 -1813
rect 20513 -1847 20529 -1813
rect 20463 -1863 20529 -1847
rect 20852 -1923 20886 -1799
rect 21805 -1855 21817 -1784
rect 21888 -1855 21901 -1784
rect 21805 -1865 21901 -1855
rect 22090 -1572 22218 -1564
rect 22090 -1640 22159 -1572
rect 22216 -1640 22226 -1572
rect 22090 -1648 22218 -1640
rect 19986 -1935 20032 -1923
rect 19986 -2111 19992 -1935
rect 20026 -2111 20032 -1935
rect 19986 -2123 20032 -2111
rect 20104 -1935 20224 -1923
rect 20104 -2111 20110 -1935
rect 20144 -2111 20184 -1935
rect 20104 -2123 20184 -2111
rect 20110 -2490 20144 -2123
rect 20178 -2311 20184 -2123
rect 20218 -2311 20224 -1935
rect 20178 -2323 20224 -2311
rect 20296 -1935 20342 -1923
rect 20296 -2311 20302 -1935
rect 20336 -2311 20342 -1935
rect 20296 -2323 20342 -2311
rect 20414 -1935 20460 -1923
rect 20414 -2311 20420 -1935
rect 20454 -2311 20460 -1935
rect 20414 -2323 20460 -2311
rect 20532 -1935 20578 -1923
rect 20532 -2311 20538 -1935
rect 20572 -2311 20578 -1935
rect 20532 -2323 20578 -2311
rect 20650 -1935 20774 -1923
rect 20650 -2311 20656 -1935
rect 20690 -2111 20734 -1935
rect 20768 -2111 20774 -1935
rect 20690 -2123 20774 -2111
rect 20846 -1935 20892 -1923
rect 20846 -2111 20852 -1935
rect 20886 -2111 20892 -1935
rect 20846 -2123 20892 -2111
rect 20690 -2311 20696 -2123
rect 20650 -2323 20696 -2311
rect 20420 -2396 20454 -2323
rect 20405 -2412 20471 -2396
rect 20405 -2446 20421 -2412
rect 20455 -2446 20471 -2412
rect 20405 -2462 20471 -2446
rect 20734 -2490 20768 -2123
rect 20110 -2542 20768 -2490
rect 20408 -2564 20500 -2542
rect 20408 -2616 20420 -2564
rect 20486 -2616 20500 -2564
rect 20408 -2620 20500 -2616
rect 22090 -2839 22141 -1648
rect 22301 -1753 22336 -1243
rect 22391 -1289 22483 -1276
rect 22391 -1352 22403 -1289
rect 22474 -1352 22483 -1289
rect 22391 -1361 22483 -1352
rect 23476 -1289 23568 -1279
rect 23476 -1351 23488 -1289
rect 23558 -1351 23568 -1289
rect 23476 -1364 23568 -1351
rect 24864 -1344 24899 -990
rect 23723 -1406 23788 -1403
rect 23723 -1409 23792 -1406
rect 23723 -1469 23729 -1409
rect 23788 -1469 23798 -1409
rect 23723 -1473 23792 -1469
rect 23723 -1475 23788 -1473
rect 24864 -1490 25344 -1344
rect 23358 -1572 23450 -1564
rect 23358 -1637 23370 -1572
rect 23438 -1637 23450 -1572
rect 23358 -1649 23450 -1637
rect 24864 -1752 24899 -1490
rect 22301 -1800 23673 -1753
rect 23995 -1799 24899 -1752
rect 25240 -1777 25344 -1767
rect 23135 -1923 23169 -1800
rect 23607 -1813 23673 -1800
rect 23607 -1847 23623 -1813
rect 23657 -1847 23673 -1813
rect 23607 -1863 23673 -1847
rect 23996 -1923 24030 -1799
rect 25197 -1847 25207 -1777
rect 25266 -1847 25344 -1777
rect 25240 -1855 25344 -1847
rect 23130 -1935 23176 -1923
rect 23130 -2111 23136 -1935
rect 23170 -2111 23176 -1935
rect 23130 -2123 23176 -2111
rect 23248 -1935 23368 -1923
rect 23248 -2111 23254 -1935
rect 23288 -2111 23328 -1935
rect 23248 -2123 23328 -2111
rect 23254 -2490 23288 -2123
rect 23322 -2311 23328 -2123
rect 23362 -2311 23368 -1935
rect 23322 -2323 23368 -2311
rect 23440 -1935 23486 -1923
rect 23440 -2311 23446 -1935
rect 23480 -2311 23486 -1935
rect 23440 -2323 23486 -2311
rect 23558 -1935 23604 -1923
rect 23558 -2311 23564 -1935
rect 23598 -2311 23604 -1935
rect 23558 -2323 23604 -2311
rect 23676 -1935 23722 -1923
rect 23676 -2311 23682 -1935
rect 23716 -2311 23722 -1935
rect 23676 -2323 23722 -2311
rect 23794 -1935 23918 -1923
rect 23794 -2311 23800 -1935
rect 23834 -2111 23878 -1935
rect 23912 -2111 23918 -1935
rect 23834 -2123 23918 -2111
rect 23990 -1935 24036 -1923
rect 23990 -2111 23996 -1935
rect 24030 -2111 24036 -1935
rect 25195 -1969 25344 -1956
rect 25195 -2032 25206 -1969
rect 25267 -2032 25344 -1969
rect 25195 -2042 25344 -2032
rect 23990 -2123 24036 -2111
rect 23834 -2311 23840 -2123
rect 23794 -2323 23840 -2311
rect 23564 -2396 23598 -2323
rect 23549 -2412 23615 -2396
rect 23549 -2446 23565 -2412
rect 23599 -2446 23615 -2412
rect 23549 -2462 23615 -2446
rect 23878 -2490 23912 -2123
rect 25193 -2189 25344 -2172
rect 25193 -2255 25205 -2189
rect 25267 -2255 25344 -2189
rect 25193 -2267 25344 -2255
rect 25195 -2385 25345 -2368
rect 25195 -2443 25205 -2385
rect 25268 -2443 25345 -2385
rect 25195 -2454 25345 -2443
rect 23254 -2542 23912 -2490
rect 23552 -2564 23644 -2542
rect 23552 -2616 23564 -2564
rect 23630 -2616 23644 -2564
rect 23552 -2620 23644 -2616
rect 25193 -2728 25346 -2710
rect 25193 -2789 25204 -2728
rect 25268 -2789 25346 -2728
rect 25193 -2800 25346 -2789
rect 18906 -2900 21891 -2839
rect 20386 -3138 20396 -3078
rect 20476 -3138 20486 -3078
rect 20386 -3178 20486 -3138
rect 19589 -3235 21392 -3178
rect 19589 -3322 19623 -3235
rect 20764 -3322 20798 -3235
rect 19583 -3334 19629 -3322
rect 19583 -3522 19589 -3334
rect 19142 -3534 19188 -3522
rect 19142 -3710 19148 -3534
rect 19182 -3710 19188 -3534
rect 19142 -3722 19188 -3710
rect 19260 -3534 19306 -3522
rect 19260 -3710 19266 -3534
rect 19300 -3710 19306 -3534
rect 19260 -3722 19306 -3710
rect 19378 -3534 19424 -3522
rect 19378 -3710 19384 -3534
rect 19418 -3710 19424 -3534
rect 19378 -3722 19424 -3710
rect 19496 -3534 19589 -3522
rect 19496 -3710 19502 -3534
rect 19536 -3710 19589 -3534
rect 19623 -3710 19629 -3334
rect 19496 -3722 19629 -3710
rect 19701 -3334 19747 -3322
rect 19701 -3710 19707 -3334
rect 19741 -3710 19747 -3334
rect 19701 -3722 19747 -3710
rect 19819 -3334 19865 -3322
rect 19819 -3710 19825 -3334
rect 19859 -3710 19865 -3334
rect 19819 -3722 19865 -3710
rect 19937 -3334 19983 -3322
rect 19937 -3710 19943 -3334
rect 19977 -3710 19983 -3334
rect 19937 -3722 19983 -3710
rect 20050 -3334 20096 -3322
rect 20050 -3710 20056 -3334
rect 20090 -3710 20096 -3334
rect 20050 -3722 20096 -3710
rect 20168 -3334 20214 -3322
rect 20168 -3710 20174 -3334
rect 20208 -3710 20214 -3334
rect 20168 -3722 20214 -3710
rect 20286 -3334 20332 -3322
rect 20286 -3710 20292 -3334
rect 20326 -3710 20332 -3334
rect 20286 -3722 20332 -3710
rect 20404 -3334 20450 -3322
rect 20404 -3710 20410 -3334
rect 20444 -3710 20450 -3334
rect 20404 -3722 20450 -3710
rect 20522 -3334 20568 -3322
rect 20522 -3710 20528 -3334
rect 20562 -3710 20568 -3334
rect 20522 -3722 20568 -3710
rect 20640 -3334 20686 -3322
rect 20640 -3710 20646 -3334
rect 20680 -3710 20686 -3334
rect 20640 -3722 20686 -3710
rect 20758 -3334 20804 -3322
rect 20758 -3710 20764 -3334
rect 20798 -3710 20804 -3334
rect 20758 -3722 20804 -3710
rect 20877 -3334 20923 -3322
rect 20877 -3710 20883 -3334
rect 20917 -3710 20923 -3334
rect 20877 -3722 20923 -3710
rect 20995 -3334 21041 -3322
rect 20995 -3710 21001 -3334
rect 21035 -3710 21041 -3334
rect 20995 -3722 21041 -3710
rect 21113 -3334 21159 -3322
rect 21113 -3710 21119 -3334
rect 21153 -3710 21159 -3334
rect 21113 -3722 21159 -3710
rect 21231 -3334 21277 -3322
rect 21231 -3710 21237 -3334
rect 21271 -3710 21277 -3334
rect 21355 -3522 21392 -3235
rect 21231 -3722 21277 -3710
rect 21350 -3534 21396 -3522
rect 21350 -3710 21356 -3534
rect 21390 -3710 21396 -3534
rect 21350 -3722 21396 -3710
rect 21468 -3534 21514 -3522
rect 21468 -3710 21474 -3534
rect 21508 -3710 21514 -3534
rect 21468 -3722 21514 -3710
rect 21586 -3534 21632 -3522
rect 21586 -3710 21592 -3534
rect 21626 -3710 21632 -3534
rect 21586 -3722 21632 -3710
rect 21704 -3534 21750 -3522
rect 21704 -3710 21710 -3534
rect 21744 -3710 21750 -3534
rect 21704 -3722 21750 -3710
rect 19147 -3908 19182 -3722
rect 20056 -3806 20090 -3722
rect 21237 -3806 21271 -3722
rect 20056 -3848 21271 -3806
rect 21237 -3868 21271 -3848
rect 21237 -3884 21594 -3868
rect 19147 -3925 20284 -3908
rect 19147 -3959 20234 -3925
rect 20268 -3959 20284 -3925
rect 21237 -3918 21544 -3884
rect 21578 -3918 21594 -3884
rect 21237 -3934 21594 -3918
rect 19147 -3975 20284 -3959
rect 17437 -4142 17502 -4139
rect 17437 -4145 17506 -4142
rect 17437 -4205 17443 -4145
rect 17502 -4205 17512 -4145
rect 17437 -4209 17506 -4205
rect 17437 -4211 17502 -4209
rect 18578 -4226 18759 -4080
rect 18888 -4020 19064 -4012
rect 18888 -4088 19005 -4020
rect 19062 -4088 19072 -4020
rect 18888 -4096 19064 -4088
rect 18994 -4136 19064 -4128
rect 18994 -4204 19005 -4136
rect 19062 -4204 19072 -4136
rect 18994 -4212 19064 -4204
rect 17072 -4308 17164 -4300
rect 17072 -4373 17084 -4308
rect 17152 -4373 17164 -4308
rect 17072 -4385 17164 -4373
rect 18578 -4488 18613 -4226
rect 16015 -4536 17387 -4489
rect 17709 -4535 18613 -4488
rect 18945 -4304 19064 -4296
rect 18945 -4372 19005 -4304
rect 19062 -4372 19072 -4304
rect 18945 -4380 19064 -4372
rect 16849 -4659 16883 -4536
rect 17321 -4549 17387 -4536
rect 17321 -4583 17337 -4549
rect 17371 -4583 17387 -4549
rect 17321 -4599 17387 -4583
rect 17710 -4659 17744 -4535
rect 16844 -4671 16890 -4659
rect 16844 -4847 16850 -4671
rect 16884 -4847 16890 -4671
rect 16844 -4859 16890 -4847
rect 16962 -4671 17082 -4659
rect 16962 -4847 16968 -4671
rect 17002 -4847 17042 -4671
rect 16962 -4859 17042 -4847
rect 16968 -5226 17002 -4859
rect 17036 -5047 17042 -4859
rect 17076 -5047 17082 -4671
rect 17036 -5059 17082 -5047
rect 17154 -4671 17200 -4659
rect 17154 -5047 17160 -4671
rect 17194 -5047 17200 -4671
rect 17154 -5059 17200 -5047
rect 17272 -4671 17318 -4659
rect 17272 -5047 17278 -4671
rect 17312 -5047 17318 -4671
rect 17272 -5059 17318 -5047
rect 17390 -4671 17436 -4659
rect 17390 -5047 17396 -4671
rect 17430 -5047 17436 -4671
rect 17390 -5059 17436 -5047
rect 17508 -4671 17632 -4659
rect 17508 -5047 17514 -4671
rect 17548 -4847 17592 -4671
rect 17626 -4847 17632 -4671
rect 17548 -4859 17632 -4847
rect 17704 -4671 17750 -4659
rect 17704 -4847 17710 -4671
rect 17744 -4847 17750 -4671
rect 17704 -4859 17750 -4847
rect 17548 -5047 17554 -4859
rect 17508 -5059 17554 -5047
rect 17278 -5132 17312 -5059
rect 17263 -5148 17329 -5132
rect 17263 -5182 17279 -5148
rect 17313 -5182 17329 -5148
rect 17263 -5198 17329 -5182
rect 17592 -5226 17626 -4859
rect 16968 -5278 17626 -5226
rect 17266 -5300 17358 -5278
rect 17266 -5352 17278 -5300
rect 17344 -5352 17358 -5300
rect 17266 -5356 17358 -5352
rect 18945 -5388 18993 -4380
rect 19147 -4485 19182 -3975
rect 19237 -4021 19329 -4008
rect 19237 -4084 19249 -4021
rect 19320 -4084 19329 -4021
rect 19237 -4093 19329 -4084
rect 20322 -4021 20414 -4011
rect 20322 -4083 20334 -4021
rect 20404 -4083 20414 -4021
rect 20322 -4096 20414 -4083
rect 21710 -4076 21745 -3722
rect 21820 -4076 21891 -2900
rect 22090 -2840 23444 -2839
rect 22090 -2901 24894 -2840
rect 23530 -3138 23540 -3078
rect 23620 -3138 23630 -3078
rect 23530 -3178 23630 -3138
rect 22733 -3235 24536 -3178
rect 22733 -3322 22767 -3235
rect 23908 -3322 23942 -3235
rect 22727 -3334 22773 -3322
rect 22727 -3522 22733 -3334
rect 22286 -3534 22332 -3522
rect 22286 -3710 22292 -3534
rect 22326 -3710 22332 -3534
rect 22286 -3722 22332 -3710
rect 22404 -3534 22450 -3522
rect 22404 -3710 22410 -3534
rect 22444 -3710 22450 -3534
rect 22404 -3722 22450 -3710
rect 22522 -3534 22568 -3522
rect 22522 -3710 22528 -3534
rect 22562 -3710 22568 -3534
rect 22522 -3722 22568 -3710
rect 22640 -3534 22733 -3522
rect 22640 -3710 22646 -3534
rect 22680 -3710 22733 -3534
rect 22767 -3710 22773 -3334
rect 22640 -3722 22773 -3710
rect 22845 -3334 22891 -3322
rect 22845 -3710 22851 -3334
rect 22885 -3710 22891 -3334
rect 22845 -3722 22891 -3710
rect 22963 -3334 23009 -3322
rect 22963 -3710 22969 -3334
rect 23003 -3710 23009 -3334
rect 22963 -3722 23009 -3710
rect 23081 -3334 23127 -3322
rect 23081 -3710 23087 -3334
rect 23121 -3710 23127 -3334
rect 23081 -3722 23127 -3710
rect 23194 -3334 23240 -3322
rect 23194 -3710 23200 -3334
rect 23234 -3710 23240 -3334
rect 23194 -3722 23240 -3710
rect 23312 -3334 23358 -3322
rect 23312 -3710 23318 -3334
rect 23352 -3710 23358 -3334
rect 23312 -3722 23358 -3710
rect 23430 -3334 23476 -3322
rect 23430 -3710 23436 -3334
rect 23470 -3710 23476 -3334
rect 23430 -3722 23476 -3710
rect 23548 -3334 23594 -3322
rect 23548 -3710 23554 -3334
rect 23588 -3710 23594 -3334
rect 23548 -3722 23594 -3710
rect 23666 -3334 23712 -3322
rect 23666 -3710 23672 -3334
rect 23706 -3710 23712 -3334
rect 23666 -3722 23712 -3710
rect 23784 -3334 23830 -3322
rect 23784 -3710 23790 -3334
rect 23824 -3710 23830 -3334
rect 23784 -3722 23830 -3710
rect 23902 -3334 23948 -3322
rect 23902 -3710 23908 -3334
rect 23942 -3710 23948 -3334
rect 23902 -3722 23948 -3710
rect 24021 -3334 24067 -3322
rect 24021 -3710 24027 -3334
rect 24061 -3710 24067 -3334
rect 24021 -3722 24067 -3710
rect 24139 -3334 24185 -3322
rect 24139 -3710 24145 -3334
rect 24179 -3710 24185 -3334
rect 24139 -3722 24185 -3710
rect 24257 -3334 24303 -3322
rect 24257 -3710 24263 -3334
rect 24297 -3710 24303 -3334
rect 24257 -3722 24303 -3710
rect 24375 -3334 24421 -3322
rect 24375 -3710 24381 -3334
rect 24415 -3710 24421 -3334
rect 24499 -3522 24536 -3235
rect 24375 -3722 24421 -3710
rect 24494 -3534 24540 -3522
rect 24494 -3710 24500 -3534
rect 24534 -3710 24540 -3534
rect 24494 -3722 24540 -3710
rect 24612 -3534 24658 -3522
rect 24612 -3710 24618 -3534
rect 24652 -3710 24658 -3534
rect 24612 -3722 24658 -3710
rect 24730 -3534 24776 -3522
rect 24730 -3710 24736 -3534
rect 24770 -3710 24776 -3534
rect 24730 -3722 24776 -3710
rect 24848 -3534 24894 -2901
rect 25195 -2900 25346 -2883
rect 25195 -2960 25206 -2900
rect 25270 -2960 25346 -2900
rect 25195 -2972 25346 -2960
rect 25192 -3254 25348 -3234
rect 25192 -3315 25205 -3254
rect 25272 -3315 25348 -3254
rect 25192 -3328 25348 -3315
rect 24848 -3710 24854 -3534
rect 24888 -3710 24894 -3534
rect 24848 -3722 24894 -3710
rect 22291 -3908 22326 -3722
rect 23200 -3806 23234 -3722
rect 24381 -3806 24415 -3722
rect 23200 -3848 24415 -3806
rect 24381 -3868 24415 -3848
rect 24381 -3884 24738 -3868
rect 22291 -3925 23428 -3908
rect 22291 -3959 23378 -3925
rect 23412 -3959 23428 -3925
rect 24381 -3918 24688 -3884
rect 24722 -3918 24738 -3884
rect 24381 -3934 24738 -3918
rect 22291 -3975 23428 -3959
rect 20569 -4138 20634 -4135
rect 20569 -4141 20638 -4138
rect 20569 -4201 20575 -4141
rect 20634 -4201 20644 -4141
rect 20569 -4205 20638 -4201
rect 20569 -4207 20634 -4205
rect 21710 -4222 21891 -4076
rect 22032 -4020 22208 -4012
rect 22032 -4088 22149 -4020
rect 22206 -4088 22216 -4020
rect 22032 -4096 22208 -4088
rect 22138 -4136 22208 -4128
rect 22138 -4204 22149 -4136
rect 22206 -4204 22216 -4136
rect 22138 -4212 22208 -4204
rect 20204 -4304 20296 -4296
rect 20204 -4369 20216 -4304
rect 20284 -4369 20296 -4304
rect 20204 -4381 20296 -4369
rect 21710 -4484 21745 -4222
rect 19147 -4532 20519 -4485
rect 20841 -4531 21745 -4484
rect 22074 -4296 22138 -4295
rect 22074 -4304 22208 -4296
rect 22074 -4372 22149 -4304
rect 22206 -4372 22216 -4304
rect 22074 -4380 22208 -4372
rect 19981 -4655 20015 -4532
rect 20453 -4545 20519 -4532
rect 20453 -4579 20469 -4545
rect 20503 -4579 20519 -4545
rect 20453 -4595 20519 -4579
rect 20842 -4655 20876 -4531
rect 19976 -4667 20022 -4655
rect 19976 -4843 19982 -4667
rect 20016 -4843 20022 -4667
rect 19976 -4855 20022 -4843
rect 20094 -4667 20214 -4655
rect 20094 -4843 20100 -4667
rect 20134 -4843 20174 -4667
rect 20094 -4855 20174 -4843
rect 20100 -5222 20134 -4855
rect 20168 -5043 20174 -4855
rect 20208 -5043 20214 -4667
rect 20168 -5055 20214 -5043
rect 20286 -4667 20332 -4655
rect 20286 -5043 20292 -4667
rect 20326 -5043 20332 -4667
rect 20286 -5055 20332 -5043
rect 20404 -4667 20450 -4655
rect 20404 -5043 20410 -4667
rect 20444 -5043 20450 -4667
rect 20404 -5055 20450 -5043
rect 20522 -4667 20568 -4655
rect 20522 -5043 20528 -4667
rect 20562 -5043 20568 -4667
rect 20522 -5055 20568 -5043
rect 20640 -4667 20764 -4655
rect 20640 -5043 20646 -4667
rect 20680 -4843 20724 -4667
rect 20758 -4843 20764 -4667
rect 20680 -4855 20764 -4843
rect 20836 -4667 20882 -4655
rect 20836 -4843 20842 -4667
rect 20876 -4843 20882 -4667
rect 20836 -4855 20882 -4843
rect 20680 -5043 20686 -4855
rect 20640 -5055 20686 -5043
rect 20410 -5128 20444 -5055
rect 20395 -5144 20461 -5128
rect 20395 -5178 20411 -5144
rect 20445 -5178 20461 -5144
rect 20395 -5194 20461 -5178
rect 20724 -5222 20758 -4855
rect 20100 -5274 20758 -5222
rect 20398 -5296 20490 -5274
rect 20398 -5348 20410 -5296
rect 20476 -5348 20490 -5296
rect 20398 -5352 20490 -5348
rect 9468 -5442 12640 -5394
rect 12672 -5440 15786 -5391
rect 15814 -5392 17421 -5391
rect 15814 -5440 18909 -5392
rect 18945 -5436 21665 -5388
rect 12592 -5468 12640 -5442
rect 6308 -5518 12564 -5470
rect 12592 -5516 15710 -5468
rect 12516 -5544 12564 -5518
rect 12516 -5592 15639 -5544
rect 15591 -5623 15639 -5592
rect 15667 -5546 15710 -5516
rect 15738 -5470 15786 -5440
rect 18861 -5464 18909 -5440
rect 15738 -5518 18789 -5470
rect 18861 -5512 20922 -5464
rect 18741 -5542 18789 -5518
rect 15667 -5594 18713 -5546
rect 18741 -5590 20189 -5542
rect 18665 -5618 18713 -5594
rect 15591 -5671 18637 -5623
rect 18665 -5666 19445 -5618
rect 3176 -5754 17951 -5706
rect 32 -5863 17207 -5815
rect 16867 -5975 16877 -5961
rect 16837 -5981 16877 -5975
rect 16953 -5975 16963 -5961
rect 16953 -5981 16995 -5975
rect 804 -6042 814 -6020
rect 776 -6074 814 -6042
rect 868 -6042 878 -6020
rect 2872 -6040 2882 -6018
rect 868 -6074 910 -6042
rect 776 -6125 910 -6074
rect 2844 -6072 2882 -6040
rect 2936 -6040 2946 -6018
rect 2936 -6072 2978 -6040
rect 4941 -6042 4951 -6020
rect 2844 -6123 2978 -6072
rect 4913 -6074 4951 -6042
rect 5005 -6042 5015 -6020
rect 7009 -6040 7019 -6018
rect 5005 -6074 5047 -6042
rect 105 -6168 1578 -6125
rect 105 -6471 139 -6168
rect 471 -6271 505 -6168
rect 707 -6271 741 -6168
rect 943 -6271 977 -6168
rect 1179 -6271 1213 -6168
rect 465 -6283 511 -6271
rect -19 -6483 27 -6471
rect -19 -6659 -13 -6483
rect 21 -6659 27 -6483
rect -19 -6671 27 -6659
rect 99 -6483 145 -6471
rect 99 -6659 105 -6483
rect 139 -6659 145 -6483
rect 99 -6671 145 -6659
rect 217 -6483 263 -6471
rect 217 -6659 223 -6483
rect 257 -6659 263 -6483
rect 217 -6671 263 -6659
rect 335 -6483 381 -6471
rect 465 -6483 471 -6283
rect 335 -6659 341 -6483
rect 375 -6659 471 -6483
rect 505 -6659 511 -6283
rect 335 -6671 381 -6659
rect 465 -6671 511 -6659
rect 583 -6283 629 -6271
rect 583 -6659 589 -6283
rect 623 -6659 629 -6283
rect 583 -6671 629 -6659
rect 701 -6283 747 -6271
rect 701 -6659 707 -6283
rect 741 -6659 747 -6283
rect 701 -6671 747 -6659
rect 819 -6283 865 -6271
rect 819 -6659 825 -6283
rect 859 -6659 865 -6283
rect 819 -6671 865 -6659
rect 937 -6283 983 -6271
rect 937 -6659 943 -6283
rect 977 -6659 983 -6283
rect 937 -6671 983 -6659
rect 1055 -6283 1101 -6271
rect 1055 -6659 1061 -6283
rect 1095 -6659 1101 -6283
rect 1055 -6671 1101 -6659
rect 1173 -6283 1219 -6271
rect 1173 -6659 1179 -6283
rect 1213 -6483 1219 -6283
rect 1544 -6471 1578 -6168
rect 2173 -6166 3646 -6123
rect 4913 -6125 5047 -6074
rect 6981 -6072 7019 -6040
rect 7073 -6040 7083 -6018
rect 9078 -6040 9088 -6018
rect 7073 -6072 7115 -6040
rect 6981 -6123 7115 -6072
rect 9050 -6072 9088 -6040
rect 9142 -6040 9152 -6018
rect 11146 -6038 11156 -6016
rect 9142 -6072 9184 -6040
rect 9050 -6123 9184 -6072
rect 11118 -6070 11156 -6038
rect 11210 -6038 11220 -6016
rect 11210 -6070 11252 -6038
rect 13215 -6040 13225 -6018
rect 11118 -6121 11252 -6070
rect 13187 -6072 13225 -6040
rect 13279 -6040 13289 -6018
rect 15283 -6038 15293 -6016
rect 13279 -6072 13321 -6040
rect 2173 -6469 2207 -6166
rect 2539 -6269 2573 -6166
rect 2775 -6269 2809 -6166
rect 3011 -6269 3045 -6166
rect 3247 -6269 3281 -6166
rect 2533 -6281 2579 -6269
rect 1302 -6483 1348 -6471
rect 1213 -6659 1308 -6483
rect 1342 -6659 1348 -6483
rect 1173 -6671 1219 -6659
rect 1302 -6671 1348 -6659
rect 1420 -6483 1466 -6471
rect 1420 -6659 1426 -6483
rect 1460 -6659 1466 -6483
rect 1420 -6671 1466 -6659
rect 1538 -6483 1584 -6471
rect 1538 -6659 1544 -6483
rect 1578 -6659 1584 -6483
rect 1538 -6671 1584 -6659
rect 1656 -6483 1702 -6471
rect 1656 -6659 1662 -6483
rect 1696 -6659 1702 -6483
rect 1656 -6671 1702 -6659
rect 2049 -6481 2095 -6469
rect 2049 -6657 2055 -6481
rect 2089 -6657 2095 -6481
rect 2049 -6669 2095 -6657
rect 2167 -6481 2213 -6469
rect 2167 -6657 2173 -6481
rect 2207 -6657 2213 -6481
rect 2167 -6669 2213 -6657
rect 2285 -6481 2331 -6469
rect 2285 -6657 2291 -6481
rect 2325 -6657 2331 -6481
rect 2285 -6669 2331 -6657
rect 2403 -6481 2449 -6469
rect 2533 -6481 2539 -6281
rect 2403 -6657 2409 -6481
rect 2443 -6657 2539 -6481
rect 2573 -6657 2579 -6281
rect 2403 -6669 2449 -6657
rect 2533 -6669 2579 -6657
rect 2651 -6281 2697 -6269
rect 2651 -6657 2657 -6281
rect 2691 -6657 2697 -6281
rect 2651 -6669 2697 -6657
rect 2769 -6281 2815 -6269
rect 2769 -6657 2775 -6281
rect 2809 -6657 2815 -6281
rect 2769 -6669 2815 -6657
rect 2887 -6281 2933 -6269
rect 2887 -6657 2893 -6281
rect 2927 -6657 2933 -6281
rect 2887 -6669 2933 -6657
rect 3005 -6281 3051 -6269
rect 3005 -6657 3011 -6281
rect 3045 -6657 3051 -6281
rect 3005 -6669 3051 -6657
rect 3123 -6281 3169 -6269
rect 3123 -6657 3129 -6281
rect 3163 -6657 3169 -6281
rect 3123 -6669 3169 -6657
rect 3241 -6281 3287 -6269
rect 3241 -6657 3247 -6281
rect 3281 -6481 3287 -6281
rect 3612 -6469 3646 -6166
rect 4242 -6168 5715 -6125
rect 3370 -6481 3416 -6469
rect 3281 -6657 3376 -6481
rect 3410 -6657 3416 -6481
rect 3241 -6669 3287 -6657
rect 3370 -6669 3416 -6657
rect 3488 -6481 3534 -6469
rect 3488 -6657 3494 -6481
rect 3528 -6657 3534 -6481
rect 3488 -6669 3534 -6657
rect 3606 -6481 3652 -6469
rect 3606 -6657 3612 -6481
rect 3646 -6657 3652 -6481
rect 3606 -6669 3652 -6657
rect 3724 -6481 3770 -6469
rect 4242 -6471 4276 -6168
rect 4608 -6271 4642 -6168
rect 4844 -6271 4878 -6168
rect 5080 -6271 5114 -6168
rect 5316 -6271 5350 -6168
rect 4602 -6283 4648 -6271
rect 3724 -6657 3730 -6481
rect 3764 -6657 3770 -6481
rect 3724 -6669 3770 -6657
rect 4118 -6483 4164 -6471
rect 4118 -6659 4124 -6483
rect 4158 -6659 4164 -6483
rect -13 -6705 21 -6671
rect 589 -6705 623 -6671
rect 825 -6705 859 -6671
rect -13 -6740 146 -6705
rect 589 -6740 859 -6705
rect 1426 -6705 1460 -6671
rect 1662 -6705 1696 -6671
rect 1426 -6740 1696 -6705
rect 2055 -6703 2089 -6669
rect 2657 -6703 2691 -6669
rect 2893 -6703 2927 -6669
rect 2055 -6738 2214 -6703
rect 2657 -6738 2927 -6703
rect 3494 -6703 3528 -6669
rect 3730 -6703 3764 -6669
rect 4118 -6671 4164 -6659
rect 4236 -6483 4282 -6471
rect 4236 -6659 4242 -6483
rect 4276 -6659 4282 -6483
rect 4236 -6671 4282 -6659
rect 4354 -6483 4400 -6471
rect 4354 -6659 4360 -6483
rect 4394 -6659 4400 -6483
rect 4354 -6671 4400 -6659
rect 4472 -6483 4518 -6471
rect 4602 -6483 4608 -6283
rect 4472 -6659 4478 -6483
rect 4512 -6659 4608 -6483
rect 4642 -6659 4648 -6283
rect 4472 -6671 4518 -6659
rect 4602 -6671 4648 -6659
rect 4720 -6283 4766 -6271
rect 4720 -6659 4726 -6283
rect 4760 -6659 4766 -6283
rect 4720 -6671 4766 -6659
rect 4838 -6283 4884 -6271
rect 4838 -6659 4844 -6283
rect 4878 -6659 4884 -6283
rect 4838 -6671 4884 -6659
rect 4956 -6283 5002 -6271
rect 4956 -6659 4962 -6283
rect 4996 -6659 5002 -6283
rect 4956 -6671 5002 -6659
rect 5074 -6283 5120 -6271
rect 5074 -6659 5080 -6283
rect 5114 -6659 5120 -6283
rect 5074 -6671 5120 -6659
rect 5192 -6283 5238 -6271
rect 5192 -6659 5198 -6283
rect 5232 -6659 5238 -6283
rect 5192 -6671 5238 -6659
rect 5310 -6283 5356 -6271
rect 5310 -6659 5316 -6283
rect 5350 -6483 5356 -6283
rect 5681 -6471 5715 -6168
rect 6310 -6166 7783 -6123
rect 6310 -6469 6344 -6166
rect 6676 -6269 6710 -6166
rect 6912 -6269 6946 -6166
rect 7148 -6269 7182 -6166
rect 7384 -6269 7418 -6166
rect 6670 -6281 6716 -6269
rect 5439 -6483 5485 -6471
rect 5350 -6659 5445 -6483
rect 5479 -6659 5485 -6483
rect 5310 -6671 5356 -6659
rect 5439 -6671 5485 -6659
rect 5557 -6483 5603 -6471
rect 5557 -6659 5563 -6483
rect 5597 -6659 5603 -6483
rect 5557 -6671 5603 -6659
rect 5675 -6483 5721 -6471
rect 5675 -6659 5681 -6483
rect 5715 -6659 5721 -6483
rect 5675 -6671 5721 -6659
rect 5793 -6483 5839 -6471
rect 5793 -6659 5799 -6483
rect 5833 -6659 5839 -6483
rect 5793 -6671 5839 -6659
rect 6186 -6481 6232 -6469
rect 6186 -6657 6192 -6481
rect 6226 -6657 6232 -6481
rect 6186 -6669 6232 -6657
rect 6304 -6481 6350 -6469
rect 6304 -6657 6310 -6481
rect 6344 -6657 6350 -6481
rect 6304 -6669 6350 -6657
rect 6422 -6481 6468 -6469
rect 6422 -6657 6428 -6481
rect 6462 -6657 6468 -6481
rect 6422 -6669 6468 -6657
rect 6540 -6481 6586 -6469
rect 6670 -6481 6676 -6281
rect 6540 -6657 6546 -6481
rect 6580 -6657 6676 -6481
rect 6710 -6657 6716 -6281
rect 6540 -6669 6586 -6657
rect 6670 -6669 6716 -6657
rect 6788 -6281 6834 -6269
rect 6788 -6657 6794 -6281
rect 6828 -6657 6834 -6281
rect 6788 -6669 6834 -6657
rect 6906 -6281 6952 -6269
rect 6906 -6657 6912 -6281
rect 6946 -6657 6952 -6281
rect 6906 -6669 6952 -6657
rect 7024 -6281 7070 -6269
rect 7024 -6657 7030 -6281
rect 7064 -6657 7070 -6281
rect 7024 -6669 7070 -6657
rect 7142 -6281 7188 -6269
rect 7142 -6657 7148 -6281
rect 7182 -6657 7188 -6281
rect 7142 -6669 7188 -6657
rect 7260 -6281 7306 -6269
rect 7260 -6657 7266 -6281
rect 7300 -6657 7306 -6281
rect 7260 -6669 7306 -6657
rect 7378 -6281 7424 -6269
rect 7378 -6657 7384 -6281
rect 7418 -6481 7424 -6281
rect 7749 -6469 7783 -6166
rect 8379 -6166 9852 -6123
rect 8379 -6469 8413 -6166
rect 8745 -6269 8779 -6166
rect 8981 -6269 9015 -6166
rect 9217 -6269 9251 -6166
rect 9453 -6269 9487 -6166
rect 8739 -6281 8785 -6269
rect 7507 -6481 7553 -6469
rect 7418 -6657 7513 -6481
rect 7547 -6657 7553 -6481
rect 7378 -6669 7424 -6657
rect 7507 -6669 7553 -6657
rect 7625 -6481 7671 -6469
rect 7625 -6657 7631 -6481
rect 7665 -6657 7671 -6481
rect 7625 -6669 7671 -6657
rect 7743 -6481 7789 -6469
rect 7743 -6657 7749 -6481
rect 7783 -6657 7789 -6481
rect 7743 -6669 7789 -6657
rect 7861 -6481 7907 -6469
rect 7861 -6657 7867 -6481
rect 7901 -6657 7907 -6481
rect 7861 -6669 7907 -6657
rect 8255 -6481 8301 -6469
rect 8255 -6657 8261 -6481
rect 8295 -6657 8301 -6481
rect 8255 -6669 8301 -6657
rect 8373 -6481 8419 -6469
rect 8373 -6657 8379 -6481
rect 8413 -6657 8419 -6481
rect 8373 -6669 8419 -6657
rect 8491 -6481 8537 -6469
rect 8491 -6657 8497 -6481
rect 8531 -6657 8537 -6481
rect 8491 -6669 8537 -6657
rect 8609 -6481 8655 -6469
rect 8739 -6481 8745 -6281
rect 8609 -6657 8615 -6481
rect 8649 -6657 8745 -6481
rect 8779 -6657 8785 -6281
rect 8609 -6669 8655 -6657
rect 8739 -6669 8785 -6657
rect 8857 -6281 8903 -6269
rect 8857 -6657 8863 -6281
rect 8897 -6657 8903 -6281
rect 8857 -6669 8903 -6657
rect 8975 -6281 9021 -6269
rect 8975 -6657 8981 -6281
rect 9015 -6657 9021 -6281
rect 8975 -6669 9021 -6657
rect 9093 -6281 9139 -6269
rect 9093 -6657 9099 -6281
rect 9133 -6657 9139 -6281
rect 9093 -6669 9139 -6657
rect 9211 -6281 9257 -6269
rect 9211 -6657 9217 -6281
rect 9251 -6657 9257 -6281
rect 9211 -6669 9257 -6657
rect 9329 -6281 9375 -6269
rect 9329 -6657 9335 -6281
rect 9369 -6657 9375 -6281
rect 9329 -6669 9375 -6657
rect 9447 -6281 9493 -6269
rect 9447 -6657 9453 -6281
rect 9487 -6481 9493 -6281
rect 9818 -6469 9852 -6166
rect 10447 -6164 11920 -6121
rect 13187 -6123 13321 -6072
rect 15255 -6070 15293 -6038
rect 15347 -6038 15357 -6016
rect 16837 -6017 16863 -5981
rect 16959 -6017 16995 -5981
rect 16837 -6035 16877 -6017
rect 16953 -6035 16995 -6017
rect 15347 -6070 15389 -6038
rect 15255 -6121 15389 -6070
rect 16837 -6075 16995 -6035
rect 16713 -6121 16995 -6075
rect 10447 -6467 10481 -6164
rect 10813 -6267 10847 -6164
rect 11049 -6267 11083 -6164
rect 11285 -6267 11319 -6164
rect 11521 -6267 11555 -6164
rect 10807 -6279 10853 -6267
rect 9576 -6481 9622 -6469
rect 9487 -6657 9582 -6481
rect 9616 -6657 9622 -6481
rect 9447 -6669 9493 -6657
rect 9576 -6669 9622 -6657
rect 9694 -6481 9740 -6469
rect 9694 -6657 9700 -6481
rect 9734 -6657 9740 -6481
rect 9694 -6669 9740 -6657
rect 9812 -6481 9858 -6469
rect 9812 -6657 9818 -6481
rect 9852 -6657 9858 -6481
rect 9812 -6669 9858 -6657
rect 9930 -6481 9976 -6469
rect 9930 -6657 9936 -6481
rect 9970 -6657 9976 -6481
rect 9930 -6669 9976 -6657
rect 10323 -6479 10369 -6467
rect 10323 -6655 10329 -6479
rect 10363 -6655 10369 -6479
rect 10323 -6667 10369 -6655
rect 10441 -6479 10487 -6467
rect 10441 -6655 10447 -6479
rect 10481 -6655 10487 -6479
rect 10441 -6667 10487 -6655
rect 10559 -6479 10605 -6467
rect 10559 -6655 10565 -6479
rect 10599 -6655 10605 -6479
rect 10559 -6667 10605 -6655
rect 10677 -6479 10723 -6467
rect 10807 -6479 10813 -6279
rect 10677 -6655 10683 -6479
rect 10717 -6655 10813 -6479
rect 10847 -6655 10853 -6279
rect 10677 -6667 10723 -6655
rect 10807 -6667 10853 -6655
rect 10925 -6279 10971 -6267
rect 10925 -6655 10931 -6279
rect 10965 -6655 10971 -6279
rect 10925 -6667 10971 -6655
rect 11043 -6279 11089 -6267
rect 11043 -6655 11049 -6279
rect 11083 -6655 11089 -6279
rect 11043 -6667 11089 -6655
rect 11161 -6279 11207 -6267
rect 11161 -6655 11167 -6279
rect 11201 -6655 11207 -6279
rect 11161 -6667 11207 -6655
rect 11279 -6279 11325 -6267
rect 11279 -6655 11285 -6279
rect 11319 -6655 11325 -6279
rect 11279 -6667 11325 -6655
rect 11397 -6279 11443 -6267
rect 11397 -6655 11403 -6279
rect 11437 -6655 11443 -6279
rect 11397 -6667 11443 -6655
rect 11515 -6279 11561 -6267
rect 11515 -6655 11521 -6279
rect 11555 -6479 11561 -6279
rect 11886 -6467 11920 -6164
rect 12516 -6166 13989 -6123
rect 11644 -6479 11690 -6467
rect 11555 -6655 11650 -6479
rect 11684 -6655 11690 -6479
rect 11515 -6667 11561 -6655
rect 11644 -6667 11690 -6655
rect 11762 -6479 11808 -6467
rect 11762 -6655 11768 -6479
rect 11802 -6655 11808 -6479
rect 11762 -6667 11808 -6655
rect 11880 -6479 11926 -6467
rect 11880 -6655 11886 -6479
rect 11920 -6655 11926 -6479
rect 11880 -6667 11926 -6655
rect 11998 -6479 12044 -6467
rect 12516 -6469 12550 -6166
rect 12882 -6269 12916 -6166
rect 13118 -6269 13152 -6166
rect 13354 -6269 13388 -6166
rect 13590 -6269 13624 -6166
rect 12876 -6281 12922 -6269
rect 11998 -6655 12004 -6479
rect 12038 -6655 12044 -6479
rect 11998 -6667 12044 -6655
rect 12392 -6481 12438 -6469
rect 12392 -6657 12398 -6481
rect 12432 -6657 12438 -6481
rect 3494 -6738 3764 -6703
rect 4124 -6705 4158 -6671
rect 4726 -6705 4760 -6671
rect 4962 -6705 4996 -6671
rect -713 -6873 -703 -6813
rect -639 -6873 -629 -6813
rect -284 -6829 6 -6822
rect -703 -8445 -639 -6873
rect -290 -6882 -280 -6829
rect -220 -6882 6 -6829
rect -284 -6888 6 -6882
rect 72 -6888 82 -6822
rect -19 -7012 -9 -7010
rect -284 -7021 -9 -7012
rect -290 -7079 -280 -7021
rect -228 -7079 -9 -7021
rect -284 -7084 -9 -7079
rect -19 -7087 -9 -7084
rect 62 -7087 72 -7010
rect 112 -7524 146 -6740
rect 825 -6802 859 -6740
rect 414 -6840 1156 -6802
rect 414 -6964 448 -6840
rect 650 -6964 684 -6840
rect 886 -6964 920 -6840
rect 1122 -6964 1156 -6840
rect 1382 -6828 1460 -6822
rect 1382 -6882 1394 -6828
rect 1448 -6882 1460 -6828
rect 1382 -6888 1460 -6882
rect 408 -6976 454 -6964
rect 408 -7352 414 -6976
rect 448 -7352 454 -6976
rect 408 -7364 454 -7352
rect 526 -6976 572 -6964
rect 526 -7352 532 -6976
rect 566 -7352 572 -6976
rect 526 -7364 572 -7352
rect 644 -6976 690 -6964
rect 644 -7352 650 -6976
rect 684 -7352 690 -6976
rect 644 -7364 690 -7352
rect 762 -6976 808 -6964
rect 762 -7352 768 -6976
rect 802 -7352 808 -6976
rect 762 -7364 808 -7352
rect 880 -6976 926 -6964
rect 880 -7352 886 -6976
rect 920 -7352 926 -6976
rect 880 -7364 926 -7352
rect 998 -6976 1044 -6964
rect 998 -7352 1004 -6976
rect 1038 -7352 1044 -6976
rect 998 -7364 1044 -7352
rect 1116 -6976 1162 -6964
rect 1116 -7352 1122 -6976
rect 1156 -7352 1162 -6976
rect 1116 -7364 1162 -7352
rect 1528 -7523 1562 -6740
rect 2000 -6886 2074 -6820
rect 2140 -6886 2150 -6820
rect 2000 -7016 2140 -7010
rect 2000 -7076 2062 -7016
rect 2128 -7076 2140 -7016
rect 2000 -7082 2140 -7076
rect 1614 -7380 1740 -7374
rect 1614 -7482 1626 -7380
rect 1728 -7482 1740 -7380
rect 1614 -7488 1740 -7482
rect 1255 -7524 1562 -7523
rect 112 -7529 428 -7524
rect 1142 -7529 1562 -7524
rect 112 -7540 495 -7529
rect 112 -7567 444 -7540
rect 112 -7696 146 -7567
rect 428 -7574 444 -7567
rect 478 -7574 495 -7540
rect 428 -7580 495 -7574
rect 1075 -7540 1562 -7529
rect 1075 -7574 1092 -7540
rect 1126 -7567 1562 -7540
rect 1126 -7574 1142 -7567
rect 1255 -7568 1562 -7567
rect 1075 -7580 1142 -7574
rect 253 -7607 309 -7595
rect 253 -7641 259 -7607
rect 293 -7608 309 -7607
rect 1366 -7608 1422 -7596
rect 293 -7624 760 -7608
rect 293 -7641 710 -7624
rect 253 -7657 710 -7641
rect 694 -7658 710 -7657
rect 744 -7658 760 -7624
rect 694 -7665 760 -7658
rect 812 -7623 1382 -7608
rect 812 -7657 828 -7623
rect 862 -7642 1382 -7623
rect 1416 -7642 1422 -7608
rect 862 -7657 1422 -7642
rect 812 -7667 879 -7657
rect 1366 -7658 1422 -7657
rect 1528 -7696 1562 -7568
rect 106 -7708 152 -7696
rect 106 -7884 112 -7708
rect 146 -7884 152 -7708
rect 106 -7896 152 -7884
rect 224 -7708 270 -7696
rect 224 -7884 230 -7708
rect 264 -7884 270 -7708
rect 224 -7896 270 -7884
rect 526 -7708 572 -7696
rect 229 -8190 263 -7896
rect 526 -8084 532 -7708
rect 566 -8084 572 -7708
rect 526 -8096 572 -8084
rect 644 -7708 690 -7696
rect 644 -8084 650 -7708
rect 684 -8084 690 -7708
rect 644 -8096 690 -8084
rect 762 -7708 808 -7696
rect 762 -8084 768 -7708
rect 802 -8084 808 -7708
rect 762 -8096 808 -8084
rect 880 -7708 926 -7696
rect 880 -8084 886 -7708
rect 920 -8084 926 -7708
rect 880 -8096 926 -8084
rect 998 -7708 1044 -7696
rect 998 -8084 1004 -7708
rect 1038 -8084 1044 -7708
rect 1404 -7708 1450 -7696
rect 1404 -7884 1410 -7708
rect 1444 -7884 1450 -7708
rect 1404 -7896 1450 -7884
rect 1522 -7708 1568 -7696
rect 1522 -7884 1528 -7708
rect 1562 -7884 1568 -7708
rect 1522 -7896 1568 -7884
rect 998 -8096 1044 -8084
rect 886 -8190 920 -8096
rect 1410 -8190 1443 -7896
rect 229 -8222 1443 -8190
rect 722 -8244 854 -8222
rect 722 -8302 756 -8244
rect 818 -8302 854 -8244
rect 722 -8307 854 -8302
rect 2000 -8445 2064 -7082
rect 2180 -7522 2214 -6738
rect 2893 -6800 2927 -6738
rect 2482 -6838 3224 -6800
rect 2482 -6962 2516 -6838
rect 2718 -6962 2752 -6838
rect 2954 -6962 2988 -6838
rect 3190 -6962 3224 -6838
rect 3450 -6826 3528 -6820
rect 3450 -6880 3462 -6826
rect 3516 -6880 3528 -6826
rect 3450 -6886 3528 -6880
rect 2476 -6974 2522 -6962
rect 2476 -7350 2482 -6974
rect 2516 -7350 2522 -6974
rect 2476 -7362 2522 -7350
rect 2594 -6974 2640 -6962
rect 2594 -7350 2600 -6974
rect 2634 -7350 2640 -6974
rect 2594 -7362 2640 -7350
rect 2712 -6974 2758 -6962
rect 2712 -7350 2718 -6974
rect 2752 -7350 2758 -6974
rect 2712 -7362 2758 -7350
rect 2830 -6974 2876 -6962
rect 2830 -7350 2836 -6974
rect 2870 -7350 2876 -6974
rect 2830 -7362 2876 -7350
rect 2948 -6974 2994 -6962
rect 2948 -7350 2954 -6974
rect 2988 -7350 2994 -6974
rect 2948 -7362 2994 -7350
rect 3066 -6974 3112 -6962
rect 3066 -7350 3072 -6974
rect 3106 -7350 3112 -6974
rect 3066 -7362 3112 -7350
rect 3184 -6974 3230 -6962
rect 3184 -7350 3190 -6974
rect 3224 -7350 3230 -6974
rect 3184 -7362 3230 -7350
rect 3596 -7521 3630 -6738
rect 4124 -6740 4283 -6705
rect 4726 -6740 4996 -6705
rect 5563 -6705 5597 -6671
rect 5799 -6705 5833 -6671
rect 5563 -6740 5833 -6705
rect 6192 -6703 6226 -6669
rect 6794 -6703 6828 -6669
rect 7030 -6703 7064 -6669
rect 6192 -6738 6351 -6703
rect 6794 -6738 7064 -6703
rect 7631 -6703 7665 -6669
rect 7867 -6703 7901 -6669
rect 7631 -6738 7901 -6703
rect 8261 -6703 8295 -6669
rect 8863 -6703 8897 -6669
rect 9099 -6703 9133 -6669
rect 8261 -6738 8420 -6703
rect 8863 -6738 9133 -6703
rect 9700 -6703 9734 -6669
rect 9936 -6703 9970 -6669
rect 9700 -6738 9970 -6703
rect 10329 -6701 10363 -6667
rect 10931 -6701 10965 -6667
rect 11167 -6701 11201 -6667
rect 10329 -6736 10488 -6701
rect 10931 -6736 11201 -6701
rect 11768 -6701 11802 -6667
rect 12004 -6701 12038 -6667
rect 12392 -6669 12438 -6657
rect 12510 -6481 12556 -6469
rect 12510 -6657 12516 -6481
rect 12550 -6657 12556 -6481
rect 12510 -6669 12556 -6657
rect 12628 -6481 12674 -6469
rect 12628 -6657 12634 -6481
rect 12668 -6657 12674 -6481
rect 12628 -6669 12674 -6657
rect 12746 -6481 12792 -6469
rect 12876 -6481 12882 -6281
rect 12746 -6657 12752 -6481
rect 12786 -6657 12882 -6481
rect 12916 -6657 12922 -6281
rect 12746 -6669 12792 -6657
rect 12876 -6669 12922 -6657
rect 12994 -6281 13040 -6269
rect 12994 -6657 13000 -6281
rect 13034 -6657 13040 -6281
rect 12994 -6669 13040 -6657
rect 13112 -6281 13158 -6269
rect 13112 -6657 13118 -6281
rect 13152 -6657 13158 -6281
rect 13112 -6669 13158 -6657
rect 13230 -6281 13276 -6269
rect 13230 -6657 13236 -6281
rect 13270 -6657 13276 -6281
rect 13230 -6669 13276 -6657
rect 13348 -6281 13394 -6269
rect 13348 -6657 13354 -6281
rect 13388 -6657 13394 -6281
rect 13348 -6669 13394 -6657
rect 13466 -6281 13512 -6269
rect 13466 -6657 13472 -6281
rect 13506 -6657 13512 -6281
rect 13466 -6669 13512 -6657
rect 13584 -6281 13630 -6269
rect 13584 -6657 13590 -6281
rect 13624 -6481 13630 -6281
rect 13955 -6469 13989 -6166
rect 14584 -6164 16057 -6121
rect 14584 -6467 14618 -6164
rect 14950 -6267 14984 -6164
rect 15186 -6267 15220 -6164
rect 15422 -6267 15456 -6164
rect 15658 -6267 15692 -6164
rect 14944 -6279 14990 -6267
rect 13713 -6481 13759 -6469
rect 13624 -6657 13719 -6481
rect 13753 -6657 13759 -6481
rect 13584 -6669 13630 -6657
rect 13713 -6669 13759 -6657
rect 13831 -6481 13877 -6469
rect 13831 -6657 13837 -6481
rect 13871 -6657 13877 -6481
rect 13831 -6669 13877 -6657
rect 13949 -6481 13995 -6469
rect 13949 -6657 13955 -6481
rect 13989 -6657 13995 -6481
rect 13949 -6669 13995 -6657
rect 14067 -6481 14113 -6469
rect 14067 -6657 14073 -6481
rect 14107 -6657 14113 -6481
rect 14067 -6669 14113 -6657
rect 14460 -6479 14506 -6467
rect 14460 -6655 14466 -6479
rect 14500 -6655 14506 -6479
rect 14460 -6667 14506 -6655
rect 14578 -6479 14624 -6467
rect 14578 -6655 14584 -6479
rect 14618 -6655 14624 -6479
rect 14578 -6667 14624 -6655
rect 14696 -6479 14742 -6467
rect 14696 -6655 14702 -6479
rect 14736 -6655 14742 -6479
rect 14696 -6667 14742 -6655
rect 14814 -6479 14860 -6467
rect 14944 -6479 14950 -6279
rect 14814 -6655 14820 -6479
rect 14854 -6655 14950 -6479
rect 14984 -6655 14990 -6279
rect 14814 -6667 14860 -6655
rect 14944 -6667 14990 -6655
rect 15062 -6279 15108 -6267
rect 15062 -6655 15068 -6279
rect 15102 -6655 15108 -6279
rect 15062 -6667 15108 -6655
rect 15180 -6279 15226 -6267
rect 15180 -6655 15186 -6279
rect 15220 -6655 15226 -6279
rect 15180 -6667 15226 -6655
rect 15298 -6279 15344 -6267
rect 15298 -6655 15304 -6279
rect 15338 -6655 15344 -6279
rect 15298 -6667 15344 -6655
rect 15416 -6279 15462 -6267
rect 15416 -6655 15422 -6279
rect 15456 -6655 15462 -6279
rect 15416 -6667 15462 -6655
rect 15534 -6279 15580 -6267
rect 15534 -6655 15540 -6279
rect 15574 -6655 15580 -6279
rect 15534 -6667 15580 -6655
rect 15652 -6279 15698 -6267
rect 15652 -6655 15658 -6279
rect 15692 -6479 15698 -6279
rect 16023 -6467 16057 -6164
rect 16713 -6167 16759 -6121
rect 16713 -6343 16719 -6167
rect 16753 -6343 16759 -6167
rect 16713 -6355 16759 -6343
rect 16831 -6167 16877 -6155
rect 16831 -6343 16837 -6167
rect 16871 -6343 16877 -6167
rect 16831 -6355 16877 -6343
rect 16949 -6167 16995 -6121
rect 16949 -6343 16955 -6167
rect 16989 -6343 16995 -6167
rect 16949 -6355 16995 -6343
rect 17067 -6167 17113 -6155
rect 17067 -6343 17073 -6167
rect 17107 -6343 17113 -6167
rect 17067 -6345 17113 -6343
rect 17067 -6432 17115 -6345
rect 17143 -6432 17207 -5863
rect 17605 -5977 17615 -5963
rect 17575 -5983 17615 -5977
rect 17691 -5977 17701 -5963
rect 17691 -5983 17733 -5977
rect 17575 -6019 17601 -5983
rect 17697 -6019 17733 -5983
rect 17575 -6037 17615 -6019
rect 17691 -6037 17733 -6019
rect 17575 -6077 17733 -6037
rect 17451 -6123 17733 -6077
rect 17451 -6163 17497 -6123
rect 17451 -6339 17457 -6163
rect 17491 -6339 17497 -6163
rect 17451 -6351 17497 -6339
rect 17569 -6163 17615 -6151
rect 17569 -6339 17575 -6163
rect 17609 -6339 17615 -6163
rect 17569 -6351 17615 -6339
rect 17687 -6163 17733 -6123
rect 17687 -6339 17693 -6163
rect 17727 -6339 17733 -6163
rect 17687 -6351 17733 -6339
rect 17805 -6163 17851 -6151
rect 17805 -6339 17811 -6163
rect 17845 -6339 17851 -6163
rect 17805 -6347 17851 -6339
rect 17805 -6430 17853 -6347
rect 17887 -6430 17951 -5754
rect 18589 -5727 18637 -5671
rect 18589 -5755 18676 -5727
rect 18343 -5977 18353 -5963
rect 18313 -5983 18353 -5977
rect 18429 -5977 18439 -5963
rect 18429 -5983 18471 -5977
rect 18313 -6019 18339 -5983
rect 18435 -6019 18471 -5983
rect 18313 -6037 18353 -6019
rect 18429 -6037 18471 -6019
rect 18313 -6077 18471 -6037
rect 18189 -6123 18471 -6077
rect 18189 -6167 18235 -6123
rect 18189 -6343 18195 -6167
rect 18229 -6343 18235 -6167
rect 18189 -6355 18235 -6343
rect 18307 -6167 18353 -6155
rect 18307 -6343 18313 -6167
rect 18347 -6343 18353 -6167
rect 18307 -6355 18353 -6343
rect 18425 -6167 18471 -6123
rect 18425 -6343 18431 -6167
rect 18465 -6343 18471 -6167
rect 18425 -6355 18471 -6343
rect 18543 -6167 18589 -6155
rect 18543 -6343 18549 -6167
rect 18583 -6343 18589 -6167
rect 18543 -6347 18589 -6343
rect 18543 -6428 18591 -6347
rect 18628 -6428 18676 -5755
rect 19085 -5977 19095 -5963
rect 19055 -5983 19095 -5977
rect 19171 -5977 19181 -5963
rect 19171 -5983 19213 -5977
rect 19055 -6019 19081 -5983
rect 19177 -6019 19213 -5983
rect 19055 -6037 19095 -6019
rect 19171 -6037 19213 -6019
rect 19055 -6077 19213 -6037
rect 18931 -6123 19213 -6077
rect 18931 -6169 18977 -6123
rect 18931 -6345 18937 -6169
rect 18971 -6345 18977 -6169
rect 18931 -6357 18977 -6345
rect 19049 -6169 19095 -6157
rect 19049 -6345 19055 -6169
rect 19089 -6345 19095 -6169
rect 19049 -6357 19095 -6345
rect 19167 -6169 19213 -6123
rect 19167 -6345 19173 -6169
rect 19207 -6345 19213 -6169
rect 19167 -6357 19213 -6345
rect 19285 -6169 19331 -6157
rect 19285 -6345 19291 -6169
rect 19325 -6345 19331 -6169
rect 19285 -6347 19331 -6345
rect 16864 -6449 16941 -6443
rect 15781 -6479 15827 -6467
rect 15692 -6655 15787 -6479
rect 15821 -6655 15827 -6479
rect 15652 -6667 15698 -6655
rect 15781 -6667 15827 -6655
rect 15899 -6479 15945 -6467
rect 15899 -6655 15905 -6479
rect 15939 -6655 15945 -6479
rect 15899 -6667 15945 -6655
rect 16017 -6479 16063 -6467
rect 16017 -6655 16023 -6479
rect 16057 -6655 16063 -6479
rect 16017 -6667 16063 -6655
rect 16135 -6479 16181 -6467
rect 16135 -6655 16141 -6479
rect 16175 -6655 16181 -6479
rect 16864 -6483 16895 -6449
rect 16929 -6483 16941 -6449
rect 16864 -6489 16941 -6483
rect 17063 -6493 17207 -6432
rect 17593 -6451 17679 -6445
rect 17593 -6485 17633 -6451
rect 17667 -6485 17679 -6451
rect 17593 -6491 17679 -6485
rect 17067 -6537 17115 -6493
rect 17801 -6494 17951 -6430
rect 18338 -6451 18417 -6445
rect 18338 -6485 18371 -6451
rect 18405 -6485 18417 -6451
rect 18338 -6491 18417 -6485
rect 18539 -6490 18676 -6428
rect 19285 -6429 19333 -6347
rect 19381 -6429 19445 -5666
rect 19825 -5977 19835 -5963
rect 19795 -5983 19835 -5977
rect 19911 -5977 19921 -5963
rect 19911 -5983 19953 -5977
rect 19795 -6019 19821 -5983
rect 19917 -6019 19953 -5983
rect 19795 -6037 19835 -6019
rect 19911 -6037 19953 -6019
rect 19795 -6077 19953 -6037
rect 19671 -6123 19953 -6077
rect 19671 -6169 19717 -6123
rect 19671 -6345 19677 -6169
rect 19711 -6345 19717 -6169
rect 19671 -6357 19717 -6345
rect 19789 -6169 19835 -6157
rect 19789 -6345 19795 -6169
rect 19829 -6345 19835 -6169
rect 19789 -6357 19835 -6345
rect 19907 -6169 19953 -6123
rect 19907 -6345 19913 -6169
rect 19947 -6345 19953 -6169
rect 19907 -6357 19953 -6345
rect 20025 -6169 20071 -6157
rect 20025 -6345 20031 -6169
rect 20065 -6345 20071 -6169
rect 20025 -6347 20071 -6345
rect 20025 -6429 20073 -6347
rect 20125 -6429 20189 -5590
rect 20563 -5977 20573 -5963
rect 20533 -5983 20573 -5977
rect 20649 -5977 20659 -5963
rect 20649 -5983 20691 -5977
rect 20533 -6019 20559 -5983
rect 20655 -6019 20691 -5983
rect 20533 -6037 20573 -6019
rect 20649 -6037 20691 -6019
rect 20533 -6077 20691 -6037
rect 20409 -6123 20691 -6077
rect 20409 -6169 20455 -6123
rect 20409 -6345 20415 -6169
rect 20449 -6345 20455 -6169
rect 20409 -6357 20455 -6345
rect 20527 -6169 20573 -6157
rect 20527 -6345 20533 -6169
rect 20567 -6345 20573 -6169
rect 20527 -6357 20573 -6345
rect 20645 -6169 20691 -6123
rect 20645 -6345 20651 -6169
rect 20685 -6345 20691 -6169
rect 20645 -6357 20691 -6345
rect 20763 -6169 20809 -6157
rect 20763 -6345 20769 -6169
rect 20803 -6345 20809 -6169
rect 20763 -6347 20809 -6345
rect 20763 -6429 20811 -6347
rect 20858 -6429 20922 -5512
rect 21301 -5977 21311 -5963
rect 21271 -5983 21311 -5977
rect 21387 -5977 21397 -5963
rect 21387 -5983 21429 -5977
rect 21271 -6019 21297 -5983
rect 21393 -6019 21429 -5983
rect 21271 -6037 21311 -6019
rect 21387 -6037 21429 -6019
rect 21271 -6077 21429 -6037
rect 21147 -6123 21429 -6077
rect 21147 -6169 21193 -6123
rect 21147 -6345 21153 -6169
rect 21187 -6345 21193 -6169
rect 21147 -6357 21193 -6345
rect 21265 -6169 21311 -6157
rect 21265 -6345 21271 -6169
rect 21305 -6345 21311 -6169
rect 21265 -6357 21311 -6345
rect 21383 -6169 21429 -6123
rect 21383 -6345 21389 -6169
rect 21423 -6345 21429 -6169
rect 21383 -6357 21429 -6345
rect 21501 -6169 21547 -6157
rect 21501 -6345 21507 -6169
rect 21541 -6345 21547 -6169
rect 21501 -6347 21547 -6345
rect 19079 -6451 19159 -6445
rect 19079 -6485 19113 -6451
rect 19147 -6485 19159 -6451
rect 16135 -6667 16181 -6655
rect 16831 -6553 16877 -6541
rect 11768 -6736 12038 -6701
rect 12398 -6703 12432 -6669
rect 13000 -6703 13034 -6669
rect 13236 -6703 13270 -6669
rect 4069 -6888 4143 -6822
rect 4209 -6888 4219 -6822
rect 4034 -7018 4209 -7012
rect 4034 -7078 4131 -7018
rect 4197 -7078 4209 -7018
rect 4034 -7084 4209 -7078
rect 3682 -7378 3808 -7372
rect 3682 -7480 3694 -7378
rect 3796 -7480 3808 -7378
rect 3682 -7486 3808 -7480
rect 3323 -7522 3630 -7521
rect 2180 -7527 2496 -7522
rect 3210 -7527 3630 -7522
rect 2180 -7538 2563 -7527
rect 2180 -7565 2512 -7538
rect 2180 -7694 2214 -7565
rect 2496 -7572 2512 -7565
rect 2546 -7572 2563 -7538
rect 2496 -7578 2563 -7572
rect 3143 -7538 3630 -7527
rect 3143 -7572 3160 -7538
rect 3194 -7565 3630 -7538
rect 3194 -7572 3210 -7565
rect 3323 -7566 3630 -7565
rect 3143 -7578 3210 -7572
rect 2321 -7605 2377 -7593
rect 2321 -7639 2327 -7605
rect 2361 -7606 2377 -7605
rect 3434 -7606 3490 -7594
rect 2361 -7622 2828 -7606
rect 2361 -7639 2778 -7622
rect 2321 -7655 2778 -7639
rect 2762 -7656 2778 -7655
rect 2812 -7656 2828 -7622
rect 2762 -7663 2828 -7656
rect 2880 -7621 3450 -7606
rect 2880 -7655 2896 -7621
rect 2930 -7640 3450 -7621
rect 3484 -7640 3490 -7606
rect 2930 -7655 3490 -7640
rect 2880 -7665 2947 -7655
rect 3434 -7656 3490 -7655
rect 3596 -7694 3630 -7566
rect 2174 -7706 2220 -7694
rect 2174 -7882 2180 -7706
rect 2214 -7882 2220 -7706
rect 2174 -7894 2220 -7882
rect 2292 -7706 2338 -7694
rect 2292 -7882 2298 -7706
rect 2332 -7882 2338 -7706
rect 2292 -7894 2338 -7882
rect 2594 -7706 2640 -7694
rect 2297 -8188 2331 -7894
rect 2594 -8082 2600 -7706
rect 2634 -8082 2640 -7706
rect 2594 -8094 2640 -8082
rect 2712 -7706 2758 -7694
rect 2712 -8082 2718 -7706
rect 2752 -8082 2758 -7706
rect 2712 -8094 2758 -8082
rect 2830 -7706 2876 -7694
rect 2830 -8082 2836 -7706
rect 2870 -8082 2876 -7706
rect 2830 -8094 2876 -8082
rect 2948 -7706 2994 -7694
rect 2948 -8082 2954 -7706
rect 2988 -8082 2994 -7706
rect 2948 -8094 2994 -8082
rect 3066 -7706 3112 -7694
rect 3066 -8082 3072 -7706
rect 3106 -8082 3112 -7706
rect 3472 -7706 3518 -7694
rect 3472 -7882 3478 -7706
rect 3512 -7882 3518 -7706
rect 3472 -7894 3518 -7882
rect 3590 -7706 3636 -7694
rect 3590 -7882 3596 -7706
rect 3630 -7882 3636 -7706
rect 3590 -7894 3636 -7882
rect 3066 -8094 3112 -8082
rect 2954 -8188 2988 -8094
rect 3478 -8188 3511 -7894
rect 2297 -8220 3511 -8188
rect 2790 -8242 2922 -8220
rect 2790 -8300 2824 -8242
rect 2886 -8300 2922 -8242
rect 2790 -8305 2922 -8300
rect -703 -8509 2065 -8445
rect -703 -8510 -398 -8509
rect 2000 -8653 2064 -8509
rect 1995 -8659 2070 -8653
rect 1995 -8710 2007 -8659
rect 2058 -8710 2070 -8659
rect 1995 -8716 2070 -8710
rect 4034 -8756 4098 -7084
rect 4249 -7524 4283 -6740
rect 4962 -6802 4996 -6740
rect 4551 -6840 5293 -6802
rect 4551 -6964 4585 -6840
rect 4787 -6964 4821 -6840
rect 5023 -6964 5057 -6840
rect 5259 -6964 5293 -6840
rect 5519 -6828 5597 -6822
rect 5519 -6882 5531 -6828
rect 5585 -6882 5597 -6828
rect 5519 -6888 5597 -6882
rect 4545 -6976 4591 -6964
rect 4545 -7352 4551 -6976
rect 4585 -7352 4591 -6976
rect 4545 -7364 4591 -7352
rect 4663 -6976 4709 -6964
rect 4663 -7352 4669 -6976
rect 4703 -7352 4709 -6976
rect 4663 -7364 4709 -7352
rect 4781 -6976 4827 -6964
rect 4781 -7352 4787 -6976
rect 4821 -7352 4827 -6976
rect 4781 -7364 4827 -7352
rect 4899 -6976 4945 -6964
rect 4899 -7352 4905 -6976
rect 4939 -7352 4945 -6976
rect 4899 -7364 4945 -7352
rect 5017 -6976 5063 -6964
rect 5017 -7352 5023 -6976
rect 5057 -7352 5063 -6976
rect 5017 -7364 5063 -7352
rect 5135 -6976 5181 -6964
rect 5135 -7352 5141 -6976
rect 5175 -7352 5181 -6976
rect 5135 -7364 5181 -7352
rect 5253 -6976 5299 -6964
rect 5253 -7352 5259 -6976
rect 5293 -7352 5299 -6976
rect 5253 -7364 5299 -7352
rect 5665 -7523 5699 -6740
rect 6137 -6886 6211 -6820
rect 6277 -6886 6287 -6820
rect 6080 -7016 6277 -7010
rect 6080 -7076 6199 -7016
rect 6265 -7076 6277 -7016
rect 6080 -7082 6277 -7076
rect 5751 -7380 5877 -7374
rect 5751 -7482 5763 -7380
rect 5865 -7482 5877 -7380
rect 5751 -7488 5877 -7482
rect 5392 -7524 5699 -7523
rect 4249 -7529 4565 -7524
rect 5279 -7529 5699 -7524
rect 4249 -7540 4632 -7529
rect 4249 -7567 4581 -7540
rect 4249 -7696 4283 -7567
rect 4565 -7574 4581 -7567
rect 4615 -7574 4632 -7540
rect 4565 -7580 4632 -7574
rect 5212 -7540 5699 -7529
rect 5212 -7574 5229 -7540
rect 5263 -7567 5699 -7540
rect 5263 -7574 5279 -7567
rect 5392 -7568 5699 -7567
rect 5212 -7580 5279 -7574
rect 4390 -7607 4446 -7595
rect 4390 -7641 4396 -7607
rect 4430 -7608 4446 -7607
rect 5503 -7608 5559 -7596
rect 4430 -7624 4897 -7608
rect 4430 -7641 4847 -7624
rect 4390 -7657 4847 -7641
rect 4831 -7658 4847 -7657
rect 4881 -7658 4897 -7624
rect 4831 -7665 4897 -7658
rect 4949 -7623 5519 -7608
rect 4949 -7657 4965 -7623
rect 4999 -7642 5519 -7623
rect 5553 -7642 5559 -7608
rect 4999 -7657 5559 -7642
rect 4949 -7667 5016 -7657
rect 5503 -7658 5559 -7657
rect 5665 -7696 5699 -7568
rect 4243 -7708 4289 -7696
rect 4243 -7884 4249 -7708
rect 4283 -7884 4289 -7708
rect 4243 -7896 4289 -7884
rect 4361 -7708 4407 -7696
rect 4361 -7884 4367 -7708
rect 4401 -7884 4407 -7708
rect 4361 -7896 4407 -7884
rect 4663 -7708 4709 -7696
rect 4366 -8190 4400 -7896
rect 4663 -8084 4669 -7708
rect 4703 -8084 4709 -7708
rect 4663 -8096 4709 -8084
rect 4781 -7708 4827 -7696
rect 4781 -8084 4787 -7708
rect 4821 -8084 4827 -7708
rect 4781 -8096 4827 -8084
rect 4899 -7708 4945 -7696
rect 4899 -8084 4905 -7708
rect 4939 -8084 4945 -7708
rect 4899 -8096 4945 -8084
rect 5017 -7708 5063 -7696
rect 5017 -8084 5023 -7708
rect 5057 -8084 5063 -7708
rect 5017 -8096 5063 -8084
rect 5135 -7708 5181 -7696
rect 5135 -8084 5141 -7708
rect 5175 -8084 5181 -7708
rect 5541 -7708 5587 -7696
rect 5541 -7884 5547 -7708
rect 5581 -7884 5587 -7708
rect 5541 -7896 5587 -7884
rect 5659 -7708 5705 -7696
rect 5659 -7884 5665 -7708
rect 5699 -7884 5705 -7708
rect 5659 -7896 5705 -7884
rect 5135 -8096 5181 -8084
rect 5023 -8190 5057 -8096
rect 5547 -8190 5580 -7896
rect 4366 -8222 5580 -8190
rect 4859 -8244 4991 -8222
rect 4859 -8302 4893 -8244
rect 4955 -8302 4991 -8244
rect 4859 -8307 4991 -8302
rect -933 -8764 4098 -8756
rect -933 -8818 4042 -8764
rect 4089 -8818 4098 -8764
rect -933 -8837 4098 -8818
rect 6080 -8865 6144 -7082
rect 6317 -7522 6351 -6738
rect 7030 -6800 7064 -6738
rect 6619 -6838 7361 -6800
rect 6619 -6962 6653 -6838
rect 6855 -6962 6889 -6838
rect 7091 -6962 7125 -6838
rect 7327 -6962 7361 -6838
rect 7587 -6826 7665 -6820
rect 7587 -6880 7599 -6826
rect 7653 -6880 7665 -6826
rect 7587 -6886 7665 -6880
rect 6613 -6974 6659 -6962
rect 6613 -7350 6619 -6974
rect 6653 -7350 6659 -6974
rect 6613 -7362 6659 -7350
rect 6731 -6974 6777 -6962
rect 6731 -7350 6737 -6974
rect 6771 -7350 6777 -6974
rect 6731 -7362 6777 -7350
rect 6849 -6974 6895 -6962
rect 6849 -7350 6855 -6974
rect 6889 -7350 6895 -6974
rect 6849 -7362 6895 -7350
rect 6967 -6974 7013 -6962
rect 6967 -7350 6973 -6974
rect 7007 -7350 7013 -6974
rect 6967 -7362 7013 -7350
rect 7085 -6974 7131 -6962
rect 7085 -7350 7091 -6974
rect 7125 -7350 7131 -6974
rect 7085 -7362 7131 -7350
rect 7203 -6974 7249 -6962
rect 7203 -7350 7209 -6974
rect 7243 -7350 7249 -6974
rect 7203 -7362 7249 -7350
rect 7321 -6974 7367 -6962
rect 7321 -7350 7327 -6974
rect 7361 -7350 7367 -6974
rect 7321 -7362 7367 -7350
rect 7733 -7521 7767 -6738
rect 8206 -6886 8280 -6820
rect 8346 -6886 8356 -6820
rect 8170 -7016 8346 -7010
rect 8170 -7076 8268 -7016
rect 8334 -7076 8346 -7016
rect 8170 -7082 8346 -7076
rect 7819 -7378 7945 -7372
rect 7819 -7480 7831 -7378
rect 7933 -7480 7945 -7378
rect 7819 -7486 7945 -7480
rect 7460 -7522 7767 -7521
rect 6317 -7527 6633 -7522
rect 7347 -7527 7767 -7522
rect 6317 -7538 6700 -7527
rect 6317 -7565 6649 -7538
rect 6317 -7694 6351 -7565
rect 6633 -7572 6649 -7565
rect 6683 -7572 6700 -7538
rect 6633 -7578 6700 -7572
rect 7280 -7538 7767 -7527
rect 7280 -7572 7297 -7538
rect 7331 -7565 7767 -7538
rect 7331 -7572 7347 -7565
rect 7460 -7566 7767 -7565
rect 7280 -7578 7347 -7572
rect 6458 -7605 6514 -7593
rect 6458 -7639 6464 -7605
rect 6498 -7606 6514 -7605
rect 7571 -7606 7627 -7594
rect 6498 -7622 6965 -7606
rect 6498 -7639 6915 -7622
rect 6458 -7655 6915 -7639
rect 6899 -7656 6915 -7655
rect 6949 -7656 6965 -7622
rect 6899 -7663 6965 -7656
rect 7017 -7621 7587 -7606
rect 7017 -7655 7033 -7621
rect 7067 -7640 7587 -7621
rect 7621 -7640 7627 -7606
rect 7067 -7655 7627 -7640
rect 7017 -7665 7084 -7655
rect 7571 -7656 7627 -7655
rect 7733 -7694 7767 -7566
rect 6311 -7706 6357 -7694
rect 6311 -7882 6317 -7706
rect 6351 -7882 6357 -7706
rect 6311 -7894 6357 -7882
rect 6429 -7706 6475 -7694
rect 6429 -7882 6435 -7706
rect 6469 -7882 6475 -7706
rect 6429 -7894 6475 -7882
rect 6731 -7706 6777 -7694
rect 6434 -8188 6468 -7894
rect 6731 -8082 6737 -7706
rect 6771 -8082 6777 -7706
rect 6731 -8094 6777 -8082
rect 6849 -7706 6895 -7694
rect 6849 -8082 6855 -7706
rect 6889 -8082 6895 -7706
rect 6849 -8094 6895 -8082
rect 6967 -7706 7013 -7694
rect 6967 -8082 6973 -7706
rect 7007 -8082 7013 -7706
rect 6967 -8094 7013 -8082
rect 7085 -7706 7131 -7694
rect 7085 -8082 7091 -7706
rect 7125 -8082 7131 -7706
rect 7085 -8094 7131 -8082
rect 7203 -7706 7249 -7694
rect 7203 -8082 7209 -7706
rect 7243 -8082 7249 -7706
rect 7609 -7706 7655 -7694
rect 7609 -7882 7615 -7706
rect 7649 -7882 7655 -7706
rect 7609 -7894 7655 -7882
rect 7727 -7706 7773 -7694
rect 7727 -7882 7733 -7706
rect 7767 -7882 7773 -7706
rect 7727 -7894 7773 -7882
rect 7203 -8094 7249 -8082
rect 7091 -8188 7125 -8094
rect 7615 -8188 7648 -7894
rect 6434 -8220 7648 -8188
rect 6927 -8242 7059 -8220
rect 6927 -8300 6961 -8242
rect 7023 -8300 7059 -8242
rect 6927 -8305 7059 -8300
rect -1130 -8867 6144 -8865
rect -1130 -8921 6089 -8867
rect 6136 -8921 6144 -8867
rect -1130 -8957 6144 -8921
rect 8170 -8965 8234 -7082
rect 8386 -7522 8420 -6738
rect 9099 -6800 9133 -6738
rect 8688 -6838 9430 -6800
rect 8688 -6962 8722 -6838
rect 8924 -6962 8958 -6838
rect 9160 -6962 9194 -6838
rect 9396 -6962 9430 -6838
rect 9656 -6826 9734 -6820
rect 9656 -6880 9668 -6826
rect 9722 -6880 9734 -6826
rect 9656 -6886 9734 -6880
rect 8682 -6974 8728 -6962
rect 8682 -7350 8688 -6974
rect 8722 -7350 8728 -6974
rect 8682 -7362 8728 -7350
rect 8800 -6974 8846 -6962
rect 8800 -7350 8806 -6974
rect 8840 -7350 8846 -6974
rect 8800 -7362 8846 -7350
rect 8918 -6974 8964 -6962
rect 8918 -7350 8924 -6974
rect 8958 -7350 8964 -6974
rect 8918 -7362 8964 -7350
rect 9036 -6974 9082 -6962
rect 9036 -7350 9042 -6974
rect 9076 -7350 9082 -6974
rect 9036 -7362 9082 -7350
rect 9154 -6974 9200 -6962
rect 9154 -7350 9160 -6974
rect 9194 -7350 9200 -6974
rect 9154 -7362 9200 -7350
rect 9272 -6974 9318 -6962
rect 9272 -7350 9278 -6974
rect 9312 -7350 9318 -6974
rect 9272 -7362 9318 -7350
rect 9390 -6974 9436 -6962
rect 9390 -7350 9396 -6974
rect 9430 -7350 9436 -6974
rect 9390 -7362 9436 -7350
rect 9802 -7521 9836 -6738
rect 10274 -6884 10348 -6818
rect 10414 -6884 10424 -6818
rect 10244 -7014 10414 -7008
rect 10244 -7074 10336 -7014
rect 10402 -7074 10414 -7014
rect 10244 -7080 10414 -7074
rect 9888 -7378 10014 -7372
rect 9888 -7480 9900 -7378
rect 10002 -7480 10014 -7378
rect 9888 -7486 10014 -7480
rect 9529 -7522 9836 -7521
rect 8386 -7527 8702 -7522
rect 9416 -7527 9836 -7522
rect 8386 -7538 8769 -7527
rect 8386 -7565 8718 -7538
rect 8386 -7694 8420 -7565
rect 8702 -7572 8718 -7565
rect 8752 -7572 8769 -7538
rect 8702 -7578 8769 -7572
rect 9349 -7538 9836 -7527
rect 9349 -7572 9366 -7538
rect 9400 -7565 9836 -7538
rect 9400 -7572 9416 -7565
rect 9529 -7566 9836 -7565
rect 9349 -7578 9416 -7572
rect 8527 -7605 8583 -7593
rect 8527 -7639 8533 -7605
rect 8567 -7606 8583 -7605
rect 9640 -7606 9696 -7594
rect 8567 -7622 9034 -7606
rect 8567 -7639 8984 -7622
rect 8527 -7655 8984 -7639
rect 8968 -7656 8984 -7655
rect 9018 -7656 9034 -7622
rect 8968 -7663 9034 -7656
rect 9086 -7621 9656 -7606
rect 9086 -7655 9102 -7621
rect 9136 -7640 9656 -7621
rect 9690 -7640 9696 -7606
rect 9136 -7655 9696 -7640
rect 9086 -7665 9153 -7655
rect 9640 -7656 9696 -7655
rect 9802 -7694 9836 -7566
rect 8380 -7706 8426 -7694
rect 8380 -7882 8386 -7706
rect 8420 -7882 8426 -7706
rect 8380 -7894 8426 -7882
rect 8498 -7706 8544 -7694
rect 8498 -7882 8504 -7706
rect 8538 -7882 8544 -7706
rect 8498 -7894 8544 -7882
rect 8800 -7706 8846 -7694
rect 8503 -8188 8537 -7894
rect 8800 -8082 8806 -7706
rect 8840 -8082 8846 -7706
rect 8800 -8094 8846 -8082
rect 8918 -7706 8964 -7694
rect 8918 -8082 8924 -7706
rect 8958 -8082 8964 -7706
rect 8918 -8094 8964 -8082
rect 9036 -7706 9082 -7694
rect 9036 -8082 9042 -7706
rect 9076 -8082 9082 -7706
rect 9036 -8094 9082 -8082
rect 9154 -7706 9200 -7694
rect 9154 -8082 9160 -7706
rect 9194 -8082 9200 -7706
rect 9154 -8094 9200 -8082
rect 9272 -7706 9318 -7694
rect 9272 -8082 9278 -7706
rect 9312 -8082 9318 -7706
rect 9678 -7706 9724 -7694
rect 9678 -7882 9684 -7706
rect 9718 -7882 9724 -7706
rect 9678 -7894 9724 -7882
rect 9796 -7706 9842 -7694
rect 9796 -7882 9802 -7706
rect 9836 -7882 9842 -7706
rect 9796 -7894 9842 -7882
rect 9272 -8094 9318 -8082
rect 9160 -8188 9194 -8094
rect 9684 -8188 9717 -7894
rect 8503 -8220 9717 -8188
rect 8996 -8242 9128 -8220
rect 8996 -8300 9030 -8242
rect 9092 -8300 9128 -8242
rect 8996 -8305 9128 -8300
rect 8170 -8977 8235 -8965
rect -1333 -8985 -1170 -8984
rect 8170 -8985 8179 -8977
rect -1333 -9028 8179 -8985
rect 8229 -8985 8235 -8977
rect 8229 -9028 8263 -8985
rect -1333 -9065 8263 -9028
rect -1333 -9066 -1170 -9065
rect 10244 -9072 10308 -7080
rect 10454 -7520 10488 -6736
rect 11167 -6798 11201 -6736
rect 10756 -6836 11498 -6798
rect 10756 -6960 10790 -6836
rect 10992 -6960 11026 -6836
rect 11228 -6960 11262 -6836
rect 11464 -6960 11498 -6836
rect 11724 -6824 11802 -6818
rect 11724 -6878 11736 -6824
rect 11790 -6878 11802 -6824
rect 11724 -6884 11802 -6878
rect 10750 -6972 10796 -6960
rect 10750 -7348 10756 -6972
rect 10790 -7348 10796 -6972
rect 10750 -7360 10796 -7348
rect 10868 -6972 10914 -6960
rect 10868 -7348 10874 -6972
rect 10908 -7348 10914 -6972
rect 10868 -7360 10914 -7348
rect 10986 -6972 11032 -6960
rect 10986 -7348 10992 -6972
rect 11026 -7348 11032 -6972
rect 10986 -7360 11032 -7348
rect 11104 -6972 11150 -6960
rect 11104 -7348 11110 -6972
rect 11144 -7348 11150 -6972
rect 11104 -7360 11150 -7348
rect 11222 -6972 11268 -6960
rect 11222 -7348 11228 -6972
rect 11262 -7348 11268 -6972
rect 11222 -7360 11268 -7348
rect 11340 -6972 11386 -6960
rect 11340 -7348 11346 -6972
rect 11380 -7348 11386 -6972
rect 11340 -7360 11386 -7348
rect 11458 -6972 11504 -6960
rect 11458 -7348 11464 -6972
rect 11498 -7348 11504 -6972
rect 11458 -7360 11504 -7348
rect 11870 -7519 11904 -6736
rect 12398 -6738 12557 -6703
rect 13000 -6738 13270 -6703
rect 13837 -6703 13871 -6669
rect 14073 -6703 14107 -6669
rect 13837 -6738 14107 -6703
rect 14466 -6701 14500 -6667
rect 15068 -6701 15102 -6667
rect 15304 -6701 15338 -6667
rect 14466 -6736 14625 -6701
rect 15068 -6736 15338 -6701
rect 15905 -6701 15939 -6667
rect 16141 -6701 16175 -6667
rect 15905 -6736 16175 -6701
rect 16831 -6729 16837 -6553
rect 16871 -6729 16877 -6553
rect 12343 -6886 12417 -6820
rect 12483 -6886 12493 -6820
rect 12343 -7016 12483 -7010
rect 12343 -7076 12405 -7016
rect 12471 -7076 12483 -7016
rect 12343 -7082 12483 -7076
rect 11956 -7376 12082 -7370
rect 11956 -7478 11968 -7376
rect 12070 -7478 12082 -7376
rect 11956 -7484 12082 -7478
rect 11597 -7520 11904 -7519
rect 10454 -7525 10770 -7520
rect 11484 -7525 11904 -7520
rect 10454 -7536 10837 -7525
rect 10454 -7563 10786 -7536
rect 10454 -7692 10488 -7563
rect 10770 -7570 10786 -7563
rect 10820 -7570 10837 -7536
rect 10770 -7576 10837 -7570
rect 11417 -7536 11904 -7525
rect 11417 -7570 11434 -7536
rect 11468 -7563 11904 -7536
rect 11468 -7570 11484 -7563
rect 11597 -7564 11904 -7563
rect 11417 -7576 11484 -7570
rect 10595 -7603 10651 -7591
rect 10595 -7637 10601 -7603
rect 10635 -7604 10651 -7603
rect 11708 -7604 11764 -7592
rect 10635 -7620 11102 -7604
rect 10635 -7637 11052 -7620
rect 10595 -7653 11052 -7637
rect 11036 -7654 11052 -7653
rect 11086 -7654 11102 -7620
rect 11036 -7661 11102 -7654
rect 11154 -7619 11724 -7604
rect 11154 -7653 11170 -7619
rect 11204 -7638 11724 -7619
rect 11758 -7638 11764 -7604
rect 11204 -7653 11764 -7638
rect 11154 -7663 11221 -7653
rect 11708 -7654 11764 -7653
rect 11870 -7692 11904 -7564
rect 10448 -7704 10494 -7692
rect 10448 -7880 10454 -7704
rect 10488 -7880 10494 -7704
rect 10448 -7892 10494 -7880
rect 10566 -7704 10612 -7692
rect 10566 -7880 10572 -7704
rect 10606 -7880 10612 -7704
rect 10566 -7892 10612 -7880
rect 10868 -7704 10914 -7692
rect 10571 -8186 10605 -7892
rect 10868 -8080 10874 -7704
rect 10908 -8080 10914 -7704
rect 10868 -8092 10914 -8080
rect 10986 -7704 11032 -7692
rect 10986 -8080 10992 -7704
rect 11026 -8080 11032 -7704
rect 10986 -8092 11032 -8080
rect 11104 -7704 11150 -7692
rect 11104 -8080 11110 -7704
rect 11144 -8080 11150 -7704
rect 11104 -8092 11150 -8080
rect 11222 -7704 11268 -7692
rect 11222 -8080 11228 -7704
rect 11262 -8080 11268 -7704
rect 11222 -8092 11268 -8080
rect 11340 -7704 11386 -7692
rect 11340 -8080 11346 -7704
rect 11380 -8080 11386 -7704
rect 11746 -7704 11792 -7692
rect 11746 -7880 11752 -7704
rect 11786 -7880 11792 -7704
rect 11746 -7892 11792 -7880
rect 11864 -7704 11910 -7692
rect 11864 -7880 11870 -7704
rect 11904 -7880 11910 -7704
rect 11864 -7892 11910 -7880
rect 11340 -8092 11386 -8080
rect 11228 -8186 11262 -8092
rect 11752 -8186 11785 -7892
rect 10571 -8218 11785 -8186
rect 11064 -8240 11196 -8218
rect 11064 -8298 11098 -8240
rect 11160 -8298 11196 -8240
rect 11064 -8303 11196 -8298
rect 10244 -9112 10250 -9072
rect -1505 -9125 10250 -9112
rect 10301 -9112 10308 -9072
rect 10301 -9125 10309 -9112
rect -1505 -9180 10309 -9125
rect -1505 -9181 -1441 -9180
rect 12343 -9211 12407 -7082
rect 12523 -7522 12557 -6738
rect 13236 -6800 13270 -6738
rect 12825 -6838 13567 -6800
rect 12825 -6962 12859 -6838
rect 13061 -6962 13095 -6838
rect 13297 -6962 13331 -6838
rect 13533 -6962 13567 -6838
rect 13793 -6826 13871 -6820
rect 13793 -6880 13805 -6826
rect 13859 -6880 13871 -6826
rect 13793 -6886 13871 -6880
rect 12819 -6974 12865 -6962
rect 12819 -7350 12825 -6974
rect 12859 -7350 12865 -6974
rect 12819 -7362 12865 -7350
rect 12937 -6974 12983 -6962
rect 12937 -7350 12943 -6974
rect 12977 -7350 12983 -6974
rect 12937 -7362 12983 -7350
rect 13055 -6974 13101 -6962
rect 13055 -7350 13061 -6974
rect 13095 -7350 13101 -6974
rect 13055 -7362 13101 -7350
rect 13173 -6974 13219 -6962
rect 13173 -7350 13179 -6974
rect 13213 -7350 13219 -6974
rect 13173 -7362 13219 -7350
rect 13291 -6974 13337 -6962
rect 13291 -7350 13297 -6974
rect 13331 -7350 13337 -6974
rect 13291 -7362 13337 -7350
rect 13409 -6974 13455 -6962
rect 13409 -7350 13415 -6974
rect 13449 -7350 13455 -6974
rect 13409 -7362 13455 -7350
rect 13527 -6974 13573 -6962
rect 13527 -7350 13533 -6974
rect 13567 -7350 13573 -6974
rect 13527 -7362 13573 -7350
rect 13939 -7521 13973 -6738
rect 14411 -6884 14485 -6818
rect 14551 -6884 14561 -6818
rect 14414 -7008 14478 -7007
rect 14414 -7014 14551 -7008
rect 14414 -7074 14473 -7014
rect 14539 -7074 14551 -7014
rect 14414 -7080 14551 -7074
rect 14025 -7378 14151 -7372
rect 14025 -7480 14037 -7378
rect 14139 -7480 14151 -7378
rect 14025 -7486 14151 -7480
rect 13666 -7522 13973 -7521
rect 12523 -7527 12839 -7522
rect 13553 -7527 13973 -7522
rect 12523 -7538 12906 -7527
rect 12523 -7565 12855 -7538
rect 12523 -7694 12557 -7565
rect 12839 -7572 12855 -7565
rect 12889 -7572 12906 -7538
rect 12839 -7578 12906 -7572
rect 13486 -7538 13973 -7527
rect 13486 -7572 13503 -7538
rect 13537 -7565 13973 -7538
rect 13537 -7572 13553 -7565
rect 13666 -7566 13973 -7565
rect 13486 -7578 13553 -7572
rect 12664 -7605 12720 -7593
rect 12664 -7639 12670 -7605
rect 12704 -7606 12720 -7605
rect 13777 -7606 13833 -7594
rect 12704 -7622 13171 -7606
rect 12704 -7639 13121 -7622
rect 12664 -7655 13121 -7639
rect 13105 -7656 13121 -7655
rect 13155 -7656 13171 -7622
rect 13105 -7663 13171 -7656
rect 13223 -7621 13793 -7606
rect 13223 -7655 13239 -7621
rect 13273 -7640 13793 -7621
rect 13827 -7640 13833 -7606
rect 13273 -7655 13833 -7640
rect 13223 -7665 13290 -7655
rect 13777 -7656 13833 -7655
rect 13939 -7694 13973 -7566
rect 12517 -7706 12563 -7694
rect 12517 -7882 12523 -7706
rect 12557 -7882 12563 -7706
rect 12517 -7894 12563 -7882
rect 12635 -7706 12681 -7694
rect 12635 -7882 12641 -7706
rect 12675 -7882 12681 -7706
rect 12635 -7894 12681 -7882
rect 12937 -7706 12983 -7694
rect 12640 -8188 12674 -7894
rect 12937 -8082 12943 -7706
rect 12977 -8082 12983 -7706
rect 12937 -8094 12983 -8082
rect 13055 -7706 13101 -7694
rect 13055 -8082 13061 -7706
rect 13095 -8082 13101 -7706
rect 13055 -8094 13101 -8082
rect 13173 -7706 13219 -7694
rect 13173 -8082 13179 -7706
rect 13213 -8082 13219 -7706
rect 13173 -8094 13219 -8082
rect 13291 -7706 13337 -7694
rect 13291 -8082 13297 -7706
rect 13331 -8082 13337 -7706
rect 13291 -8094 13337 -8082
rect 13409 -7706 13455 -7694
rect 13409 -8082 13415 -7706
rect 13449 -8082 13455 -7706
rect 13815 -7706 13861 -7694
rect 13815 -7882 13821 -7706
rect 13855 -7882 13861 -7706
rect 13815 -7894 13861 -7882
rect 13933 -7706 13979 -7694
rect 13933 -7882 13939 -7706
rect 13973 -7882 13979 -7706
rect 13933 -7894 13979 -7882
rect 13409 -8094 13455 -8082
rect 13297 -8188 13331 -8094
rect 13821 -8188 13854 -7894
rect 12640 -8220 13854 -8188
rect 13133 -8242 13265 -8220
rect 13133 -8300 13167 -8242
rect 13229 -8300 13265 -8242
rect 13133 -8305 13265 -8300
rect -1734 -9216 12408 -9211
rect -1734 -9267 12353 -9216
rect 12397 -9267 12408 -9216
rect -1734 -9278 12408 -9267
rect -1734 -9279 -1654 -9278
rect 12343 -9279 12407 -9278
rect 14414 -9299 14478 -7080
rect 14591 -7520 14625 -6736
rect 15304 -6798 15338 -6736
rect 14893 -6836 15635 -6798
rect 14893 -6960 14927 -6836
rect 15129 -6960 15163 -6836
rect 15365 -6960 15399 -6836
rect 15601 -6960 15635 -6836
rect 15861 -6824 15939 -6818
rect 15861 -6878 15873 -6824
rect 15927 -6878 15939 -6824
rect 15861 -6884 15939 -6878
rect 14887 -6972 14933 -6960
rect 14887 -7348 14893 -6972
rect 14927 -7348 14933 -6972
rect 14887 -7360 14933 -7348
rect 15005 -6972 15051 -6960
rect 15005 -7348 15011 -6972
rect 15045 -7348 15051 -6972
rect 15005 -7360 15051 -7348
rect 15123 -6972 15169 -6960
rect 15123 -7348 15129 -6972
rect 15163 -7348 15169 -6972
rect 15123 -7360 15169 -7348
rect 15241 -6972 15287 -6960
rect 15241 -7348 15247 -6972
rect 15281 -7348 15287 -6972
rect 15241 -7360 15287 -7348
rect 15359 -6972 15405 -6960
rect 15359 -7348 15365 -6972
rect 15399 -7348 15405 -6972
rect 15359 -7360 15405 -7348
rect 15477 -6972 15523 -6960
rect 15477 -7348 15483 -6972
rect 15517 -7348 15523 -6972
rect 15477 -7360 15523 -7348
rect 15595 -6972 15641 -6960
rect 15595 -7348 15601 -6972
rect 15635 -7348 15641 -6972
rect 15595 -7360 15641 -7348
rect 16007 -7519 16041 -6736
rect 16831 -6843 16877 -6729
rect 16949 -6553 17115 -6537
rect 17805 -6539 17853 -6494
rect 18543 -6539 18591 -6490
rect 19079 -6491 19159 -6485
rect 19281 -6493 19445 -6429
rect 19819 -6451 19899 -6445
rect 19819 -6485 19853 -6451
rect 19887 -6485 19899 -6451
rect 19819 -6491 19899 -6485
rect 20021 -6493 20189 -6429
rect 20555 -6451 20637 -6445
rect 20555 -6485 20591 -6451
rect 20625 -6485 20637 -6451
rect 20555 -6491 20637 -6485
rect 20759 -6493 20922 -6429
rect 21501 -6432 21549 -6347
rect 21601 -6432 21665 -5436
rect 22074 -5760 22138 -4380
rect 22291 -4485 22326 -3975
rect 22381 -4021 22473 -4008
rect 22381 -4084 22393 -4021
rect 22464 -4084 22473 -4021
rect 22381 -4093 22473 -4084
rect 23466 -4021 23558 -4011
rect 23466 -4083 23478 -4021
rect 23548 -4083 23558 -4021
rect 23466 -4096 23558 -4083
rect 24854 -4076 24889 -3722
rect 23713 -4138 23778 -4135
rect 23713 -4141 23782 -4138
rect 23713 -4201 23719 -4141
rect 23778 -4201 23788 -4141
rect 23713 -4205 23782 -4201
rect 23713 -4207 23778 -4205
rect 24854 -4222 24890 -4076
rect 23348 -4304 23440 -4296
rect 23348 -4369 23360 -4304
rect 23428 -4369 23440 -4304
rect 23348 -4381 23440 -4369
rect 24854 -4484 24889 -4222
rect 22291 -4532 23663 -4485
rect 23985 -4531 24889 -4484
rect 23125 -4655 23159 -4532
rect 23597 -4545 23663 -4532
rect 23597 -4579 23613 -4545
rect 23647 -4579 23663 -4545
rect 23597 -4595 23663 -4579
rect 23986 -4655 24020 -4531
rect 23120 -4667 23166 -4655
rect 23120 -4843 23126 -4667
rect 23160 -4843 23166 -4667
rect 23120 -4855 23166 -4843
rect 23238 -4667 23358 -4655
rect 23238 -4843 23244 -4667
rect 23278 -4843 23318 -4667
rect 23238 -4855 23318 -4843
rect 23244 -5222 23278 -4855
rect 23312 -5043 23318 -4855
rect 23352 -5043 23358 -4667
rect 23312 -5055 23358 -5043
rect 23430 -4667 23476 -4655
rect 23430 -5043 23436 -4667
rect 23470 -5043 23476 -4667
rect 23430 -5055 23476 -5043
rect 23548 -4667 23594 -4655
rect 23548 -5043 23554 -4667
rect 23588 -5043 23594 -4667
rect 23548 -5055 23594 -5043
rect 23666 -4667 23712 -4655
rect 23666 -5043 23672 -4667
rect 23706 -5043 23712 -4667
rect 23666 -5055 23712 -5043
rect 23784 -4667 23908 -4655
rect 23784 -5043 23790 -4667
rect 23824 -4843 23868 -4667
rect 23902 -4843 23908 -4667
rect 23824 -4855 23908 -4843
rect 23980 -4667 24026 -4655
rect 23980 -4843 23986 -4667
rect 24020 -4843 24026 -4667
rect 23980 -4855 24026 -4843
rect 23824 -5043 23830 -4855
rect 23784 -5055 23830 -5043
rect 23554 -5128 23588 -5055
rect 23539 -5144 23605 -5128
rect 23539 -5178 23555 -5144
rect 23589 -5178 23605 -5144
rect 23539 -5194 23605 -5178
rect 23868 -5222 23902 -4855
rect 23244 -5274 23902 -5222
rect 23542 -5296 23634 -5274
rect 23542 -5348 23554 -5296
rect 23620 -5348 23634 -5296
rect 23542 -5352 23634 -5348
rect 22074 -5824 22405 -5760
rect 22039 -5977 22049 -5963
rect 22009 -5983 22049 -5977
rect 22125 -5977 22135 -5963
rect 22125 -5983 22167 -5977
rect 22009 -6019 22035 -5983
rect 22131 -6019 22167 -5983
rect 22009 -6037 22049 -6019
rect 22125 -6037 22167 -6019
rect 22009 -6077 22167 -6037
rect 21885 -6123 22167 -6077
rect 21885 -6169 21931 -6123
rect 21885 -6345 21891 -6169
rect 21925 -6345 21931 -6169
rect 21885 -6357 21931 -6345
rect 22003 -6169 22049 -6157
rect 22003 -6345 22009 -6169
rect 22043 -6345 22049 -6169
rect 22003 -6357 22049 -6345
rect 22121 -6169 22167 -6123
rect 22121 -6345 22127 -6169
rect 22161 -6345 22167 -6169
rect 22121 -6357 22167 -6345
rect 22239 -6169 22285 -6157
rect 22239 -6345 22245 -6169
rect 22279 -6345 22285 -6169
rect 22239 -6347 22285 -6345
rect 22239 -6429 22287 -6347
rect 22341 -6429 22405 -5824
rect 21140 -6445 21188 -6433
rect 21140 -6491 21146 -6445
rect 21182 -6451 21375 -6445
rect 21182 -6485 21329 -6451
rect 21363 -6485 21375 -6451
rect 21182 -6491 21375 -6485
rect 19285 -6539 19333 -6493
rect 20025 -6539 20073 -6493
rect 20763 -6539 20811 -6493
rect 21140 -6503 21188 -6491
rect 21494 -6496 21665 -6432
rect 21877 -6445 21927 -6433
rect 21877 -6491 21883 -6445
rect 21921 -6451 22113 -6445
rect 21921 -6485 22067 -6451
rect 22101 -6485 22113 -6451
rect 21921 -6491 22113 -6485
rect 21501 -6539 21549 -6496
rect 21877 -6503 21927 -6491
rect 22235 -6493 22405 -6429
rect 22239 -6539 22287 -6493
rect 16949 -6729 16955 -6553
rect 16989 -6567 17115 -6553
rect 17569 -6551 17615 -6539
rect 16989 -6729 16995 -6567
rect 16949 -6741 16995 -6729
rect 17569 -6727 17575 -6551
rect 17609 -6727 17615 -6551
rect 16791 -6909 16801 -6843
rect 16903 -6909 16913 -6843
rect 17569 -6845 17615 -6727
rect 17687 -6551 17853 -6539
rect 17687 -6727 17693 -6551
rect 17727 -6569 17853 -6551
rect 18307 -6555 18353 -6543
rect 17727 -6727 17733 -6569
rect 17687 -6739 17733 -6727
rect 18307 -6731 18313 -6555
rect 18347 -6731 18353 -6555
rect 18307 -6845 18353 -6731
rect 18425 -6555 18591 -6539
rect 18425 -6731 18431 -6555
rect 18465 -6569 18591 -6555
rect 19049 -6555 19095 -6543
rect 18465 -6731 18471 -6569
rect 18425 -6743 18471 -6731
rect 19049 -6731 19055 -6555
rect 19089 -6731 19095 -6555
rect 19049 -6845 19095 -6731
rect 19167 -6555 19333 -6539
rect 19167 -6731 19173 -6555
rect 19207 -6569 19333 -6555
rect 19789 -6555 19835 -6543
rect 19207 -6731 19213 -6569
rect 19167 -6743 19213 -6731
rect 19789 -6731 19795 -6555
rect 19829 -6731 19835 -6555
rect 19789 -6845 19835 -6731
rect 19907 -6555 20073 -6539
rect 19907 -6731 19913 -6555
rect 19947 -6569 20073 -6555
rect 20527 -6555 20573 -6543
rect 19947 -6731 19953 -6569
rect 19907 -6743 19953 -6731
rect 20527 -6731 20533 -6555
rect 20567 -6731 20573 -6555
rect 20527 -6845 20573 -6731
rect 20645 -6555 20811 -6539
rect 20645 -6731 20651 -6555
rect 20685 -6569 20811 -6555
rect 21265 -6551 21311 -6539
rect 20685 -6731 20691 -6569
rect 20645 -6743 20691 -6731
rect 21265 -6727 21271 -6551
rect 21305 -6727 21311 -6551
rect 21265 -6845 21311 -6727
rect 21383 -6551 21549 -6539
rect 21383 -6727 21389 -6551
rect 21423 -6569 21549 -6551
rect 22003 -6551 22049 -6539
rect 21423 -6727 21429 -6569
rect 21383 -6739 21429 -6727
rect 22003 -6727 22009 -6551
rect 22043 -6727 22049 -6551
rect 22003 -6845 22049 -6727
rect 22121 -6551 22287 -6539
rect 22121 -6727 22127 -6551
rect 22161 -6569 22287 -6551
rect 22161 -6727 22167 -6569
rect 22121 -6739 22167 -6727
rect 17529 -6911 17539 -6845
rect 17641 -6911 17651 -6845
rect 18267 -6911 18277 -6845
rect 18379 -6911 18389 -6845
rect 19009 -6911 19019 -6845
rect 19121 -6911 19131 -6845
rect 19749 -6911 19759 -6845
rect 19861 -6911 19871 -6845
rect 20487 -6911 20497 -6845
rect 20599 -6911 20609 -6845
rect 21225 -6911 21235 -6845
rect 21337 -6911 21347 -6845
rect 21963 -6911 21973 -6845
rect 22075 -6911 22085 -6845
rect 16093 -7376 16219 -7370
rect 16093 -7478 16105 -7376
rect 16207 -7478 16219 -7376
rect 16093 -7484 16219 -7478
rect 15734 -7520 16041 -7519
rect 14591 -7525 14907 -7520
rect 15621 -7525 16041 -7520
rect 14591 -7536 14974 -7525
rect 14591 -7563 14923 -7536
rect 14591 -7692 14625 -7563
rect 14907 -7570 14923 -7563
rect 14957 -7570 14974 -7536
rect 14907 -7576 14974 -7570
rect 15554 -7536 16041 -7525
rect 15554 -7570 15571 -7536
rect 15605 -7563 16041 -7536
rect 15605 -7570 15621 -7563
rect 15734 -7564 16041 -7563
rect 15554 -7576 15621 -7570
rect 14732 -7603 14788 -7591
rect 14732 -7637 14738 -7603
rect 14772 -7604 14788 -7603
rect 15845 -7604 15901 -7592
rect 14772 -7620 15239 -7604
rect 14772 -7637 15189 -7620
rect 14732 -7653 15189 -7637
rect 15173 -7654 15189 -7653
rect 15223 -7654 15239 -7620
rect 15173 -7661 15239 -7654
rect 15291 -7619 15861 -7604
rect 15291 -7653 15307 -7619
rect 15341 -7638 15861 -7619
rect 15895 -7638 15901 -7604
rect 15341 -7653 15901 -7638
rect 15291 -7663 15358 -7653
rect 15845 -7654 15901 -7653
rect 16007 -7692 16041 -7564
rect 14585 -7704 14631 -7692
rect 14585 -7880 14591 -7704
rect 14625 -7880 14631 -7704
rect 14585 -7892 14631 -7880
rect 14703 -7704 14749 -7692
rect 14703 -7880 14709 -7704
rect 14743 -7880 14749 -7704
rect 14703 -7892 14749 -7880
rect 15005 -7704 15051 -7692
rect 14708 -8186 14742 -7892
rect 15005 -8080 15011 -7704
rect 15045 -8080 15051 -7704
rect 15005 -8092 15051 -8080
rect 15123 -7704 15169 -7692
rect 15123 -8080 15129 -7704
rect 15163 -8080 15169 -7704
rect 15123 -8092 15169 -8080
rect 15241 -7704 15287 -7692
rect 15241 -8080 15247 -7704
rect 15281 -8080 15287 -7704
rect 15241 -8092 15287 -8080
rect 15359 -7704 15405 -7692
rect 15359 -8080 15365 -7704
rect 15399 -8080 15405 -7704
rect 15359 -8092 15405 -8080
rect 15477 -7704 15523 -7692
rect 15477 -8080 15483 -7704
rect 15517 -8080 15523 -7704
rect 15883 -7704 15929 -7692
rect 15883 -7880 15889 -7704
rect 15923 -7880 15929 -7704
rect 15883 -7892 15929 -7880
rect 16001 -7704 16047 -7692
rect 16001 -7880 16007 -7704
rect 16041 -7880 16047 -7704
rect 16001 -7892 16047 -7880
rect 15477 -8092 15523 -8080
rect 15365 -8186 15399 -8092
rect 15889 -8186 15922 -7892
rect 14708 -8218 15922 -8186
rect 15201 -8240 15333 -8218
rect 15201 -8298 15235 -8240
rect 15297 -8298 15333 -8240
rect 15201 -8303 15333 -8298
rect 14414 -9310 14480 -9299
rect -1987 -9311 14480 -9310
rect -1987 -9365 14421 -9311
rect 14474 -9365 14480 -9311
rect -1987 -9388 14480 -9365
<< via1 >>
rect -2478 5863 -2418 5922
rect 10304 5847 10358 5901
rect 10398 5754 10452 5808
rect -2481 5660 -2421 5722
rect -2488 5470 -2428 5532
rect -2488 5281 -2428 5350
rect -2501 5100 -2440 5163
rect -2514 4900 -2443 4972
rect -2497 3111 -2443 3166
rect -2526 2737 -2470 2791
rect -2507 -1364 -2445 -1289
rect -2506 -1691 -2444 -1616
rect 8766 5662 8820 5716
rect 8941 5567 8995 5621
rect -2237 -5618 -2182 -5557
rect -1981 -5615 -1913 -5557
rect -2237 -5910 -2182 -5849
rect -2237 -6215 -2182 -6154
rect -2237 -6376 -2182 -6315
rect -2237 -6527 -2181 -6466
rect -2237 -6687 -2182 -6626
rect -2237 -6874 -2182 -6813
rect -2237 -7080 -2182 -7019
rect 7305 5477 7359 5531
rect -1722 -5908 -1666 -5851
rect 7443 5383 7497 5437
rect 5803 5289 5857 5343
rect 5982 5195 6036 5249
rect -1504 -6212 -1443 -6159
rect 4347 5105 4401 5159
rect 4475 5010 4529 5064
rect -1329 -6374 -1259 -6316
rect 2894 4919 2948 4973
rect -1127 -6524 -1059 -6466
rect 3025 4824 3079 4878
rect 1449 4733 1503 4787
rect 1559 4640 1613 4694
rect -931 -6683 -873 -6629
rect -293 3408 -222 3467
rect 542 4061 602 4123
rect 1990 4061 2050 4123
rect 3488 4063 3548 4125
rect 4936 4063 4996 4125
rect 6456 4061 6516 4123
rect 7904 4061 7964 4123
rect 9402 4063 9462 4125
rect 10850 4063 10910 4125
rect 12536 4259 12588 4311
rect 13704 4259 13756 4311
rect -7 3307 62 3371
rect 764 2911 826 2919
rect 764 2865 770 2911
rect 770 2865 822 2911
rect 822 2865 826 2911
rect 764 2859 826 2865
rect 1766 3244 1820 3298
rect 1651 3112 1705 3167
rect 2212 2911 2274 2919
rect 2212 2865 2218 2911
rect 2218 2865 2270 2911
rect 2270 2865 2274 2911
rect 2212 2859 2274 2865
rect 3260 3243 3314 3297
rect 3149 3111 3203 3165
rect 3710 2913 3772 2921
rect 3710 2867 3716 2913
rect 3716 2867 3768 2913
rect 3768 2867 3772 2913
rect 3710 2861 3772 2867
rect -503 1356 -420 1444
rect 1508 2378 1588 2384
rect 1508 2324 1512 2378
rect 1512 2324 1584 2378
rect 1584 2324 1588 2378
rect 117 1322 174 1326
rect 117 1262 121 1322
rect 121 1262 170 1322
rect 170 1262 174 1322
rect 117 1258 174 1262
rect 117 1154 174 1158
rect 117 1094 121 1154
rect 121 1094 170 1154
rect 170 1094 174 1154
rect 117 1090 174 1094
rect 361 1437 432 1441
rect 361 1382 365 1437
rect 365 1382 425 1437
rect 425 1382 432 1437
rect 361 1378 432 1382
rect 1446 1438 1516 1441
rect 1446 1383 1450 1438
rect 1450 1383 1510 1438
rect 1510 1383 1516 1438
rect 1446 1379 1516 1383
rect 1687 1307 1746 1321
rect 1687 1273 1700 1307
rect 1700 1273 1734 1307
rect 1734 1273 1746 1307
rect 1687 1261 1746 1273
rect 4710 3246 4764 3300
rect 4597 3116 4651 3170
rect 14872 4259 14924 4311
rect 16040 4259 16092 4311
rect 5158 2913 5220 2921
rect 5158 2867 5164 2913
rect 5164 2867 5216 2913
rect 5216 2867 5220 2913
rect 5158 2861 5220 2867
rect 6229 3241 6283 3295
rect 6113 3116 6167 3170
rect 6678 2911 6740 2919
rect 6678 2865 6684 2911
rect 6684 2865 6736 2911
rect 6736 2865 6740 2911
rect 6678 2859 6740 2865
rect 7677 3248 7731 3302
rect 7565 3110 7619 3164
rect 8126 2911 8188 2919
rect 8126 2865 8132 2911
rect 8132 2865 8184 2911
rect 8184 2865 8188 2911
rect 8126 2859 8188 2865
rect 9174 3246 9228 3300
rect 9062 3116 9116 3170
rect 9624 2913 9686 2921
rect 9624 2867 9630 2913
rect 9630 2867 9682 2913
rect 9682 2867 9686 2913
rect 9624 2861 9686 2867
rect 10606 3228 10692 3316
rect 10492 3099 10578 3187
rect 11072 2913 11134 2921
rect 11072 2867 11078 2913
rect 11078 2867 11130 2913
rect 11130 2867 11134 2913
rect 11072 2861 11134 2867
rect 17214 4261 17266 4313
rect 18382 4261 18434 4313
rect 19550 4261 19602 4313
rect 20718 4261 20770 4313
rect 12065 2935 12117 2987
rect 13233 2935 13285 2987
rect 14401 2935 14453 2987
rect 15569 2935 15621 2987
rect 16743 2937 16795 2989
rect 17911 2937 17963 2989
rect 19079 2937 19131 2989
rect 20247 2937 20299 2989
rect 4652 2378 4732 2384
rect 4652 2324 4656 2378
rect 4656 2324 4728 2378
rect 4728 2324 4732 2378
rect 3261 1322 3318 1326
rect 3261 1262 3265 1322
rect 3265 1262 3314 1322
rect 3314 1262 3318 1322
rect 3261 1258 3318 1262
rect 1328 1153 1396 1158
rect 1328 1098 1332 1153
rect 1332 1098 1392 1153
rect 1392 1098 1396 1153
rect 1328 1093 1396 1098
rect 1522 120 1526 166
rect 1526 120 1584 166
rect 1584 120 1588 166
rect 1522 114 1588 120
rect 3261 1154 3318 1158
rect 3261 1094 3265 1154
rect 3265 1094 3314 1154
rect 3314 1094 3318 1154
rect 3261 1090 3318 1094
rect 3505 1437 3576 1441
rect 3505 1382 3509 1437
rect 3509 1382 3569 1437
rect 3569 1382 3576 1437
rect 3505 1378 3576 1382
rect 4590 1438 4660 1441
rect 4590 1383 4594 1438
rect 4594 1383 4654 1438
rect 4654 1383 4660 1438
rect 4590 1379 4660 1383
rect 4831 1307 4890 1321
rect 4831 1273 4844 1307
rect 4844 1273 4878 1307
rect 4878 1273 4890 1307
rect 4831 1261 4890 1273
rect 7784 2382 7864 2388
rect 7784 2328 7788 2382
rect 7788 2328 7860 2382
rect 7860 2328 7864 2382
rect 6393 1326 6450 1330
rect 6393 1266 6397 1326
rect 6397 1266 6446 1326
rect 6446 1266 6450 1326
rect 6393 1262 6450 1266
rect 4472 1153 4540 1158
rect 4472 1098 4476 1153
rect 4476 1098 4536 1153
rect 4536 1098 4540 1153
rect 4472 1093 4540 1098
rect 4666 120 4670 166
rect 4670 120 4728 166
rect 4728 120 4732 166
rect 4666 114 4732 120
rect 6393 1158 6450 1162
rect 6393 1098 6397 1158
rect 6397 1098 6446 1158
rect 6446 1098 6450 1158
rect 6393 1094 6450 1098
rect 6637 1441 6708 1445
rect 6637 1386 6641 1441
rect 6641 1386 6701 1441
rect 6701 1386 6708 1441
rect 6637 1382 6708 1386
rect 7722 1442 7792 1445
rect 7722 1387 7726 1442
rect 7726 1387 7786 1442
rect 7786 1387 7792 1442
rect 7722 1383 7792 1387
rect 7963 1311 8022 1325
rect 7963 1277 7976 1311
rect 7976 1277 8010 1311
rect 8010 1277 8022 1311
rect 7963 1265 8022 1277
rect 10928 2382 11008 2388
rect 10928 2328 10932 2382
rect 10932 2328 11004 2382
rect 11004 2328 11008 2382
rect 9537 1326 9594 1330
rect 9537 1266 9541 1326
rect 9541 1266 9590 1326
rect 9590 1266 9594 1326
rect 9537 1262 9594 1266
rect 7604 1157 7672 1162
rect 7604 1102 7608 1157
rect 7608 1102 7668 1157
rect 7668 1102 7672 1157
rect 7604 1097 7672 1102
rect 7798 124 7802 170
rect 7802 124 7860 170
rect 7860 124 7864 170
rect 7798 118 7864 124
rect 9781 1441 9852 1445
rect 9781 1386 9785 1441
rect 9785 1386 9845 1441
rect 9845 1386 9852 1441
rect 9781 1382 9852 1386
rect 10866 1442 10936 1445
rect 10866 1387 10870 1442
rect 10870 1387 10930 1442
rect 10930 1387 10936 1442
rect 10866 1383 10936 1387
rect 11107 1311 11166 1325
rect 11107 1277 11120 1311
rect 11120 1277 11154 1311
rect 11154 1277 11166 1311
rect 11107 1265 11166 1277
rect 14130 2378 14210 2384
rect 14130 2324 14134 2378
rect 14134 2324 14206 2378
rect 14206 2324 14210 2378
rect 12739 1322 12796 1326
rect 12739 1262 12743 1322
rect 12743 1262 12792 1322
rect 12792 1262 12796 1322
rect 12739 1258 12796 1262
rect 10942 124 10946 170
rect 10946 124 11004 170
rect 11004 124 11008 170
rect 10942 118 11008 124
rect 12983 1437 13054 1441
rect 12983 1382 12987 1437
rect 12987 1382 13047 1437
rect 13047 1382 13054 1437
rect 12983 1378 13054 1382
rect 14068 1438 14138 1441
rect 14068 1383 14072 1438
rect 14072 1383 14132 1438
rect 14132 1383 14138 1438
rect 14068 1379 14138 1383
rect 14309 1307 14368 1321
rect 14309 1273 14322 1307
rect 14322 1273 14356 1307
rect 14356 1273 14368 1307
rect 14309 1261 14368 1273
rect 17274 2378 17354 2384
rect 17274 2324 17278 2378
rect 17278 2324 17350 2378
rect 17350 2324 17354 2378
rect 15883 1322 15940 1326
rect 15883 1262 15887 1322
rect 15887 1262 15936 1322
rect 15936 1262 15940 1322
rect 15883 1258 15940 1262
rect 14144 120 14148 166
rect 14148 120 14206 166
rect 14206 120 14210 166
rect 14144 114 14210 120
rect 15883 1154 15940 1158
rect 15883 1094 15887 1154
rect 15887 1094 15936 1154
rect 15936 1094 15940 1154
rect 15883 1090 15940 1094
rect 16127 1437 16198 1441
rect 16127 1382 16131 1437
rect 16131 1382 16191 1437
rect 16191 1382 16198 1437
rect 16127 1378 16198 1382
rect 17212 1438 17282 1441
rect 17212 1383 17216 1438
rect 17216 1383 17276 1438
rect 17276 1383 17282 1438
rect 17212 1379 17282 1383
rect 17453 1307 17512 1321
rect 17453 1273 17466 1307
rect 17466 1273 17500 1307
rect 17500 1273 17512 1307
rect 17453 1261 17512 1273
rect 20406 2382 20486 2388
rect 20406 2328 20410 2382
rect 20410 2328 20482 2382
rect 20482 2328 20486 2382
rect 19015 1326 19072 1330
rect 19015 1266 19019 1326
rect 19019 1266 19068 1326
rect 19068 1266 19072 1326
rect 19015 1262 19072 1266
rect 17094 1153 17162 1158
rect 17094 1098 17098 1153
rect 17098 1098 17158 1153
rect 17158 1098 17162 1153
rect 17094 1093 17162 1098
rect 17288 120 17292 166
rect 17292 120 17350 166
rect 17350 120 17354 166
rect 17288 114 17354 120
rect 19015 1158 19072 1162
rect 19015 1098 19019 1158
rect 19019 1098 19068 1158
rect 19068 1098 19072 1158
rect 19015 1094 19072 1098
rect 19259 1441 19330 1445
rect 19259 1386 19263 1441
rect 19263 1386 19323 1441
rect 19323 1386 19330 1441
rect 19259 1382 19330 1386
rect 20344 1442 20414 1445
rect 20344 1387 20348 1442
rect 20348 1387 20408 1442
rect 20408 1387 20414 1442
rect 20344 1383 20414 1387
rect 20585 1311 20644 1325
rect 20585 1277 20598 1311
rect 20598 1277 20632 1311
rect 20632 1277 20644 1311
rect 20585 1265 20644 1277
rect 23550 2382 23630 2388
rect 23550 2328 23554 2382
rect 23554 2328 23626 2382
rect 23626 2328 23630 2382
rect 22159 1326 22216 1330
rect 22159 1266 22163 1326
rect 22163 1266 22212 1326
rect 22212 1266 22216 1326
rect 22159 1262 22216 1266
rect 20226 1157 20294 1162
rect 20226 1102 20230 1157
rect 20230 1102 20290 1157
rect 20290 1102 20294 1157
rect 20226 1097 20294 1102
rect 20420 124 20424 170
rect 20424 124 20482 170
rect 20482 124 20486 170
rect 20420 118 20486 124
rect 22159 1158 22216 1162
rect 22159 1098 22163 1158
rect 22163 1098 22212 1158
rect 22212 1098 22216 1158
rect 22159 1094 22216 1098
rect 22403 1441 22474 1445
rect 22403 1386 22407 1441
rect 22407 1386 22467 1441
rect 22467 1386 22474 1441
rect 22403 1382 22474 1386
rect 23488 1442 23558 1445
rect 23488 1387 23492 1442
rect 23492 1387 23552 1442
rect 23552 1387 23558 1442
rect 23488 1383 23558 1387
rect 23729 1311 23788 1325
rect 23729 1277 23742 1311
rect 23742 1277 23776 1311
rect 23776 1277 23788 1311
rect 23729 1265 23788 1277
rect 23370 1157 23438 1162
rect 23370 1102 23374 1157
rect 23374 1102 23434 1157
rect 23434 1102 23438 1157
rect 23370 1097 23438 1102
rect 23564 124 23568 170
rect 23568 124 23626 170
rect 23626 124 23630 170
rect 23564 118 23630 124
rect 1508 -356 1588 -350
rect 1508 -410 1512 -356
rect 1512 -410 1584 -356
rect 1584 -410 1588 -356
rect 117 -1412 174 -1408
rect 117 -1472 121 -1412
rect 121 -1472 170 -1412
rect 170 -1472 174 -1412
rect 117 -1476 174 -1472
rect -496 -1685 -429 -1615
rect 117 -1580 174 -1576
rect 117 -1640 121 -1580
rect 121 -1640 170 -1580
rect 170 -1640 174 -1580
rect 117 -1644 174 -1640
rect 361 -1297 432 -1293
rect 361 -1352 365 -1297
rect 365 -1352 425 -1297
rect 425 -1352 432 -1297
rect 361 -1356 432 -1352
rect 1446 -1296 1516 -1293
rect 1446 -1351 1450 -1296
rect 1450 -1351 1510 -1296
rect 1510 -1351 1516 -1296
rect 1446 -1355 1516 -1351
rect 1687 -1427 1746 -1413
rect 1687 -1461 1700 -1427
rect 1700 -1461 1734 -1427
rect 1734 -1461 1746 -1427
rect 1687 -1473 1746 -1461
rect 4652 -356 4732 -350
rect 4652 -410 4656 -356
rect 4656 -410 4728 -356
rect 4728 -410 4732 -356
rect 3261 -1412 3318 -1408
rect 3261 -1472 3265 -1412
rect 3265 -1472 3314 -1412
rect 3314 -1472 3318 -1412
rect 3261 -1476 3318 -1472
rect 1328 -1581 1396 -1576
rect 1328 -1636 1332 -1581
rect 1332 -1636 1392 -1581
rect 1392 -1636 1396 -1581
rect 1328 -1641 1396 -1636
rect 3261 -1580 3318 -1576
rect 3261 -1640 3265 -1580
rect 3265 -1640 3314 -1580
rect 3314 -1640 3318 -1580
rect 3261 -1644 3318 -1640
rect 1522 -2614 1526 -2568
rect 1526 -2614 1584 -2568
rect 1584 -2614 1588 -2568
rect 1522 -2620 1588 -2614
rect 2936 -2614 3000 -2537
rect 3505 -1297 3576 -1293
rect 3505 -1352 3509 -1297
rect 3509 -1352 3569 -1297
rect 3569 -1352 3576 -1297
rect 3505 -1356 3576 -1352
rect 4590 -1296 4660 -1293
rect 4590 -1351 4594 -1296
rect 4594 -1351 4654 -1296
rect 4654 -1351 4660 -1296
rect 4590 -1355 4660 -1351
rect 4831 -1427 4890 -1413
rect 4831 -1461 4844 -1427
rect 4844 -1461 4878 -1427
rect 4878 -1461 4890 -1427
rect 4831 -1473 4890 -1461
rect 7784 -352 7864 -346
rect 7784 -406 7788 -352
rect 7788 -406 7860 -352
rect 7860 -406 7864 -352
rect 6393 -1408 6450 -1404
rect 6393 -1468 6397 -1408
rect 6397 -1468 6446 -1408
rect 6446 -1468 6450 -1408
rect 6393 -1472 6450 -1468
rect 4472 -1581 4540 -1576
rect 4472 -1636 4476 -1581
rect 4476 -1636 4536 -1581
rect 4536 -1636 4540 -1581
rect 4472 -1641 4540 -1636
rect 4666 -2614 4670 -2568
rect 4670 -2614 4728 -2568
rect 4728 -2614 4732 -2568
rect 4666 -2620 4732 -2614
rect 6046 -2668 6114 -2596
rect 6393 -1576 6450 -1572
rect 6393 -1636 6397 -1576
rect 6397 -1636 6446 -1576
rect 6446 -1636 6450 -1576
rect 6393 -1640 6450 -1636
rect 6637 -1293 6708 -1289
rect 6637 -1348 6641 -1293
rect 6641 -1348 6701 -1293
rect 6701 -1348 6708 -1293
rect 6637 -1352 6708 -1348
rect 7722 -1292 7792 -1289
rect 7722 -1347 7726 -1292
rect 7726 -1347 7786 -1292
rect 7786 -1347 7792 -1292
rect 7722 -1351 7792 -1347
rect 7963 -1423 8022 -1409
rect 7963 -1457 7976 -1423
rect 7976 -1457 8010 -1423
rect 8010 -1457 8022 -1423
rect 7963 -1469 8022 -1457
rect 10928 -352 11008 -346
rect 10928 -406 10932 -352
rect 10932 -406 11004 -352
rect 11004 -406 11008 -352
rect 9537 -1408 9594 -1404
rect 9537 -1468 9541 -1408
rect 9541 -1468 9590 -1408
rect 9590 -1468 9594 -1408
rect 9537 -1472 9594 -1468
rect 7604 -1577 7672 -1572
rect 7604 -1632 7608 -1577
rect 7608 -1632 7668 -1577
rect 7668 -1632 7672 -1577
rect 7604 -1637 7672 -1632
rect 7798 -2610 7802 -2564
rect 7802 -2610 7860 -2564
rect 7860 -2610 7864 -2564
rect 7798 -2616 7864 -2610
rect 9182 -2790 9249 -2722
rect 9537 -1576 9594 -1572
rect 9537 -1636 9541 -1576
rect 9541 -1636 9590 -1576
rect 9590 -1636 9594 -1576
rect 9537 -1640 9594 -1636
rect 9781 -1293 9852 -1289
rect 9781 -1348 9785 -1293
rect 9785 -1348 9845 -1293
rect 9845 -1348 9852 -1293
rect 9781 -1352 9852 -1348
rect 10866 -1292 10936 -1289
rect 10866 -1347 10870 -1292
rect 10870 -1347 10930 -1292
rect 10930 -1347 10936 -1292
rect 10866 -1351 10936 -1347
rect 11107 -1423 11166 -1409
rect 11107 -1457 11120 -1423
rect 11120 -1457 11154 -1423
rect 11154 -1457 11166 -1423
rect 11107 -1469 11166 -1457
rect 14130 -356 14210 -350
rect 14130 -410 14134 -356
rect 14134 -410 14206 -356
rect 14206 -410 14210 -356
rect 12739 -1412 12796 -1408
rect 12739 -1472 12743 -1412
rect 12743 -1472 12792 -1412
rect 12792 -1472 12796 -1412
rect 12739 -1476 12796 -1472
rect 10748 -1577 10816 -1572
rect 10748 -1632 10752 -1577
rect 10752 -1632 10812 -1577
rect 10812 -1632 10816 -1577
rect 10748 -1637 10816 -1632
rect 12329 -2447 12407 -2378
rect 12739 -1580 12796 -1576
rect 12739 -1640 12743 -1580
rect 12743 -1640 12792 -1580
rect 12792 -1640 12796 -1580
rect 12739 -1644 12796 -1640
rect 10942 -2610 10946 -2564
rect 10946 -2610 11004 -2564
rect 11004 -2610 11008 -2564
rect 10942 -2616 11008 -2610
rect 12983 -1297 13054 -1293
rect 12983 -1352 12987 -1297
rect 12987 -1352 13047 -1297
rect 13047 -1352 13054 -1297
rect 12983 -1356 13054 -1352
rect 14068 -1296 14138 -1293
rect 14068 -1351 14072 -1296
rect 14072 -1351 14132 -1296
rect 14132 -1351 14138 -1296
rect 14068 -1355 14138 -1351
rect 14309 -1427 14368 -1413
rect 14309 -1461 14322 -1427
rect 14322 -1461 14356 -1427
rect 14356 -1461 14368 -1427
rect 14309 -1473 14368 -1461
rect 17274 -356 17354 -350
rect 17274 -410 17278 -356
rect 17278 -410 17350 -356
rect 17350 -410 17354 -356
rect 15883 -1296 15940 -1292
rect 15883 -1356 15887 -1296
rect 15887 -1356 15936 -1296
rect 15936 -1356 15940 -1296
rect 15883 -1360 15940 -1356
rect 15883 -1412 15940 -1408
rect 15883 -1472 15887 -1412
rect 15887 -1472 15936 -1412
rect 15936 -1472 15940 -1412
rect 15883 -1476 15940 -1472
rect 13950 -1581 14018 -1576
rect 13950 -1636 13954 -1581
rect 13954 -1636 14014 -1581
rect 14014 -1636 14018 -1581
rect 13950 -1641 14018 -1636
rect 15883 -1580 15940 -1576
rect 15883 -1640 15887 -1580
rect 15887 -1640 15936 -1580
rect 15936 -1640 15940 -1580
rect 15883 -1644 15940 -1640
rect 15529 -2269 15625 -2174
rect 14144 -2614 14148 -2568
rect 14148 -2614 14206 -2568
rect 14206 -2614 14210 -2568
rect 14144 -2620 14210 -2614
rect 16127 -1297 16198 -1293
rect 16127 -1352 16131 -1297
rect 16131 -1352 16191 -1297
rect 16191 -1352 16198 -1297
rect 16127 -1356 16198 -1352
rect 17212 -1296 17282 -1293
rect 17212 -1351 17216 -1296
rect 17216 -1351 17276 -1296
rect 17276 -1351 17282 -1296
rect 17212 -1355 17282 -1351
rect 17453 -1427 17512 -1413
rect 17453 -1461 17466 -1427
rect 17466 -1461 17500 -1427
rect 17500 -1461 17512 -1427
rect 17453 -1473 17512 -1461
rect 20406 -352 20486 -346
rect 20406 -406 20410 -352
rect 20410 -406 20482 -352
rect 20482 -406 20486 -352
rect 19015 -1408 19072 -1404
rect 19015 -1468 19019 -1408
rect 19019 -1468 19068 -1408
rect 19068 -1468 19072 -1408
rect 19015 -1472 19072 -1468
rect 17094 -1581 17162 -1576
rect 17094 -1636 17098 -1581
rect 17098 -1636 17158 -1581
rect 17158 -1636 17162 -1581
rect 17094 -1641 17162 -1636
rect 18688 -2036 18758 -1943
rect 19015 -1576 19072 -1572
rect 19015 -1636 19019 -1576
rect 19019 -1636 19068 -1576
rect 19068 -1636 19072 -1576
rect 19015 -1640 19072 -1636
rect 17288 -2614 17292 -2568
rect 17292 -2614 17350 -2568
rect 17350 -2614 17354 -2568
rect 17288 -2620 17354 -2614
rect 1498 -3088 1578 -3082
rect 1498 -3142 1502 -3088
rect 1502 -3142 1574 -3088
rect 1574 -3142 1578 -3088
rect 107 -4028 164 -4024
rect 107 -4088 111 -4028
rect 111 -4088 160 -4028
rect 160 -4088 164 -4028
rect 107 -4092 164 -4088
rect 107 -4144 164 -4140
rect 107 -4204 111 -4144
rect 111 -4204 160 -4144
rect 160 -4204 164 -4144
rect 107 -4208 164 -4204
rect 107 -4312 164 -4308
rect 107 -4372 111 -4312
rect 111 -4372 160 -4312
rect 160 -4372 164 -4312
rect 107 -4376 164 -4372
rect 351 -4029 422 -4025
rect 351 -4084 355 -4029
rect 355 -4084 415 -4029
rect 415 -4084 422 -4029
rect 351 -4088 422 -4084
rect 1436 -4028 1506 -4025
rect 1436 -4083 1440 -4028
rect 1440 -4083 1500 -4028
rect 1500 -4083 1506 -4028
rect 1436 -4087 1506 -4083
rect 4642 -3088 4722 -3082
rect 4642 -3142 4646 -3088
rect 4646 -3142 4718 -3088
rect 4718 -3142 4722 -3088
rect 1677 -4159 1736 -4145
rect 1677 -4193 1690 -4159
rect 1690 -4193 1724 -4159
rect 1724 -4193 1736 -4159
rect 1677 -4205 1736 -4193
rect 3251 -4028 3308 -4024
rect 3251 -4088 3255 -4028
rect 3255 -4088 3304 -4028
rect 3304 -4088 3308 -4028
rect 3251 -4092 3308 -4088
rect 3251 -4144 3308 -4140
rect 3251 -4204 3255 -4144
rect 3255 -4204 3304 -4144
rect 3304 -4204 3308 -4144
rect 3251 -4208 3308 -4204
rect 1318 -4313 1386 -4308
rect 1318 -4368 1322 -4313
rect 1322 -4368 1382 -4313
rect 1382 -4368 1386 -4313
rect 1318 -4373 1386 -4368
rect 3251 -4312 3308 -4308
rect 3251 -4372 3255 -4312
rect 3255 -4372 3304 -4312
rect 3304 -4372 3308 -4312
rect 3251 -4376 3308 -4372
rect 1512 -5346 1516 -5300
rect 1516 -5346 1574 -5300
rect 1574 -5346 1578 -5300
rect 1512 -5352 1578 -5346
rect 3495 -4029 3566 -4025
rect 3495 -4084 3499 -4029
rect 3499 -4084 3559 -4029
rect 3559 -4084 3566 -4029
rect 3495 -4088 3566 -4084
rect 4580 -4028 4650 -4025
rect 4580 -4083 4584 -4028
rect 4584 -4083 4644 -4028
rect 4644 -4083 4650 -4028
rect 4580 -4087 4650 -4083
rect 7774 -3084 7854 -3078
rect 7774 -3138 7778 -3084
rect 7778 -3138 7850 -3084
rect 7850 -3138 7854 -3084
rect 4821 -4159 4880 -4145
rect 4821 -4193 4834 -4159
rect 4834 -4193 4868 -4159
rect 4868 -4193 4880 -4159
rect 4821 -4205 4880 -4193
rect 6383 -4024 6440 -4020
rect 6383 -4084 6387 -4024
rect 6387 -4084 6436 -4024
rect 6436 -4084 6440 -4024
rect 6383 -4088 6440 -4084
rect 6383 -4140 6440 -4136
rect 6383 -4200 6387 -4140
rect 6387 -4200 6436 -4140
rect 6436 -4200 6440 -4140
rect 6383 -4204 6440 -4200
rect 4462 -4313 4530 -4308
rect 4462 -4368 4466 -4313
rect 4466 -4368 4526 -4313
rect 4526 -4368 4530 -4313
rect 4462 -4373 4530 -4368
rect 6383 -4308 6440 -4304
rect 6383 -4368 6387 -4308
rect 6387 -4368 6436 -4308
rect 6436 -4368 6440 -4308
rect 6383 -4372 6440 -4368
rect 4656 -5346 4660 -5300
rect 4660 -5346 4718 -5300
rect 4718 -5346 4722 -5300
rect 4656 -5352 4722 -5346
rect 6627 -4025 6698 -4021
rect 6627 -4080 6631 -4025
rect 6631 -4080 6691 -4025
rect 6691 -4080 6698 -4025
rect 6627 -4084 6698 -4080
rect 7712 -4024 7782 -4021
rect 7712 -4079 7716 -4024
rect 7716 -4079 7776 -4024
rect 7776 -4079 7782 -4024
rect 7712 -4083 7782 -4079
rect 10918 -3084 10998 -3078
rect 10918 -3138 10922 -3084
rect 10922 -3138 10994 -3084
rect 10994 -3138 10998 -3084
rect 7953 -4155 8012 -4141
rect 7953 -4189 7966 -4155
rect 7966 -4189 8000 -4155
rect 8000 -4189 8012 -4155
rect 7953 -4201 8012 -4189
rect 9527 -4024 9584 -4020
rect 9527 -4084 9531 -4024
rect 9531 -4084 9580 -4024
rect 9580 -4084 9584 -4024
rect 9527 -4088 9584 -4084
rect 9527 -4140 9584 -4136
rect 9527 -4200 9531 -4140
rect 9531 -4200 9580 -4140
rect 9580 -4200 9584 -4140
rect 9527 -4204 9584 -4200
rect 7594 -4309 7662 -4304
rect 7594 -4364 7598 -4309
rect 7598 -4364 7658 -4309
rect 7658 -4364 7662 -4309
rect 7594 -4369 7662 -4364
rect 9527 -4308 9584 -4304
rect 9527 -4368 9531 -4308
rect 9531 -4368 9580 -4308
rect 9580 -4368 9584 -4308
rect 9527 -4372 9584 -4368
rect 7788 -5342 7792 -5296
rect 7792 -5342 7850 -5296
rect 7850 -5342 7854 -5296
rect 7788 -5348 7854 -5342
rect 9771 -4025 9842 -4021
rect 9771 -4080 9775 -4025
rect 9775 -4080 9835 -4025
rect 9835 -4080 9842 -4025
rect 9771 -4084 9842 -4080
rect 10856 -4024 10926 -4021
rect 10856 -4079 10860 -4024
rect 10860 -4079 10920 -4024
rect 10920 -4079 10926 -4024
rect 10856 -4083 10926 -4079
rect 14120 -3088 14200 -3082
rect 14120 -3142 14124 -3088
rect 14124 -3142 14196 -3088
rect 14196 -3142 14200 -3088
rect 17264 -3088 17344 -3082
rect 17264 -3142 17268 -3088
rect 17268 -3142 17340 -3088
rect 17340 -3142 17344 -3088
rect 11097 -4155 11156 -4141
rect 11097 -4189 11110 -4155
rect 11110 -4189 11144 -4155
rect 11144 -4189 11156 -4155
rect 11097 -4201 11156 -4189
rect 12729 -4028 12786 -4024
rect 12729 -4088 12733 -4028
rect 12733 -4088 12782 -4028
rect 12782 -4088 12786 -4028
rect 12729 -4092 12786 -4088
rect 12729 -4144 12786 -4140
rect 12729 -4204 12733 -4144
rect 12733 -4204 12782 -4144
rect 12782 -4204 12786 -4144
rect 12729 -4208 12786 -4204
rect 10738 -4309 10806 -4304
rect 10738 -4364 10742 -4309
rect 10742 -4364 10802 -4309
rect 10802 -4364 10806 -4309
rect 10738 -4369 10806 -4364
rect 12729 -4312 12786 -4308
rect 12729 -4372 12733 -4312
rect 12733 -4372 12782 -4312
rect 12782 -4372 12786 -4312
rect 12729 -4376 12786 -4372
rect 10932 -5342 10936 -5296
rect 10936 -5342 10994 -5296
rect 10994 -5342 10998 -5296
rect 10932 -5348 10998 -5342
rect 12973 -4029 13044 -4025
rect 12973 -4084 12977 -4029
rect 12977 -4084 13037 -4029
rect 13037 -4084 13044 -4029
rect 12973 -4088 13044 -4084
rect 14058 -4028 14128 -4025
rect 14058 -4083 14062 -4028
rect 14062 -4083 14122 -4028
rect 14122 -4083 14128 -4028
rect 14058 -4087 14128 -4083
rect 14299 -4159 14358 -4145
rect 14299 -4193 14312 -4159
rect 14312 -4193 14346 -4159
rect 14346 -4193 14358 -4159
rect 14299 -4205 14358 -4193
rect 13940 -4313 14008 -4308
rect 13940 -4368 13944 -4313
rect 13944 -4368 14004 -4313
rect 14004 -4368 14008 -4313
rect 13940 -4373 14008 -4368
rect 15873 -4028 15930 -4024
rect 15873 -4088 15877 -4028
rect 15877 -4088 15926 -4028
rect 15926 -4088 15930 -4028
rect 15873 -4092 15930 -4088
rect 15873 -4144 15930 -4140
rect 15873 -4204 15877 -4144
rect 15877 -4204 15926 -4144
rect 15926 -4204 15930 -4144
rect 15873 -4208 15930 -4204
rect 15873 -4312 15930 -4308
rect 15873 -4372 15877 -4312
rect 15877 -4372 15926 -4312
rect 15926 -4372 15930 -4312
rect 15873 -4376 15930 -4372
rect 14134 -5346 14138 -5300
rect 14138 -5346 14196 -5300
rect 14196 -5346 14200 -5300
rect 14134 -5352 14200 -5346
rect 16117 -4029 16188 -4025
rect 16117 -4084 16121 -4029
rect 16121 -4084 16181 -4029
rect 16181 -4084 16188 -4029
rect 16117 -4088 16188 -4084
rect 17202 -4028 17272 -4025
rect 17202 -4083 17206 -4028
rect 17206 -4083 17266 -4028
rect 17266 -4083 17272 -4028
rect 17202 -4087 17272 -4083
rect 19259 -1293 19330 -1289
rect 19259 -1348 19263 -1293
rect 19263 -1348 19323 -1293
rect 19323 -1348 19330 -1293
rect 19259 -1352 19330 -1348
rect 20344 -1292 20414 -1289
rect 20344 -1347 20348 -1292
rect 20348 -1347 20408 -1292
rect 20408 -1347 20414 -1292
rect 20344 -1351 20414 -1347
rect 20585 -1423 20644 -1409
rect 20585 -1457 20598 -1423
rect 20598 -1457 20632 -1423
rect 20632 -1457 20644 -1423
rect 20585 -1469 20644 -1457
rect 23550 -352 23630 -346
rect 23550 -406 23554 -352
rect 23554 -406 23626 -352
rect 23626 -406 23630 -352
rect 22159 -1408 22216 -1404
rect 22159 -1468 22163 -1408
rect 22163 -1468 22212 -1408
rect 22212 -1468 22216 -1408
rect 22159 -1472 22216 -1468
rect 20226 -1577 20294 -1572
rect 20226 -1632 20230 -1577
rect 20230 -1632 20290 -1577
rect 20290 -1632 20294 -1577
rect 20226 -1637 20294 -1632
rect 21817 -1855 21888 -1784
rect 22159 -1576 22216 -1572
rect 22159 -1636 22163 -1576
rect 22163 -1636 22212 -1576
rect 22212 -1636 22216 -1576
rect 22159 -1640 22216 -1636
rect 20420 -2610 20424 -2564
rect 20424 -2610 20482 -2564
rect 20482 -2610 20486 -2564
rect 20420 -2616 20486 -2610
rect 22403 -1293 22474 -1289
rect 22403 -1348 22407 -1293
rect 22407 -1348 22467 -1293
rect 22467 -1348 22474 -1293
rect 22403 -1352 22474 -1348
rect 23488 -1292 23558 -1289
rect 23488 -1347 23492 -1292
rect 23492 -1347 23552 -1292
rect 23552 -1347 23558 -1292
rect 23488 -1351 23558 -1347
rect 23729 -1423 23788 -1409
rect 23729 -1457 23742 -1423
rect 23742 -1457 23776 -1423
rect 23776 -1457 23788 -1423
rect 23729 -1469 23788 -1457
rect 23370 -1577 23438 -1572
rect 23370 -1632 23374 -1577
rect 23374 -1632 23434 -1577
rect 23434 -1632 23438 -1577
rect 23370 -1637 23438 -1632
rect 25207 -1847 25266 -1777
rect 25206 -2032 25267 -1969
rect 25205 -2255 25267 -2189
rect 25205 -2443 25268 -2385
rect 23564 -2610 23568 -2564
rect 23568 -2610 23626 -2564
rect 23626 -2610 23630 -2564
rect 23564 -2616 23630 -2610
rect 25204 -2789 25268 -2728
rect 20396 -3084 20476 -3078
rect 20396 -3138 20400 -3084
rect 20400 -3138 20472 -3084
rect 20472 -3138 20476 -3084
rect 17443 -4159 17502 -4145
rect 17443 -4193 17456 -4159
rect 17456 -4193 17490 -4159
rect 17490 -4193 17502 -4159
rect 17443 -4205 17502 -4193
rect 19005 -4024 19062 -4020
rect 19005 -4084 19009 -4024
rect 19009 -4084 19058 -4024
rect 19058 -4084 19062 -4024
rect 19005 -4088 19062 -4084
rect 19005 -4140 19062 -4136
rect 19005 -4200 19009 -4140
rect 19009 -4200 19058 -4140
rect 19058 -4200 19062 -4140
rect 19005 -4204 19062 -4200
rect 17084 -4313 17152 -4308
rect 17084 -4368 17088 -4313
rect 17088 -4368 17148 -4313
rect 17148 -4368 17152 -4313
rect 17084 -4373 17152 -4368
rect 19005 -4308 19062 -4304
rect 19005 -4368 19009 -4308
rect 19009 -4368 19058 -4308
rect 19058 -4368 19062 -4308
rect 19005 -4372 19062 -4368
rect 17278 -5346 17282 -5300
rect 17282 -5346 17340 -5300
rect 17340 -5346 17344 -5300
rect 17278 -5352 17344 -5346
rect 19249 -4025 19320 -4021
rect 19249 -4080 19253 -4025
rect 19253 -4080 19313 -4025
rect 19313 -4080 19320 -4025
rect 19249 -4084 19320 -4080
rect 20334 -4024 20404 -4021
rect 20334 -4079 20338 -4024
rect 20338 -4079 20398 -4024
rect 20398 -4079 20404 -4024
rect 20334 -4083 20404 -4079
rect 23540 -3084 23620 -3078
rect 23540 -3138 23544 -3084
rect 23544 -3138 23616 -3084
rect 23616 -3138 23620 -3084
rect 25206 -2960 25270 -2900
rect 25205 -3315 25272 -3254
rect 20575 -4155 20634 -4141
rect 20575 -4189 20588 -4155
rect 20588 -4189 20622 -4155
rect 20622 -4189 20634 -4155
rect 20575 -4201 20634 -4189
rect 22149 -4024 22206 -4020
rect 22149 -4084 22153 -4024
rect 22153 -4084 22202 -4024
rect 22202 -4084 22206 -4024
rect 22149 -4088 22206 -4084
rect 22149 -4140 22206 -4136
rect 22149 -4200 22153 -4140
rect 22153 -4200 22202 -4140
rect 22202 -4200 22206 -4140
rect 22149 -4204 22206 -4200
rect 20216 -4309 20284 -4304
rect 20216 -4364 20220 -4309
rect 20220 -4364 20280 -4309
rect 20280 -4364 20284 -4309
rect 20216 -4369 20284 -4364
rect 22149 -4308 22206 -4304
rect 22149 -4368 22153 -4308
rect 22153 -4368 22202 -4308
rect 22202 -4368 22206 -4308
rect 22149 -4372 22206 -4368
rect 20410 -5342 20414 -5296
rect 20414 -5342 20472 -5296
rect 20472 -5342 20476 -5296
rect 20410 -5348 20476 -5342
rect 16877 -5981 16953 -5961
rect 814 -6028 868 -6020
rect 814 -6066 824 -6028
rect 824 -6066 862 -6028
rect 862 -6066 868 -6028
rect 2882 -6026 2936 -6018
rect 814 -6074 868 -6066
rect 2882 -6064 2892 -6026
rect 2892 -6064 2930 -6026
rect 2930 -6064 2936 -6026
rect 2882 -6072 2936 -6064
rect 4951 -6028 5005 -6020
rect 4951 -6066 4961 -6028
rect 4961 -6066 4999 -6028
rect 4999 -6066 5005 -6028
rect 7019 -6026 7073 -6018
rect 4951 -6074 5005 -6066
rect 7019 -6064 7029 -6026
rect 7029 -6064 7067 -6026
rect 7067 -6064 7073 -6026
rect 9088 -6026 9142 -6018
rect 7019 -6072 7073 -6064
rect 9088 -6064 9098 -6026
rect 9098 -6064 9136 -6026
rect 9136 -6064 9142 -6026
rect 11156 -6024 11210 -6016
rect 9088 -6072 9142 -6064
rect 11156 -6062 11166 -6024
rect 11166 -6062 11204 -6024
rect 11204 -6062 11210 -6024
rect 11156 -6070 11210 -6062
rect 13225 -6026 13279 -6018
rect 13225 -6064 13235 -6026
rect 13235 -6064 13273 -6026
rect 13273 -6064 13279 -6026
rect 15293 -6024 15347 -6016
rect 13225 -6072 13279 -6064
rect 15293 -6062 15303 -6024
rect 15303 -6062 15341 -6024
rect 15341 -6062 15347 -6024
rect 16877 -6017 16953 -5981
rect 16877 -6035 16953 -6017
rect 15293 -6070 15347 -6062
rect -703 -6873 -639 -6813
rect -280 -6882 -220 -6829
rect 6 -6888 72 -6822
rect -9 -7018 62 -7010
rect -280 -7079 -228 -7021
rect -9 -7078 -6 -7018
rect -6 -7078 60 -7018
rect 60 -7078 62 -7018
rect -9 -7087 62 -7078
rect 1394 -6882 1448 -6828
rect 2074 -6886 2140 -6820
rect 756 -8250 818 -8244
rect 756 -8292 762 -8250
rect 762 -8292 812 -8250
rect 812 -8292 818 -8250
rect 756 -8302 818 -8292
rect 3462 -6880 3516 -6826
rect 17615 -5983 17691 -5963
rect 17615 -6019 17691 -5983
rect 17615 -6037 17691 -6019
rect 18353 -5983 18429 -5963
rect 18353 -6019 18429 -5983
rect 18353 -6037 18429 -6019
rect 19095 -5983 19171 -5963
rect 19095 -6019 19171 -5983
rect 19095 -6037 19171 -6019
rect 19835 -5983 19911 -5963
rect 19835 -6019 19911 -5983
rect 19835 -6037 19911 -6019
rect 20573 -5983 20649 -5963
rect 20573 -6019 20649 -5983
rect 20573 -6037 20649 -6019
rect 21311 -5983 21387 -5963
rect 21311 -6019 21387 -5983
rect 21311 -6037 21387 -6019
rect 4143 -6888 4209 -6822
rect 2824 -8248 2886 -8242
rect 2824 -8290 2830 -8248
rect 2830 -8290 2880 -8248
rect 2880 -8290 2886 -8248
rect 2824 -8300 2886 -8290
rect 5531 -6882 5585 -6828
rect 6211 -6886 6277 -6820
rect 4893 -8250 4955 -8244
rect 4893 -8292 4899 -8250
rect 4899 -8292 4949 -8250
rect 4949 -8292 4955 -8250
rect 4893 -8302 4955 -8292
rect 7599 -6880 7653 -6826
rect 8280 -6886 8346 -6820
rect 6961 -8248 7023 -8242
rect 6961 -8290 6967 -8248
rect 6967 -8290 7017 -8248
rect 7017 -8290 7023 -8248
rect 6961 -8300 7023 -8290
rect 9668 -6880 9722 -6826
rect 10348 -6884 10414 -6818
rect 9030 -8248 9092 -8242
rect 9030 -8290 9036 -8248
rect 9036 -8290 9086 -8248
rect 9086 -8290 9092 -8248
rect 9030 -8300 9092 -8290
rect 11736 -6878 11790 -6824
rect 12417 -6886 12483 -6820
rect 11098 -8246 11160 -8240
rect 11098 -8288 11104 -8246
rect 11104 -8288 11154 -8246
rect 11154 -8288 11160 -8246
rect 11098 -8298 11160 -8288
rect 13805 -6880 13859 -6826
rect 14485 -6884 14551 -6818
rect 13167 -8248 13229 -8242
rect 13167 -8290 13173 -8248
rect 13173 -8290 13223 -8248
rect 13223 -8290 13229 -8248
rect 13167 -8300 13229 -8290
rect 15873 -6878 15927 -6824
rect 22393 -4025 22464 -4021
rect 22393 -4080 22397 -4025
rect 22397 -4080 22457 -4025
rect 22457 -4080 22464 -4025
rect 22393 -4084 22464 -4080
rect 23478 -4024 23548 -4021
rect 23478 -4079 23482 -4024
rect 23482 -4079 23542 -4024
rect 23542 -4079 23548 -4024
rect 23478 -4083 23548 -4079
rect 23719 -4155 23778 -4141
rect 23719 -4189 23732 -4155
rect 23732 -4189 23766 -4155
rect 23766 -4189 23778 -4155
rect 23719 -4201 23778 -4189
rect 23360 -4309 23428 -4304
rect 23360 -4364 23364 -4309
rect 23364 -4364 23424 -4309
rect 23424 -4364 23428 -4309
rect 23360 -4369 23428 -4364
rect 23554 -5342 23558 -5296
rect 23558 -5342 23616 -5296
rect 23616 -5342 23620 -5296
rect 23554 -5348 23620 -5342
rect 22049 -5983 22125 -5963
rect 22049 -6019 22125 -5983
rect 22049 -6037 22125 -6019
rect 16801 -6849 16903 -6843
rect 16801 -6903 16813 -6849
rect 16813 -6903 16891 -6849
rect 16891 -6903 16903 -6849
rect 16801 -6909 16903 -6903
rect 17539 -6851 17641 -6845
rect 17539 -6905 17551 -6851
rect 17551 -6905 17629 -6851
rect 17629 -6905 17641 -6851
rect 17539 -6911 17641 -6905
rect 18277 -6851 18379 -6845
rect 18277 -6905 18289 -6851
rect 18289 -6905 18367 -6851
rect 18367 -6905 18379 -6851
rect 18277 -6911 18379 -6905
rect 19019 -6851 19121 -6845
rect 19019 -6905 19031 -6851
rect 19031 -6905 19109 -6851
rect 19109 -6905 19121 -6851
rect 19019 -6911 19121 -6905
rect 19759 -6851 19861 -6845
rect 19759 -6905 19771 -6851
rect 19771 -6905 19849 -6851
rect 19849 -6905 19861 -6851
rect 19759 -6911 19861 -6905
rect 20497 -6851 20599 -6845
rect 20497 -6905 20509 -6851
rect 20509 -6905 20587 -6851
rect 20587 -6905 20599 -6851
rect 20497 -6911 20599 -6905
rect 21235 -6851 21337 -6845
rect 21235 -6905 21247 -6851
rect 21247 -6905 21325 -6851
rect 21325 -6905 21337 -6851
rect 21235 -6911 21337 -6905
rect 21973 -6851 22075 -6845
rect 21973 -6905 21985 -6851
rect 21985 -6905 22063 -6851
rect 22063 -6905 22075 -6851
rect 21973 -6911 22075 -6905
rect 15235 -8246 15297 -8240
rect 15235 -8288 15241 -8246
rect 15241 -8288 15291 -8246
rect 15291 -8288 15297 -8246
rect 15235 -8298 15297 -8288
<< metal2 >>
rect -2478 5922 -2418 5932
rect -2418 5901 10358 5911
rect -2418 5863 10304 5901
rect -2478 5853 -2418 5863
rect 10304 5837 10358 5847
rect -2481 5725 -2421 5732
rect 8766 5725 8820 5726
rect -2481 5722 8823 5725
rect -2421 5716 8823 5722
rect -2421 5662 8766 5716
rect 8820 5662 8823 5716
rect -2421 5660 8823 5662
rect -2481 5650 -2421 5660
rect -2488 5536 -2428 5542
rect 7305 5536 7359 5541
rect -2488 5532 7360 5536
rect -2428 5531 7360 5532
rect -2428 5477 7305 5531
rect 7359 5477 7360 5531
rect -2428 5470 7360 5477
rect -2488 5460 -2428 5470
rect -2488 5350 -2428 5360
rect 5803 5350 5857 5353
rect -2428 5343 5857 5350
rect -2428 5289 5803 5343
rect -2428 5281 5857 5289
rect -2488 5271 -2428 5281
rect 5802 5279 5857 5281
rect -2501 5163 -2440 5173
rect 4347 5163 4401 5169
rect -2440 5159 4401 5163
rect -2440 5105 4347 5159
rect -2440 5100 4401 5105
rect -2501 5090 -2440 5100
rect -2514 4972 -2443 4982
rect 2894 4973 2948 4983
rect -2443 4919 2894 4972
rect -2443 4900 2948 4919
rect -2514 4890 -2443 4900
rect 1449 4787 1503 4797
rect 542 4123 602 4133
rect 542 4051 602 4061
rect -293 3467 -222 3477
rect -293 3398 -222 3408
rect -7 3371 62 3381
rect -7 3297 62 3307
rect -2497 3166 -2443 3176
rect 1449 3168 1503 4733
rect 1559 4702 1613 4704
rect 1558 4694 1613 4702
rect 1558 4640 1559 4694
rect 1558 3298 1613 4640
rect 1990 4123 2050 4133
rect 1990 4051 2050 4061
rect 1766 3298 1820 3308
rect 1558 3244 1766 3298
rect 1766 3234 1820 3244
rect 1640 3185 1716 3195
rect -2022 3167 1510 3168
rect -2239 3166 1640 3167
rect -2443 3112 1640 3166
rect -2443 3111 1510 3112
rect -2497 3101 -2443 3111
rect 2894 3165 2948 4900
rect 3025 4878 3079 4888
rect 3025 3297 3079 4824
rect 3488 4125 3548 4135
rect 3488 4053 3548 4063
rect 3260 3297 3314 3307
rect 3025 3243 3260 3297
rect 3260 3233 3314 3243
rect 3142 3177 3206 3187
rect 2894 3111 3142 3165
rect 4347 3170 4401 5100
rect 4475 5064 4529 5074
rect 4475 3300 4529 5010
rect 4936 4125 4996 4135
rect 4936 4053 4996 4063
rect 4686 3300 4764 3310
rect 4475 3246 4710 3300
rect 4475 3245 4764 3246
rect 4686 3236 4764 3245
rect 4591 3183 4658 3193
rect 4347 3116 4591 3170
rect 5802 3170 5856 5279
rect 5982 5249 6036 5259
rect 5982 3295 6036 5195
rect 6456 4123 6516 4133
rect 6456 4051 6516 4061
rect 6229 3295 6283 3305
rect 5982 3241 6229 3295
rect 6229 3231 6283 3241
rect 6110 3181 6170 3191
rect 5802 3116 6110 3170
rect 1640 3088 1716 3098
rect 3142 3093 3206 3103
rect 4591 3095 4658 3105
rect 7305 3164 7359 5470
rect 7443 5437 7497 5447
rect 7443 3303 7497 5383
rect 7904 4123 7964 4133
rect 7904 4051 7964 4061
rect 7677 3303 7731 3312
rect 7443 3302 7731 3303
rect 7443 3248 7677 3302
rect 7677 3238 7731 3248
rect 7560 3174 7620 3184
rect 7305 3110 7560 3164
rect 8766 3170 8820 5660
rect 8941 5621 8995 5631
rect 8941 3390 8995 5567
rect 9402 4125 9462 4135
rect 9402 4053 9462 4063
rect 8941 3336 9228 3390
rect 9174 3300 9228 3336
rect 9174 3236 9228 3246
rect 9059 3183 9120 3193
rect 8766 3116 9059 3170
rect 6110 3096 6170 3106
rect 7560 3096 7620 3106
rect 9059 3094 9120 3104
rect 10307 3187 10357 5837
rect 10398 5808 10452 5818
rect 10398 5744 10452 5754
rect 10400 3407 10450 5744
rect 12514 4332 12604 4342
rect 12514 4231 12604 4241
rect 13682 4332 13772 4342
rect 13682 4231 13772 4241
rect 14850 4332 14940 4342
rect 14850 4231 14940 4241
rect 16018 4332 16108 4342
rect 16018 4231 16108 4241
rect 17192 4334 17282 4344
rect 17192 4233 17282 4243
rect 18360 4334 18450 4344
rect 18360 4233 18450 4243
rect 19528 4334 19618 4344
rect 19528 4233 19618 4243
rect 20696 4334 20786 4344
rect 20696 4233 20786 4243
rect 10850 4125 10910 4135
rect 10850 4053 10910 4063
rect 10400 3357 10678 3407
rect 10627 3326 10677 3357
rect 10606 3316 10692 3326
rect 10606 3218 10692 3228
rect 10493 3197 10578 3198
rect 10492 3188 10578 3197
rect 10492 3187 10493 3188
rect 10307 3099 10492 3187
rect 10492 3098 10493 3099
rect 10492 3089 10578 3098
rect 10493 3088 10578 3089
rect 12049 3005 12139 3015
rect 3710 2929 3772 2931
rect 5158 2929 5220 2931
rect 9624 2929 9686 2931
rect 11072 2929 11134 2931
rect 764 2927 826 2929
rect 2212 2927 2274 2929
rect 764 2919 828 2927
rect 826 2917 828 2919
rect 764 2845 828 2855
rect 2212 2919 2276 2927
rect 2274 2917 2276 2919
rect 2212 2845 2276 2855
rect 3710 2921 3774 2929
rect 3772 2919 3774 2921
rect 3710 2847 3774 2857
rect 5158 2921 5222 2929
rect 5220 2919 5222 2921
rect 5158 2847 5222 2857
rect 6678 2927 6740 2929
rect 8126 2927 8188 2929
rect 6678 2919 6742 2927
rect 6740 2917 6742 2919
rect 6678 2845 6742 2855
rect 8126 2919 8190 2927
rect 8188 2917 8190 2919
rect 8126 2845 8190 2855
rect 9624 2921 9688 2929
rect 9686 2919 9688 2921
rect 9624 2847 9688 2857
rect 11072 2921 11136 2929
rect 11134 2919 11136 2921
rect 12049 2904 12139 2914
rect 13217 3005 13307 3015
rect 13217 2904 13307 2914
rect 14385 3005 14475 3015
rect 14385 2904 14475 2914
rect 15553 3005 15643 3015
rect 15553 2904 15643 2914
rect 16727 3007 16817 3017
rect 16727 2906 16817 2916
rect 17895 3007 17985 3017
rect 17895 2906 17985 2916
rect 19063 3007 19153 3017
rect 19063 2906 19153 2916
rect 20231 3007 20321 3017
rect 20231 2906 20321 2916
rect 11072 2847 11136 2857
rect -2527 2792 -2469 2802
rect -2527 2726 -2469 2736
rect 1496 2412 1596 2422
rect 1496 2310 1596 2320
rect 4640 2412 4740 2422
rect 4640 2310 4740 2320
rect 7772 2416 7872 2426
rect 7772 2314 7872 2324
rect 10916 2416 11016 2426
rect 10916 2314 11016 2324
rect 14118 2412 14218 2422
rect 14118 2310 14218 2320
rect 17262 2412 17362 2422
rect 17262 2310 17362 2320
rect 20394 2416 20494 2426
rect 20394 2314 20494 2324
rect 23538 2416 23638 2426
rect 23538 2314 23638 2324
rect 6626 1455 6719 1457
rect 9770 1455 9863 1457
rect 19248 1455 19341 1457
rect 22392 1455 22485 1457
rect 350 1451 443 1453
rect 3494 1451 3587 1453
rect 6382 1451 7801 1455
rect 9526 1451 10945 1455
rect 12972 1451 13065 1453
rect 16116 1451 16209 1453
rect 19004 1451 20423 1455
rect 22148 1451 23567 1455
rect -519 1445 23567 1451
rect -519 1444 6637 1445
rect -519 1367 -503 1444
rect -420 1441 6637 1444
rect -420 1378 361 1441
rect 432 1379 1446 1441
rect 1516 1379 3505 1441
rect 432 1378 3505 1379
rect 3576 1379 4590 1441
rect 4660 1382 6637 1441
rect 6708 1383 7722 1445
rect 7792 1383 9781 1445
rect 6708 1382 9781 1383
rect 9852 1383 10866 1445
rect 10936 1441 19259 1445
rect 10936 1383 12983 1441
rect 9852 1382 12983 1383
rect 4660 1379 12983 1382
rect 3576 1378 12983 1379
rect 13054 1379 14068 1441
rect 14138 1379 16127 1441
rect 13054 1378 16127 1379
rect 16198 1379 17212 1441
rect 17282 1382 19259 1441
rect 19330 1383 20344 1445
rect 20414 1383 22403 1445
rect 19330 1382 22403 1383
rect 22474 1383 23488 1445
rect 23558 1383 23567 1445
rect 22474 1382 23567 1383
rect 17282 1379 23567 1382
rect 16198 1378 23567 1379
rect -420 1367 23567 1378
rect -503 1346 -420 1356
rect 3261 1334 3318 1336
rect 106 1331 202 1334
rect 3250 1331 3346 1334
rect 106 1326 1746 1331
rect 106 1258 117 1326
rect 174 1321 1746 1326
rect 174 1261 1687 1321
rect 174 1258 1746 1261
rect 106 1252 1746 1258
rect 106 1249 202 1252
rect 1687 1251 1746 1252
rect 3250 1326 4890 1331
rect 3250 1258 3261 1326
rect 3318 1321 4890 1326
rect 3318 1261 4831 1321
rect 3318 1258 4890 1261
rect 3250 1252 4890 1258
rect 6382 1330 8022 1335
rect 6382 1262 6393 1330
rect 6450 1325 8022 1330
rect 6450 1265 7963 1325
rect 6450 1262 8022 1265
rect 6382 1256 8022 1262
rect 7963 1255 8022 1256
rect 9526 1330 11166 1335
rect 9526 1262 9537 1330
rect 9594 1325 11166 1330
rect 9594 1265 11107 1325
rect 9594 1262 11166 1265
rect 9526 1256 11166 1262
rect 9526 1253 9622 1256
rect 11107 1255 11166 1256
rect 12728 1331 12824 1334
rect 15872 1331 15968 1334
rect 12728 1326 14368 1331
rect 12728 1258 12739 1326
rect 12796 1321 14368 1326
rect 12796 1261 14309 1321
rect 12796 1258 14368 1261
rect 9537 1252 9594 1253
rect 12728 1252 14368 1258
rect 3250 1249 3346 1252
rect 4831 1251 4890 1252
rect 12728 1249 12824 1252
rect 14309 1251 14368 1252
rect 15872 1326 17512 1331
rect 15872 1258 15883 1326
rect 15940 1321 17512 1326
rect 15940 1261 17453 1321
rect 15940 1258 17512 1261
rect 15872 1252 17512 1258
rect 19004 1330 20644 1335
rect 19004 1262 19015 1330
rect 19072 1325 20644 1330
rect 19072 1265 20585 1325
rect 19072 1262 20644 1265
rect 19004 1256 20644 1262
rect 19004 1253 19100 1256
rect 20585 1255 20644 1256
rect 22148 1330 23788 1335
rect 22148 1262 22159 1330
rect 22216 1325 23788 1330
rect 22216 1265 23729 1325
rect 22216 1262 23788 1265
rect 22148 1256 23788 1262
rect 22148 1253 22244 1256
rect 23729 1255 23788 1256
rect 19015 1252 19072 1253
rect 22159 1252 22216 1253
rect 15872 1249 15968 1252
rect 17453 1251 17512 1252
rect 117 1248 174 1249
rect 3261 1248 3318 1249
rect 12739 1248 12796 1249
rect 15883 1248 15940 1249
rect 6393 1171 6450 1172
rect 19015 1171 19072 1172
rect 22159 1171 22216 1172
rect 6382 1170 6478 1171
rect 19004 1170 19100 1171
rect 22148 1170 22244 1171
rect 117 1167 174 1168
rect 3261 1167 3318 1168
rect 106 1166 202 1167
rect 3250 1166 3346 1167
rect 106 1158 1407 1166
rect 106 1090 117 1158
rect 174 1093 1328 1158
rect 1396 1093 1407 1158
rect 174 1090 1407 1093
rect 106 1082 1407 1090
rect 3250 1158 4551 1166
rect 3250 1090 3261 1158
rect 3318 1093 4472 1158
rect 4540 1093 4551 1158
rect 3318 1090 4551 1093
rect 3250 1082 4551 1090
rect 6382 1162 7683 1170
rect 15883 1167 15940 1168
rect 6382 1094 6393 1162
rect 6450 1097 7604 1162
rect 7672 1097 7683 1162
rect 6450 1094 7683 1097
rect 6382 1086 7683 1094
rect 15872 1166 15968 1167
rect 15872 1158 17173 1166
rect 15872 1090 15883 1158
rect 15940 1093 17094 1158
rect 17162 1093 17173 1158
rect 15940 1090 17173 1093
rect 6393 1084 6450 1086
rect 15872 1082 17173 1090
rect 19004 1162 20305 1170
rect 19004 1094 19015 1162
rect 19072 1097 20226 1162
rect 20294 1097 20305 1162
rect 19072 1094 20305 1097
rect 19004 1086 20305 1094
rect 22148 1162 23449 1170
rect 22148 1094 22159 1162
rect 22216 1097 23370 1162
rect 23438 1097 23449 1162
rect 22216 1094 23449 1097
rect 22148 1086 23449 1094
rect 19015 1084 19072 1086
rect 22159 1084 22216 1086
rect 117 1080 174 1082
rect 3261 1080 3318 1082
rect 15883 1080 15940 1082
rect 1516 168 1592 178
rect 1516 100 1592 110
rect 4660 168 4736 178
rect 4660 100 4736 110
rect 7792 172 7868 182
rect 7792 104 7868 114
rect 10936 172 11012 182
rect 10936 104 11012 114
rect 14138 168 14214 178
rect 14138 100 14214 110
rect 17282 168 17358 178
rect 17282 100 17358 110
rect 20414 172 20490 182
rect 20414 104 20490 114
rect 23558 172 23634 182
rect 23558 104 23634 114
rect 1496 -322 1596 -312
rect 1496 -424 1596 -414
rect 4640 -322 4740 -312
rect 4640 -424 4740 -414
rect 7772 -318 7872 -308
rect 7772 -420 7872 -410
rect 10916 -318 11016 -308
rect 10916 -420 11016 -410
rect 14118 -322 14218 -312
rect 14118 -424 14218 -414
rect 17262 -322 17362 -312
rect 17262 -424 17362 -414
rect 20394 -318 20494 -308
rect 20394 -420 20494 -410
rect 23538 -318 23638 -308
rect 23538 -420 23638 -410
rect 9770 -1279 9863 -1277
rect 19248 -1279 19341 -1277
rect 22392 -1279 22485 -1277
rect -2507 -1283 -2445 -1279
rect 6385 -1280 10945 -1279
rect 19007 -1280 20423 -1279
rect 22151 -1280 23567 -1279
rect 350 -1283 443 -1281
rect 3494 -1283 3587 -1281
rect 6382 -1283 10945 -1280
rect 12972 -1283 13065 -1281
rect 16116 -1283 16209 -1281
rect 17229 -1283 23567 -1280
rect -2512 -1284 10945 -1283
rect 12731 -1284 14147 -1283
rect 15875 -1284 23567 -1283
rect -2512 -1285 14147 -1284
rect 15872 -1285 23567 -1284
rect -2512 -1289 23567 -1285
rect -2512 -1364 -2507 -1289
rect -2445 -1293 6637 -1289
rect -2445 -1356 361 -1293
rect 432 -1355 1446 -1293
rect 1516 -1355 3505 -1293
rect 432 -1356 3505 -1355
rect 3576 -1355 4590 -1293
rect 4660 -1352 6637 -1293
rect 6708 -1351 7722 -1289
rect 7792 -1351 9781 -1289
rect 6708 -1352 9781 -1351
rect 9852 -1351 10866 -1289
rect 10936 -1292 19259 -1289
rect 10936 -1293 15883 -1292
rect 10936 -1351 12983 -1293
rect 9852 -1352 12983 -1351
rect 4660 -1355 12983 -1352
rect 3576 -1356 12983 -1355
rect 13054 -1355 14068 -1293
rect 14138 -1355 15883 -1293
rect 13054 -1356 15883 -1355
rect -2445 -1360 15883 -1356
rect 15940 -1293 19259 -1292
rect 15940 -1356 16127 -1293
rect 16198 -1355 17212 -1293
rect 17282 -1352 19259 -1293
rect 19330 -1351 20344 -1289
rect 20414 -1351 22403 -1289
rect 19330 -1352 22403 -1351
rect 22474 -1351 23488 -1289
rect 23558 -1351 23567 -1289
rect 22474 -1352 23567 -1351
rect 17282 -1355 23567 -1352
rect 16198 -1356 23567 -1355
rect 15940 -1360 23567 -1356
rect -2445 -1363 23567 -1360
rect -2445 -1364 6460 -1363
rect -2512 -1366 6450 -1364
rect -2512 -1367 6413 -1366
rect 12728 -1367 19036 -1363
rect -2512 -1368 16 -1367
rect -2507 -1374 -2445 -1368
rect 9537 -1396 9594 -1394
rect 22159 -1396 22216 -1394
rect 117 -1400 174 -1398
rect 3261 -1400 3318 -1398
rect 9526 -1399 9622 -1396
rect 106 -1403 202 -1400
rect 3250 -1403 3346 -1400
rect 106 -1408 1746 -1403
rect 106 -1476 117 -1408
rect 174 -1413 1746 -1408
rect 174 -1473 1687 -1413
rect 174 -1476 1746 -1473
rect 106 -1482 1746 -1476
rect 106 -1485 202 -1482
rect 1687 -1483 1746 -1482
rect 3250 -1408 4890 -1403
rect 3250 -1476 3261 -1408
rect 3318 -1413 4890 -1408
rect 3318 -1473 4831 -1413
rect 3318 -1476 4890 -1473
rect 3250 -1482 4890 -1476
rect 6382 -1404 8022 -1399
rect 6382 -1472 6393 -1404
rect 6450 -1409 8022 -1404
rect 6450 -1469 7963 -1409
rect 6450 -1472 8022 -1469
rect 6382 -1478 8022 -1472
rect 6382 -1481 6478 -1478
rect 7963 -1479 8022 -1478
rect 9526 -1404 11166 -1399
rect 15883 -1400 15940 -1398
rect 22148 -1399 22244 -1396
rect 9526 -1472 9537 -1404
rect 9594 -1409 11166 -1404
rect 9594 -1469 11107 -1409
rect 9594 -1472 11166 -1469
rect 9526 -1478 11166 -1472
rect 9526 -1481 9622 -1478
rect 11107 -1479 11166 -1478
rect 12728 -1403 12824 -1400
rect 15872 -1403 15968 -1400
rect 12728 -1408 14368 -1403
rect 12728 -1476 12739 -1408
rect 12796 -1413 14368 -1408
rect 12796 -1473 14309 -1413
rect 12796 -1476 14368 -1473
rect 6393 -1482 6450 -1481
rect 9537 -1482 9594 -1481
rect 12728 -1482 14368 -1476
rect 3250 -1485 3346 -1482
rect 4831 -1483 4890 -1482
rect 12728 -1485 12824 -1482
rect 14309 -1483 14368 -1482
rect 15872 -1408 17512 -1403
rect 15872 -1476 15883 -1408
rect 15940 -1413 17512 -1408
rect 15940 -1473 17453 -1413
rect 15940 -1476 17512 -1473
rect 15872 -1482 17512 -1476
rect 19004 -1404 20644 -1399
rect 19004 -1472 19015 -1404
rect 19072 -1409 20644 -1404
rect 19072 -1469 20585 -1409
rect 19072 -1472 20644 -1469
rect 19004 -1478 20644 -1472
rect 19004 -1481 19100 -1478
rect 20585 -1479 20644 -1478
rect 22148 -1404 23788 -1399
rect 22148 -1472 22159 -1404
rect 22216 -1409 23788 -1404
rect 22216 -1469 23729 -1409
rect 22216 -1472 23788 -1469
rect 22148 -1478 23788 -1472
rect 22148 -1481 22244 -1478
rect 23729 -1479 23788 -1478
rect 19015 -1482 19072 -1481
rect 22159 -1482 22216 -1481
rect 15872 -1485 15968 -1482
rect 17453 -1483 17512 -1482
rect 117 -1486 174 -1485
rect 3261 -1486 3318 -1485
rect 12739 -1486 12796 -1485
rect 15883 -1486 15940 -1485
rect 6393 -1563 6450 -1562
rect 9537 -1563 9594 -1562
rect 19015 -1563 19072 -1562
rect 22159 -1563 22216 -1562
rect 6382 -1564 6478 -1563
rect 9526 -1564 9622 -1563
rect 19004 -1564 19100 -1563
rect 22148 -1564 22244 -1563
rect 117 -1567 174 -1566
rect 3261 -1567 3318 -1566
rect 106 -1568 202 -1567
rect 3250 -1568 3346 -1567
rect 106 -1576 1407 -1568
rect -2506 -1608 -2444 -1606
rect -496 -1608 -429 -1605
rect -2506 -1610 -409 -1608
rect -2511 -1615 -409 -1610
rect -2511 -1616 -496 -1615
rect -2511 -1691 -2506 -1616
rect -2444 -1685 -496 -1616
rect -429 -1685 -409 -1615
rect 106 -1644 117 -1576
rect 174 -1641 1328 -1576
rect 1396 -1641 1407 -1576
rect 174 -1644 1407 -1641
rect 106 -1652 1407 -1644
rect 3250 -1576 4551 -1568
rect 3250 -1644 3261 -1576
rect 3318 -1641 4472 -1576
rect 4540 -1641 4551 -1576
rect 3318 -1644 4551 -1641
rect 3250 -1652 4551 -1644
rect 6382 -1572 7683 -1564
rect 6382 -1640 6393 -1572
rect 6450 -1637 7604 -1572
rect 7672 -1637 7683 -1572
rect 6450 -1640 7683 -1637
rect 6382 -1648 7683 -1640
rect 9526 -1572 10827 -1564
rect 12739 -1567 12796 -1566
rect 15883 -1567 15940 -1566
rect 9526 -1640 9537 -1572
rect 9594 -1637 10748 -1572
rect 10816 -1637 10827 -1572
rect 9594 -1640 10827 -1637
rect 9526 -1648 10827 -1640
rect 12728 -1568 12824 -1567
rect 15872 -1568 15968 -1567
rect 12728 -1576 14029 -1568
rect 12728 -1644 12739 -1576
rect 12796 -1641 13950 -1576
rect 14018 -1641 14029 -1576
rect 12796 -1644 14029 -1641
rect 6393 -1650 6450 -1648
rect 9537 -1650 9594 -1648
rect 12728 -1652 14029 -1644
rect 15872 -1576 17173 -1568
rect 15872 -1644 15883 -1576
rect 15940 -1641 17094 -1576
rect 17162 -1641 17173 -1576
rect 15940 -1644 17173 -1641
rect 15872 -1652 17173 -1644
rect 19004 -1572 20305 -1564
rect 19004 -1640 19015 -1572
rect 19072 -1637 20226 -1572
rect 20294 -1637 20305 -1572
rect 19072 -1640 20305 -1637
rect 19004 -1648 20305 -1640
rect 22148 -1572 23449 -1564
rect 22148 -1640 22159 -1572
rect 22216 -1637 23370 -1572
rect 23438 -1637 23449 -1572
rect 22216 -1640 23449 -1637
rect 22148 -1648 23449 -1640
rect 19015 -1650 19072 -1648
rect 22159 -1650 22216 -1648
rect 117 -1654 174 -1652
rect 3261 -1654 3318 -1652
rect 12739 -1654 12796 -1652
rect 15883 -1654 15940 -1652
rect -2444 -1691 -409 -1685
rect -2511 -1694 -409 -1691
rect -2511 -1695 -2420 -1694
rect -496 -1695 -429 -1694
rect -2506 -1701 -2444 -1695
rect 21817 -1777 25266 -1767
rect 21817 -1784 25207 -1777
rect 21888 -1847 25207 -1784
rect 21888 -1855 25266 -1847
rect 21817 -1865 21888 -1855
rect 25207 -1857 25266 -1855
rect 18688 -1943 18758 -1933
rect 18758 -1969 25268 -1956
rect 18758 -2032 25206 -1969
rect 25267 -2032 25268 -1969
rect 18758 -2036 25268 -2032
rect 18688 -2042 25268 -2036
rect 18688 -2046 18758 -2042
rect 15529 -2172 15625 -2164
rect 15529 -2174 25268 -2172
rect 15625 -2189 25268 -2174
rect 15625 -2255 25205 -2189
rect 25267 -2255 25268 -2189
rect 15625 -2266 25268 -2255
rect 15529 -2279 15625 -2269
rect 12329 -2378 25269 -2368
rect 12407 -2385 25269 -2378
rect 12407 -2443 25205 -2385
rect 25268 -2443 25269 -2385
rect 12407 -2447 25269 -2443
rect 12329 -2454 25269 -2447
rect 12329 -2457 12407 -2454
rect 2936 -2530 3000 -2527
rect 2926 -2537 3011 -2530
rect 1516 -2566 1592 -2556
rect 1516 -2634 1592 -2624
rect 2926 -2614 2936 -2537
rect 3000 -2614 3011 -2537
rect 1486 -3054 1586 -3044
rect 1486 -3156 1586 -3146
rect 2926 -3235 3011 -2614
rect 4660 -2566 4736 -2556
rect 7792 -2562 7868 -2552
rect 6046 -2596 6114 -2586
rect 4660 -2634 4736 -2624
rect 6037 -2668 6046 -2608
rect 6114 -2668 6124 -2608
rect 7792 -2630 7868 -2620
rect 10936 -2562 11012 -2552
rect 10936 -2630 11012 -2620
rect 14138 -2566 14214 -2556
rect 14138 -2634 14214 -2624
rect 17282 -2566 17358 -2556
rect 17282 -2634 17358 -2624
rect 20414 -2562 20490 -2552
rect 20414 -2630 20490 -2620
rect 23558 -2562 23634 -2552
rect 23558 -2630 23634 -2620
rect 6037 -2884 6124 -2668
rect 9184 -2712 25269 -2711
rect 9182 -2722 25269 -2712
rect 9249 -2728 25269 -2722
rect 9249 -2789 25204 -2728
rect 25268 -2789 25269 -2728
rect 9249 -2790 25269 -2789
rect 9182 -2800 25269 -2790
rect 6037 -2900 25272 -2884
rect 6037 -2960 25206 -2900
rect 25270 -2960 25272 -2900
rect 6037 -2971 25272 -2960
rect 4630 -3054 4730 -3044
rect 4630 -3156 4730 -3146
rect 7762 -3050 7862 -3040
rect 7762 -3152 7862 -3142
rect 10906 -3050 11006 -3040
rect 10906 -3152 11006 -3142
rect 14108 -3054 14208 -3044
rect 14108 -3156 14208 -3146
rect 17252 -3054 17352 -3044
rect 17252 -3156 17352 -3146
rect 20384 -3050 20484 -3040
rect 20384 -3152 20484 -3142
rect 23528 -3050 23628 -3040
rect 23528 -3152 23628 -3142
rect 2926 -3254 25272 -3235
rect 2926 -3315 25205 -3254
rect 2926 -3327 25272 -3315
rect 2926 -3328 3011 -3327
rect 6383 -4011 6440 -4010
rect 6616 -4011 6709 -4009
rect 9527 -4011 9584 -4010
rect 9760 -4011 9853 -4009
rect 19005 -4011 19062 -4010
rect 19238 -4011 19331 -4009
rect 22149 -4011 22206 -4010
rect 22382 -4011 22475 -4009
rect 6375 -4012 7791 -4011
rect 9519 -4012 10935 -4011
rect 18997 -4012 20413 -4011
rect 22141 -4012 23557 -4011
rect 107 -4015 164 -4014
rect 340 -4015 433 -4013
rect 3251 -4015 3308 -4014
rect 3484 -4015 3577 -4013
rect 6372 -4015 7791 -4012
rect 9516 -4015 10935 -4012
rect 12729 -4015 12786 -4014
rect 12962 -4015 13055 -4013
rect 15873 -4015 15930 -4014
rect 16106 -4015 16199 -4013
rect 18994 -4015 20413 -4012
rect 22138 -4015 23557 -4012
rect 96 -4020 23557 -4015
rect 96 -4024 6383 -4020
rect 96 -4092 107 -4024
rect 164 -4025 3251 -4024
rect 164 -4088 351 -4025
rect 422 -4087 1436 -4025
rect 1506 -4087 3251 -4025
rect 422 -4088 3251 -4087
rect 164 -4092 3251 -4088
rect 3308 -4025 6383 -4024
rect 3308 -4088 3495 -4025
rect 3566 -4087 4580 -4025
rect 4650 -4087 6383 -4025
rect 3566 -4088 6383 -4087
rect 6440 -4021 9527 -4020
rect 6440 -4084 6627 -4021
rect 6698 -4083 7712 -4021
rect 7782 -4083 9527 -4021
rect 6698 -4084 9527 -4083
rect 6440 -4088 9527 -4084
rect 9584 -4021 19005 -4020
rect 9584 -4084 9771 -4021
rect 9842 -4083 10856 -4021
rect 10926 -4024 19005 -4021
rect 10926 -4083 12729 -4024
rect 9842 -4084 12729 -4083
rect 9584 -4088 12729 -4084
rect 3308 -4092 12729 -4088
rect 12786 -4025 15873 -4024
rect 12786 -4088 12973 -4025
rect 13044 -4087 14058 -4025
rect 14128 -4087 15873 -4025
rect 13044 -4088 15873 -4087
rect 12786 -4092 15873 -4088
rect 15930 -4025 19005 -4024
rect 15930 -4088 16117 -4025
rect 16188 -4087 17202 -4025
rect 17272 -4087 19005 -4025
rect 16188 -4088 19005 -4087
rect 19062 -4021 22149 -4020
rect 19062 -4084 19249 -4021
rect 19320 -4083 20334 -4021
rect 20404 -4083 22149 -4021
rect 19320 -4084 22149 -4083
rect 19062 -4088 22149 -4084
rect 22206 -4021 23557 -4020
rect 22206 -4084 22393 -4021
rect 22464 -4083 23478 -4021
rect 23548 -4083 23557 -4021
rect 22464 -4084 23557 -4083
rect 22206 -4088 23557 -4084
rect 15930 -4092 23557 -4088
rect 96 -4100 23557 -4092
rect 107 -4102 164 -4100
rect 3251 -4102 3308 -4100
rect 12729 -4102 12786 -4100
rect 15873 -4102 15930 -4100
rect 107 -4132 164 -4130
rect 3251 -4132 3308 -4130
rect 96 -4135 192 -4132
rect 3240 -4135 3336 -4132
rect 96 -4140 1736 -4135
rect 96 -4208 107 -4140
rect 164 -4145 1736 -4140
rect 164 -4205 1677 -4145
rect 164 -4208 1736 -4205
rect 96 -4214 1736 -4208
rect 96 -4217 192 -4214
rect 1677 -4215 1736 -4214
rect 3240 -4140 4880 -4135
rect 3240 -4208 3251 -4140
rect 3308 -4145 4880 -4140
rect 3308 -4205 4821 -4145
rect 3308 -4208 4880 -4205
rect 3240 -4214 4880 -4208
rect 6372 -4136 8012 -4131
rect 6372 -4204 6383 -4136
rect 6440 -4141 8012 -4136
rect 6440 -4201 7953 -4141
rect 6440 -4204 8012 -4201
rect 6372 -4210 8012 -4204
rect 6372 -4213 6468 -4210
rect 7953 -4211 8012 -4210
rect 9516 -4136 11156 -4131
rect 12729 -4132 12786 -4130
rect 15873 -4132 15930 -4130
rect 9516 -4204 9527 -4136
rect 9584 -4141 11156 -4136
rect 9584 -4201 11097 -4141
rect 9584 -4204 11156 -4201
rect 9516 -4210 11156 -4204
rect 9516 -4213 9612 -4210
rect 11097 -4211 11156 -4210
rect 12718 -4135 12814 -4132
rect 15862 -4135 15958 -4132
rect 12718 -4140 14358 -4135
rect 12718 -4208 12729 -4140
rect 12786 -4145 14358 -4140
rect 12786 -4205 14299 -4145
rect 12786 -4208 14358 -4205
rect 6383 -4214 6440 -4213
rect 9527 -4214 9584 -4213
rect 12718 -4214 14358 -4208
rect 3240 -4217 3336 -4214
rect 4821 -4215 4880 -4214
rect 12718 -4217 12814 -4214
rect 14299 -4215 14358 -4214
rect 15862 -4140 17502 -4135
rect 15862 -4208 15873 -4140
rect 15930 -4145 17502 -4140
rect 15930 -4205 17443 -4145
rect 15930 -4208 17502 -4205
rect 15862 -4214 17502 -4208
rect 18994 -4136 20634 -4131
rect 18994 -4204 19005 -4136
rect 19062 -4141 20634 -4136
rect 19062 -4201 20575 -4141
rect 19062 -4204 20634 -4201
rect 18994 -4210 20634 -4204
rect 18994 -4213 19090 -4210
rect 20575 -4211 20634 -4210
rect 22138 -4136 23778 -4131
rect 22138 -4204 22149 -4136
rect 22206 -4141 23778 -4136
rect 22206 -4201 23719 -4141
rect 22206 -4204 23778 -4201
rect 22138 -4210 23778 -4204
rect 22138 -4213 22234 -4210
rect 23719 -4211 23778 -4210
rect 19005 -4214 19062 -4213
rect 22149 -4214 22206 -4213
rect 15862 -4217 15958 -4214
rect 17443 -4215 17502 -4214
rect 107 -4218 164 -4217
rect 3251 -4218 3308 -4217
rect 12729 -4218 12786 -4217
rect 15873 -4218 15930 -4217
rect 6383 -4295 6440 -4294
rect 9527 -4295 9584 -4294
rect 19005 -4295 19062 -4294
rect 22149 -4295 22206 -4294
rect 6372 -4296 6468 -4295
rect 9516 -4296 9612 -4295
rect 18994 -4296 19090 -4295
rect 22138 -4296 22234 -4295
rect 107 -4299 164 -4298
rect 3251 -4299 3308 -4298
rect 96 -4300 192 -4299
rect 3240 -4300 3336 -4299
rect 96 -4308 1397 -4300
rect 96 -4376 107 -4308
rect 164 -4373 1318 -4308
rect 1386 -4373 1397 -4308
rect 164 -4376 1397 -4373
rect 96 -4384 1397 -4376
rect 3240 -4308 4541 -4300
rect 3240 -4376 3251 -4308
rect 3308 -4373 4462 -4308
rect 4530 -4373 4541 -4308
rect 3308 -4376 4541 -4373
rect 3240 -4384 4541 -4376
rect 6372 -4304 7673 -4296
rect 6372 -4372 6383 -4304
rect 6440 -4369 7594 -4304
rect 7662 -4369 7673 -4304
rect 6440 -4372 7673 -4369
rect 6372 -4380 7673 -4372
rect 9516 -4304 10817 -4296
rect 12729 -4299 12786 -4298
rect 15873 -4299 15930 -4298
rect 9516 -4372 9527 -4304
rect 9584 -4369 10738 -4304
rect 10806 -4369 10817 -4304
rect 9584 -4372 10817 -4369
rect 9516 -4380 10817 -4372
rect 12718 -4300 12814 -4299
rect 15862 -4300 15958 -4299
rect 12718 -4308 14019 -4300
rect 12718 -4376 12729 -4308
rect 12786 -4373 13940 -4308
rect 14008 -4373 14019 -4308
rect 12786 -4376 14019 -4373
rect 6383 -4382 6440 -4380
rect 9527 -4382 9584 -4380
rect 12718 -4384 14019 -4376
rect 15862 -4308 17163 -4300
rect 15862 -4376 15873 -4308
rect 15930 -4373 17084 -4308
rect 17152 -4373 17163 -4308
rect 15930 -4376 17163 -4373
rect 15862 -4384 17163 -4376
rect 18994 -4304 20295 -4296
rect 18994 -4372 19005 -4304
rect 19062 -4369 20216 -4304
rect 20284 -4369 20295 -4304
rect 19062 -4372 20295 -4369
rect 18994 -4380 20295 -4372
rect 22138 -4304 23439 -4296
rect 22138 -4372 22149 -4304
rect 22206 -4369 23360 -4304
rect 23428 -4369 23439 -4304
rect 22206 -4372 23439 -4369
rect 22138 -4380 23439 -4372
rect 19005 -4382 19062 -4380
rect 22149 -4382 22206 -4380
rect 107 -4386 164 -4384
rect 3251 -4386 3308 -4384
rect 12729 -4386 12786 -4384
rect 15873 -4386 15930 -4384
rect 1506 -5298 1582 -5288
rect 1506 -5366 1582 -5356
rect 4650 -5298 4726 -5288
rect 4650 -5366 4726 -5356
rect 7782 -5294 7858 -5284
rect 7782 -5362 7858 -5352
rect 10926 -5294 11002 -5284
rect 10926 -5362 11002 -5352
rect 14128 -5298 14204 -5288
rect 14128 -5366 14204 -5356
rect 17272 -5298 17348 -5288
rect 17272 -5366 17348 -5356
rect 20404 -5294 20480 -5284
rect 20404 -5362 20480 -5352
rect 23548 -5294 23624 -5284
rect 23548 -5362 23624 -5352
rect -2237 -5556 -2182 -5547
rect -1981 -5556 -1913 -5547
rect -2237 -5557 -1909 -5556
rect -2182 -5615 -1981 -5557
rect -1913 -5615 -1909 -5557
rect -2182 -5618 -1909 -5615
rect -2237 -5628 -2182 -5618
rect -1981 -5625 -1913 -5618
rect -2237 -5848 -2182 -5839
rect -2237 -5849 -2167 -5848
rect -1722 -5849 -1666 -5841
rect -2182 -5851 -1655 -5849
rect -2182 -5908 -1722 -5851
rect -1666 -5908 -1655 -5851
rect -2182 -5910 -1655 -5908
rect -2237 -5920 -2182 -5910
rect -1722 -5918 -1666 -5910
rect 16869 -5951 16963 -5941
rect 802 -6012 880 -6002
rect 802 -6092 880 -6082
rect 2870 -6010 2948 -6000
rect 2870 -6090 2948 -6080
rect 4939 -6012 5017 -6002
rect 4939 -6092 5017 -6082
rect 7007 -6010 7085 -6000
rect 7007 -6090 7085 -6080
rect 9076 -6010 9154 -6000
rect 9076 -6090 9154 -6080
rect 11144 -6008 11222 -5998
rect 11144 -6088 11222 -6078
rect 13213 -6010 13291 -6000
rect 13213 -6090 13291 -6080
rect 15281 -6008 15359 -5998
rect 16869 -6045 16963 -6035
rect 17607 -5953 17701 -5943
rect 17607 -6047 17701 -6037
rect 18345 -5953 18439 -5943
rect 18345 -6047 18439 -6037
rect 19087 -5953 19181 -5943
rect 19087 -6047 19181 -6037
rect 19827 -5953 19921 -5943
rect 19827 -6047 19921 -6037
rect 20565 -5953 20659 -5943
rect 20565 -6047 20659 -6037
rect 21303 -5953 21397 -5943
rect 21303 -6047 21397 -6037
rect 22041 -5953 22135 -5943
rect 22041 -6047 22135 -6037
rect 15281 -6088 15359 -6078
rect -2237 -6153 -2182 -6144
rect -2237 -6154 -2167 -6153
rect -1504 -6154 -1443 -6149
rect -2182 -6159 -1441 -6154
rect -2182 -6212 -1504 -6159
rect -1443 -6212 -1441 -6159
rect -2182 -6215 -1441 -6212
rect -2237 -6225 -2182 -6215
rect -1504 -6222 -1443 -6215
rect -2237 -6314 -2182 -6305
rect -2237 -6315 -2167 -6314
rect -1329 -6315 -1259 -6306
rect -2182 -6316 -1254 -6315
rect -2182 -6374 -1329 -6316
rect -1259 -6374 -1254 -6316
rect -2182 -6376 -1254 -6374
rect -2237 -6386 -2182 -6376
rect -1329 -6384 -1259 -6376
rect -2237 -6465 -2181 -6456
rect -2237 -6466 -2180 -6465
rect -1127 -6466 -1059 -6456
rect -2181 -6524 -1127 -6466
rect -1059 -6524 -1056 -6466
rect -2181 -6527 -1056 -6524
rect -2237 -6537 -2181 -6527
rect -1127 -6534 -1059 -6527
rect -2237 -6625 -2182 -6616
rect -2237 -6626 -2167 -6625
rect -931 -6626 -873 -6619
rect -2182 -6629 -869 -6626
rect -2182 -6683 -931 -6629
rect -873 -6683 -869 -6629
rect -2182 -6687 -869 -6683
rect -2237 -6697 -2182 -6687
rect -931 -6693 -873 -6687
rect -2237 -6812 -2182 -6803
rect -703 -6812 -639 -6803
rect 2069 -6804 2144 -6794
rect -2237 -6813 -638 -6812
rect -2182 -6873 -703 -6813
rect -639 -6873 -638 -6813
rect -2182 -6874 -638 -6873
rect -282 -6828 -216 -6818
rect -2237 -6884 -2182 -6874
rect -703 -6883 -639 -6874
rect -282 -6895 -216 -6885
rect 0 -6888 6 -6822
rect 72 -6828 1448 -6822
rect 72 -6882 1394 -6828
rect 72 -6888 1448 -6882
rect 2068 -6886 2069 -6820
rect 2144 -6826 3516 -6820
rect 4140 -6822 4209 -6812
rect 6212 -6820 6276 -6811
rect 8280 -6818 8347 -6808
rect 10343 -6818 10408 -6808
rect 14478 -6809 14561 -6799
rect 2144 -6880 3462 -6826
rect 2144 -6886 3516 -6880
rect 4137 -6888 4140 -6822
rect 4209 -6828 5585 -6822
rect 4209 -6882 5531 -6828
rect 4209 -6888 5585 -6882
rect 6205 -6886 6211 -6820
rect 6277 -6826 7653 -6820
rect 6277 -6880 7599 -6826
rect 6277 -6886 7653 -6880
rect 8274 -6886 8280 -6820
rect 8347 -6826 9722 -6820
rect 8347 -6880 9668 -6826
rect 8347 -6886 9722 -6880
rect 10342 -6884 10343 -6818
rect 10414 -6824 11790 -6818
rect 12414 -6820 12481 -6811
rect 10414 -6878 11736 -6824
rect 10414 -6884 11790 -6878
rect 12411 -6821 12417 -6820
rect 12411 -6885 12414 -6821
rect 12483 -6826 13859 -6820
rect 12483 -6880 13805 -6826
rect 12411 -6886 12417 -6885
rect 12483 -6886 13859 -6880
rect 14561 -6824 15927 -6818
rect 14561 -6878 15873 -6824
rect 14561 -6884 15927 -6878
rect 16801 -6839 16903 -6833
rect 16801 -6843 16905 -6839
rect 2069 -6900 2144 -6890
rect 4140 -6898 4209 -6888
rect 6212 -6896 6276 -6886
rect 8280 -6897 8347 -6887
rect 10343 -6896 10408 -6886
rect 12414 -6895 12481 -6886
rect 14478 -6899 14561 -6889
rect 16903 -6909 16905 -6843
rect 16801 -6917 16905 -6909
rect 17539 -6841 17641 -6835
rect 18277 -6841 18379 -6835
rect 19019 -6841 19121 -6835
rect 19759 -6841 19861 -6835
rect 20497 -6841 20599 -6835
rect 21235 -6841 21337 -6835
rect 21973 -6841 22075 -6835
rect 17539 -6845 17643 -6841
rect 17641 -6911 17643 -6845
rect 16801 -6919 16903 -6917
rect 17539 -6919 17643 -6911
rect 18277 -6845 18381 -6841
rect 18379 -6911 18381 -6845
rect 18277 -6919 18381 -6911
rect 19019 -6845 19123 -6841
rect 19121 -6911 19123 -6845
rect 19019 -6919 19123 -6911
rect 19759 -6845 19863 -6841
rect 19861 -6911 19863 -6845
rect 19759 -6919 19863 -6911
rect 20497 -6845 20601 -6841
rect 20599 -6911 20601 -6845
rect 20497 -6919 20601 -6911
rect 21235 -6845 21339 -6841
rect 21337 -6911 21339 -6845
rect 21235 -6919 21339 -6911
rect 21973 -6845 22077 -6841
rect 22075 -6911 22077 -6845
rect 21973 -6919 22077 -6911
rect 17539 -6921 17641 -6919
rect 18277 -6921 18379 -6919
rect 19019 -6921 19121 -6919
rect 19759 -6921 19861 -6919
rect 20497 -6921 20599 -6919
rect 21235 -6921 21337 -6919
rect 21973 -6921 22075 -6919
rect -2237 -7019 -2182 -7009
rect -9 -7010 62 -7000
rect -280 -7020 -228 -7011
rect -2182 -7021 -228 -7020
rect -2182 -7079 -280 -7021
rect -2237 -7090 -2182 -7080
rect -280 -7089 -228 -7079
rect -9 -7097 62 -7087
rect 750 -8242 822 -8232
rect 750 -8322 822 -8312
rect 2818 -8240 2890 -8230
rect 2818 -8320 2890 -8310
rect 4887 -8242 4959 -8232
rect 4887 -8322 4959 -8312
rect 6955 -8240 7027 -8230
rect 6955 -8320 7027 -8310
rect 9024 -8240 9096 -8230
rect 9024 -8320 9096 -8310
rect 11092 -8238 11164 -8228
rect 11092 -8318 11164 -8308
rect 13161 -8240 13233 -8230
rect 13161 -8320 13233 -8310
rect 15229 -8238 15301 -8228
rect 15229 -8318 15301 -8308
<< via2 >>
rect 542 4061 602 4123
rect -293 3408 -222 3467
rect -7 3307 62 3371
rect 1990 4061 2050 4123
rect 1640 3167 1716 3185
rect 1640 3112 1651 3167
rect 1651 3112 1705 3167
rect 1705 3112 1716 3167
rect 1640 3098 1716 3112
rect 3488 4063 3548 4125
rect 3142 3165 3206 3177
rect 3142 3111 3149 3165
rect 3149 3111 3203 3165
rect 3203 3111 3206 3165
rect 4936 4063 4996 4125
rect 4591 3170 4658 3183
rect 4591 3116 4597 3170
rect 4597 3116 4651 3170
rect 4651 3116 4658 3170
rect 6456 4061 6516 4123
rect 6110 3170 6170 3181
rect 6110 3116 6113 3170
rect 6113 3116 6167 3170
rect 6167 3116 6170 3170
rect 3142 3103 3206 3111
rect 4591 3105 4658 3116
rect 6110 3106 6170 3116
rect 7904 4061 7964 4123
rect 7560 3164 7620 3174
rect 7560 3110 7565 3164
rect 7565 3110 7619 3164
rect 7619 3110 7620 3164
rect 9402 4063 9462 4125
rect 9059 3170 9120 3183
rect 9059 3116 9062 3170
rect 9062 3116 9116 3170
rect 9116 3116 9120 3170
rect 7560 3106 7620 3110
rect 9059 3104 9120 3116
rect 12514 4311 12604 4332
rect 12514 4259 12536 4311
rect 12536 4259 12588 4311
rect 12588 4259 12604 4311
rect 12514 4241 12604 4259
rect 13682 4311 13772 4332
rect 13682 4259 13704 4311
rect 13704 4259 13756 4311
rect 13756 4259 13772 4311
rect 13682 4241 13772 4259
rect 14850 4311 14940 4332
rect 14850 4259 14872 4311
rect 14872 4259 14924 4311
rect 14924 4259 14940 4311
rect 14850 4241 14940 4259
rect 16018 4311 16108 4332
rect 16018 4259 16040 4311
rect 16040 4259 16092 4311
rect 16092 4259 16108 4311
rect 16018 4241 16108 4259
rect 17192 4313 17282 4334
rect 17192 4261 17214 4313
rect 17214 4261 17266 4313
rect 17266 4261 17282 4313
rect 17192 4243 17282 4261
rect 18360 4313 18450 4334
rect 18360 4261 18382 4313
rect 18382 4261 18434 4313
rect 18434 4261 18450 4313
rect 18360 4243 18450 4261
rect 19528 4313 19618 4334
rect 19528 4261 19550 4313
rect 19550 4261 19602 4313
rect 19602 4261 19618 4313
rect 19528 4243 19618 4261
rect 20696 4313 20786 4334
rect 20696 4261 20718 4313
rect 20718 4261 20770 4313
rect 20770 4261 20786 4313
rect 20696 4243 20786 4261
rect 10850 4063 10910 4125
rect 10493 3187 10578 3188
rect 10493 3099 10578 3187
rect 10493 3098 10578 3099
rect 12049 2987 12139 3005
rect 12049 2935 12065 2987
rect 12065 2935 12117 2987
rect 12117 2935 12139 2987
rect 764 2859 826 2917
rect 826 2859 828 2917
rect 764 2855 828 2859
rect 2212 2859 2274 2917
rect 2274 2859 2276 2917
rect 2212 2855 2276 2859
rect 3710 2861 3772 2919
rect 3772 2861 3774 2919
rect 3710 2857 3774 2861
rect 5158 2861 5220 2919
rect 5220 2861 5222 2919
rect 5158 2857 5222 2861
rect 6678 2859 6740 2917
rect 6740 2859 6742 2917
rect 6678 2855 6742 2859
rect 8126 2859 8188 2917
rect 8188 2859 8190 2917
rect 8126 2855 8190 2859
rect 9624 2861 9686 2919
rect 9686 2861 9688 2919
rect 9624 2857 9688 2861
rect 11072 2861 11134 2919
rect 11134 2861 11136 2919
rect 12049 2914 12139 2935
rect 13217 2987 13307 3005
rect 13217 2935 13233 2987
rect 13233 2935 13285 2987
rect 13285 2935 13307 2987
rect 13217 2914 13307 2935
rect 14385 2987 14475 3005
rect 14385 2935 14401 2987
rect 14401 2935 14453 2987
rect 14453 2935 14475 2987
rect 14385 2914 14475 2935
rect 15553 2987 15643 3005
rect 15553 2935 15569 2987
rect 15569 2935 15621 2987
rect 15621 2935 15643 2987
rect 15553 2914 15643 2935
rect 16727 2989 16817 3007
rect 16727 2937 16743 2989
rect 16743 2937 16795 2989
rect 16795 2937 16817 2989
rect 16727 2916 16817 2937
rect 17895 2989 17985 3007
rect 17895 2937 17911 2989
rect 17911 2937 17963 2989
rect 17963 2937 17985 2989
rect 17895 2916 17985 2937
rect 19063 2989 19153 3007
rect 19063 2937 19079 2989
rect 19079 2937 19131 2989
rect 19131 2937 19153 2989
rect 19063 2916 19153 2937
rect 20231 2989 20321 3007
rect 20231 2937 20247 2989
rect 20247 2937 20299 2989
rect 20299 2937 20321 2989
rect 20231 2916 20321 2937
rect 11072 2857 11136 2861
rect -2527 2791 -2469 2792
rect -2527 2737 -2526 2791
rect -2526 2737 -2470 2791
rect -2470 2737 -2469 2791
rect -2527 2736 -2469 2737
rect 1496 2384 1596 2412
rect 1496 2324 1508 2384
rect 1508 2324 1588 2384
rect 1588 2324 1596 2384
rect 1496 2320 1596 2324
rect 4640 2384 4740 2412
rect 4640 2324 4652 2384
rect 4652 2324 4732 2384
rect 4732 2324 4740 2384
rect 4640 2320 4740 2324
rect 7772 2388 7872 2416
rect 7772 2328 7784 2388
rect 7784 2328 7864 2388
rect 7864 2328 7872 2388
rect 7772 2324 7872 2328
rect 10916 2388 11016 2416
rect 10916 2328 10928 2388
rect 10928 2328 11008 2388
rect 11008 2328 11016 2388
rect 10916 2324 11016 2328
rect 14118 2384 14218 2412
rect 14118 2324 14130 2384
rect 14130 2324 14210 2384
rect 14210 2324 14218 2384
rect 14118 2320 14218 2324
rect 17262 2384 17362 2412
rect 17262 2324 17274 2384
rect 17274 2324 17354 2384
rect 17354 2324 17362 2384
rect 17262 2320 17362 2324
rect 20394 2388 20494 2416
rect 20394 2328 20406 2388
rect 20406 2328 20486 2388
rect 20486 2328 20494 2388
rect 20394 2324 20494 2328
rect 23538 2388 23638 2416
rect 23538 2328 23550 2388
rect 23550 2328 23630 2388
rect 23630 2328 23638 2388
rect 23538 2324 23638 2328
rect 1516 166 1592 168
rect 1516 114 1522 166
rect 1522 114 1588 166
rect 1588 114 1592 166
rect 1516 110 1592 114
rect 4660 166 4736 168
rect 4660 114 4666 166
rect 4666 114 4732 166
rect 4732 114 4736 166
rect 4660 110 4736 114
rect 7792 170 7868 172
rect 7792 118 7798 170
rect 7798 118 7864 170
rect 7864 118 7868 170
rect 7792 114 7868 118
rect 10936 170 11012 172
rect 10936 118 10942 170
rect 10942 118 11008 170
rect 11008 118 11012 170
rect 10936 114 11012 118
rect 14138 166 14214 168
rect 14138 114 14144 166
rect 14144 114 14210 166
rect 14210 114 14214 166
rect 14138 110 14214 114
rect 17282 166 17358 168
rect 17282 114 17288 166
rect 17288 114 17354 166
rect 17354 114 17358 166
rect 17282 110 17358 114
rect 20414 170 20490 172
rect 20414 118 20420 170
rect 20420 118 20486 170
rect 20486 118 20490 170
rect 20414 114 20490 118
rect 23558 170 23634 172
rect 23558 118 23564 170
rect 23564 118 23630 170
rect 23630 118 23634 170
rect 23558 114 23634 118
rect 1496 -350 1596 -322
rect 1496 -410 1508 -350
rect 1508 -410 1588 -350
rect 1588 -410 1596 -350
rect 1496 -414 1596 -410
rect 4640 -350 4740 -322
rect 4640 -410 4652 -350
rect 4652 -410 4732 -350
rect 4732 -410 4740 -350
rect 4640 -414 4740 -410
rect 7772 -346 7872 -318
rect 7772 -406 7784 -346
rect 7784 -406 7864 -346
rect 7864 -406 7872 -346
rect 7772 -410 7872 -406
rect 10916 -346 11016 -318
rect 10916 -406 10928 -346
rect 10928 -406 11008 -346
rect 11008 -406 11016 -346
rect 10916 -410 11016 -406
rect 14118 -350 14218 -322
rect 14118 -410 14130 -350
rect 14130 -410 14210 -350
rect 14210 -410 14218 -350
rect 14118 -414 14218 -410
rect 17262 -350 17362 -322
rect 17262 -410 17274 -350
rect 17274 -410 17354 -350
rect 17354 -410 17362 -350
rect 17262 -414 17362 -410
rect 20394 -346 20494 -318
rect 20394 -406 20406 -346
rect 20406 -406 20486 -346
rect 20486 -406 20494 -346
rect 20394 -410 20494 -406
rect 23538 -346 23638 -318
rect 23538 -406 23550 -346
rect 23550 -406 23630 -346
rect 23630 -406 23638 -346
rect 23538 -410 23638 -406
rect 1516 -2568 1592 -2566
rect 1516 -2620 1522 -2568
rect 1522 -2620 1588 -2568
rect 1588 -2620 1592 -2568
rect 1516 -2624 1592 -2620
rect 1486 -3082 1586 -3054
rect 1486 -3142 1498 -3082
rect 1498 -3142 1578 -3082
rect 1578 -3142 1586 -3082
rect 1486 -3146 1586 -3142
rect 4660 -2568 4736 -2566
rect 4660 -2620 4666 -2568
rect 4666 -2620 4732 -2568
rect 4732 -2620 4736 -2568
rect 7792 -2564 7868 -2562
rect 4660 -2624 4736 -2620
rect 7792 -2616 7798 -2564
rect 7798 -2616 7864 -2564
rect 7864 -2616 7868 -2564
rect 7792 -2620 7868 -2616
rect 10936 -2564 11012 -2562
rect 10936 -2616 10942 -2564
rect 10942 -2616 11008 -2564
rect 11008 -2616 11012 -2564
rect 10936 -2620 11012 -2616
rect 14138 -2568 14214 -2566
rect 14138 -2620 14144 -2568
rect 14144 -2620 14210 -2568
rect 14210 -2620 14214 -2568
rect 14138 -2624 14214 -2620
rect 17282 -2568 17358 -2566
rect 17282 -2620 17288 -2568
rect 17288 -2620 17354 -2568
rect 17354 -2620 17358 -2568
rect 17282 -2624 17358 -2620
rect 20414 -2564 20490 -2562
rect 20414 -2616 20420 -2564
rect 20420 -2616 20486 -2564
rect 20486 -2616 20490 -2564
rect 20414 -2620 20490 -2616
rect 23558 -2564 23634 -2562
rect 23558 -2616 23564 -2564
rect 23564 -2616 23630 -2564
rect 23630 -2616 23634 -2564
rect 23558 -2620 23634 -2616
rect 4630 -3082 4730 -3054
rect 4630 -3142 4642 -3082
rect 4642 -3142 4722 -3082
rect 4722 -3142 4730 -3082
rect 4630 -3146 4730 -3142
rect 7762 -3078 7862 -3050
rect 7762 -3138 7774 -3078
rect 7774 -3138 7854 -3078
rect 7854 -3138 7862 -3078
rect 7762 -3142 7862 -3138
rect 10906 -3078 11006 -3050
rect 10906 -3138 10918 -3078
rect 10918 -3138 10998 -3078
rect 10998 -3138 11006 -3078
rect 10906 -3142 11006 -3138
rect 14108 -3082 14208 -3054
rect 14108 -3142 14120 -3082
rect 14120 -3142 14200 -3082
rect 14200 -3142 14208 -3082
rect 14108 -3146 14208 -3142
rect 17252 -3082 17352 -3054
rect 17252 -3142 17264 -3082
rect 17264 -3142 17344 -3082
rect 17344 -3142 17352 -3082
rect 17252 -3146 17352 -3142
rect 20384 -3078 20484 -3050
rect 20384 -3138 20396 -3078
rect 20396 -3138 20476 -3078
rect 20476 -3138 20484 -3078
rect 20384 -3142 20484 -3138
rect 23528 -3078 23628 -3050
rect 23528 -3138 23540 -3078
rect 23540 -3138 23620 -3078
rect 23620 -3138 23628 -3078
rect 23528 -3142 23628 -3138
rect 1506 -5300 1582 -5298
rect 1506 -5352 1512 -5300
rect 1512 -5352 1578 -5300
rect 1578 -5352 1582 -5300
rect 1506 -5356 1582 -5352
rect 4650 -5300 4726 -5298
rect 4650 -5352 4656 -5300
rect 4656 -5352 4722 -5300
rect 4722 -5352 4726 -5300
rect 4650 -5356 4726 -5352
rect 7782 -5296 7858 -5294
rect 7782 -5348 7788 -5296
rect 7788 -5348 7854 -5296
rect 7854 -5348 7858 -5296
rect 7782 -5352 7858 -5348
rect 10926 -5296 11002 -5294
rect 10926 -5348 10932 -5296
rect 10932 -5348 10998 -5296
rect 10998 -5348 11002 -5296
rect 10926 -5352 11002 -5348
rect 14128 -5300 14204 -5298
rect 14128 -5352 14134 -5300
rect 14134 -5352 14200 -5300
rect 14200 -5352 14204 -5300
rect 14128 -5356 14204 -5352
rect 17272 -5300 17348 -5298
rect 17272 -5352 17278 -5300
rect 17278 -5352 17344 -5300
rect 17344 -5352 17348 -5300
rect 17272 -5356 17348 -5352
rect 20404 -5296 20480 -5294
rect 20404 -5348 20410 -5296
rect 20410 -5348 20476 -5296
rect 20476 -5348 20480 -5296
rect 20404 -5352 20480 -5348
rect 23548 -5296 23624 -5294
rect 23548 -5348 23554 -5296
rect 23554 -5348 23620 -5296
rect 23620 -5348 23624 -5296
rect 23548 -5352 23624 -5348
rect 16869 -5961 16963 -5951
rect 802 -6020 880 -6012
rect 802 -6074 814 -6020
rect 814 -6074 868 -6020
rect 868 -6074 880 -6020
rect 802 -6082 880 -6074
rect 2870 -6018 2948 -6010
rect 2870 -6072 2882 -6018
rect 2882 -6072 2936 -6018
rect 2936 -6072 2948 -6018
rect 2870 -6080 2948 -6072
rect 4939 -6020 5017 -6012
rect 4939 -6074 4951 -6020
rect 4951 -6074 5005 -6020
rect 5005 -6074 5017 -6020
rect 4939 -6082 5017 -6074
rect 7007 -6018 7085 -6010
rect 7007 -6072 7019 -6018
rect 7019 -6072 7073 -6018
rect 7073 -6072 7085 -6018
rect 7007 -6080 7085 -6072
rect 9076 -6018 9154 -6010
rect 9076 -6072 9088 -6018
rect 9088 -6072 9142 -6018
rect 9142 -6072 9154 -6018
rect 9076 -6080 9154 -6072
rect 11144 -6016 11222 -6008
rect 11144 -6070 11156 -6016
rect 11156 -6070 11210 -6016
rect 11210 -6070 11222 -6016
rect 11144 -6078 11222 -6070
rect 13213 -6018 13291 -6010
rect 13213 -6072 13225 -6018
rect 13225 -6072 13279 -6018
rect 13279 -6072 13291 -6018
rect 13213 -6080 13291 -6072
rect 15281 -6016 15359 -6008
rect 15281 -6070 15293 -6016
rect 15293 -6070 15347 -6016
rect 15347 -6070 15359 -6016
rect 16869 -6035 16877 -5961
rect 16877 -6035 16953 -5961
rect 16953 -6035 16963 -5961
rect 17607 -5963 17701 -5953
rect 17607 -6037 17615 -5963
rect 17615 -6037 17691 -5963
rect 17691 -6037 17701 -5963
rect 18345 -5963 18439 -5953
rect 18345 -6037 18353 -5963
rect 18353 -6037 18429 -5963
rect 18429 -6037 18439 -5963
rect 19087 -5963 19181 -5953
rect 19087 -6037 19095 -5963
rect 19095 -6037 19171 -5963
rect 19171 -6037 19181 -5963
rect 19827 -5963 19921 -5953
rect 19827 -6037 19835 -5963
rect 19835 -6037 19911 -5963
rect 19911 -6037 19921 -5963
rect 20565 -5963 20659 -5953
rect 20565 -6037 20573 -5963
rect 20573 -6037 20649 -5963
rect 20649 -6037 20659 -5963
rect 21303 -5963 21397 -5953
rect 21303 -6037 21311 -5963
rect 21311 -6037 21387 -5963
rect 21387 -6037 21397 -5963
rect 22041 -5963 22135 -5953
rect 22041 -6037 22049 -5963
rect 22049 -6037 22125 -5963
rect 22125 -6037 22135 -5963
rect 15281 -6078 15359 -6070
rect 2069 -6820 2144 -6804
rect -282 -6829 -216 -6828
rect -282 -6882 -280 -6829
rect -280 -6882 -220 -6829
rect -220 -6882 -216 -6829
rect -282 -6885 -216 -6882
rect 2069 -6886 2074 -6820
rect 2074 -6886 2140 -6820
rect 2140 -6886 2144 -6820
rect 8280 -6820 8347 -6818
rect 2069 -6890 2144 -6886
rect 4140 -6888 4143 -6822
rect 4143 -6888 4209 -6822
rect 6212 -6886 6276 -6821
rect 8280 -6886 8346 -6820
rect 8346 -6886 8347 -6820
rect 10343 -6884 10348 -6818
rect 10348 -6884 10408 -6818
rect 14478 -6818 14561 -6809
rect 10343 -6886 10408 -6884
rect 12414 -6885 12417 -6821
rect 12417 -6885 12481 -6821
rect 14478 -6884 14485 -6818
rect 14485 -6884 14551 -6818
rect 14551 -6884 14561 -6818
rect 8280 -6887 8347 -6886
rect 14478 -6889 14561 -6884
rect 16817 -6907 16883 -6849
rect 17555 -6909 17621 -6851
rect 18293 -6909 18359 -6851
rect 19035 -6909 19101 -6851
rect 19775 -6909 19841 -6851
rect 20513 -6909 20579 -6851
rect 21251 -6909 21317 -6851
rect 21989 -6909 22055 -6851
rect -9 -7087 62 -7010
rect 750 -8244 822 -8242
rect 750 -8302 756 -8244
rect 756 -8302 818 -8244
rect 818 -8302 822 -8244
rect 750 -8312 822 -8302
rect 2818 -8242 2890 -8240
rect 2818 -8300 2824 -8242
rect 2824 -8300 2886 -8242
rect 2886 -8300 2890 -8242
rect 2818 -8310 2890 -8300
rect 4887 -8244 4959 -8242
rect 4887 -8302 4893 -8244
rect 4893 -8302 4955 -8244
rect 4955 -8302 4959 -8244
rect 4887 -8312 4959 -8302
rect 6955 -8242 7027 -8240
rect 6955 -8300 6961 -8242
rect 6961 -8300 7023 -8242
rect 7023 -8300 7027 -8242
rect 6955 -8310 7027 -8300
rect 9024 -8242 9096 -8240
rect 9024 -8300 9030 -8242
rect 9030 -8300 9092 -8242
rect 9092 -8300 9096 -8242
rect 9024 -8310 9096 -8300
rect 11092 -8240 11164 -8238
rect 11092 -8298 11098 -8240
rect 11098 -8298 11160 -8240
rect 11160 -8298 11164 -8240
rect 11092 -8308 11164 -8298
rect 13161 -8242 13233 -8240
rect 13161 -8300 13167 -8242
rect 13167 -8300 13229 -8242
rect 13229 -8300 13233 -8242
rect 13161 -8310 13233 -8300
rect 15229 -8240 15301 -8238
rect 15229 -8298 15235 -8240
rect 15235 -8298 15297 -8240
rect 15297 -8298 15301 -8240
rect 15229 -8308 15301 -8298
<< metal3 >>
rect 12486 4226 12496 4346
rect 12618 4226 12628 4346
rect 13654 4332 13796 4346
rect 13654 4241 13682 4332
rect 13772 4241 13796 4332
rect 13654 4226 13796 4241
rect 14822 4332 14964 4346
rect 14822 4241 14850 4332
rect 14940 4241 14964 4332
rect 14822 4226 14964 4241
rect 15990 4332 16132 4346
rect 15990 4241 16018 4332
rect 16108 4241 16132 4332
rect 15990 4226 16132 4241
rect 17164 4334 17306 4348
rect 17164 4243 17192 4334
rect 17282 4243 17306 4334
rect 17164 4228 17306 4243
rect 18332 4334 18474 4348
rect 18332 4243 18360 4334
rect 18450 4243 18474 4334
rect 18332 4228 18474 4243
rect 19500 4334 19642 4348
rect 19500 4243 19528 4334
rect 19618 4243 19642 4334
rect 19500 4228 19642 4243
rect 20668 4334 20810 4348
rect 20668 4243 20696 4334
rect 20786 4243 20810 4334
rect 20668 4228 20810 4243
rect 526 4127 624 4145
rect 526 4055 536 4127
rect 606 4055 624 4127
rect 526 4047 624 4055
rect 1974 4127 2072 4145
rect 1974 4055 1984 4127
rect 2054 4055 2072 4127
rect 1974 4047 2072 4055
rect 3472 4129 3570 4147
rect 3472 4057 3482 4129
rect 3552 4057 3570 4129
rect 3472 4049 3570 4057
rect 4920 4129 5018 4147
rect 4920 4057 4930 4129
rect 5000 4057 5018 4129
rect 4920 4049 5018 4057
rect 6440 4127 6538 4145
rect 6440 4055 6450 4127
rect 6520 4055 6538 4127
rect 6440 4047 6538 4055
rect 7888 4127 7986 4145
rect 7888 4055 7898 4127
rect 7968 4055 7986 4127
rect 7888 4047 7986 4055
rect 9386 4129 9484 4147
rect 9386 4057 9396 4129
rect 9466 4057 9484 4129
rect 9386 4049 9484 4057
rect 10834 4129 10932 4147
rect 10834 4057 10844 4129
rect 10914 4057 10932 4129
rect 10834 4049 10932 4057
rect -293 3472 -221 3477
rect -303 3467 -212 3472
rect -303 3408 -293 3467
rect -222 3408 -212 3467
rect -303 3403 -212 3408
rect -2537 2795 -2459 2797
rect -293 2795 -221 3403
rect -17 3371 72 3376
rect -17 3307 -7 3371
rect 62 3307 72 3371
rect -17 3302 72 3307
rect -2537 2792 -221 2795
rect -2537 2736 -2527 2792
rect -2469 2736 -221 2792
rect -2537 2733 -221 2736
rect -2537 2731 -2459 2733
rect -293 -6823 -221 2733
rect -293 -6828 -206 -6823
rect -293 -6885 -282 -6828
rect -216 -6885 -206 -6828
rect -293 -6890 -206 -6885
rect -293 -6899 -221 -6890
rect -9 -6965 63 3302
rect 1630 3185 2116 3197
rect 9049 3189 9910 3191
rect 1630 3098 1640 3185
rect 1716 3098 2116 3185
rect 1630 3092 2116 3098
rect 3129 3177 4194 3188
rect 3129 3103 3142 3177
rect 3206 3103 4194 3177
rect 3129 3097 4194 3103
rect 744 2923 846 2939
rect 744 2855 758 2923
rect 832 2855 846 2923
rect 744 2841 846 2855
rect 1486 2412 1606 2417
rect 1486 2318 1496 2412
rect 1596 2318 1606 2412
rect 1486 2315 1606 2318
rect 1476 168 1642 176
rect 1476 100 1510 168
rect 1594 100 1642 168
rect 1476 96 1642 100
rect 1486 -322 1606 -317
rect 1486 -416 1496 -322
rect 1596 -416 1606 -322
rect 1486 -419 1606 -416
rect 1476 -2566 1642 -2558
rect 1476 -2634 1510 -2566
rect 1594 -2634 1642 -2566
rect 1476 -2638 1642 -2634
rect 1476 -3054 1596 -3049
rect 1476 -3148 1486 -3054
rect 1586 -3148 1596 -3054
rect 1476 -3151 1596 -3148
rect 1466 -5298 1632 -5290
rect 1466 -5366 1500 -5298
rect 1584 -5366 1632 -5298
rect 1466 -5370 1632 -5366
rect 732 -6010 946 -6006
rect 732 -6082 802 -6010
rect 878 -6012 946 -6010
rect 880 -6082 946 -6012
rect 732 -6084 946 -6082
rect 792 -6087 890 -6084
rect 2051 -6799 2116 3092
rect 2192 2923 2294 2939
rect 2192 2855 2206 2923
rect 2280 2855 2294 2923
rect 2192 2841 2294 2855
rect 3690 2925 3792 2941
rect 3690 2857 3704 2925
rect 3778 2857 3792 2925
rect 3690 2843 3792 2857
rect 2800 -6008 3014 -6004
rect 2800 -6080 2870 -6008
rect 2946 -6010 3014 -6008
rect 2948 -6080 3014 -6010
rect 2800 -6082 3014 -6080
rect 2860 -6085 2958 -6082
rect 2051 -6804 2154 -6799
rect 2051 -6890 2069 -6804
rect 2144 -6890 2154 -6804
rect 2051 -6895 2154 -6890
rect 4130 -6817 4194 3097
rect 4581 3183 4668 3188
rect 6350 3186 6416 3187
rect 4581 3105 4591 3183
rect 4658 3105 4668 3183
rect 4581 2968 4668 3105
rect 6100 3181 6416 3186
rect 6100 3106 6110 3181
rect 6170 3106 6416 3181
rect 9049 3183 9965 3189
rect 7627 3179 8645 3180
rect 6100 3102 6416 3106
rect 6100 3101 6180 3102
rect 4582 2767 4668 2968
rect 5138 2925 5240 2941
rect 5138 2857 5152 2925
rect 5226 2857 5240 2925
rect 5138 2843 5240 2857
rect 4582 2695 6268 2767
rect 4630 2412 4750 2417
rect 4630 2318 4640 2412
rect 4740 2318 4750 2412
rect 4630 2315 4750 2318
rect 4620 168 4786 176
rect 4620 100 4654 168
rect 4738 100 4786 168
rect 4620 96 4786 100
rect 4630 -322 4750 -317
rect 4630 -416 4640 -322
rect 4740 -416 4750 -322
rect 4630 -419 4750 -416
rect 4620 -2566 4786 -2558
rect 4620 -2634 4654 -2566
rect 4738 -2634 4786 -2566
rect 4620 -2638 4786 -2634
rect 4620 -3054 4740 -3049
rect 4620 -3148 4630 -3054
rect 4730 -3148 4740 -3054
rect 4620 -3151 4740 -3148
rect 4610 -5298 4776 -5290
rect 4610 -5366 4644 -5298
rect 4728 -5366 4776 -5298
rect 4610 -5370 4776 -5366
rect 4869 -6010 5083 -6006
rect 4869 -6082 4939 -6010
rect 5015 -6012 5083 -6010
rect 5017 -6082 5083 -6012
rect 4869 -6084 5083 -6082
rect 4929 -6087 5027 -6084
rect 6201 -6816 6268 2695
rect 6350 2737 6416 3102
rect 7550 3174 8645 3179
rect 7550 3106 7560 3174
rect 7620 3106 8645 3174
rect 7550 3102 8645 3106
rect 7550 3101 7630 3102
rect 6658 2923 6760 2939
rect 6658 2855 6672 2923
rect 6746 2855 6760 2923
rect 6658 2841 6760 2855
rect 8106 2923 8208 2939
rect 8106 2855 8120 2923
rect 8194 2855 8208 2923
rect 8106 2841 8208 2855
rect 8563 2746 8645 3102
rect 9049 3104 9059 3183
rect 9120 3104 9965 3183
rect 9049 3099 9965 3104
rect 9902 2953 9965 3099
rect 10483 3188 10588 3193
rect 10483 3098 10493 3188
rect 10578 3180 10588 3188
rect 13851 3180 13936 3181
rect 10578 3103 13936 3180
rect 10578 3098 10588 3103
rect 10483 3093 10588 3098
rect 10398 2953 10834 2954
rect 9604 2925 9706 2941
rect 9604 2857 9618 2925
rect 9692 2857 9706 2925
rect 9902 2868 10834 2953
rect 9604 2843 9706 2857
rect 10773 2762 10834 2868
rect 11052 2925 11154 2941
rect 11052 2857 11066 2925
rect 11140 2857 11154 2925
rect 12029 2904 12039 3015
rect 12149 2904 12159 3015
rect 13197 2904 13207 3015
rect 13317 2904 13327 3015
rect 11052 2843 11154 2857
rect 10332 2746 10398 2748
rect 8271 2737 8345 2738
rect 6350 2662 8345 2737
rect 6350 2661 6416 2662
rect 7762 2416 7882 2421
rect 7762 2322 7772 2416
rect 7872 2322 7882 2416
rect 7762 2319 7882 2322
rect 7752 172 7918 180
rect 7752 104 7786 172
rect 7870 104 7918 172
rect 7752 100 7918 104
rect 7762 -318 7882 -313
rect 7762 -412 7772 -318
rect 7872 -412 7882 -318
rect 7762 -415 7882 -412
rect 7752 -2562 7918 -2554
rect 7752 -2630 7786 -2562
rect 7870 -2630 7918 -2562
rect 7752 -2634 7918 -2630
rect 7752 -3050 7872 -3045
rect 7752 -3144 7762 -3050
rect 7862 -3144 7872 -3050
rect 7752 -3147 7872 -3144
rect 7742 -5294 7908 -5286
rect 7742 -5362 7776 -5294
rect 7860 -5362 7908 -5294
rect 7742 -5366 7908 -5362
rect 6937 -6008 7151 -6004
rect 6937 -6080 7007 -6008
rect 7083 -6010 7151 -6008
rect 7085 -6080 7151 -6010
rect 6937 -6082 7151 -6080
rect 6997 -6085 7095 -6082
rect 8271 -6813 8345 2662
rect 8563 2657 10402 2746
rect 10773 2702 12084 2762
rect 8563 2655 8645 2657
rect 9006 -6008 9220 -6004
rect 9006 -6080 9076 -6008
rect 9152 -6010 9220 -6008
rect 9154 -6080 9220 -6010
rect 9006 -6082 9220 -6080
rect 9066 -6085 9164 -6082
rect 10332 -6813 10398 2657
rect 10906 2416 11026 2421
rect 10906 2322 10916 2416
rect 11016 2322 11026 2416
rect 10906 2319 11026 2322
rect 10896 172 11062 180
rect 10896 104 10930 172
rect 11014 104 11062 172
rect 10896 100 11062 104
rect 10906 -318 11026 -313
rect 10906 -412 10916 -318
rect 11016 -412 11026 -318
rect 10906 -415 11026 -412
rect 10896 -2562 11062 -2554
rect 10896 -2630 10930 -2562
rect 11014 -2630 11062 -2562
rect 10896 -2634 11062 -2630
rect 10896 -3050 11016 -3045
rect 10896 -3144 10906 -3050
rect 11006 -3144 11016 -3050
rect 10896 -3147 11016 -3144
rect 10886 -5294 11052 -5286
rect 10886 -5362 10920 -5294
rect 11004 -5362 11052 -5294
rect 10886 -5366 11052 -5362
rect 11074 -6006 11288 -6002
rect 11074 -6078 11144 -6006
rect 11220 -6008 11288 -6006
rect 11222 -6078 11288 -6008
rect 11074 -6080 11288 -6078
rect 11134 -6083 11232 -6080
rect 4130 -6822 4219 -6817
rect 4130 -6888 4140 -6822
rect 4209 -6888 4219 -6822
rect 4130 -6893 4219 -6888
rect 6201 -6821 6286 -6816
rect 6201 -6886 6212 -6821
rect 6276 -6886 6286 -6821
rect 6201 -6891 6286 -6886
rect 8270 -6818 8357 -6813
rect 8270 -6887 8280 -6818
rect 8347 -6887 8357 -6818
rect 2051 -6909 2116 -6895
rect 4130 -6900 4194 -6893
rect 6201 -6899 6268 -6891
rect 8270 -6892 8357 -6887
rect 10332 -6818 10418 -6813
rect 10332 -6886 10343 -6818
rect 10408 -6886 10418 -6818
rect 10332 -6891 10418 -6886
rect 12019 -6815 12084 2702
rect 13851 2671 13936 3103
rect 14365 2904 14375 3015
rect 14485 2904 14495 3015
rect 15533 2904 15543 3015
rect 15653 2904 15663 3015
rect 16707 2906 16717 3017
rect 16827 2906 16837 3017
rect 17875 2906 17885 3017
rect 17995 2906 18005 3017
rect 19043 2906 19053 3017
rect 19163 2906 19173 3017
rect 20211 2906 20221 3017
rect 20331 2906 20341 3017
rect 13851 2666 14440 2671
rect 13852 2601 14440 2666
rect 14108 2412 14228 2417
rect 14108 2318 14118 2412
rect 14218 2318 14228 2412
rect 14108 2315 14228 2318
rect 14098 168 14264 176
rect 14098 100 14132 168
rect 14216 100 14264 168
rect 14098 96 14264 100
rect 14108 -322 14228 -317
rect 14108 -416 14118 -322
rect 14218 -416 14228 -322
rect 14108 -419 14228 -416
rect 14098 -2566 14264 -2558
rect 14098 -2634 14132 -2566
rect 14216 -2634 14264 -2566
rect 14098 -2638 14264 -2634
rect 14098 -3054 14218 -3049
rect 14098 -3148 14108 -3054
rect 14208 -3148 14218 -3054
rect 14098 -3151 14218 -3148
rect 14088 -5298 14254 -5290
rect 14088 -5366 14122 -5298
rect 14206 -5366 14254 -5298
rect 14088 -5370 14254 -5366
rect 13143 -6008 13357 -6004
rect 13143 -6080 13213 -6008
rect 13289 -6010 13357 -6008
rect 13291 -6080 13357 -6010
rect 13143 -6082 13357 -6080
rect 13203 -6085 13301 -6082
rect 14367 -6804 14438 2601
rect 17252 2412 17372 2417
rect 17252 2318 17262 2412
rect 17362 2318 17372 2412
rect 20384 2416 20504 2421
rect 20384 2322 20394 2416
rect 20494 2322 20504 2416
rect 20384 2319 20504 2322
rect 23528 2416 23648 2421
rect 23528 2322 23538 2416
rect 23638 2322 23648 2416
rect 23528 2319 23648 2322
rect 17252 2315 17372 2318
rect 17242 168 17408 176
rect 17242 100 17276 168
rect 17360 100 17408 168
rect 20374 172 20540 180
rect 20374 104 20408 172
rect 20492 104 20540 172
rect 20374 100 20540 104
rect 23518 172 23684 180
rect 23518 104 23552 172
rect 23636 104 23684 172
rect 23518 100 23684 104
rect 17242 96 17408 100
rect 17252 -322 17372 -317
rect 17252 -416 17262 -322
rect 17362 -416 17372 -322
rect 20384 -318 20504 -313
rect 20384 -412 20394 -318
rect 20494 -412 20504 -318
rect 20384 -415 20504 -412
rect 23528 -318 23648 -313
rect 23528 -412 23538 -318
rect 23638 -412 23648 -318
rect 23528 -415 23648 -412
rect 17252 -419 17372 -416
rect 17242 -2566 17408 -2558
rect 17242 -2634 17276 -2566
rect 17360 -2634 17408 -2566
rect 20374 -2562 20540 -2554
rect 20374 -2630 20408 -2562
rect 20492 -2630 20540 -2562
rect 20374 -2634 20540 -2630
rect 23518 -2562 23684 -2554
rect 23518 -2630 23552 -2562
rect 23636 -2630 23684 -2562
rect 23518 -2634 23684 -2630
rect 17242 -2638 17408 -2634
rect 17242 -3054 17362 -3049
rect 17242 -3148 17252 -3054
rect 17352 -3148 17362 -3054
rect 20374 -3050 20494 -3045
rect 20374 -3144 20384 -3050
rect 20484 -3144 20494 -3050
rect 20374 -3147 20494 -3144
rect 23518 -3050 23638 -3045
rect 23518 -3144 23528 -3050
rect 23628 -3144 23638 -3050
rect 23518 -3147 23638 -3144
rect 17242 -3151 17362 -3148
rect 17232 -5298 17398 -5290
rect 17232 -5366 17266 -5298
rect 17350 -5366 17398 -5298
rect 20364 -5294 20530 -5286
rect 20364 -5362 20398 -5294
rect 20482 -5362 20530 -5294
rect 20364 -5366 20530 -5362
rect 23508 -5294 23674 -5286
rect 23508 -5362 23542 -5294
rect 23626 -5362 23674 -5294
rect 23508 -5366 23674 -5362
rect 17232 -5370 17398 -5366
rect 16713 -5937 17107 -5931
rect 15211 -6006 15425 -6002
rect 15211 -6078 15281 -6006
rect 15357 -6008 15425 -6006
rect 15359 -6078 15425 -6008
rect 15211 -6080 15425 -6078
rect 16713 -6045 16861 -5937
rect 16971 -6045 17107 -5937
rect 15271 -6083 15369 -6080
rect 16713 -6081 17107 -6045
rect 17451 -5939 17845 -5933
rect 17451 -6047 17599 -5939
rect 17709 -6047 17845 -5939
rect 17451 -6083 17845 -6047
rect 18189 -5939 18583 -5933
rect 18189 -6047 18337 -5939
rect 18447 -6047 18583 -5939
rect 18189 -6083 18583 -6047
rect 18931 -5939 19325 -5933
rect 18931 -6047 19079 -5939
rect 19189 -6047 19325 -5939
rect 18931 -6083 19325 -6047
rect 19671 -5939 20065 -5933
rect 19671 -6047 19819 -5939
rect 19929 -6047 20065 -5939
rect 19671 -6083 20065 -6047
rect 20409 -5939 20803 -5933
rect 20409 -6047 20557 -5939
rect 20667 -6047 20803 -5939
rect 20409 -6083 20803 -6047
rect 21147 -5939 21541 -5933
rect 21147 -6047 21295 -5939
rect 21405 -6047 21541 -5939
rect 21147 -6083 21541 -6047
rect 21885 -5939 22279 -5933
rect 21885 -6047 22033 -5939
rect 22143 -6047 22279 -5939
rect 21885 -6083 22279 -6047
rect 14367 -6809 14571 -6804
rect 12019 -6816 12439 -6815
rect 12019 -6821 12491 -6816
rect 12019 -6885 12414 -6821
rect 12481 -6885 12491 -6821
rect 12019 -6889 12491 -6885
rect 12019 -6890 12084 -6889
rect 12304 -6890 12491 -6889
rect 14367 -6889 14478 -6809
rect 14561 -6889 14571 -6809
rect 16771 -6829 16931 -6827
rect 16771 -6839 16801 -6829
rect 8271 -6904 8345 -6892
rect 10332 -6900 10398 -6891
rect 14367 -6902 14571 -6889
rect 16769 -6921 16801 -6839
rect 16771 -6929 16801 -6921
rect 16903 -6929 16931 -6829
rect 17509 -6831 17669 -6829
rect 17509 -6841 17539 -6831
rect 17507 -6923 17539 -6841
rect 16771 -6935 16931 -6929
rect 17509 -6931 17539 -6923
rect 17641 -6931 17669 -6831
rect 18247 -6831 18407 -6829
rect 18247 -6841 18277 -6831
rect 18245 -6923 18277 -6841
rect 17509 -6937 17669 -6931
rect 18247 -6931 18277 -6923
rect 18379 -6931 18407 -6831
rect 18989 -6831 19149 -6829
rect 18989 -6841 19019 -6831
rect 18987 -6923 19019 -6841
rect 18247 -6937 18407 -6931
rect 18989 -6931 19019 -6923
rect 19121 -6931 19149 -6831
rect 19729 -6831 19889 -6829
rect 19729 -6841 19759 -6831
rect 19727 -6923 19759 -6841
rect 18989 -6937 19149 -6931
rect 19729 -6931 19759 -6923
rect 19861 -6931 19889 -6831
rect 20467 -6831 20627 -6829
rect 20467 -6841 20497 -6831
rect 20465 -6923 20497 -6841
rect 19729 -6937 19889 -6931
rect 20467 -6931 20497 -6923
rect 20599 -6931 20627 -6831
rect 21205 -6831 21365 -6829
rect 21205 -6841 21235 -6831
rect 21203 -6923 21235 -6841
rect 20467 -6937 20627 -6931
rect 21205 -6931 21235 -6923
rect 21337 -6931 21365 -6831
rect 21943 -6831 22103 -6829
rect 21943 -6841 21973 -6831
rect 21941 -6923 21973 -6841
rect 21205 -6937 21365 -6931
rect 21943 -6931 21973 -6923
rect 22075 -6931 22103 -6831
rect 21943 -6937 22103 -6931
rect -29 -7010 81 -6965
rect -29 -7087 -9 -7010
rect 62 -7087 81 -7010
rect -29 -7107 81 -7087
rect 11054 -8224 11206 -8222
rect 15191 -8224 15343 -8222
rect 2780 -8226 2932 -8224
rect 6917 -8226 7069 -8224
rect 8986 -8226 9138 -8224
rect 712 -8228 864 -8226
rect 710 -8232 864 -8228
rect 710 -8320 740 -8232
rect 834 -8320 864 -8232
rect 710 -8326 864 -8320
rect 2778 -8230 2932 -8226
rect 4849 -8228 5001 -8226
rect 2778 -8318 2808 -8230
rect 2902 -8318 2932 -8230
rect 2778 -8324 2932 -8318
rect 712 -8336 864 -8326
rect 2780 -8334 2932 -8324
rect 4847 -8232 5001 -8228
rect 4847 -8320 4877 -8232
rect 4971 -8320 5001 -8232
rect 4847 -8326 5001 -8320
rect 6915 -8230 7069 -8226
rect 6915 -8318 6945 -8230
rect 7039 -8318 7069 -8230
rect 6915 -8324 7069 -8318
rect 8984 -8230 9138 -8226
rect 8984 -8318 9014 -8230
rect 9108 -8318 9138 -8230
rect 8984 -8324 9138 -8318
rect 11052 -8228 11206 -8224
rect 13123 -8226 13275 -8224
rect 11052 -8316 11082 -8228
rect 11176 -8316 11206 -8228
rect 11052 -8322 11206 -8316
rect 4849 -8336 5001 -8326
rect 6917 -8334 7069 -8324
rect 8986 -8334 9138 -8324
rect 11054 -8332 11206 -8322
rect 13121 -8230 13275 -8226
rect 13121 -8318 13151 -8230
rect 13245 -8318 13275 -8230
rect 13121 -8324 13275 -8318
rect 15189 -8228 15343 -8224
rect 15189 -8316 15219 -8228
rect 15313 -8316 15343 -8228
rect 15189 -8322 15343 -8316
rect 13123 -8334 13275 -8324
rect 15191 -8332 15343 -8322
<< via3 >>
rect 12496 4332 12618 4346
rect 12496 4241 12514 4332
rect 12514 4241 12604 4332
rect 12604 4241 12618 4332
rect 12496 4226 12618 4241
rect 13698 4254 13762 4318
rect 14866 4254 14930 4318
rect 16036 4256 16100 4320
rect 17208 4256 17272 4320
rect 18376 4254 18440 4318
rect 19544 4256 19608 4320
rect 20712 4256 20776 4320
rect 536 4123 606 4127
rect 536 4061 542 4123
rect 542 4061 602 4123
rect 602 4061 606 4123
rect 536 4055 606 4061
rect 1984 4123 2054 4127
rect 1984 4061 1990 4123
rect 1990 4061 2050 4123
rect 2050 4061 2054 4123
rect 1984 4055 2054 4061
rect 3482 4125 3552 4129
rect 3482 4063 3488 4125
rect 3488 4063 3548 4125
rect 3548 4063 3552 4125
rect 3482 4057 3552 4063
rect 4930 4125 5000 4129
rect 4930 4063 4936 4125
rect 4936 4063 4996 4125
rect 4996 4063 5000 4125
rect 4930 4057 5000 4063
rect 6450 4123 6520 4127
rect 6450 4061 6456 4123
rect 6456 4061 6516 4123
rect 6516 4061 6520 4123
rect 6450 4055 6520 4061
rect 7898 4123 7968 4127
rect 7898 4061 7904 4123
rect 7904 4061 7964 4123
rect 7964 4061 7968 4123
rect 7898 4055 7968 4061
rect 9396 4125 9466 4129
rect 9396 4063 9402 4125
rect 9402 4063 9462 4125
rect 9462 4063 9466 4125
rect 9396 4057 9466 4063
rect 10844 4125 10914 4129
rect 10844 4063 10850 4125
rect 10850 4063 10910 4125
rect 10910 4063 10914 4125
rect 10844 4057 10914 4063
rect 758 2917 832 2923
rect 758 2855 764 2917
rect 764 2855 828 2917
rect 828 2855 832 2917
rect 1496 2320 1596 2410
rect 1496 2318 1596 2320
rect 1510 110 1516 168
rect 1516 110 1592 168
rect 1592 110 1594 168
rect 1510 100 1594 110
rect 1496 -414 1596 -324
rect 1496 -416 1596 -414
rect 1510 -2624 1516 -2566
rect 1516 -2624 1592 -2566
rect 1592 -2624 1594 -2566
rect 1510 -2634 1594 -2624
rect 1486 -3146 1586 -3056
rect 1486 -3148 1586 -3146
rect 1500 -5356 1506 -5298
rect 1506 -5356 1582 -5298
rect 1582 -5356 1584 -5298
rect 1500 -5366 1584 -5356
rect 802 -6012 878 -6010
rect 802 -6076 878 -6012
rect 2206 2917 2280 2923
rect 2206 2855 2212 2917
rect 2212 2855 2276 2917
rect 2276 2855 2280 2917
rect 3704 2919 3778 2925
rect 3704 2857 3710 2919
rect 3710 2857 3774 2919
rect 3774 2857 3778 2919
rect 2870 -6010 2946 -6008
rect 2870 -6074 2946 -6010
rect 5152 2919 5226 2925
rect 5152 2857 5158 2919
rect 5158 2857 5222 2919
rect 5222 2857 5226 2919
rect 4640 2320 4740 2410
rect 4640 2318 4740 2320
rect 4654 110 4660 168
rect 4660 110 4736 168
rect 4736 110 4738 168
rect 4654 100 4738 110
rect 4640 -414 4740 -324
rect 4640 -416 4740 -414
rect 4654 -2624 4660 -2566
rect 4660 -2624 4736 -2566
rect 4736 -2624 4738 -2566
rect 4654 -2634 4738 -2624
rect 4630 -3146 4730 -3056
rect 4630 -3148 4730 -3146
rect 4644 -5356 4650 -5298
rect 4650 -5356 4726 -5298
rect 4726 -5356 4728 -5298
rect 4644 -5366 4728 -5356
rect 4939 -6012 5015 -6010
rect 4939 -6076 5015 -6012
rect 6672 2917 6746 2923
rect 6672 2855 6678 2917
rect 6678 2855 6742 2917
rect 6742 2855 6746 2917
rect 8120 2917 8194 2923
rect 8120 2855 8126 2917
rect 8126 2855 8190 2917
rect 8190 2855 8194 2917
rect 9618 2919 9692 2925
rect 9618 2857 9624 2919
rect 9624 2857 9688 2919
rect 9688 2857 9692 2919
rect 11066 2919 11140 2925
rect 11066 2857 11072 2919
rect 11072 2857 11136 2919
rect 11136 2857 11140 2919
rect 12039 3005 12149 3015
rect 12039 2914 12049 3005
rect 12049 2914 12139 3005
rect 12139 2914 12149 3005
rect 12039 2904 12149 2914
rect 13207 3005 13317 3015
rect 13207 2914 13217 3005
rect 13217 2914 13307 3005
rect 13307 2914 13317 3005
rect 13207 2904 13317 2914
rect 7772 2324 7872 2414
rect 7772 2322 7872 2324
rect 7786 114 7792 172
rect 7792 114 7868 172
rect 7868 114 7870 172
rect 7786 104 7870 114
rect 7772 -410 7872 -320
rect 7772 -412 7872 -410
rect 7786 -2620 7792 -2562
rect 7792 -2620 7868 -2562
rect 7868 -2620 7870 -2562
rect 7786 -2630 7870 -2620
rect 7762 -3142 7862 -3052
rect 7762 -3144 7862 -3142
rect 7776 -5352 7782 -5294
rect 7782 -5352 7858 -5294
rect 7858 -5352 7860 -5294
rect 7776 -5362 7860 -5352
rect 7007 -6010 7083 -6008
rect 7007 -6074 7083 -6010
rect 9076 -6010 9152 -6008
rect 9076 -6074 9152 -6010
rect 10916 2324 11016 2414
rect 10916 2322 11016 2324
rect 10930 114 10936 172
rect 10936 114 11012 172
rect 11012 114 11014 172
rect 10930 104 11014 114
rect 10916 -410 11016 -320
rect 10916 -412 11016 -410
rect 10930 -2620 10936 -2562
rect 10936 -2620 11012 -2562
rect 11012 -2620 11014 -2562
rect 10930 -2630 11014 -2620
rect 10906 -3142 11006 -3052
rect 10906 -3144 11006 -3142
rect 10920 -5352 10926 -5294
rect 10926 -5352 11002 -5294
rect 11002 -5352 11004 -5294
rect 10920 -5362 11004 -5352
rect 11144 -6008 11220 -6006
rect 11144 -6072 11220 -6008
rect 14375 3005 14485 3015
rect 14375 2914 14385 3005
rect 14385 2914 14475 3005
rect 14475 2914 14485 3005
rect 14375 2904 14485 2914
rect 15543 3005 15653 3015
rect 15543 2914 15553 3005
rect 15553 2914 15643 3005
rect 15643 2914 15653 3005
rect 15543 2904 15653 2914
rect 16717 3007 16827 3017
rect 16717 2916 16727 3007
rect 16727 2916 16817 3007
rect 16817 2916 16827 3007
rect 16717 2906 16827 2916
rect 17885 3007 17995 3017
rect 17885 2916 17895 3007
rect 17895 2916 17985 3007
rect 17985 2916 17995 3007
rect 17885 2906 17995 2916
rect 19053 3007 19163 3017
rect 19053 2916 19063 3007
rect 19063 2916 19153 3007
rect 19153 2916 19163 3007
rect 19053 2906 19163 2916
rect 20221 3007 20331 3017
rect 20221 2916 20231 3007
rect 20231 2916 20321 3007
rect 20321 2916 20331 3007
rect 20221 2906 20331 2916
rect 14118 2320 14218 2410
rect 14118 2318 14218 2320
rect 14132 110 14138 168
rect 14138 110 14214 168
rect 14214 110 14216 168
rect 14132 100 14216 110
rect 14118 -414 14218 -324
rect 14118 -416 14218 -414
rect 14132 -2624 14138 -2566
rect 14138 -2624 14214 -2566
rect 14214 -2624 14216 -2566
rect 14132 -2634 14216 -2624
rect 14108 -3146 14208 -3056
rect 14108 -3148 14208 -3146
rect 14122 -5356 14128 -5298
rect 14128 -5356 14204 -5298
rect 14204 -5356 14206 -5298
rect 14122 -5366 14206 -5356
rect 13213 -6010 13289 -6008
rect 13213 -6074 13289 -6010
rect 17262 2320 17362 2410
rect 17262 2318 17362 2320
rect 20394 2324 20494 2414
rect 20394 2322 20494 2324
rect 23538 2324 23638 2414
rect 23538 2322 23638 2324
rect 17276 110 17282 168
rect 17282 110 17358 168
rect 17358 110 17360 168
rect 17276 100 17360 110
rect 20408 114 20414 172
rect 20414 114 20490 172
rect 20490 114 20492 172
rect 20408 104 20492 114
rect 23552 114 23558 172
rect 23558 114 23634 172
rect 23634 114 23636 172
rect 23552 104 23636 114
rect 17262 -414 17362 -324
rect 17262 -416 17362 -414
rect 20394 -410 20494 -320
rect 20394 -412 20494 -410
rect 23538 -410 23638 -320
rect 23538 -412 23638 -410
rect 17276 -2624 17282 -2566
rect 17282 -2624 17358 -2566
rect 17358 -2624 17360 -2566
rect 17276 -2634 17360 -2624
rect 20408 -2620 20414 -2562
rect 20414 -2620 20490 -2562
rect 20490 -2620 20492 -2562
rect 20408 -2630 20492 -2620
rect 23552 -2620 23558 -2562
rect 23558 -2620 23634 -2562
rect 23634 -2620 23636 -2562
rect 23552 -2630 23636 -2620
rect 17252 -3146 17352 -3056
rect 17252 -3148 17352 -3146
rect 20384 -3142 20484 -3052
rect 20384 -3144 20484 -3142
rect 23528 -3142 23628 -3052
rect 23528 -3144 23628 -3142
rect 17266 -5356 17272 -5298
rect 17272 -5356 17348 -5298
rect 17348 -5356 17350 -5298
rect 17266 -5366 17350 -5356
rect 20398 -5352 20404 -5294
rect 20404 -5352 20480 -5294
rect 20480 -5352 20482 -5294
rect 20398 -5362 20482 -5352
rect 23542 -5352 23548 -5294
rect 23548 -5352 23624 -5294
rect 23624 -5352 23626 -5294
rect 23542 -5362 23626 -5352
rect 15281 -6008 15357 -6006
rect 15281 -6072 15357 -6008
rect 16861 -5951 16971 -5937
rect 16861 -6035 16869 -5951
rect 16869 -6035 16963 -5951
rect 16963 -6035 16971 -5951
rect 16861 -6045 16971 -6035
rect 17599 -5953 17709 -5939
rect 17599 -6037 17607 -5953
rect 17607 -6037 17701 -5953
rect 17701 -6037 17709 -5953
rect 17599 -6047 17709 -6037
rect 18337 -5953 18447 -5939
rect 18337 -6037 18345 -5953
rect 18345 -6037 18439 -5953
rect 18439 -6037 18447 -5953
rect 18337 -6047 18447 -6037
rect 19079 -5953 19189 -5939
rect 19079 -6037 19087 -5953
rect 19087 -6037 19181 -5953
rect 19181 -6037 19189 -5953
rect 19079 -6047 19189 -6037
rect 19819 -5953 19929 -5939
rect 19819 -6037 19827 -5953
rect 19827 -6037 19921 -5953
rect 19921 -6037 19929 -5953
rect 19819 -6047 19929 -6037
rect 20557 -5953 20667 -5939
rect 20557 -6037 20565 -5953
rect 20565 -6037 20659 -5953
rect 20659 -6037 20667 -5953
rect 20557 -6047 20667 -6037
rect 21295 -5953 21405 -5939
rect 21295 -6037 21303 -5953
rect 21303 -6037 21397 -5953
rect 21397 -6037 21405 -5953
rect 21295 -6047 21405 -6037
rect 22033 -5953 22143 -5939
rect 22033 -6037 22041 -5953
rect 22041 -6037 22135 -5953
rect 22135 -6037 22143 -5953
rect 22033 -6047 22143 -6037
rect 16801 -6849 16903 -6829
rect 16801 -6907 16817 -6849
rect 16817 -6907 16883 -6849
rect 16883 -6907 16903 -6849
rect 16801 -6929 16903 -6907
rect 17539 -6851 17641 -6831
rect 17539 -6909 17555 -6851
rect 17555 -6909 17621 -6851
rect 17621 -6909 17641 -6851
rect 17539 -6931 17641 -6909
rect 18277 -6851 18379 -6831
rect 18277 -6909 18293 -6851
rect 18293 -6909 18359 -6851
rect 18359 -6909 18379 -6851
rect 18277 -6931 18379 -6909
rect 19019 -6851 19121 -6831
rect 19019 -6909 19035 -6851
rect 19035 -6909 19101 -6851
rect 19101 -6909 19121 -6851
rect 19019 -6931 19121 -6909
rect 19759 -6851 19861 -6831
rect 19759 -6909 19775 -6851
rect 19775 -6909 19841 -6851
rect 19841 -6909 19861 -6851
rect 19759 -6931 19861 -6909
rect 20497 -6851 20599 -6831
rect 20497 -6909 20513 -6851
rect 20513 -6909 20579 -6851
rect 20579 -6909 20599 -6851
rect 20497 -6931 20599 -6909
rect 21235 -6851 21337 -6831
rect 21235 -6909 21251 -6851
rect 21251 -6909 21317 -6851
rect 21317 -6909 21337 -6851
rect 21235 -6931 21337 -6909
rect 21973 -6851 22075 -6831
rect 21973 -6909 21989 -6851
rect 21989 -6909 22055 -6851
rect 22055 -6909 22075 -6851
rect 21973 -6931 22075 -6909
rect 740 -8242 834 -8232
rect 740 -8312 750 -8242
rect 750 -8312 822 -8242
rect 822 -8312 834 -8242
rect 740 -8320 834 -8312
rect 2808 -8240 2902 -8230
rect 2808 -8310 2818 -8240
rect 2818 -8310 2890 -8240
rect 2890 -8310 2902 -8240
rect 2808 -8318 2902 -8310
rect 4877 -8242 4971 -8232
rect 4877 -8312 4887 -8242
rect 4887 -8312 4959 -8242
rect 4959 -8312 4971 -8242
rect 4877 -8320 4971 -8312
rect 6945 -8240 7039 -8230
rect 6945 -8310 6955 -8240
rect 6955 -8310 7027 -8240
rect 7027 -8310 7039 -8240
rect 6945 -8318 7039 -8310
rect 9014 -8240 9108 -8230
rect 9014 -8310 9024 -8240
rect 9024 -8310 9096 -8240
rect 9096 -8310 9108 -8240
rect 9014 -8318 9108 -8310
rect 11082 -8238 11176 -8228
rect 11082 -8308 11092 -8238
rect 11092 -8308 11164 -8238
rect 11164 -8308 11176 -8238
rect 11082 -8316 11176 -8308
rect 13151 -8240 13245 -8230
rect 13151 -8310 13161 -8240
rect 13161 -8310 13233 -8240
rect 13233 -8310 13245 -8240
rect 13151 -8318 13245 -8310
rect 15219 -8238 15313 -8228
rect 15219 -8308 15229 -8238
rect 15229 -8308 15301 -8238
rect 15301 -8308 15313 -8238
rect 15219 -8316 15313 -8308
<< metal4 >>
rect 11131 4346 20908 4412
rect 11131 4226 12496 4346
rect 12618 4320 20908 4346
rect 12618 4318 16036 4320
rect 12618 4254 13698 4318
rect 13762 4254 14866 4318
rect 14930 4256 16036 4318
rect 16100 4256 17208 4320
rect 17272 4318 19544 4320
rect 17272 4256 18376 4318
rect 14930 4254 18376 4256
rect 18440 4256 19544 4318
rect 19608 4256 20712 4320
rect 20776 4256 20908 4320
rect 18440 4254 20908 4256
rect 12618 4226 20908 4254
rect 11131 4216 20908 4226
rect 11131 4185 11987 4216
rect 75 4129 11987 4185
rect 75 4127 3482 4129
rect 75 4055 536 4127
rect 606 4055 1984 4127
rect 2054 4057 3482 4127
rect 3552 4057 4930 4129
rect 5000 4127 9396 4129
rect 5000 4057 6450 4127
rect 2054 4055 6450 4057
rect 6520 4055 7898 4127
rect 7968 4057 9396 4127
rect 9466 4057 10844 4129
rect 10914 4057 11987 4129
rect 7968 4055 11987 4057
rect 75 4028 11987 4055
rect 75 4027 11314 4028
rect 75 2517 391 4027
rect 640 2517 24570 2520
rect 70 2414 24570 2517
rect 70 2410 7772 2414
rect 70 2374 1496 2410
rect 62 2318 1496 2374
rect 1596 2318 4640 2410
rect 4740 2322 7772 2410
rect 7872 2322 10916 2414
rect 11016 2410 20394 2414
rect 11016 2322 14118 2410
rect 4740 2318 14118 2322
rect 14218 2318 17262 2410
rect 17362 2322 20394 2410
rect 20494 2322 23538 2414
rect 23638 2322 24570 2414
rect 17362 2318 24570 2322
rect 62 2286 24570 2318
rect 62 2284 751 2286
rect 62 -216 350 2284
rect 640 -216 24570 -214
rect 62 -320 24570 -216
rect 62 -324 7772 -320
rect 62 -416 1496 -324
rect 1596 -416 4640 -324
rect 4740 -412 7772 -324
rect 7872 -412 10916 -320
rect 11016 -324 20394 -320
rect 11016 -412 14118 -324
rect 4740 -416 14118 -412
rect 14218 -416 17262 -324
rect 17362 -412 20394 -324
rect 20494 -412 23538 -320
rect 23638 -412 24570 -320
rect 17362 -416 24570 -412
rect 62 -448 24570 -416
rect 62 -451 861 -448
rect 62 -2939 350 -451
rect 62 -2946 825 -2939
rect 62 -3052 24560 -2946
rect 62 -3056 7762 -3052
rect 62 -3148 1486 -3056
rect 1586 -3148 4630 -3056
rect 4730 -3144 7762 -3056
rect 7862 -3144 10906 -3052
rect 11006 -3056 20384 -3052
rect 11006 -3144 14108 -3056
rect 4730 -3148 14108 -3144
rect 14208 -3148 17252 -3056
rect 17352 -3144 20384 -3056
rect 20484 -3144 23528 -3052
rect 23628 -3144 24560 -3052
rect 17352 -3148 24560 -3144
rect 62 -3174 24560 -3148
rect 62 -5874 350 -3174
rect 630 -3180 24560 -3174
rect 15976 -5863 16734 -5862
rect 15976 -5874 22331 -5863
rect -42 -5937 22331 -5874
rect -42 -6006 16861 -5937
rect -42 -6008 11144 -6006
rect -42 -6010 2870 -6008
rect -42 -6076 802 -6010
rect 878 -6074 2870 -6010
rect 2946 -6010 7007 -6008
rect 2946 -6074 4939 -6010
rect 878 -6076 4939 -6074
rect 5015 -6074 7007 -6010
rect 7083 -6074 9076 -6008
rect 9152 -6072 11144 -6008
rect 11220 -6008 15281 -6006
rect 11220 -6072 13213 -6008
rect 9152 -6074 13213 -6072
rect 13289 -6072 15281 -6008
rect 15357 -6045 16861 -6006
rect 16971 -5939 22331 -5937
rect 16971 -6045 17599 -5939
rect 15357 -6047 17599 -6045
rect 17709 -6047 18337 -5939
rect 18447 -6047 19079 -5939
rect 19189 -6047 19819 -5939
rect 19929 -6047 20557 -5939
rect 20667 -6047 21295 -5939
rect 21405 -6047 22033 -5939
rect 22143 -6047 22331 -5939
rect 15357 -6053 22331 -6047
rect 15357 -6072 16734 -6053
rect 13289 -6074 16734 -6072
rect 5015 -6076 16734 -6074
rect -42 -6118 16734 -6076
rect 62 -6127 350 -6118
rect 15976 -6120 16734 -6118
rect 16714 -6963 16732 -6773
rect 16968 -6963 16975 -6773
rect 17453 -6963 17466 -6773
rect 17702 -6963 17715 -6773
rect 18191 -6963 18214 -6773
rect 18450 -6963 18451 -6773
rect 18933 -6963 18955 -6773
rect 19191 -6963 19194 -6773
rect 19673 -6963 19686 -6773
rect 19922 -6963 19935 -6773
rect 20411 -6963 20425 -6773
rect 20661 -6963 20672 -6773
rect 21148 -6963 21171 -6773
rect 21407 -6963 21409 -6773
rect 21885 -6963 21898 -6773
rect 22134 -6963 22147 -6773
rect 665 -8416 671 -8226
rect 907 -8416 917 -8226
rect 2732 -8416 2738 -8224
rect 2974 -8416 2984 -8224
rect 4800 -8416 4811 -8226
rect 5047 -8416 5055 -8226
rect 6869 -8416 6879 -8224
rect 7115 -8416 7123 -8224
rect 8937 -8416 8952 -8224
rect 9188 -8416 9190 -8224
rect 11004 -8416 11016 -8222
rect 11252 -8416 11260 -8222
rect 13074 -8416 13079 -8224
rect 13315 -8416 13328 -8224
rect 15142 -8416 15152 -8222
rect 15388 -8416 15397 -8222
<< via4 >>
rect 679 2923 915 3016
rect 679 2855 758 2923
rect 758 2855 832 2923
rect 832 2855 915 2923
rect 679 2780 915 2855
rect 2128 2923 2364 3001
rect 2128 2855 2206 2923
rect 2206 2855 2280 2923
rect 2280 2855 2364 2923
rect 2128 2765 2364 2855
rect 3623 2925 3859 3010
rect 3623 2857 3704 2925
rect 3704 2857 3778 2925
rect 3778 2857 3859 2925
rect 3623 2774 3859 2857
rect 5072 2925 5308 3005
rect 5072 2857 5152 2925
rect 5152 2857 5226 2925
rect 5226 2857 5308 2925
rect 5072 2769 5308 2857
rect 6591 2923 6827 3005
rect 6591 2855 6672 2923
rect 6672 2855 6746 2923
rect 6746 2855 6827 2923
rect 6591 2769 6827 2855
rect 8039 2923 8275 3001
rect 8039 2855 8120 2923
rect 8120 2855 8194 2923
rect 8194 2855 8275 2923
rect 8039 2765 8275 2855
rect 9534 2925 9770 3016
rect 11970 3015 12206 3032
rect 9534 2857 9618 2925
rect 9618 2857 9692 2925
rect 9692 2857 9770 2925
rect 9534 2780 9770 2857
rect 10983 2925 11219 3010
rect 10983 2857 11066 2925
rect 11066 2857 11140 2925
rect 11140 2857 11219 2925
rect 10983 2774 11219 2857
rect 11970 2904 12039 3015
rect 12039 2904 12149 3015
rect 12149 2904 12206 3015
rect 11970 2796 12206 2904
rect 13142 3015 13378 3045
rect 13142 2904 13207 3015
rect 13207 2904 13317 3015
rect 13317 2904 13378 3015
rect 13142 2809 13378 2904
rect 14316 3015 14552 3032
rect 14316 2904 14375 3015
rect 14375 2904 14485 3015
rect 14485 2904 14552 3015
rect 14316 2796 14552 2904
rect 15480 3015 15716 3074
rect 15480 2904 15543 3015
rect 15543 2904 15653 3015
rect 15653 2904 15716 3015
rect 15480 2838 15716 2904
rect 16650 3017 16886 3072
rect 16650 2906 16717 3017
rect 16717 2906 16827 3017
rect 16827 2906 16886 3017
rect 16650 2836 16886 2906
rect 17819 3017 18055 3038
rect 17819 2906 17885 3017
rect 17885 2906 17995 3017
rect 17995 2906 18055 3017
rect 17819 2802 18055 2906
rect 18997 3017 19233 3050
rect 18997 2906 19053 3017
rect 19053 2906 19163 3017
rect 19163 2906 19233 3017
rect 18997 2814 19233 2906
rect 20162 3017 20398 3034
rect 20162 2906 20221 3017
rect 20221 2906 20331 3017
rect 20331 2906 20398 3017
rect 20162 2798 20398 2906
rect 1438 168 1674 208
rect 1438 100 1510 168
rect 1510 100 1594 168
rect 1594 100 1674 168
rect 1438 -28 1674 100
rect 4575 168 4811 194
rect 4575 100 4654 168
rect 4654 100 4738 168
rect 4738 100 4811 168
rect 4575 -42 4811 100
rect 7711 172 7947 212
rect 7711 104 7786 172
rect 7786 104 7870 172
rect 7870 104 7947 172
rect 7711 -24 7947 104
rect 10862 172 11098 203
rect 10862 104 10930 172
rect 10930 104 11014 172
rect 11014 104 11098 172
rect 10862 -33 11098 104
rect 14052 168 14288 216
rect 14052 100 14132 168
rect 14132 100 14216 168
rect 14216 100 14288 168
rect 14052 -20 14288 100
rect 17198 168 17434 212
rect 17198 100 17276 168
rect 17276 100 17360 168
rect 17360 100 17434 168
rect 17198 -24 17434 100
rect 20316 172 20552 221
rect 20316 104 20408 172
rect 20408 104 20492 172
rect 20492 104 20552 172
rect 20316 -15 20552 104
rect 23471 172 23707 194
rect 23471 104 23552 172
rect 23552 104 23636 172
rect 23636 104 23707 172
rect 23471 -42 23707 104
rect 1449 -2566 1685 -2507
rect 1449 -2634 1510 -2566
rect 1510 -2634 1594 -2566
rect 1594 -2634 1685 -2566
rect 1449 -2743 1685 -2634
rect 4589 -2566 4825 -2521
rect 4589 -2634 4654 -2566
rect 4654 -2634 4738 -2566
rect 4738 -2634 4825 -2566
rect 4589 -2757 4825 -2634
rect 7711 -2562 7947 -2529
rect 7711 -2630 7786 -2562
rect 7786 -2630 7870 -2562
rect 7870 -2630 7947 -2562
rect 7711 -2765 7947 -2630
rect 10867 -2562 11103 -2525
rect 10867 -2630 10930 -2562
rect 10930 -2630 11014 -2562
rect 11014 -2630 11103 -2562
rect 10867 -2761 11103 -2630
rect 14064 -2566 14300 -2529
rect 14064 -2634 14132 -2566
rect 14132 -2634 14216 -2566
rect 14216 -2634 14300 -2566
rect 14064 -2765 14300 -2634
rect 17197 -2566 17433 -2529
rect 17197 -2634 17276 -2566
rect 17276 -2634 17360 -2566
rect 17360 -2634 17433 -2566
rect 17197 -2765 17433 -2634
rect 20330 -2562 20566 -2520
rect 20330 -2630 20408 -2562
rect 20408 -2630 20492 -2562
rect 20492 -2630 20566 -2562
rect 20330 -2756 20566 -2630
rect 23462 -2562 23698 -2529
rect 23462 -2630 23552 -2562
rect 23552 -2630 23636 -2562
rect 23636 -2630 23698 -2562
rect 23462 -2765 23698 -2630
rect 1425 -5298 1661 -5258
rect 1425 -5366 1500 -5298
rect 1500 -5366 1584 -5298
rect 1584 -5366 1661 -5298
rect 1425 -5494 1661 -5366
rect 4579 -5298 4815 -5267
rect 4579 -5366 4644 -5298
rect 4644 -5366 4728 -5298
rect 4728 -5366 4815 -5298
rect 4579 -5503 4815 -5366
rect 7710 -5294 7946 -5267
rect 7710 -5362 7776 -5294
rect 7776 -5362 7860 -5294
rect 7860 -5362 7946 -5294
rect 7710 -5503 7946 -5362
rect 10841 -5294 11077 -5267
rect 10841 -5362 10920 -5294
rect 10920 -5362 11004 -5294
rect 11004 -5362 11077 -5294
rect 10841 -5503 11077 -5362
rect 14050 -5298 14286 -5272
rect 14050 -5366 14122 -5298
rect 14122 -5366 14206 -5298
rect 14206 -5366 14286 -5298
rect 14050 -5508 14286 -5366
rect 17191 -5298 17427 -5253
rect 17191 -5366 17266 -5298
rect 17266 -5366 17350 -5298
rect 17350 -5366 17427 -5298
rect 17191 -5489 17427 -5366
rect 20326 -5294 20562 -5267
rect 20326 -5362 20398 -5294
rect 20398 -5362 20482 -5294
rect 20482 -5362 20562 -5294
rect 20326 -5503 20562 -5362
rect 23466 -5294 23702 -5249
rect 23466 -5362 23542 -5294
rect 23542 -5362 23626 -5294
rect 23626 -5362 23702 -5294
rect 23466 -5485 23702 -5362
rect 16732 -6829 16968 -6754
rect 16732 -6929 16801 -6829
rect 16801 -6929 16903 -6829
rect 16903 -6929 16968 -6829
rect 16732 -6990 16968 -6929
rect 17466 -6831 17702 -6756
rect 17466 -6931 17539 -6831
rect 17539 -6931 17641 -6831
rect 17641 -6931 17702 -6831
rect 17466 -6992 17702 -6931
rect 18214 -6831 18450 -6758
rect 18214 -6931 18277 -6831
rect 18277 -6931 18379 -6831
rect 18379 -6931 18450 -6831
rect 18214 -6994 18450 -6931
rect 18955 -6831 19191 -6763
rect 18955 -6931 19019 -6831
rect 19019 -6931 19121 -6831
rect 19121 -6931 19191 -6831
rect 18955 -6999 19191 -6931
rect 19686 -6831 19922 -6752
rect 19686 -6931 19759 -6831
rect 19759 -6931 19861 -6831
rect 19861 -6931 19922 -6831
rect 19686 -6988 19922 -6931
rect 20425 -6831 20661 -6752
rect 20425 -6931 20497 -6831
rect 20497 -6931 20599 -6831
rect 20599 -6931 20661 -6831
rect 20425 -6988 20661 -6931
rect 21171 -6831 21407 -6754
rect 21171 -6931 21235 -6831
rect 21235 -6931 21337 -6831
rect 21337 -6931 21407 -6831
rect 21171 -6990 21407 -6931
rect 21898 -6831 22134 -6756
rect 21898 -6931 21973 -6831
rect 21973 -6931 22075 -6831
rect 22075 -6931 22134 -6831
rect 21898 -6992 22134 -6931
rect 671 -8232 907 -8199
rect 671 -8320 740 -8232
rect 740 -8320 834 -8232
rect 834 -8320 907 -8232
rect 671 -8435 907 -8320
rect 2738 -8230 2974 -8190
rect 2738 -8318 2808 -8230
rect 2808 -8318 2902 -8230
rect 2902 -8318 2974 -8230
rect 2738 -8426 2974 -8318
rect 4811 -8232 5047 -8185
rect 4811 -8320 4877 -8232
rect 4877 -8320 4971 -8232
rect 4971 -8320 5047 -8232
rect 4811 -8421 5047 -8320
rect 6879 -8230 7115 -8192
rect 6879 -8318 6945 -8230
rect 6945 -8318 7039 -8230
rect 7039 -8318 7115 -8230
rect 6879 -8428 7115 -8318
rect 8952 -8230 9188 -8199
rect 8952 -8318 9014 -8230
rect 9014 -8318 9108 -8230
rect 9108 -8318 9188 -8230
rect 8952 -8435 9188 -8318
rect 11016 -8228 11252 -8195
rect 11016 -8316 11082 -8228
rect 11082 -8316 11176 -8228
rect 11176 -8316 11252 -8228
rect 11016 -8431 11252 -8316
rect 13079 -8230 13315 -8195
rect 13079 -8318 13151 -8230
rect 13151 -8318 13245 -8230
rect 13245 -8318 13315 -8230
rect 13079 -8431 13315 -8318
rect 15152 -8228 15388 -8183
rect 15152 -8316 15219 -8228
rect 15219 -8316 15313 -8228
rect 15313 -8316 15388 -8228
rect 15152 -8419 15388 -8316
<< metal5 >>
rect 495 3074 23948 3241
rect 495 3045 15480 3074
rect 495 3032 13142 3045
rect 495 3016 11970 3032
rect 495 2780 679 3016
rect 915 3010 9534 3016
rect 915 3001 3623 3010
rect 915 2780 2128 3001
rect 495 2765 2128 2780
rect 2364 2774 3623 3001
rect 3859 3005 9534 3010
rect 3859 2774 5072 3005
rect 2364 2769 5072 2774
rect 5308 2769 6591 3005
rect 6827 3001 9534 3005
rect 6827 2769 8039 3001
rect 2364 2765 8039 2769
rect 8275 2780 9534 3001
rect 9770 3010 11970 3016
rect 9770 2780 10983 3010
rect 8275 2774 10983 2780
rect 11219 2796 11970 3010
rect 12206 2809 13142 3032
rect 13378 3032 15480 3045
rect 13378 2809 14316 3032
rect 12206 2796 14316 2809
rect 14552 2838 15480 3032
rect 15716 3072 23948 3074
rect 15716 2838 16650 3072
rect 14552 2836 16650 2838
rect 16886 3050 23948 3072
rect 16886 3038 18997 3050
rect 16886 2836 17819 3038
rect 14552 2802 17819 2836
rect 18055 2814 18997 3038
rect 19233 3034 23948 3050
rect 19233 2814 20162 3034
rect 18055 2802 20162 2814
rect 14552 2798 20162 2802
rect 20398 2798 23948 3034
rect 14552 2796 23948 2798
rect 11219 2774 23948 2796
rect 8275 2765 23948 2774
rect 495 221 23948 2765
rect 495 216 20316 221
rect 495 212 14052 216
rect 495 208 7711 212
rect 495 -28 1438 208
rect 1674 194 7711 208
rect 1674 -28 4575 194
rect 495 -42 4575 -28
rect 4811 -24 7711 194
rect 7947 203 14052 212
rect 7947 -24 10862 203
rect 4811 -33 10862 -24
rect 11098 -20 14052 203
rect 14288 212 20316 216
rect 14288 -20 17198 212
rect 11098 -24 17198 -20
rect 17434 -15 20316 212
rect 20552 194 23948 221
rect 20552 -15 23471 194
rect 17434 -24 23471 -15
rect 11098 -33 23471 -24
rect 4811 -42 23471 -33
rect 23707 -42 23948 194
rect 495 -2507 23948 -42
rect 495 -2743 1449 -2507
rect 1685 -2520 23948 -2507
rect 1685 -2521 20330 -2520
rect 1685 -2743 4589 -2521
rect 495 -2757 4589 -2743
rect 4825 -2525 20330 -2521
rect 4825 -2529 10867 -2525
rect 4825 -2757 7711 -2529
rect 495 -2765 7711 -2757
rect 7947 -2761 10867 -2529
rect 11103 -2529 20330 -2525
rect 11103 -2761 14064 -2529
rect 7947 -2765 14064 -2761
rect 14300 -2765 17197 -2529
rect 17433 -2756 20330 -2529
rect 20566 -2529 23948 -2520
rect 20566 -2756 23462 -2529
rect 17433 -2765 23462 -2756
rect 23698 -2765 23948 -2529
rect 495 -5249 23948 -2765
rect 495 -5253 23466 -5249
rect 495 -5258 17191 -5253
rect 495 -5494 1425 -5258
rect 1661 -5267 17191 -5258
rect 1661 -5494 4579 -5267
rect 495 -5503 4579 -5494
rect 4815 -5503 7710 -5267
rect 7946 -5503 10841 -5267
rect 11077 -5272 17191 -5267
rect 11077 -5503 14050 -5272
rect 495 -5508 14050 -5503
rect 14286 -5489 17191 -5272
rect 17427 -5267 23466 -5253
rect 17427 -5489 20326 -5267
rect 14286 -5503 20326 -5489
rect 20562 -5485 23466 -5267
rect 23702 -5485 23948 -5249
rect 20562 -5503 23948 -5485
rect 14286 -5508 23948 -5503
rect 495 -6752 23948 -5508
rect 495 -6754 19686 -6752
rect 495 -6990 16732 -6754
rect 16968 -6756 19686 -6754
rect 16968 -6990 17466 -6756
rect 495 -6992 17466 -6990
rect 17702 -6758 19686 -6756
rect 17702 -6992 18214 -6758
rect 495 -6994 18214 -6992
rect 18450 -6763 19686 -6758
rect 18450 -6994 18955 -6763
rect 495 -6999 18955 -6994
rect 19191 -6988 19686 -6763
rect 19922 -6988 20425 -6752
rect 20661 -6754 23948 -6752
rect 20661 -6988 21171 -6754
rect 19191 -6990 21171 -6988
rect 21407 -6756 23948 -6754
rect 21407 -6990 21898 -6756
rect 19191 -6992 21898 -6990
rect 22134 -6992 23948 -6756
rect 19191 -6999 23948 -6992
rect 495 -8183 23948 -6999
rect 495 -8185 15152 -8183
rect 495 -8190 4811 -8185
rect 495 -8199 2738 -8190
rect 495 -8435 671 -8199
rect 907 -8426 2738 -8199
rect 2974 -8421 4811 -8190
rect 5047 -8192 15152 -8185
rect 5047 -8421 6879 -8192
rect 2974 -8426 6879 -8421
rect 907 -8428 6879 -8426
rect 7115 -8195 15152 -8192
rect 7115 -8199 11016 -8195
rect 7115 -8428 8952 -8199
rect 907 -8435 8952 -8428
rect 9188 -8431 11016 -8199
rect 11252 -8431 13079 -8195
rect 13315 -8419 15152 -8195
rect 15388 -8419 23948 -8183
rect 13315 -8431 23948 -8419
rect 9188 -8435 23948 -8431
rect 495 -8882 23948 -8435
<< labels >>
flabel metal5 17354 -8713 19521 -7975 1 FreeSerif 3200 0 0 0 VSS
port 27 n
flabel metal4 11192 4053 11897 4378 1 FreeSerif 1600 0 0 0 VDD
port 28 n
flabel metal1 -2300 -7075 -2258 -7026 1 FreeSerif 640 0 0 0 A[0]
port 30 n
flabel metal1 -2302 -6869 -2253 -6816 1 FreeSerif 640 0 0 0 A[1]
port 31 n
flabel metal1 -2298 -6681 -2240 -6627 1 FreeSerif 640 0 0 0 A[2]
port 32 n
flabel metal1 -2300 -6374 -2241 -6318 1 FreeSerif 640 0 0 0 A[4]
port 16 n
flabel metal1 -2302 -6525 -2238 -6471 1 FreeSerif 640 0 0 0 A[3]
port 33 n
flabel metal1 -2302 -6214 -2240 -6156 1 FreeSerif 640 0 0 0 A[5]
port 17 n
flabel metal1 -2300 -5905 -2243 -5853 1 FreeSerif 720 0 0 0 A[6]
port 18 n
flabel metal1 -2300 -5614 -2240 -5561 1 FreeSerif 720 0 0 0 A[7]
port 34 n
flabel metal1 -2580 2740 -2542 2788 1 FreeSerif 720 0 0 0 B[0]
port 35 n
flabel metal1 -2579 3115 -2518 3161 1 FreeSerif 720 0 0 0 B[1]
port 36 n
flabel metal1 -2580 4905 -2520 4964 1 FreeSerif 720 0 0 0 B[2]
port 37 n
flabel metal1 -2581 5102 -2521 5161 1 FreeSerif 720 0 0 0 B[3]
port 38 n
flabel metal1 -2579 5286 -2519 5345 1 FreeSerif 720 0 0 0 B[4]
port 39 n
flabel metal1 -2579 5473 -2519 5532 1 FreeSerif 720 0 0 0 B[5]
port 40 n
flabel metal1 -2578 5663 -2518 5722 1 FreeSerif 720 0 0 0 B[6]
port 41 n
flabel metal1 -2577 5865 -2518 5920 1 FreeSerif 720 0 0 0 B[7]
port 42 n
flabel metal1 -2605 -1361 -2535 -1289 1 FreeSerif 720 0 0 0 opcode[1]
port 43 n
flabel metal1 -2607 -1687 -2529 -1619 1 FreeSerif 720 0 0 0 opcode[0]
port 44 n
flabel metal1 25246 -1483 25335 -1353 1 FreeSerif 720 0 0 0 Y[7]
port 45 n
flabel metal1 25288 -1842 25336 -1780 1 FreeSerif 720 0 0 0 Y[6]
port 46 n
flabel metal1 25283 -2033 25336 -1971 1 FreeSerif 720 0 0 0 Y[5]
port 7 n
flabel metal1 25283 -2255 25334 -2193 1 FreeSerif 720 0 0 0 Y[4]
port 6 n
flabel metal1 25278 -2446 25333 -2382 1 FreeSerif 720 0 0 0 Y[3]
port 5 n
flabel metal1 25278 -2787 25334 -2723 1 FreeSerif 720 0 0 0 Y[2]
port 4 n
flabel metal1 25282 -2959 25335 -2898 1 FreeSerif 720 0 0 0 Y[1]
port 3 n
flabel metal1 25282 -3319 25340 -3254 1 FreeSerif 720 0 0 0 Y[0]
port 47 n
<< end >>
