** sch_path: /home/ume/Desktop/designFinal/xschem/arithmetic_unit.sch
**.subckt arithmetic_unit A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7]
*+ B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7] opcode[0],opcode[1] Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7] Cout VSS VDD
*.ipin A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7]
*.ipin B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7]
*.ipin opcode[0],opcode[1]
*.opin Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7]
*.opin Cout
*.iopin VSS
*.iopin VDD
x1 sub[0] opcode[0] VDD VSS B[0] xor2
x2 sub[1] opcode[0] VDD VSS B[1] xor2
x3 sub[2] opcode[0] VDD VSS B[2] xor2
x4 sub[3] opcode[0] VDD VSS B[3] xor2
x5 sub[4] opcode[0] VDD VSS B[4] xor2
x6 sub[5] opcode[0] VDD VSS B[5] xor2
x7 sub[6] opcode[0] VDD VSS B[6] xor2
x8 sub[7] opcode[0] VDD VSS B[7] xor2
x9 VSS VDD opcode[1] adder[0] multi[0] Y[0] 2x1_mux
x10 VSS VDD opcode[1] adder[1] multi[1] Y[1] 2x1_mux
x11 VSS VDD opcode[1] adder[2] multi[2] Y[2] 2x1_mux
x12 VSS VDD opcode[1] adder[3] multi[3] Y[3] 2x1_mux
x13 VSS VDD opcode[1] adder[4] multi[4] Y[4] 2x1_mux
x14 VSS VDD opcode[1] adder[5] multi[5] Y[5] 2x1_mux
x15 VSS VDD opcode[1] adder[6] multi[6] Y[6] 2x1_mux
x16 VSS VDD opcode[1] adder[7] multi[7] Y[7] 2x1_mux
x18 A[3] A[4] A[5] A[6] B[3] B[4] B[5] B[6] VDD VSS multi[0] multi[1] multi[2] multi[3] multi[4]
+ multi[5] multi[6] multi[7] array_multiplier
x17 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] sub[0] sub[1] sub[2] sub[3] sub[4] sub[5] sub[6] sub[7]
+ opcode[0] VDD VSS adder[0] adder[1] adder[2] adder[3] adder[4] adder[5] adder[6] adder[7] Cout
+ carry_ripple_adder
**.ends

* expanding   symbol:  xor2.sym # of pins=5
** sym_path: /home/ume/Desktop/designFinal/xschem/xor2.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/xor2.sch
.subckt xor2  Y A VDD VSS B
*.opin Y
*.ipin A
*.iopin VDD
*.iopin VSS
*.ipin B
XM7 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Y inv_B net1 VDD sky130_fd_pr__pfet_01v8 L=0.30 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Y inv_A net1 VDD sky130_fd_pr__pfet_01v8 L=0.30 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Y A net2 VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y inv_A net3 VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 inv_B VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 inv_B B VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 inv_B B VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 inv_A A VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 inv_A A VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  2x1_mux.sym # of pins=6
** sym_path: /home/ume/Desktop/designFinal/xschem/2x1_mux.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/2x1_mux.sch
.subckt 2x1_mux  VSS VDD S D0 D1 OUT
*.iopin VSS
*.iopin VDD
*.ipin S
*.ipin D0
*.ipin D1
*.opin OUT
XM2 net1 S_BAR net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 D1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 D0 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 S_BAR net4 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 D1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net4 S VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 S_BAR S VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 S_BAR S VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 S net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 D0 net4 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  array_multiplier.sym # of pins=5
** sym_path: /home/ume/Desktop/designFinal/xschem/array_multiplier.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/array_multiplier.sch
.subckt array_multiplier  A[0] A[1] A[2] A[3] B[0] B[1] B[2] B[3] VDD VSS Y[0] Y[1] Y[2] Y[3] Y[4]
+ Y[5] Y[6] Y[7]
*.ipin A[0],A[1],A[2],A[3]
*.ipin B[0],B[1],B[2],B[3]
*.iopin VDD
*.iopin VSS
*.opin Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7]
x1 VSS A[1] B[1] VDD net1 and2
x2 VSS A[2] B[0] VDD net2 and2
x3 VSS A[2] B[1] VDD net3 and2
x4 VSS A[3] B[0] VDD net4 and2
x5 net1 net2 net30 net24 net5 VDD VSS fulladder
x6 net3 net4 net5 net7 net10 VDD VSS fulladder
x7 VSS A[1] B[2] VDD net6 and2
x8 net7 net6 net31 net26 net8 VDD VSS fulladder
x9 VSS A[3] B[1] VDD net9 and2
x10 net10 net9 net8 net12 net13 VDD VSS fulladder
x11 VSS A[2] B[2] VDD net11 and2
x12 net12 net11 net32 net20 net15 VDD VSS fulladder
x13 VSS A[3] B[2] VDD net14 and2
x14 VSS A[2] B[3] VDD net17 and2
x15 VSS A[1] B[3] VDD net19 and2
x17 VSS A[0] B[1] VDD net21 and2
x18 VSS A[1] B[0] VDD net22 and2
x19 VSS A[0] B[2] VDD net23 and2
x20 VSS A[0] B[3] VDD net25 and2
x21 VSS A[3] B[3] VDD net28 and2
x22 net16 net17 net18 Y[5] net29 VDD VSS fulladder
x23 net20 net19 Y[4] net18 VDD VSS half_adder
x16 net13 net14 net15 net16 net27 VDD VSS fulladder
x24 net24 net23 Y[2] net31 VDD VSS half_adder
x25 net21 net22 Y[1] net30 VDD VSS half_adder
x26 VSS A[0] B[0] VDD Y[0] and2
x27 net26 net25 Y[3] net32 VDD VSS half_adder
x28 net27 net28 net29 Y[6] Y[7] VDD VSS fulladder
.ends


* expanding   symbol:  carry_ripple_adder.sym # of pins=7
** sym_path: /home/ume/Desktop/designFinal/xschem/carry_ripple_adder.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/carry_ripple_adder.sch
.subckt carry_ripple_adder  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4] B[5]
+ B[6] B[7] carry_in VDD VSS Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] carry_out
*.ipin A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7]
*.ipin B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7]
*.ipin carry_in
*.iopin VDD
*.iopin VSS
*.opin Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7]
*.opin carry_out
x1 A[0] B[0] carry_in Y[0] net1 VDD VSS fulladder
x2 A[1] B[1] net1 Y[1] net2 VDD VSS fulladder
x3 A[2] B[2] net2 Y[2] net3 VDD VSS fulladder
x4 A[3] B[3] net3 Y[3] net4 VDD VSS fulladder
x5 A[4] B[4] net4 Y[4] net5 VDD VSS fulladder
x6 A[5] B[5] net5 Y[5] net6 VDD VSS fulladder
x7 A[6] B[6] net6 Y[6] net7 VDD VSS fulladder
x8 A[7] B[7] net7 Y[7] carry_out VDD VSS fulladder
.ends


* expanding   symbol:  and2.sym # of pins=5
** sym_path: /home/ume/Desktop/designFinal/xschem/and2.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/and2.sch
.subckt and2  VSS A B VDD OUT
*.iopin VSS
*.ipin A
*.ipin B
*.iopin VDD
*.opin OUT
XM2 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A net2 VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  fulladder.sym # of pins=7
** sym_path: /home/ume/Desktop/designFinal/xschem/fulladder.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/fulladder.sch
.subckt fulladder  A B carry_in Y carry_out VDD VSS
*.ipin A
*.ipin B
*.ipin carry_in
*.opin Y
*.opin carry_out
*.iopin VDD
*.iopin VSS
x1 VSS A B VDD net1 and2
x2 VSS B carry_in VDD net2 and2
x3 VSS A carry_in VDD net3 and2
x4 VDD net1 net3 net2 carry_out VSS or3
x5 VDD A Y B carry_in VSS xor3
.ends


* expanding   symbol:  half_adder.sym # of pins=6
** sym_path: /home/ume/Desktop/designFinal/xschem/half_adder.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/half_adder.sch
.subckt half_adder  A B Y carry_out VDD VSS
*.ipin A
*.ipin B
*.opin Y
*.opin carry_out
*.iopin VDD
*.iopin VSS
x1 Y A VDD VSS B xor2
x2 VSS A B VDD carry_out and2
.ends


* expanding   symbol:  or3.sym # of pins=6
** sym_path: /home/ume/Desktop/designFinal/xschem/or3.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/or3.sch
.subckt or3  VDD A B C OUT VSS
*.ipin A
*.ipin B
*.iopin VSS
*.iopin VDD
*.opin OUT
*.ipin C
XM4 net1 A net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 C VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 B net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 C VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xor3.sym # of pins=6
** sym_path: /home/ume/Desktop/designFinal/xschem/xor3.sym
** sch_path: /home/ume/Desktop/designFinal/xschem/xor3.sch
.subckt xor3  VDD A OUT B C VSS
*.ipin C
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
*.iopin VDD
x1 net1 A VDD VSS B xor2
x2 OUT net1 VDD VSS C xor2
.ends

.end
