magic
tech sky130B
magscale 1 2
timestamp 1733691381
<< error_p >>
rect -324 181 -266 187
rect -206 181 -148 187
rect -88 181 -30 187
rect 30 181 88 187
rect 148 181 206 187
rect 266 181 324 187
rect -324 147 -312 181
rect -206 147 -194 181
rect -88 147 -76 181
rect 30 147 42 181
rect 148 147 160 181
rect 266 147 278 181
rect -324 141 -266 147
rect -206 141 -148 147
rect -88 141 -30 147
rect 30 141 88 147
rect 148 141 206 147
rect 266 141 324 147
rect -324 -147 -266 -141
rect -206 -147 -148 -141
rect -88 -147 -30 -141
rect 30 -147 88 -141
rect 148 -147 206 -141
rect 266 -147 324 -141
rect -324 -181 -312 -147
rect -206 -181 -194 -147
rect -88 -181 -76 -147
rect 30 -181 42 -147
rect 148 -181 160 -147
rect 266 -181 278 -147
rect -324 -187 -266 -181
rect -206 -187 -148 -181
rect -88 -187 -30 -181
rect 30 -187 88 -181
rect 148 -187 206 -181
rect 266 -187 324 -181
<< nwell >>
rect -419 -200 419 200
<< pmos >>
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
<< pdiff >>
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
<< pdiffc >>
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
<< poly >>
rect -328 181 -262 197
rect -328 147 -312 181
rect -278 147 -262 181
rect -328 131 -262 147
rect -210 181 -144 197
rect -210 147 -194 181
rect -160 147 -144 181
rect -210 131 -144 147
rect -92 181 -26 197
rect -92 147 -76 181
rect -42 147 -26 181
rect -92 131 -26 147
rect 26 181 92 197
rect 26 147 42 181
rect 76 147 92 181
rect 26 131 92 147
rect 144 181 210 197
rect 144 147 160 181
rect 194 147 210 181
rect 144 131 210 147
rect 262 181 328 197
rect 262 147 278 181
rect 312 147 328 181
rect 262 131 328 147
rect -325 100 -265 131
rect -207 100 -147 131
rect -89 100 -29 131
rect 29 100 89 131
rect 147 100 207 131
rect 265 100 325 131
rect -325 -131 -265 -100
rect -207 -131 -147 -100
rect -89 -131 -29 -100
rect 29 -131 89 -100
rect 147 -131 207 -100
rect 265 -131 325 -100
rect -328 -147 -262 -131
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -328 -197 -262 -181
rect -210 -147 -144 -131
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -210 -197 -144 -181
rect -92 -147 -26 -131
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect -92 -197 -26 -181
rect 26 -147 92 -131
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 26 -197 92 -181
rect 144 -147 210 -131
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 144 -197 210 -181
rect 262 -147 328 -131
rect 262 -181 278 -147
rect 312 -181 328 -147
rect 262 -197 328 -181
<< polycont >>
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
<< locali >>
rect -328 147 -312 181
rect -278 147 -262 181
rect -210 147 -194 181
rect -160 147 -144 181
rect -92 147 -76 181
rect -42 147 -26 181
rect 26 147 42 181
rect 76 147 92 181
rect 144 147 160 181
rect 194 147 210 181
rect 262 147 278 181
rect 312 147 328 181
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 262 -181 278 -147
rect 312 -181 328 -147
<< viali >>
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
<< metal1 >>
rect -324 181 -266 187
rect -324 147 -312 181
rect -278 147 -266 181
rect -324 141 -266 147
rect -206 181 -148 187
rect -206 147 -194 181
rect -160 147 -148 181
rect -206 141 -148 147
rect -88 181 -30 187
rect -88 147 -76 181
rect -42 147 -30 181
rect -88 141 -30 147
rect 30 181 88 187
rect 30 147 42 181
rect 76 147 88 181
rect 30 141 88 147
rect 148 181 206 187
rect 148 147 160 181
rect 194 147 206 181
rect 148 141 206 147
rect 266 181 324 187
rect 266 147 278 181
rect 312 147 324 181
rect 266 141 324 147
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect -324 -147 -266 -141
rect -324 -181 -312 -147
rect -278 -181 -266 -147
rect -324 -187 -266 -181
rect -206 -147 -148 -141
rect -206 -181 -194 -147
rect -160 -181 -148 -147
rect -206 -187 -148 -181
rect -88 -147 -30 -141
rect -88 -181 -76 -147
rect -42 -181 -30 -147
rect -88 -187 -30 -181
rect 30 -147 88 -141
rect 30 -181 42 -147
rect 76 -181 88 -147
rect 30 -187 88 -181
rect 148 -147 206 -141
rect 148 -181 160 -147
rect 194 -181 206 -147
rect 148 -187 206 -181
rect 266 -147 324 -141
rect 266 -181 278 -147
rect 312 -181 324 -147
rect 266 -187 324 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
