* NGSPICE file created from logic_and_pex.ext - technology: sky130B

.subckt logic_and A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3]
+ Y[4] Y[5] Y[6] Y[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
X0 a_155_68.t5 A[0].t0 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 a_155_68.t4 A[0].t1 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 VDD.t5 B[0].t0 a_155_68.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 VDD.t89 B[5].t0 a_7517_68.t4 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4 a_10463_70.t5 B[7].t0 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 VDD.t7 A[7].t0 a_10463_70.t0 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 a_4549_70.t5 A[3].t0 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7 Y[0].t2 a_155_68.t7 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 VDD.t45 A[1].t0 a_1603_68.t5 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 VDD.t75 B[4].t0 a_6069_68.t2 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 VDD.t65 B[6].t0 a_9015_70.t4 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X11 a_3338_n567.t1 A[2].t0 a_3101_70.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 Y[6].t3 a_9015_70.t7 VSS.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 a_6069_68.t3 A[4].t0 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X14 Y[5].t2 a_7517_68.t7 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 VDD.t49 B[7].t1 a_10463_70.t4 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 VSS.t5 B[6].t1 a_9252_n567.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 VDD.t137 a_10463_70.t7 Y[7].t2 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X18 VDD.t57 B[3].t0 a_4549_70.t1 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X19 Y[4].t2 a_6069_68.t7 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X20 Y[1].t3 a_1603_68.t7 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X21 a_9015_70.t3 B[6].t2 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X22 a_10700_n567.t1 A[7].t1 a_10463_70.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 VDD.t15 a_155_68.t8 Y[0].t1 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X24 a_1603_68.t2 B[1].t0 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 VDD.t91 a_1603_68.t8 Y[1].t2 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VDD.t19 A[2].t1 a_3101_70.t5 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 VDD.t107 B[3].t1 a_4549_70.t6 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 VDD.t143 B[4].t1 a_6069_68.t1 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 VSS.t6 B[5].t1 a_7754_n569.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X30 VDD.t101 a_7517_68.t8 Y[5].t1 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 VDD.t119 A[6].t0 a_9015_70.t6 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 Y[7].t1 a_10463_70.t8 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X33 a_4549_70.t0 B[3].t2 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 VDD.t109 a_6069_68.t8 Y[4].t1 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X35 a_7517_68.t5 A[5].t0 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X36 Y[6].t2 a_9015_70.t8 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X37 Y[1].t1 a_1603_68.t9 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X38 Y[5].t0 a_7517_68.t9 VDD.t127 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X39 VDD.t141 B[6].t3 a_9015_70.t2 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X40 VDD.t11 B[1].t1 a_1603_68.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 a_3101_70.t4 A[2].t2 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X42 Y[3].t2 a_4549_70.t7 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 a_6069_68.t0 B[4].t2 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X44 VSS.t9 B[3].t3 a_4786_n567.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X45 a_9015_70.t5 A[6].t1 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 a_1840_n569.t1 A[1].t1 a_1603_68.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X47 a_7517_68.t3 B[5].t2 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X48 Y[7].t0 a_10463_70.t9 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X49 Y[0].t3 a_155_68.t9 VSS.t10 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 Y[4].t3 a_6069_68.t9 VSS.t8 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 Y[2].t2 a_3101_70.t7 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X52 Y[4].t0 a_6069_68.t10 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X53 VSS.t14 B[0].t1 a_392_n569.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 Y[5].t3 a_7517_68.t10 VSS.t12 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X55 VDD.t113 a_4549_70.t8 Y[3].t1 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 VDD.t83 A[5].t1 a_7517_68.t1 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 Y[6].t1 a_9015_70.t9 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X58 VSS.t2 B[4].t3 a_6306_n569.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X59 VDD.t25 B[0].t2 a_155_68.t2 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X60 Y[1].t0 a_1603_68.t10 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 VDD.t3 B[2].t0 a_3101_70.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 a_10463_70.t6 A[7].t2 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_3101_70.t3 A[2].t3 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X64 VSS.t7 B[7].t2 a_10700_n567.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X65 a_1603_68.t4 A[1].t2 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 Y[2].t3 a_3101_70.t8 VSS.t15 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 a_9252_n567.t0 A[6].t2 a_9015_70.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X68 a_3101_70.t1 B[2].t1 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 VDD.t27 a_3101_70.t9 Y[2].t1 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X70 a_4549_70.t4 A[3].t1 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 a_7517_68.t0 A[5].t2 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X72 Y[3].t3 a_4549_70.t9 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 a_155_68.t1 B[0].t3 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X74 Y[3].t0 a_4549_70.t10 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 a_6069_68.t4 A[4].t1 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 VDD.t33 a_9015_70.t10 Y[6].t0 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 VSS.t4 B[2].t2 a_3338_n567.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X78 VDD.t59 A[0].t2 a_155_68.t3 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 Y[0].t0 a_155_68.t10 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_10463_70.t1 A[7].t3 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X81 VDD.t121 B[7].t3 a_10463_70.t3 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X82 a_4786_n567.t0 A[3].t2 a_4549_70.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X83 VDD.t73 A[3].t3 a_4549_70.t3 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 VDD.t17 B[5].t3 a_7517_68.t2 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 a_9015_70.t0 A[6].t3 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X86 a_7754_n569.t1 A[5].t3 a_7517_68.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 Y[7].t3 a_10463_70.t10 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X88 a_1603_68.t3 A[1].t3 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 VDD.t97 B[1].t2 a_1603_68.t1 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X90 Y[2].t0 a_3101_70.t10 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X91 a_392_n569.t0 A[0].t3 a_155_68.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X92 VSS.t11 B[1].t3 a_1840_n569.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 a_6306_n569.t0 A[4].t2 a_6069_68.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X94 VDD.t99 B[2].t3 a_3101_70.t6 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X95 VDD.t115 A[4].t3 a_6069_68.t6 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 A[0].t3 A[0].t1 437.233
R1 A[0] A[0].t3 216.701
R2 A[0].n0 A[0].t0 214.686
R3 A[0].t1 A[0].n0 214.686
R4 A[0].n0 A[0].t2 80.333
R5 VDD.t90 VDD.t130 196.666
R6 VDD.t52 VDD.t90 196.666
R7 VDD.t10 VDD.t52 196.666
R8 VDD.t116 VDD.t10 196.666
R9 VDD.t96 VDD.t116 196.666
R10 VDD.t66 VDD.t44 196.666
R11 VDD.t44 VDD.t46 196.666
R12 VDD.t108 VDD.t128 196.666
R13 VDD.t38 VDD.t108 196.666
R14 VDD.t74 VDD.t38 196.666
R15 VDD.t50 VDD.t74 196.666
R16 VDD.t142 VDD.t50 196.666
R17 VDD.t68 VDD.t114 196.666
R18 VDD.t114 VDD.t80 196.666
R19 VDD.t100 VDD.t126 196.666
R20 VDD.t94 VDD.t100 196.666
R21 VDD.t88 VDD.t94 196.666
R22 VDD.t122 VDD.t88 196.666
R23 VDD.t16 VDD.t122 196.666
R24 VDD.t70 VDD.t82 196.666
R25 VDD.t82 VDD.t104 196.666
R26 VDD.t32 VDD.t34 196.666
R27 VDD.t86 VDD.t32 196.666
R28 VDD.t140 VDD.t86 196.666
R29 VDD.t40 VDD.t140 196.666
R30 VDD.t64 VDD.t40 196.666
R31 VDD.t102 VDD.t118 196.666
R32 VDD.t118 VDD.t0 196.666
R33 VDD.t136 VDD.t76 196.666
R34 VDD.t36 VDD.t136 196.666
R35 VDD.t48 VDD.t36 196.666
R36 VDD.t78 VDD.t48 196.666
R37 VDD.t120 VDD.t78 196.666
R38 VDD.t92 VDD.t6 196.666
R39 VDD.t6 VDD.t42 196.666
R40 VDD.t26 VDD.t28 196.666
R41 VDD.t132 VDD.t26 196.666
R42 VDD.t98 VDD.t132 196.666
R43 VDD.t12 VDD.t98 196.666
R44 VDD.t2 VDD.t12 196.666
R45 VDD.t134 VDD.t18 196.666
R46 VDD.t18 VDD.t30 196.666
R47 VDD.t112 VDD.t124 196.666
R48 VDD.t20 VDD.t112 196.666
R49 VDD.t106 VDD.t20 196.666
R50 VDD.t8 VDD.t106 196.666
R51 VDD.t56 VDD.t8 196.666
R52 VDD.t84 VDD.t72 196.666
R53 VDD.t72 VDD.t54 196.666
R54 VDD.t14 VDD.t110 196.666
R55 VDD.t138 VDD.t14 196.666
R56 VDD.t4 VDD.t138 196.666
R57 VDD.t22 VDD.t4 196.666
R58 VDD.t24 VDD.t22 196.666
R59 VDD.t60 VDD.t58 196.666
R60 VDD.t58 VDD.t62 196.666
R61 VDD.n59 VDD.t47 30.163
R62 VDD.n7 VDD.t81 30.163
R63 VDD.n15 VDD.t105 30.163
R64 VDD.n23 VDD.t1 30.163
R65 VDD.n31 VDD.t43 30.163
R66 VDD.n51 VDD.t31 30.163
R67 VDD.n43 VDD.t55 30.163
R68 VDD.n67 VDD.t63 30.163
R69 VDD.n58 VDD.t67 28.565
R70 VDD.n58 VDD.t45 28.565
R71 VDD.n53 VDD.t131 28.565
R72 VDD.n53 VDD.t91 28.565
R73 VDD.n54 VDD.t53 28.565
R74 VDD.n54 VDD.t11 28.565
R75 VDD.n56 VDD.t117 28.565
R76 VDD.n56 VDD.t97 28.565
R77 VDD.n6 VDD.t69 28.565
R78 VDD.n6 VDD.t115 28.565
R79 VDD.n1 VDD.t129 28.565
R80 VDD.n1 VDD.t109 28.565
R81 VDD.n2 VDD.t39 28.565
R82 VDD.n2 VDD.t75 28.565
R83 VDD.n4 VDD.t51 28.565
R84 VDD.n4 VDD.t143 28.565
R85 VDD.n14 VDD.t71 28.565
R86 VDD.n14 VDD.t83 28.565
R87 VDD.n9 VDD.t127 28.565
R88 VDD.n9 VDD.t101 28.565
R89 VDD.n10 VDD.t95 28.565
R90 VDD.n10 VDD.t89 28.565
R91 VDD.n12 VDD.t123 28.565
R92 VDD.n12 VDD.t17 28.565
R93 VDD.n22 VDD.t103 28.565
R94 VDD.n22 VDD.t119 28.565
R95 VDD.n17 VDD.t35 28.565
R96 VDD.n17 VDD.t33 28.565
R97 VDD.n18 VDD.t87 28.565
R98 VDD.n18 VDD.t141 28.565
R99 VDD.n20 VDD.t41 28.565
R100 VDD.n20 VDD.t65 28.565
R101 VDD.n30 VDD.t93 28.565
R102 VDD.n30 VDD.t7 28.565
R103 VDD.n25 VDD.t77 28.565
R104 VDD.n25 VDD.t137 28.565
R105 VDD.n26 VDD.t37 28.565
R106 VDD.n26 VDD.t49 28.565
R107 VDD.n28 VDD.t79 28.565
R108 VDD.n28 VDD.t121 28.565
R109 VDD.n50 VDD.t135 28.565
R110 VDD.n50 VDD.t19 28.565
R111 VDD.n45 VDD.t29 28.565
R112 VDD.n45 VDD.t27 28.565
R113 VDD.n46 VDD.t133 28.565
R114 VDD.n46 VDD.t99 28.565
R115 VDD.n48 VDD.t13 28.565
R116 VDD.n48 VDD.t3 28.565
R117 VDD.n42 VDD.t85 28.565
R118 VDD.n42 VDD.t73 28.565
R119 VDD.n37 VDD.t125 28.565
R120 VDD.n37 VDD.t113 28.565
R121 VDD.n38 VDD.t21 28.565
R122 VDD.n38 VDD.t107 28.565
R123 VDD.n40 VDD.t9 28.565
R124 VDD.n40 VDD.t57 28.565
R125 VDD.n66 VDD.t61 28.565
R126 VDD.n66 VDD.t59 28.565
R127 VDD.n61 VDD.t111 28.565
R128 VDD.n61 VDD.t15 28.565
R129 VDD.n62 VDD.t139 28.565
R130 VDD.n62 VDD.t5 28.565
R131 VDD.n64 VDD.t23 28.565
R132 VDD.n64 VDD.t25 28.565
R133 VDD.n52 VDD.t66 23.317
R134 VDD.n0 VDD.t68 23.317
R135 VDD.n8 VDD.t70 23.317
R136 VDD.n16 VDD.t102 23.317
R137 VDD.n24 VDD.t92 23.317
R138 VDD.n44 VDD.t134 23.317
R139 VDD.n36 VDD.t84 23.317
R140 VDD.n60 VDD.t60 23.317
R141 VDD.n60 VDD.t24 20.186
R142 VDD.n52 VDD.t96 20.183
R143 VDD.n0 VDD.t142 20.183
R144 VDD.n8 VDD.t16 20.183
R145 VDD.n16 VDD.t64 20.183
R146 VDD.n24 VDD.t120 20.183
R147 VDD.n44 VDD.t2 20.183
R148 VDD.n36 VDD.t56 20.183
R149 VDD.n55 VDD.n53 1.564
R150 VDD.n3 VDD.n1 1.564
R151 VDD.n11 VDD.n9 1.564
R152 VDD.n19 VDD.n17 1.564
R153 VDD.n27 VDD.n25 1.564
R154 VDD.n47 VDD.n45 1.564
R155 VDD.n39 VDD.n37 1.564
R156 VDD.n63 VDD.n61 1.564
R157 VDD.n57 VDD.n55 0.85
R158 VDD.n5 VDD.n3 0.85
R159 VDD.n13 VDD.n11 0.85
R160 VDD.n21 VDD.n19 0.85
R161 VDD.n29 VDD.n27 0.85
R162 VDD.n49 VDD.n47 0.85
R163 VDD.n41 VDD.n39 0.85
R164 VDD.n65 VDD.n63 0.85
R165 VDD.n59 VDD.n58 0.747
R166 VDD.n55 VDD.n54 0.747
R167 VDD.n57 VDD.n56 0.747
R168 VDD.n7 VDD.n6 0.747
R169 VDD.n3 VDD.n2 0.747
R170 VDD.n5 VDD.n4 0.747
R171 VDD.n15 VDD.n14 0.747
R172 VDD.n11 VDD.n10 0.747
R173 VDD.n13 VDD.n12 0.747
R174 VDD.n23 VDD.n22 0.747
R175 VDD.n19 VDD.n18 0.747
R176 VDD.n21 VDD.n20 0.747
R177 VDD.n31 VDD.n30 0.747
R178 VDD.n27 VDD.n26 0.747
R179 VDD.n29 VDD.n28 0.747
R180 VDD.n51 VDD.n50 0.747
R181 VDD.n47 VDD.n46 0.747
R182 VDD.n49 VDD.n48 0.747
R183 VDD.n43 VDD.n42 0.747
R184 VDD.n39 VDD.n38 0.747
R185 VDD.n41 VDD.n40 0.747
R186 VDD.n67 VDD.n66 0.747
R187 VDD.n63 VDD.n62 0.747
R188 VDD.n65 VDD.n64 0.747
R189 VDD.n70 VDD.n69 0.446
R190 VDD.n34 VDD.n33 0.446
R191 VDD.n69 VDD.n68 0.431
R192 VDD.n71 VDD.n70 0.431
R193 VDD.n33 VDD.n32 0.431
R194 VDD.n35 VDD.n34 0.431
R195 VDD VDD.n71 0.223
R196 VDD.n69 VDD.n59 0.208
R197 VDD.n35 VDD.n7 0.208
R198 VDD.n34 VDD.n15 0.208
R199 VDD.n33 VDD.n23 0.208
R200 VDD.n32 VDD.n31 0.208
R201 VDD.n70 VDD.n51 0.208
R202 VDD.n71 VDD.n43 0.208
R203 VDD.n68 VDD.n67 0.208
R204 VDD VDD.n35 0.198
R205 VDD.n69 VDD.n57 0.195
R206 VDD.n35 VDD.n5 0.195
R207 VDD.n34 VDD.n13 0.195
R208 VDD.n33 VDD.n21 0.195
R209 VDD.n32 VDD.n29 0.195
R210 VDD.n70 VDD.n49 0.195
R211 VDD.n71 VDD.n41 0.195
R212 VDD.n68 VDD.n65 0.195
R213 VDD.n68 VDD.n60 0.001
R214 VDD.n69 VDD.n52 0.001
R215 VDD.n35 VDD.n0 0.001
R216 VDD.n34 VDD.n8 0.001
R217 VDD.n33 VDD.n16 0.001
R218 VDD.n32 VDD.n24 0.001
R219 VDD.n70 VDD.n44 0.001
R220 VDD.n71 VDD.n36 0.001
R221 a_155_68.n4 a_155_68.t10 214.335
R222 a_155_68.t7 a_155_68.n4 214.335
R223 a_155_68.n5 a_155_68.t7 143.851
R224 a_155_68.n5 a_155_68.t9 135.658
R225 a_155_68.n4 a_155_68.t8 80.333
R226 a_155_68.n0 a_155_68.t3 28.565
R227 a_155_68.n0 a_155_68.t5 28.565
R228 a_155_68.n2 a_155_68.t2 28.565
R229 a_155_68.n2 a_155_68.t4 28.565
R230 a_155_68.t0 a_155_68.n7 28.565
R231 a_155_68.n7 a_155_68.t1 28.565
R232 a_155_68.n1 a_155_68.t6 9.714
R233 a_155_68.n1 a_155_68.n0 1.003
R234 a_155_68.n6 a_155_68.n3 0.833
R235 a_155_68.n3 a_155_68.n2 0.653
R236 a_155_68.n7 a_155_68.n6 0.653
R237 a_155_68.n3 a_155_68.n1 0.341
R238 a_155_68.n6 a_155_68.n5 0.032
R239 B[0].t1 B[0].t2 415.315
R240 B[0] B[0].t1 217.493
R241 B[0].n0 B[0].t0 214.335
R242 B[0].t2 B[0].n0 214.335
R243 B[0].n0 B[0].t3 80.333
R244 B[5].t1 B[5].t3 415.315
R245 B[5] B[5].t1 217.491
R246 B[5].n0 B[5].t0 214.335
R247 B[5].t3 B[5].n0 214.335
R248 B[5].n0 B[5].t2 80.333
R249 a_7517_68.n2 a_7517_68.t9 214.335
R250 a_7517_68.t7 a_7517_68.n2 214.335
R251 a_7517_68.n3 a_7517_68.t7 143.851
R252 a_7517_68.n3 a_7517_68.t10 135.658
R253 a_7517_68.n2 a_7517_68.t8 80.333
R254 a_7517_68.n4 a_7517_68.t4 28.565
R255 a_7517_68.n4 a_7517_68.t3 28.565
R256 a_7517_68.n0 a_7517_68.t1 28.565
R257 a_7517_68.n0 a_7517_68.t5 28.565
R258 a_7517_68.n7 a_7517_68.t2 28.565
R259 a_7517_68.t0 a_7517_68.n7 28.565
R260 a_7517_68.n1 a_7517_68.t6 9.714
R261 a_7517_68.n1 a_7517_68.n0 1.003
R262 a_7517_68.n6 a_7517_68.n5 0.833
R263 a_7517_68.n5 a_7517_68.n4 0.653
R264 a_7517_68.n7 a_7517_68.n6 0.653
R265 a_7517_68.n6 a_7517_68.n1 0.341
R266 a_7517_68.n5 a_7517_68.n3 0.032
R267 B[7].t2 B[7].t3 415.315
R268 B[7] B[7].t2 217.493
R269 B[7].n0 B[7].t1 214.335
R270 B[7].t3 B[7].n0 214.335
R271 B[7].n0 B[7].t0 80.333
R272 a_10463_70.n0 a_10463_70.t8 214.335
R273 a_10463_70.t9 a_10463_70.n0 214.335
R274 a_10463_70.n1 a_10463_70.t9 143.851
R275 a_10463_70.n1 a_10463_70.t10 135.658
R276 a_10463_70.n0 a_10463_70.t7 80.333
R277 a_10463_70.n2 a_10463_70.t4 28.565
R278 a_10463_70.n2 a_10463_70.t5 28.565
R279 a_10463_70.n4 a_10463_70.t3 28.565
R280 a_10463_70.n4 a_10463_70.t6 28.565
R281 a_10463_70.t0 a_10463_70.n7 28.565
R282 a_10463_70.n7 a_10463_70.t1 28.565
R283 a_10463_70.n6 a_10463_70.t2 9.714
R284 a_10463_70.n7 a_10463_70.n6 1.003
R285 a_10463_70.n5 a_10463_70.n3 0.833
R286 a_10463_70.n3 a_10463_70.n2 0.653
R287 a_10463_70.n5 a_10463_70.n4 0.653
R288 a_10463_70.n6 a_10463_70.n5 0.341
R289 a_10463_70.n3 a_10463_70.n1 0.032
R290 A[7].t1 A[7].t2 437.233
R291 A[7] A[7].t1 216.696
R292 A[7].n0 A[7].t3 214.686
R293 A[7].t2 A[7].n0 214.686
R294 A[7].n0 A[7].t0 80.333
R295 A[3].t2 A[3].t0 437.233
R296 A[3] A[3].t2 216.696
R297 A[3].n0 A[3].t1 214.686
R298 A[3].t0 A[3].n0 214.686
R299 A[3].n0 A[3].t3 80.333
R300 a_4549_70.n4 a_4549_70.t10 214.335
R301 a_4549_70.t7 a_4549_70.n4 214.335
R302 a_4549_70.n5 a_4549_70.t7 143.851
R303 a_4549_70.n5 a_4549_70.t9 135.658
R304 a_4549_70.n4 a_4549_70.t8 80.333
R305 a_4549_70.n0 a_4549_70.t3 28.565
R306 a_4549_70.n0 a_4549_70.t4 28.565
R307 a_4549_70.n2 a_4549_70.t1 28.565
R308 a_4549_70.n2 a_4549_70.t5 28.565
R309 a_4549_70.n7 a_4549_70.t6 28.565
R310 a_4549_70.t0 a_4549_70.n7 28.565
R311 a_4549_70.n1 a_4549_70.t2 9.714
R312 a_4549_70.n1 a_4549_70.n0 1.003
R313 a_4549_70.n6 a_4549_70.n3 0.833
R314 a_4549_70.n3 a_4549_70.n2 0.653
R315 a_4549_70.n7 a_4549_70.n6 0.653
R316 a_4549_70.n3 a_4549_70.n1 0.341
R317 a_4549_70.n6 a_4549_70.n5 0.032
R318 Y[0].n1 Y[0].n0 192.754
R319 Y[0].n1 Y[0].t0 28.568
R320 Y[0].n0 Y[0].t1 28.565
R321 Y[0].n0 Y[0].t2 28.565
R322 Y[0].n2 Y[0].t3 18.726
R323 Y[0].n2 Y[0].n1 1.123
R324 Y[0] Y[0].n2 0.009
R325 A[1].t1 A[1].t2 437.233
R326 A[1] A[1].t1 216.694
R327 A[1].n0 A[1].t3 214.686
R328 A[1].t2 A[1].n0 214.686
R329 A[1].n0 A[1].t0 80.333
R330 a_1603_68.n4 a_1603_68.t9 214.335
R331 a_1603_68.t10 a_1603_68.n4 214.335
R332 a_1603_68.n5 a_1603_68.t10 143.851
R333 a_1603_68.n5 a_1603_68.t7 135.658
R334 a_1603_68.n4 a_1603_68.t8 80.333
R335 a_1603_68.n0 a_1603_68.t5 28.565
R336 a_1603_68.n0 a_1603_68.t3 28.565
R337 a_1603_68.n2 a_1603_68.t1 28.565
R338 a_1603_68.n2 a_1603_68.t4 28.565
R339 a_1603_68.t0 a_1603_68.n7 28.565
R340 a_1603_68.n7 a_1603_68.t2 28.565
R341 a_1603_68.n1 a_1603_68.t6 9.714
R342 a_1603_68.n1 a_1603_68.n0 1.003
R343 a_1603_68.n6 a_1603_68.n3 0.833
R344 a_1603_68.n3 a_1603_68.n2 0.653
R345 a_1603_68.n7 a_1603_68.n6 0.653
R346 a_1603_68.n3 a_1603_68.n1 0.341
R347 a_1603_68.n6 a_1603_68.n5 0.032
R348 B[4].t3 B[4].t1 415.315
R349 B[4] B[4].t3 217.493
R350 B[4].n0 B[4].t0 214.335
R351 B[4].t1 B[4].n0 214.335
R352 B[4].n0 B[4].t2 80.333
R353 a_6069_68.n2 a_6069_68.t10 214.335
R354 a_6069_68.t7 a_6069_68.n2 214.335
R355 a_6069_68.n3 a_6069_68.t7 143.851
R356 a_6069_68.n3 a_6069_68.t9 135.658
R357 a_6069_68.n2 a_6069_68.t8 80.333
R358 a_6069_68.n4 a_6069_68.t2 28.565
R359 a_6069_68.n4 a_6069_68.t0 28.565
R360 a_6069_68.n0 a_6069_68.t6 28.565
R361 a_6069_68.n0 a_6069_68.t4 28.565
R362 a_6069_68.n7 a_6069_68.t1 28.565
R363 a_6069_68.t3 a_6069_68.n7 28.565
R364 a_6069_68.n1 a_6069_68.t5 9.714
R365 a_6069_68.n1 a_6069_68.n0 1.003
R366 a_6069_68.n6 a_6069_68.n5 0.833
R367 a_6069_68.n5 a_6069_68.n4 0.653
R368 a_6069_68.n7 a_6069_68.n6 0.653
R369 a_6069_68.n6 a_6069_68.n1 0.341
R370 a_6069_68.n5 a_6069_68.n3 0.032
R371 B[6].t1 B[6].t0 415.315
R372 B[6] B[6].t1 217.493
R373 B[6].n0 B[6].t3 214.335
R374 B[6].t0 B[6].n0 214.335
R375 B[6].n0 B[6].t2 80.333
R376 a_9015_70.n0 a_9015_70.t8 214.335
R377 a_9015_70.t9 a_9015_70.n0 214.335
R378 a_9015_70.n1 a_9015_70.t9 143.851
R379 a_9015_70.n1 a_9015_70.t7 135.658
R380 a_9015_70.n0 a_9015_70.t10 80.333
R381 a_9015_70.n2 a_9015_70.t2 28.565
R382 a_9015_70.n2 a_9015_70.t3 28.565
R383 a_9015_70.n4 a_9015_70.t4 28.565
R384 a_9015_70.n4 a_9015_70.t5 28.565
R385 a_9015_70.n7 a_9015_70.t6 28.565
R386 a_9015_70.t0 a_9015_70.n7 28.565
R387 a_9015_70.n6 a_9015_70.t1 9.714
R388 a_9015_70.n7 a_9015_70.n6 1.003
R389 a_9015_70.n5 a_9015_70.n3 0.833
R390 a_9015_70.n3 a_9015_70.n2 0.653
R391 a_9015_70.n5 a_9015_70.n4 0.653
R392 a_9015_70.n6 a_9015_70.n5 0.341
R393 a_9015_70.n3 a_9015_70.n1 0.032
R394 A[2].t0 A[2].t2 437.233
R395 A[2] A[2].t0 216.699
R396 A[2].n0 A[2].t3 214.686
R397 A[2].t2 A[2].n0 214.686
R398 A[2].n0 A[2].t1 80.333
R399 a_3101_70.n2 a_3101_70.t10 214.335
R400 a_3101_70.t7 a_3101_70.n2 214.335
R401 a_3101_70.n3 a_3101_70.t7 143.851
R402 a_3101_70.n3 a_3101_70.t8 135.658
R403 a_3101_70.n2 a_3101_70.t9 80.333
R404 a_3101_70.n4 a_3101_70.t6 28.565
R405 a_3101_70.n4 a_3101_70.t1 28.565
R406 a_3101_70.n0 a_3101_70.t5 28.565
R407 a_3101_70.n0 a_3101_70.t3 28.565
R408 a_3101_70.t0 a_3101_70.n7 28.565
R409 a_3101_70.n7 a_3101_70.t4 28.565
R410 a_3101_70.n1 a_3101_70.t2 9.714
R411 a_3101_70.n1 a_3101_70.n0 1.003
R412 a_3101_70.n6 a_3101_70.n5 0.833
R413 a_3101_70.n5 a_3101_70.n4 0.653
R414 a_3101_70.n7 a_3101_70.n6 0.653
R415 a_3101_70.n6 a_3101_70.n1 0.341
R416 a_3101_70.n5 a_3101_70.n3 0.032
R417 a_3338_n567.t0 a_3338_n567.t1 17.4
R418 VSS.n5 VSS.t8 18.178
R419 VSS.n3 VSS.t12 18.178
R420 VSS.n12 VSS.t13 18.178
R421 VSS.n10 VSS.t15 18.178
R422 VSS.n8 VSS.t0 18.178
R423 VSS.n7 VSS.t10 18.178
R424 VSS.n1 VSS.t1 18.178
R425 VSS.n0 VSS.t3 18.178
R426 VSS.n5 VSS.t2 9.319
R427 VSS.n3 VSS.t6 9.319
R428 VSS.n12 VSS.t9 9.319
R429 VSS.n10 VSS.t4 9.319
R430 VSS.n8 VSS.t11 9.319
R431 VSS.n7 VSS.t14 9.319
R432 VSS.n1 VSS.t5 9.319
R433 VSS.n0 VSS.t7 9.319
R434 VSS.n9 VSS.n7 0.815
R435 VSS.n2 VSS.n0 0.813
R436 VSS.n11 VSS.n9 0.524
R437 VSS.n4 VSS.n2 0.524
R438 VSS.n6 VSS.n4 0.507
R439 VSS.n13 VSS.n11 0.505
R440 VSS VSS.n6 0.329
R441 VSS.n6 VSS.n5 0.309
R442 VSS.n4 VSS.n3 0.309
R443 VSS.n13 VSS.n12 0.309
R444 VSS.n11 VSS.n10 0.309
R445 VSS.n9 VSS.n8 0.309
R446 VSS.n2 VSS.n1 0.309
R447 VSS VSS.n13 0.162
R448 Y[6].n1 Y[6].n0 192.754
R449 Y[6].n1 Y[6].t2 28.568
R450 Y[6].n0 Y[6].t0 28.565
R451 Y[6].n0 Y[6].t1 28.565
R452 Y[6].n2 Y[6].t3 18.726
R453 Y[6].n2 Y[6].n1 1.123
R454 Y[6] Y[6].n2 0.016
R455 A[4].t2 A[4].t0 437.233
R456 A[4] A[4].t2 216.701
R457 A[4].n0 A[4].t1 214.686
R458 A[4].t0 A[4].n0 214.686
R459 A[4].n0 A[4].t3 80.333
R460 Y[5].n1 Y[5].n0 192.754
R461 Y[5].n1 Y[5].t0 28.568
R462 Y[5].n0 Y[5].t1 28.565
R463 Y[5].n0 Y[5].t2 28.565
R464 Y[5].n2 Y[5].t3 18.726
R465 Y[5].n2 Y[5].n1 1.123
R466 Y[5] Y[5].n2 0.004
R467 a_9252_n567.t0 a_9252_n567.t1 17.4
R468 Y[7].n1 Y[7].n0 192.754
R469 Y[7].n1 Y[7].t1 28.568
R470 Y[7].n0 Y[7].t2 28.565
R471 Y[7].n0 Y[7].t0 28.565
R472 Y[7].n2 Y[7].t3 18.726
R473 Y[7].n2 Y[7].n1 1.123
R474 Y[7] Y[7].n2 0.009
R475 B[3].t3 B[3].t0 415.315
R476 B[3] B[3].t3 217.491
R477 B[3].n0 B[3].t1 214.335
R478 B[3].t0 B[3].n0 214.335
R479 B[3].n0 B[3].t2 80.333
R480 Y[4].n1 Y[4].n0 192.754
R481 Y[4].n1 Y[4].t0 28.568
R482 Y[4].n0 Y[4].t1 28.565
R483 Y[4].n0 Y[4].t2 28.565
R484 Y[4].n2 Y[4].t3 18.726
R485 Y[4].n2 Y[4].n1 1.123
R486 Y[4] Y[4].n2 0.002
R487 Y[1].n1 Y[1].n0 192.754
R488 Y[1].n1 Y[1].t1 28.568
R489 Y[1].n0 Y[1].t2 28.565
R490 Y[1].n0 Y[1].t0 28.565
R491 Y[1].n2 Y[1].t3 18.726
R492 Y[1].n2 Y[1].n1 1.123
R493 Y[1] Y[1].n2 0.004
R494 a_10700_n567.t0 a_10700_n567.t1 17.4
R495 B[1].t3 B[1].t2 415.315
R496 B[1] B[1].t3 217.493
R497 B[1].n0 B[1].t1 214.335
R498 B[1].t2 B[1].n0 214.335
R499 B[1].n0 B[1].t0 80.333
R500 a_7754_n569.t0 a_7754_n569.t1 17.4
R501 A[6].t2 A[6].t1 437.233
R502 A[6] A[6].t2 216.696
R503 A[6].n0 A[6].t3 214.686
R504 A[6].t1 A[6].n0 214.686
R505 A[6].n0 A[6].t0 80.333
R506 A[5].t3 A[5].t2 437.233
R507 A[5] A[5].t3 216.706
R508 A[5].n0 A[5].t0 214.686
R509 A[5].t2 A[5].n0 214.686
R510 A[5].n0 A[5].t1 80.333
R511 Y[3].n1 Y[3].n0 192.754
R512 Y[3].n1 Y[3].t0 28.568
R513 Y[3].n0 Y[3].t1 28.565
R514 Y[3].n0 Y[3].t2 28.565
R515 Y[3].n2 Y[3].t3 18.726
R516 Y[3].n2 Y[3].n1 1.123
R517 Y[3] Y[3].n2 0.007
R518 a_4786_n567.t0 a_4786_n567.t1 17.4
R519 a_1840_n569.t0 a_1840_n569.t1 17.4
R520 Y[2].n1 Y[2].n0 192.754
R521 Y[2].n1 Y[2].t0 28.568
R522 Y[2].n0 Y[2].t1 28.565
R523 Y[2].n0 Y[2].t2 28.565
R524 Y[2].n2 Y[2].t3 18.726
R525 Y[2].n2 Y[2].n1 1.123
R526 Y[2] Y[2].n2 0.004
R527 a_392_n569.t0 a_392_n569.t1 17.4
R528 a_6306_n569.t0 a_6306_n569.t1 17.4
R529 B[2].t2 B[2].t0 415.315
R530 B[2] B[2].t2 217.488
R531 B[2].n0 B[2].t3 214.335
R532 B[2].t0 B[2].n0 214.335
R533 B[2].n0 B[2].t1 80.333
C0 A[1] A[0] 0.00fF
C1 Y[5] B[4] 0.00fF
C2 A[1] B[0] 0.00fF
C3 B[3] B[2] 0.00fF
C4 Y[2] B[2] 0.01fF
C5 A[1] VDD 0.18fF
C6 A[6] B[6] 0.80fF
C7 VDD A[6] 0.18fF
C8 A[7] Y[6] 0.02fF
C9 Y[1] B[1] 0.01fF
C10 B[0] A[0] 0.80fF
C11 VDD A[0] 0.16fF
C12 Y[6] Y[7] 0.01fF
C13 A[3] B[2] 0.00fF
C14 B[0] VDD 0.19fF
C15 A[2] B[2] 0.80fF
C16 VDD B[6] 0.19fF
C17 A[4] VDD 0.18fF
C18 Y[5] A[5] 0.01fF
C19 Y[4] B[5] 0.01fF
C20 Y[0] B[1] 0.01fF
C21 Y[4] Y[3] 0.00fF
C22 VDD B[4] 0.19fF
C23 A[4] B[4] 0.80fF
C24 A[7] A[6] 0.00fF
C25 Y[1] Y[0] 0.01fF
C26 A[1] B[2] 0.00fF
C27 A[5] A[6] 0.00fF
C28 Y[3] B[3] 0.01fF
C29 Y[2] Y[3] 0.01fF
C30 A[7] B[6] 0.00fF
C31 A[7] VDD 0.17fF
C32 Y[7] B[6] 0.00fF
C33 VDD Y[7] 0.69fF
C34 Y[3] A[3] 0.01fF
C35 Y[2] Y[1] 0.00fF
C36 A[5] B[6] 0.00fF
C37 A[2] B[1] 0.00fF
C38 VDD A[5] 0.18fF
C39 VDD B[2] 0.19fF
C40 Y[5] B[5] 0.01fF
C41 A[4] A[5] 0.00fF
C42 B[7] Y[6] 0.01fF
C43 Y[1] A[2] 0.02fF
C44 A[5] B[4] 0.00fF
C45 B[5] A[6] 0.00fF
C46 A[7] Y[7] 0.01fF
C47 B[1] A[1] 0.80fF
C48 B[1] A[0] 0.00fF
C49 Y[2] B[3] 0.01fF
C50 B[5] B[6] 0.00fF
C51 VDD B[5] 0.19fF
C52 B[1] B[0] 0.00fF
C53 A[4] B[5] 0.00fF
C54 Y[1] A[1] 0.01fF
C55 B[1] VDD 0.19fF
C56 Y[5] Y[4] 0.01fF
C57 B[7] A[6] 0.00fF
C58 Y[3] VDD 0.76fF
C59 Y[2] A[3] 0.02fF
C60 B[3] A[3] 0.80fF
C61 A[4] Y[3] 0.02fF
C62 Y[2] A[2] 0.01fF
C63 B[3] A[2] 0.00fF
C64 Y[1] B[0] 0.00fF
C65 B[5] B[4] 0.00fF
C66 Y[1] VDD 0.78fF
C67 B[7] B[6] 0.00fF
C68 B[7] VDD 0.18fF
C69 A[3] A[2] 0.00fF
C70 Y[3] B[4] 0.01fF
C71 Y[0] A[1] 0.02fF
C72 Y[5] Y[6] 0.00fF
C73 Y[0] A[0] 0.01fF
C74 Y[0] B[0] 0.01fF
C75 B[5] A[5] 0.80fF
C76 Y[0] VDD 0.78fF
C77 Y[4] VDD 0.78fF
C78 Y[4] A[4] 0.01fF
C79 B[1] B[2] 0.00fF
C80 Y[3] B[2] 0.00fF
C81 B[7] A[7] 0.80fF
C82 B[7] Y[7] 0.01fF
C83 A[2] A[1] 0.00fF
C84 B[3] VDD 0.19fF
C85 Y[2] VDD 0.78fF
C86 Y[6] A[6] 0.01fF
C87 Y[4] B[4] 0.01fF
C88 A[4] B[3] 0.00fF
C89 Y[1] B[2] 0.01fF
C90 Y[5] A[6] 0.02fF
C91 A[3] VDD 0.18fF
C92 Y[6] B[6] 0.01fF
C93 Y[6] VDD 0.78fF
C94 A[2] VDD 0.18fF
C95 A[4] A[3] 0.00fF
C96 B[3] B[4] 0.00fF
C97 Y[5] B[6] 0.01fF
C98 Y[5] VDD 0.78fF
C99 A[3] B[4] 0.00fF
C100 Y[4] A[5] 0.02fF
.ends

