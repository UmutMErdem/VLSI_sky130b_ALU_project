magic
tech sky130B
magscale 1 2
timestamp 1735737881
<< nwell >>
rect 2563 677 2791 1167
rect 359 477 1197 677
rect 2257 477 3095 677
rect -125 153 3578 477
rect 302 -540 1140 153
rect 2200 -540 3038 153
<< nmos >>
rect 94 -1010 154 -810
rect 514 -1210 574 -810
rect 632 -1210 692 -810
rect 750 -1210 810 -810
rect 868 -1210 928 -810
rect 1392 -1010 1452 -810
rect 1992 -1010 2052 -810
rect 2412 -1210 2472 -810
rect 2530 -1210 2590 -810
rect 2648 -1210 2708 -810
rect 2766 -1210 2826 -810
rect 3290 -1010 3350 -810
<< pmos >>
rect -31 215 29 415
rect 87 215 147 415
rect 205 215 265 415
rect 453 215 513 615
rect 571 215 631 615
rect 689 215 749 615
rect 807 215 867 615
rect 925 215 985 615
rect 1043 215 1103 615
rect 1290 215 1350 415
rect 1408 215 1468 415
rect 1526 215 1586 415
rect 1867 215 1927 415
rect 1985 215 2045 415
rect 2103 215 2163 415
rect 2351 215 2411 615
rect 2469 215 2529 615
rect 2587 215 2647 615
rect 2705 215 2765 615
rect 2823 215 2883 615
rect 2941 215 3001 615
rect 3188 215 3248 415
rect 3306 215 3366 415
rect 3424 215 3484 415
rect 396 -478 456 -78
rect 514 -478 574 -78
rect 632 -478 692 -78
rect 750 -478 810 -78
rect 868 -478 928 -78
rect 986 -478 1046 -78
rect 2294 -478 2354 -78
rect 2412 -478 2472 -78
rect 2530 -478 2590 -78
rect 2648 -478 2708 -78
rect 2766 -478 2826 -78
rect 2884 -478 2944 -78
<< ndiff >>
rect 36 -822 94 -810
rect 36 -998 48 -822
rect 82 -998 94 -822
rect 36 -1010 94 -998
rect 154 -822 212 -810
rect 154 -998 166 -822
rect 200 -998 212 -822
rect 154 -1010 212 -998
rect 456 -822 514 -810
rect 456 -1198 468 -822
rect 502 -1198 514 -822
rect 456 -1210 514 -1198
rect 574 -822 632 -810
rect 574 -1198 586 -822
rect 620 -1198 632 -822
rect 574 -1210 632 -1198
rect 692 -822 750 -810
rect 692 -1198 704 -822
rect 738 -1198 750 -822
rect 692 -1210 750 -1198
rect 810 -822 868 -810
rect 810 -1198 822 -822
rect 856 -1198 868 -822
rect 810 -1210 868 -1198
rect 928 -822 986 -810
rect 928 -1198 940 -822
rect 974 -1198 986 -822
rect 1334 -822 1392 -810
rect 1334 -998 1346 -822
rect 1380 -998 1392 -822
rect 1334 -1010 1392 -998
rect 1452 -822 1510 -810
rect 1452 -998 1464 -822
rect 1498 -998 1510 -822
rect 1452 -1010 1510 -998
rect 1934 -822 1992 -810
rect 1934 -998 1946 -822
rect 1980 -998 1992 -822
rect 1934 -1010 1992 -998
rect 2052 -822 2110 -810
rect 2052 -998 2064 -822
rect 2098 -998 2110 -822
rect 2052 -1010 2110 -998
rect 2354 -822 2412 -810
rect 928 -1210 986 -1198
rect 2354 -1198 2366 -822
rect 2400 -1198 2412 -822
rect 2354 -1210 2412 -1198
rect 2472 -822 2530 -810
rect 2472 -1198 2484 -822
rect 2518 -1198 2530 -822
rect 2472 -1210 2530 -1198
rect 2590 -822 2648 -810
rect 2590 -1198 2602 -822
rect 2636 -1198 2648 -822
rect 2590 -1210 2648 -1198
rect 2708 -822 2766 -810
rect 2708 -1198 2720 -822
rect 2754 -1198 2766 -822
rect 2708 -1210 2766 -1198
rect 2826 -822 2884 -810
rect 2826 -1198 2838 -822
rect 2872 -1198 2884 -822
rect 3232 -822 3290 -810
rect 3232 -998 3244 -822
rect 3278 -998 3290 -822
rect 3232 -1010 3290 -998
rect 3350 -822 3408 -810
rect 3350 -998 3362 -822
rect 3396 -998 3408 -822
rect 3350 -1010 3408 -998
rect 2826 -1210 2884 -1198
<< pdiff >>
rect 395 603 453 615
rect -89 403 -31 415
rect -89 227 -77 403
rect -43 227 -31 403
rect -89 215 -31 227
rect 29 403 87 415
rect 29 227 41 403
rect 75 227 87 403
rect 29 215 87 227
rect 147 403 205 415
rect 147 227 159 403
rect 193 227 205 403
rect 147 215 205 227
rect 265 403 323 415
rect 265 227 277 403
rect 311 227 323 403
rect 265 215 323 227
rect 395 227 407 603
rect 441 227 453 603
rect 395 215 453 227
rect 513 603 571 615
rect 513 227 525 603
rect 559 227 571 603
rect 513 215 571 227
rect 631 603 689 615
rect 631 227 643 603
rect 677 227 689 603
rect 631 215 689 227
rect 749 603 807 615
rect 749 227 761 603
rect 795 227 807 603
rect 749 215 807 227
rect 867 603 925 615
rect 867 227 879 603
rect 913 227 925 603
rect 867 215 925 227
rect 985 603 1043 615
rect 985 227 997 603
rect 1031 227 1043 603
rect 985 215 1043 227
rect 1103 603 1161 615
rect 1103 227 1115 603
rect 1149 227 1161 603
rect 2293 603 2351 615
rect 1103 215 1161 227
rect 1232 403 1290 415
rect 1232 227 1244 403
rect 1278 227 1290 403
rect 1232 215 1290 227
rect 1350 403 1408 415
rect 1350 227 1362 403
rect 1396 227 1408 403
rect 1350 215 1408 227
rect 1468 403 1526 415
rect 1468 227 1480 403
rect 1514 227 1526 403
rect 1468 215 1526 227
rect 1586 403 1644 415
rect 1586 227 1598 403
rect 1632 227 1644 403
rect 1586 215 1644 227
rect 1809 403 1867 415
rect 1809 227 1821 403
rect 1855 227 1867 403
rect 1809 215 1867 227
rect 1927 403 1985 415
rect 1927 227 1939 403
rect 1973 227 1985 403
rect 1927 215 1985 227
rect 2045 403 2103 415
rect 2045 227 2057 403
rect 2091 227 2103 403
rect 2045 215 2103 227
rect 2163 403 2221 415
rect 2163 227 2175 403
rect 2209 227 2221 403
rect 2163 215 2221 227
rect 2293 227 2305 603
rect 2339 227 2351 603
rect 2293 215 2351 227
rect 2411 603 2469 615
rect 2411 227 2423 603
rect 2457 227 2469 603
rect 2411 215 2469 227
rect 2529 603 2587 615
rect 2529 227 2541 603
rect 2575 227 2587 603
rect 2529 215 2587 227
rect 2647 603 2705 615
rect 2647 227 2659 603
rect 2693 227 2705 603
rect 2647 215 2705 227
rect 2765 603 2823 615
rect 2765 227 2777 603
rect 2811 227 2823 603
rect 2765 215 2823 227
rect 2883 603 2941 615
rect 2883 227 2895 603
rect 2929 227 2941 603
rect 2883 215 2941 227
rect 3001 603 3059 615
rect 3001 227 3013 603
rect 3047 227 3059 603
rect 3001 215 3059 227
rect 3130 403 3188 415
rect 3130 227 3142 403
rect 3176 227 3188 403
rect 3130 215 3188 227
rect 3248 403 3306 415
rect 3248 227 3260 403
rect 3294 227 3306 403
rect 3248 215 3306 227
rect 3366 403 3424 415
rect 3366 227 3378 403
rect 3412 227 3424 403
rect 3366 215 3424 227
rect 3484 403 3542 415
rect 3484 227 3496 403
rect 3530 227 3542 403
rect 3484 215 3542 227
rect 338 -90 396 -78
rect 338 -466 350 -90
rect 384 -466 396 -90
rect 338 -478 396 -466
rect 456 -90 514 -78
rect 456 -466 468 -90
rect 502 -466 514 -90
rect 456 -478 514 -466
rect 574 -90 632 -78
rect 574 -466 586 -90
rect 620 -466 632 -90
rect 574 -478 632 -466
rect 692 -90 750 -78
rect 692 -466 704 -90
rect 738 -466 750 -90
rect 692 -478 750 -466
rect 810 -90 868 -78
rect 810 -466 822 -90
rect 856 -466 868 -90
rect 810 -478 868 -466
rect 928 -90 986 -78
rect 928 -466 940 -90
rect 974 -466 986 -90
rect 928 -478 986 -466
rect 1046 -90 1104 -78
rect 1046 -466 1058 -90
rect 1092 -466 1104 -90
rect 1046 -478 1104 -466
rect 2236 -90 2294 -78
rect 2236 -466 2248 -90
rect 2282 -466 2294 -90
rect 2236 -478 2294 -466
rect 2354 -90 2412 -78
rect 2354 -466 2366 -90
rect 2400 -466 2412 -90
rect 2354 -478 2412 -466
rect 2472 -90 2530 -78
rect 2472 -466 2484 -90
rect 2518 -466 2530 -90
rect 2472 -478 2530 -466
rect 2590 -90 2648 -78
rect 2590 -466 2602 -90
rect 2636 -466 2648 -90
rect 2590 -478 2648 -466
rect 2708 -90 2766 -78
rect 2708 -466 2720 -90
rect 2754 -466 2766 -90
rect 2708 -478 2766 -466
rect 2826 -90 2884 -78
rect 2826 -466 2838 -90
rect 2872 -466 2884 -90
rect 2826 -478 2884 -466
rect 2944 -90 3002 -78
rect 2944 -466 2956 -90
rect 2990 -466 3002 -90
rect 2944 -478 3002 -466
<< ndiffc >>
rect 48 -998 82 -822
rect 166 -998 200 -822
rect 468 -1198 502 -822
rect 586 -1198 620 -822
rect 704 -1198 738 -822
rect 822 -1198 856 -822
rect 940 -1198 974 -822
rect 1346 -998 1380 -822
rect 1464 -998 1498 -822
rect 1946 -998 1980 -822
rect 2064 -998 2098 -822
rect 2366 -1198 2400 -822
rect 2484 -1198 2518 -822
rect 2602 -1198 2636 -822
rect 2720 -1198 2754 -822
rect 2838 -1198 2872 -822
rect 3244 -998 3278 -822
rect 3362 -998 3396 -822
<< pdiffc >>
rect -77 227 -43 403
rect 41 227 75 403
rect 159 227 193 403
rect 277 227 311 403
rect 407 227 441 603
rect 525 227 559 603
rect 643 227 677 603
rect 761 227 795 603
rect 879 227 913 603
rect 997 227 1031 603
rect 1115 227 1149 603
rect 1244 227 1278 403
rect 1362 227 1396 403
rect 1480 227 1514 403
rect 1598 227 1632 403
rect 1821 227 1855 403
rect 1939 227 1973 403
rect 2057 227 2091 403
rect 2175 227 2209 403
rect 2305 227 2339 603
rect 2423 227 2457 603
rect 2541 227 2575 603
rect 2659 227 2693 603
rect 2777 227 2811 603
rect 2895 227 2929 603
rect 3013 227 3047 603
rect 3142 227 3176 403
rect 3260 227 3294 403
rect 3378 227 3412 403
rect 3496 227 3530 403
rect 350 -466 384 -90
rect 468 -466 502 -90
rect 586 -466 620 -90
rect 704 -466 738 -90
rect 822 -466 856 -90
rect 940 -466 974 -90
rect 1058 -466 1092 -90
rect 2248 -466 2282 -90
rect 2366 -466 2400 -90
rect 2484 -466 2518 -90
rect 2602 -466 2636 -90
rect 2720 -466 2754 -90
rect 2838 -466 2872 -90
rect 2956 -466 2990 -90
<< psubdiff >>
rect 647 -1507 802 -1461
rect 647 -1670 678 -1507
rect 768 -1670 802 -1507
rect 647 -1695 802 -1670
<< nsubdiff >>
rect 2601 1091 2754 1131
rect 2601 942 2644 1091
rect 2711 942 2754 1091
rect 2601 873 2754 942
<< psubdiffcont >>
rect 678 -1670 768 -1507
<< nsubdiffcont >>
rect 2644 942 2711 1091
<< poly >>
rect 453 630 749 681
rect 453 615 513 630
rect 571 615 631 630
rect 689 615 749 630
rect 807 615 867 641
rect 925 615 985 641
rect 1043 615 1103 641
rect 2351 630 2647 681
rect 2351 615 2411 630
rect 2469 615 2529 630
rect 2587 615 2647 630
rect 2705 615 2765 641
rect 2823 615 2883 641
rect 2941 615 3001 641
rect -31 415 29 441
rect 87 415 147 441
rect 205 415 265 441
rect 1290 432 1586 483
rect 1290 415 1350 432
rect 1408 415 1468 432
rect 1526 415 1586 432
rect 1867 415 1927 441
rect 1985 415 2045 441
rect 2103 415 2163 441
rect 3188 432 3484 483
rect 3188 415 3248 432
rect 3306 415 3366 432
rect 3424 415 3484 432
rect -31 198 29 215
rect 87 198 147 215
rect 205 198 265 215
rect 453 198 513 215
rect -31 147 513 198
rect 571 189 631 215
rect 689 189 749 215
rect 807 196 867 215
rect 925 196 985 215
rect 1043 196 1103 215
rect 1290 196 1350 215
rect 1408 196 1468 215
rect 94 63 154 147
rect 807 145 1350 196
rect 1392 189 1468 196
rect 1526 189 1586 215
rect 1867 198 1927 215
rect 1985 198 2045 215
rect 2103 198 2163 215
rect 2351 198 2411 215
rect 1392 145 1467 189
rect 1867 147 2411 198
rect 2469 189 2529 215
rect 2587 189 2647 215
rect 2705 196 2765 215
rect 2823 196 2883 215
rect 2941 196 3001 215
rect 3188 196 3248 215
rect 3306 196 3366 215
rect 1392 63 1452 145
rect 94 -5 203 63
rect 94 -705 154 -5
rect 396 -55 692 5
rect 396 -78 456 -55
rect 514 -78 574 -55
rect 632 -78 692 -55
rect 750 -54 1046 6
rect 1343 -5 1452 63
rect 750 -78 810 -54
rect 868 -78 928 -54
rect 986 -78 1046 -54
rect 396 -504 456 -478
rect 364 -645 431 -638
rect 514 -645 574 -478
rect 632 -504 692 -478
rect 750 -504 810 -478
rect 364 -654 574 -645
rect 364 -688 380 -654
rect 414 -688 574 -654
rect 364 -704 574 -688
rect 94 -721 245 -705
rect 94 -755 195 -721
rect 229 -755 245 -721
rect 94 -771 245 -755
rect 94 -810 154 -771
rect 514 -810 574 -704
rect 868 -645 928 -478
rect 986 -504 1046 -478
rect 1011 -645 1078 -638
rect 868 -654 1078 -645
rect 868 -688 1028 -654
rect 1062 -688 1078 -654
rect 868 -704 1078 -688
rect 630 -738 696 -722
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 630 -788 696 -772
rect 748 -737 814 -722
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 748 -787 814 -771
rect 632 -810 692 -788
rect 750 -810 810 -787
rect 868 -810 928 -704
rect 1392 -706 1452 -5
rect 1302 -722 1452 -706
rect 1302 -756 1318 -722
rect 1352 -756 1452 -722
rect 1302 -772 1452 -756
rect 1392 -810 1452 -772
rect 1992 -511 2052 147
rect 2705 145 3248 196
rect 3290 189 3366 196
rect 3424 189 3484 215
rect 3290 145 3365 189
rect 3290 63 3350 145
rect 2294 -55 2590 5
rect 2294 -78 2354 -55
rect 2412 -78 2472 -55
rect 2530 -78 2590 -55
rect 2648 -54 2944 6
rect 3241 -5 3350 63
rect 2648 -78 2708 -54
rect 2766 -78 2826 -54
rect 2884 -78 2944 -54
rect 2294 -504 2354 -478
rect 1992 -527 2059 -511
rect 1992 -561 2008 -527
rect 2042 -561 2059 -527
rect 1992 -577 2059 -561
rect 1992 -705 2052 -577
rect 2262 -645 2329 -638
rect 2412 -645 2472 -478
rect 2530 -504 2590 -478
rect 2648 -504 2708 -478
rect 2262 -654 2472 -645
rect 2262 -688 2278 -654
rect 2312 -688 2472 -654
rect 2262 -704 2472 -688
rect 1992 -721 2143 -705
rect 1992 -755 2093 -721
rect 2127 -755 2143 -721
rect 1992 -771 2143 -755
rect 1992 -810 2052 -771
rect 2412 -810 2472 -704
rect 2766 -645 2826 -478
rect 2884 -504 2944 -478
rect 2909 -645 2976 -638
rect 2766 -654 2976 -645
rect 2766 -688 2926 -654
rect 2960 -688 2976 -654
rect 2766 -704 2976 -688
rect 2528 -738 2594 -722
rect 2528 -772 2544 -738
rect 2578 -772 2594 -738
rect 2528 -788 2594 -772
rect 2646 -737 2712 -722
rect 2646 -771 2662 -737
rect 2696 -771 2712 -737
rect 2646 -787 2712 -771
rect 2530 -810 2590 -788
rect 2648 -810 2708 -787
rect 2766 -810 2826 -704
rect 3290 -706 3350 -5
rect 3200 -722 3350 -706
rect 3200 -756 3216 -722
rect 3250 -756 3350 -722
rect 3200 -772 3350 -756
rect 3290 -810 3350 -772
rect 94 -1036 154 -1010
rect 1392 -1036 1452 -1010
rect 1992 -1036 2052 -1010
rect 3290 -1036 3350 -1010
rect 514 -1236 574 -1210
rect 632 -1236 692 -1210
rect 750 -1236 810 -1210
rect 868 -1236 928 -1210
rect 2412 -1236 2472 -1210
rect 2530 -1236 2590 -1210
rect 2648 -1236 2708 -1210
rect 2766 -1236 2826 -1210
<< polycont >>
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1028 -688 1062 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
rect 2008 -561 2042 -527
rect 2278 -688 2312 -654
rect 2093 -755 2127 -721
rect 2926 -688 2960 -654
rect 2544 -772 2578 -738
rect 2662 -771 2696 -737
rect 3216 -756 3250 -722
<< locali >>
rect 2565 1091 2790 1167
rect 2565 942 2644 1091
rect 2711 942 2790 1091
rect 2565 836 2790 942
rect 761 656 1031 691
rect 407 603 441 619
rect -77 457 193 492
rect -77 403 -43 457
rect -77 211 -43 227
rect 41 403 75 419
rect 41 211 75 227
rect 159 403 193 457
rect 159 211 193 227
rect 277 403 311 419
rect 277 211 311 227
rect 407 211 441 227
rect 525 603 559 619
rect 525 211 559 227
rect 643 603 677 619
rect 643 211 677 227
rect 761 603 795 656
rect 761 211 795 227
rect 879 603 913 619
rect 879 211 913 227
rect 997 603 1031 656
rect 2659 656 2929 691
rect 997 211 1031 227
rect 1115 603 1149 619
rect 2305 603 2339 619
rect 1821 457 2091 492
rect 1115 211 1149 227
rect 1244 403 1278 419
rect 1244 211 1278 227
rect 1362 403 1396 419
rect 1362 211 1396 227
rect 1480 403 1514 419
rect 1480 211 1514 227
rect 1598 403 1632 419
rect 1598 211 1632 227
rect 1821 403 1855 457
rect 1821 211 1855 227
rect 1939 403 1973 419
rect 1939 211 1973 227
rect 2057 403 2091 457
rect 2057 211 2091 227
rect 2175 403 2209 419
rect 2175 211 2209 227
rect 2305 211 2339 227
rect 2423 603 2457 619
rect 2423 211 2457 227
rect 2541 603 2575 619
rect 2541 211 2575 227
rect 2659 603 2693 656
rect 2659 211 2693 227
rect 2777 603 2811 619
rect 2777 211 2811 227
rect 2895 603 2929 656
rect 2895 211 2929 227
rect 3013 603 3047 619
rect 3013 211 3047 227
rect 3142 403 3176 419
rect 3142 211 3176 227
rect 3260 403 3294 419
rect 3260 211 3294 227
rect 3378 403 3412 419
rect 3378 211 3412 227
rect 3496 403 3530 419
rect 3496 211 3530 227
rect 350 -90 384 -74
rect 468 -90 502 -74
rect 350 -482 384 -466
rect 467 -466 468 -419
rect 586 -90 620 -74
rect 502 -466 503 -419
rect 467 -524 503 -466
rect 704 -90 738 -74
rect 586 -482 620 -466
rect 702 -466 704 -419
rect 702 -524 738 -466
rect 822 -90 856 -74
rect 822 -482 856 -466
rect 940 -90 974 -74
rect 1058 -90 1092 -74
rect 974 -466 976 -420
rect 940 -524 976 -466
rect 1058 -482 1092 -466
rect 2248 -90 2282 -74
rect 2366 -90 2400 -74
rect 2248 -482 2282 -466
rect 2365 -466 2366 -419
rect 2484 -90 2518 -74
rect 2400 -466 2401 -419
rect 1563 -524 2060 -506
rect 467 -527 2060 -524
rect 467 -561 2008 -527
rect 2042 -561 2060 -527
rect 467 -564 2060 -561
rect 2365 -524 2401 -466
rect 2602 -90 2636 -74
rect 2484 -482 2518 -466
rect 2600 -466 2602 -419
rect 2600 -524 2636 -466
rect 2720 -90 2754 -74
rect 2720 -482 2754 -466
rect 2838 -90 2872 -74
rect 2956 -90 2990 -74
rect 2872 -466 2874 -420
rect 2838 -524 2874 -466
rect 2956 -482 2990 -466
rect 3461 -524 3561 -494
rect 2365 -564 3561 -524
rect 486 -565 2060 -564
rect 2384 -565 3561 -564
rect 364 -654 431 -638
rect 364 -688 380 -654
rect 414 -688 431 -654
rect 364 -704 431 -688
rect 195 -721 229 -705
rect 195 -771 229 -755
rect 541 -806 575 -565
rect 1563 -582 2060 -565
rect 1011 -654 1078 -638
rect 1011 -688 1028 -654
rect 1062 -688 1078 -654
rect 1011 -704 1078 -688
rect 2262 -654 2329 -638
rect 2262 -688 2278 -654
rect 2312 -688 2329 -654
rect 2262 -704 2329 -688
rect 1318 -722 1352 -706
rect 630 -772 646 -738
rect 680 -772 696 -738
rect 748 -771 764 -737
rect 798 -771 814 -737
rect 1318 -772 1352 -756
rect 2093 -721 2127 -705
rect 2093 -771 2127 -755
rect 2439 -806 2473 -565
rect 3461 -594 3561 -565
rect 2909 -654 2976 -638
rect 2909 -688 2926 -654
rect 2960 -688 2976 -654
rect 2909 -704 2976 -688
rect 3216 -722 3250 -706
rect 2528 -772 2544 -738
rect 2578 -772 2594 -738
rect 2646 -771 2662 -737
rect 2696 -771 2712 -737
rect 3216 -772 3250 -756
rect 48 -822 82 -806
rect 48 -1014 82 -998
rect 166 -822 200 -806
rect 166 -1014 200 -998
rect 468 -822 502 -806
rect 541 -822 620 -806
rect 541 -852 586 -822
rect 468 -1265 503 -1198
rect 586 -1214 620 -1198
rect 704 -822 738 -806
rect 704 -1214 738 -1198
rect 822 -822 856 -806
rect 940 -822 974 -806
rect 1346 -822 1380 -806
rect 1346 -1014 1380 -998
rect 1464 -822 1498 -806
rect 1464 -1014 1498 -998
rect 1946 -822 1980 -806
rect 1946 -1014 1980 -998
rect 2064 -822 2098 -806
rect 2064 -1014 2098 -998
rect 2366 -822 2400 -806
rect 822 -1214 856 -1198
rect 939 -1265 974 -1198
rect 468 -1300 974 -1265
rect 2439 -822 2518 -806
rect 2439 -852 2484 -822
rect 2366 -1265 2401 -1198
rect 2484 -1214 2518 -1198
rect 2602 -822 2636 -806
rect 2602 -1214 2636 -1198
rect 2720 -822 2754 -806
rect 2838 -822 2872 -806
rect 3244 -822 3278 -806
rect 3244 -1014 3278 -998
rect 3362 -822 3396 -806
rect 3362 -1014 3396 -998
rect 2720 -1214 2754 -1198
rect 2837 -1265 2872 -1198
rect 2366 -1300 2872 -1265
rect 639 -1507 811 -1460
rect 639 -1670 678 -1507
rect 768 -1670 811 -1507
rect 639 -1710 811 -1670
<< viali >>
rect -77 227 -43 403
rect 41 227 75 403
rect 159 227 193 403
rect 277 227 311 403
rect 407 227 441 603
rect 525 227 559 603
rect 643 227 677 603
rect 761 227 795 603
rect 879 227 913 603
rect 997 227 1031 603
rect 1115 227 1149 603
rect 1244 227 1278 403
rect 1362 227 1396 403
rect 1480 227 1514 403
rect 1598 227 1632 403
rect 1821 227 1855 403
rect 1939 227 1973 403
rect 2057 227 2091 403
rect 2175 227 2209 403
rect 2305 227 2339 603
rect 2423 227 2457 603
rect 2541 227 2575 603
rect 2659 227 2693 603
rect 2777 227 2811 603
rect 2895 227 2929 603
rect 3013 227 3047 603
rect 3142 227 3176 403
rect 3260 227 3294 403
rect 3378 227 3412 403
rect 3496 227 3530 403
rect 350 -466 384 -90
rect 468 -466 502 -90
rect 586 -466 620 -90
rect 704 -466 738 -90
rect 822 -466 856 -90
rect 940 -466 974 -90
rect 1058 -466 1092 -90
rect 2248 -466 2282 -90
rect 2366 -466 2400 -90
rect 2484 -466 2518 -90
rect 2602 -466 2636 -90
rect 2720 -466 2754 -90
rect 2838 -466 2872 -90
rect 2956 -466 2990 -90
rect 380 -688 414 -654
rect 195 -755 229 -721
rect 1028 -688 1062 -654
rect 2278 -688 2312 -654
rect 646 -772 680 -738
rect 764 -771 798 -737
rect 1318 -756 1352 -722
rect 2093 -755 2127 -721
rect 2926 -688 2960 -654
rect 2544 -772 2578 -738
rect 2662 -771 2696 -737
rect 3216 -756 3250 -722
rect 48 -998 82 -822
rect 166 -998 200 -822
rect 468 -1198 502 -822
rect 586 -1198 620 -822
rect 704 -1198 738 -822
rect 822 -1198 856 -822
rect 940 -1198 974 -822
rect 1346 -998 1380 -822
rect 1464 -998 1498 -822
rect 1946 -998 1980 -822
rect 2064 -998 2098 -822
rect 2366 -1198 2400 -822
rect 2484 -1198 2518 -822
rect 2602 -1198 2636 -822
rect 2720 -1198 2754 -822
rect 2838 -1198 2872 -822
rect 3244 -998 3278 -822
rect 3362 -998 3396 -822
<< metal1 >>
rect 703 867 713 975
rect 845 867 855 975
rect 2601 867 2611 975
rect 2743 867 2753 975
rect 713 827 845 867
rect 2611 827 2743 867
rect 712 761 845 827
rect 2610 761 2743 827
rect 41 718 1514 761
rect 41 415 75 718
rect 407 615 441 718
rect 643 615 677 718
rect 879 615 913 718
rect 1115 615 1149 718
rect 401 603 447 615
rect -83 403 -37 415
rect -83 227 -77 403
rect -43 227 -37 403
rect -83 215 -37 227
rect 35 403 81 415
rect 35 227 41 403
rect 75 227 81 403
rect 35 215 81 227
rect 153 403 199 415
rect 153 227 159 403
rect 193 227 199 403
rect 153 215 199 227
rect 271 403 317 415
rect 401 403 407 603
rect 271 227 277 403
rect 311 227 407 403
rect 441 227 447 603
rect 271 215 317 227
rect 401 215 447 227
rect 519 603 565 615
rect 519 227 525 603
rect 559 227 565 603
rect 519 215 565 227
rect 637 603 683 615
rect 637 227 643 603
rect 677 227 683 603
rect 637 215 683 227
rect 755 603 801 615
rect 755 227 761 603
rect 795 227 801 603
rect 755 215 801 227
rect 873 603 919 615
rect 873 227 879 603
rect 913 227 919 603
rect 873 215 919 227
rect 991 603 1037 615
rect 991 227 997 603
rect 1031 227 1037 603
rect 991 215 1037 227
rect 1109 603 1155 615
rect 1109 227 1115 603
rect 1149 403 1155 603
rect 1480 415 1514 718
rect 1939 718 3412 761
rect 1939 415 1973 718
rect 2305 615 2339 718
rect 2541 615 2575 718
rect 2777 615 2811 718
rect 3013 615 3047 718
rect 2299 603 2345 615
rect 1238 403 1284 415
rect 1149 227 1244 403
rect 1278 227 1284 403
rect 1109 215 1155 227
rect 1238 215 1284 227
rect 1356 403 1402 415
rect 1356 227 1362 403
rect 1396 227 1402 403
rect 1356 215 1402 227
rect 1474 403 1520 415
rect 1474 227 1480 403
rect 1514 227 1520 403
rect 1474 215 1520 227
rect 1592 403 1638 415
rect 1592 227 1598 403
rect 1632 227 1638 403
rect 1592 215 1638 227
rect 1815 403 1861 415
rect 1815 227 1821 403
rect 1855 227 1861 403
rect 1815 215 1861 227
rect 1933 403 1979 415
rect 1933 227 1939 403
rect 1973 227 1979 403
rect 1933 215 1979 227
rect 2051 403 2097 415
rect 2051 227 2057 403
rect 2091 227 2097 403
rect 2051 215 2097 227
rect 2169 403 2215 415
rect 2299 403 2305 603
rect 2169 227 2175 403
rect 2209 227 2305 403
rect 2339 227 2345 603
rect 2169 215 2215 227
rect 2299 215 2345 227
rect 2417 603 2463 615
rect 2417 227 2423 603
rect 2457 227 2463 603
rect 2417 215 2463 227
rect 2535 603 2581 615
rect 2535 227 2541 603
rect 2575 227 2581 603
rect 2535 215 2581 227
rect 2653 603 2699 615
rect 2653 227 2659 603
rect 2693 227 2699 603
rect 2653 215 2699 227
rect 2771 603 2817 615
rect 2771 227 2777 603
rect 2811 227 2817 603
rect 2771 215 2817 227
rect 2889 603 2935 615
rect 2889 227 2895 603
rect 2929 227 2935 603
rect 2889 215 2935 227
rect 3007 603 3053 615
rect 3007 227 3013 603
rect 3047 403 3053 603
rect 3378 415 3412 718
rect 3136 403 3182 415
rect 3047 227 3142 403
rect 3176 227 3182 403
rect 3007 215 3053 227
rect 3136 215 3182 227
rect 3254 403 3300 415
rect 3254 227 3260 403
rect 3294 227 3300 403
rect 3254 215 3300 227
rect 3372 403 3418 415
rect 3372 227 3378 403
rect 3412 227 3418 403
rect 3372 215 3418 227
rect 3490 403 3536 415
rect 3490 227 3496 403
rect 3530 227 3536 403
rect 3490 215 3536 227
rect -77 181 -43 215
rect 525 181 559 215
rect 761 181 795 215
rect -77 146 82 181
rect 525 146 795 181
rect 1362 181 1396 215
rect 1598 181 1632 215
rect 1362 146 1632 181
rect 1821 181 1855 215
rect 2423 181 2457 215
rect 2659 181 2693 215
rect 1821 146 1980 181
rect 2423 146 2693 181
rect 3260 181 3294 215
rect 3496 181 3530 215
rect 3260 146 3530 181
rect 48 -638 82 146
rect 761 84 795 146
rect 350 46 1092 84
rect 350 -78 384 46
rect 586 -78 620 46
rect 822 -78 856 46
rect 1058 -78 1092 46
rect 344 -90 390 -78
rect 344 -466 350 -90
rect 384 -466 390 -90
rect 344 -478 390 -466
rect 462 -90 508 -78
rect 462 -466 468 -90
rect 502 -466 508 -90
rect 462 -478 508 -466
rect 580 -90 626 -78
rect 580 -466 586 -90
rect 620 -466 626 -90
rect 580 -478 626 -466
rect 698 -90 744 -78
rect 698 -466 704 -90
rect 738 -466 744 -90
rect 698 -478 744 -466
rect 816 -90 862 -78
rect 816 -466 822 -90
rect 856 -466 862 -90
rect 816 -478 862 -466
rect 934 -90 980 -78
rect 934 -466 940 -90
rect 974 -466 980 -90
rect 934 -478 980 -466
rect 1052 -90 1098 -78
rect 1052 -466 1058 -90
rect 1092 -466 1098 -90
rect 1052 -478 1098 -466
rect 1464 -637 1498 146
rect 1191 -638 1498 -637
rect 48 -643 364 -638
rect 1078 -643 1498 -638
rect 48 -654 431 -643
rect 48 -681 380 -654
rect 48 -810 82 -681
rect 364 -688 380 -681
rect 414 -688 431 -654
rect 364 -694 431 -688
rect 1011 -654 1498 -643
rect 1011 -688 1028 -654
rect 1062 -681 1498 -654
rect 1062 -688 1078 -681
rect 1191 -682 1498 -681
rect 1011 -694 1078 -688
rect 189 -721 245 -709
rect 189 -755 195 -721
rect 229 -722 245 -721
rect 1302 -722 1358 -710
rect 229 -738 696 -722
rect 229 -755 646 -738
rect 189 -771 646 -755
rect 630 -772 646 -771
rect 680 -772 696 -738
rect 630 -779 696 -772
rect 748 -737 1318 -722
rect 748 -771 764 -737
rect 798 -756 1318 -737
rect 1352 -756 1358 -722
rect 798 -771 1358 -756
rect 748 -781 815 -771
rect 1302 -772 1358 -771
rect 1464 -810 1498 -682
rect 1946 -638 1980 146
rect 2659 84 2693 146
rect 2248 46 2990 84
rect 2248 -78 2282 46
rect 2484 -78 2518 46
rect 2720 -78 2754 46
rect 2956 -78 2990 46
rect 2242 -90 2288 -78
rect 2242 -466 2248 -90
rect 2282 -466 2288 -90
rect 2242 -478 2288 -466
rect 2360 -90 2406 -78
rect 2360 -466 2366 -90
rect 2400 -466 2406 -90
rect 2360 -478 2406 -466
rect 2478 -90 2524 -78
rect 2478 -466 2484 -90
rect 2518 -466 2524 -90
rect 2478 -478 2524 -466
rect 2596 -90 2642 -78
rect 2596 -466 2602 -90
rect 2636 -466 2642 -90
rect 2596 -478 2642 -466
rect 2714 -90 2760 -78
rect 2714 -466 2720 -90
rect 2754 -466 2760 -90
rect 2714 -478 2760 -466
rect 2832 -90 2878 -78
rect 2832 -466 2838 -90
rect 2872 -466 2878 -90
rect 2832 -478 2878 -466
rect 2950 -90 2996 -78
rect 2950 -466 2956 -90
rect 2990 -466 2996 -90
rect 2950 -478 2996 -466
rect 3362 -637 3396 146
rect 3089 -638 3396 -637
rect 1946 -643 2262 -638
rect 2976 -643 3396 -638
rect 1946 -654 2329 -643
rect 1946 -681 2278 -654
rect 1946 -810 1980 -681
rect 2262 -688 2278 -681
rect 2312 -688 2329 -654
rect 2262 -694 2329 -688
rect 2909 -654 3396 -643
rect 2909 -688 2926 -654
rect 2960 -681 3396 -654
rect 2960 -688 2976 -681
rect 3089 -682 3396 -681
rect 2909 -694 2976 -688
rect 2087 -721 2143 -709
rect 2087 -755 2093 -721
rect 2127 -722 2143 -721
rect 3200 -722 3256 -710
rect 2127 -738 2594 -722
rect 2127 -755 2544 -738
rect 2087 -771 2544 -755
rect 2528 -772 2544 -771
rect 2578 -772 2594 -738
rect 2528 -779 2594 -772
rect 2646 -737 3216 -722
rect 2646 -771 2662 -737
rect 2696 -756 3216 -737
rect 3250 -756 3256 -722
rect 2696 -771 3256 -756
rect 2646 -781 2713 -771
rect 3200 -772 3256 -771
rect 3362 -810 3396 -682
rect 42 -822 88 -810
rect 42 -998 48 -822
rect 82 -998 88 -822
rect 42 -1010 88 -998
rect 160 -822 206 -810
rect 160 -998 166 -822
rect 200 -998 206 -822
rect 160 -1010 206 -998
rect 462 -822 508 -810
rect 165 -1304 199 -1010
rect 462 -1198 468 -822
rect 502 -1198 508 -822
rect 462 -1210 508 -1198
rect 580 -822 626 -810
rect 580 -1198 586 -822
rect 620 -1198 626 -822
rect 580 -1210 626 -1198
rect 698 -822 744 -810
rect 698 -1198 704 -822
rect 738 -1198 744 -822
rect 698 -1210 744 -1198
rect 816 -822 862 -810
rect 816 -1198 822 -822
rect 856 -1198 862 -822
rect 816 -1210 862 -1198
rect 934 -822 980 -810
rect 934 -1198 940 -822
rect 974 -1198 980 -822
rect 1340 -822 1386 -810
rect 1340 -998 1346 -822
rect 1380 -998 1386 -822
rect 1340 -1010 1386 -998
rect 1458 -822 1504 -810
rect 1458 -998 1464 -822
rect 1498 -998 1504 -822
rect 1458 -1010 1504 -998
rect 1940 -822 1986 -810
rect 1940 -998 1946 -822
rect 1980 -998 1986 -822
rect 1940 -1010 1986 -998
rect 2058 -822 2104 -810
rect 2058 -998 2064 -822
rect 2098 -998 2104 -822
rect 2058 -1010 2104 -998
rect 2360 -822 2406 -810
rect 934 -1210 980 -1198
rect 822 -1304 856 -1210
rect 1346 -1304 1379 -1010
rect 165 -1336 1379 -1304
rect 2063 -1304 2097 -1010
rect 2360 -1198 2366 -822
rect 2400 -1198 2406 -822
rect 2360 -1210 2406 -1198
rect 2478 -822 2524 -810
rect 2478 -1198 2484 -822
rect 2518 -1198 2524 -822
rect 2478 -1210 2524 -1198
rect 2596 -822 2642 -810
rect 2596 -1198 2602 -822
rect 2636 -1198 2642 -822
rect 2596 -1210 2642 -1198
rect 2714 -822 2760 -810
rect 2714 -1198 2720 -822
rect 2754 -1198 2760 -822
rect 2714 -1210 2760 -1198
rect 2832 -822 2878 -810
rect 2832 -1198 2838 -822
rect 2872 -1198 2878 -822
rect 3238 -822 3284 -810
rect 3238 -998 3244 -822
rect 3278 -998 3284 -822
rect 3238 -1010 3284 -998
rect 3356 -822 3402 -810
rect 3356 -998 3362 -822
rect 3396 -998 3402 -822
rect 3356 -1010 3402 -998
rect 2832 -1210 2878 -1198
rect 2720 -1304 2754 -1210
rect 3244 -1304 3277 -1010
rect 2063 -1336 3277 -1304
rect 658 -1421 790 -1336
rect 2556 -1421 2688 -1336
rect 648 -1529 658 -1421
rect 790 -1529 800 -1421
rect 2546 -1529 2556 -1421
rect 2688 -1529 2698 -1421
<< via1 >>
rect 713 867 845 975
rect 2611 867 2743 975
rect 658 -1529 790 -1421
rect 2556 -1529 2688 -1421
<< metal2 >>
rect 702 986 855 996
rect 702 847 855 857
rect 2600 986 2753 996
rect 2600 847 2753 857
rect 648 -1411 801 -1401
rect 648 -1550 801 -1540
rect 2546 -1411 2699 -1401
rect 2546 -1550 2699 -1540
<< via2 >>
rect 702 975 855 986
rect 702 867 713 975
rect 713 867 845 975
rect 845 867 855 975
rect 702 857 855 867
rect 2600 975 2753 986
rect 2600 867 2611 975
rect 2611 867 2743 975
rect 2743 867 2753 975
rect 2600 857 2753 867
rect 648 -1421 801 -1411
rect 648 -1529 658 -1421
rect 658 -1529 790 -1421
rect 790 -1529 801 -1421
rect 648 -1540 801 -1529
rect 2546 -1421 2699 -1411
rect 2546 -1529 2556 -1421
rect 2556 -1529 2688 -1421
rect 2688 -1529 2699 -1421
rect 2546 -1540 2699 -1529
<< metal3 >>
rect 670 838 680 1017
rect 879 838 889 1017
rect 2568 838 2578 1017
rect 2777 838 2787 1017
rect 614 -1571 624 -1392
rect 823 -1571 833 -1392
rect 2512 -1571 2522 -1392
rect 2721 -1571 2731 -1392
<< via3 >>
rect 680 986 879 1017
rect 680 857 702 986
rect 702 857 855 986
rect 855 857 879 986
rect 680 838 879 857
rect 2578 986 2777 1017
rect 2578 857 2600 986
rect 2600 857 2753 986
rect 2753 857 2777 986
rect 2578 838 2777 857
rect 624 -1411 823 -1392
rect 624 -1540 648 -1411
rect 648 -1540 801 -1411
rect 801 -1540 823 -1411
rect 624 -1571 823 -1540
rect 2522 -1411 2721 -1392
rect 2522 -1540 2546 -1411
rect 2546 -1540 2699 -1411
rect 2699 -1540 2721 -1411
rect 2522 -1571 2721 -1540
<< metal4 >>
rect 935 1165 2481 1166
rect 538 1017 2905 1165
rect 538 923 680 1017
rect 658 838 680 923
rect 879 922 2578 1017
rect 879 838 969 922
rect 658 835 969 838
rect 2476 838 2578 922
rect 2777 923 2905 1017
rect 2777 838 2801 923
rect 2476 835 2801 838
rect 600 -1392 845 -1389
rect 600 -1477 624 -1392
rect 496 -1571 624 -1477
rect 823 -1477 845 -1392
rect 2498 -1392 2743 -1389
rect 2498 -1477 2522 -1392
rect 823 -1528 965 -1477
rect 2394 -1528 2522 -1477
rect 823 -1571 2522 -1528
rect 2721 -1477 2743 -1392
rect 2721 -1571 2863 -1477
rect 496 -1719 2863 -1571
rect 884 -1721 2555 -1719
<< labels >>
flabel poly 107 4 192 52 1 FreeSans 240 0 0 0 A
port 6 n
flabel poly 1358 5 1443 53 1 FreeSans 240 0 0 0 B
port 7 n
flabel metal4 1212 980 2315 1147 1 FreeSans 1040 0 0 0 VDD
port 10 n
flabel metal4 1166 -1713 2269 -1546 1 FreeSans 1040 0 0 0 VSS
port 9 n
flabel poly 3256 5 3341 53 1 FreeSans 240 0 0 0 C
port 11 n
flabel locali 3469 -586 3552 -502 1 FreeSans 320 0 0 0 OUT
port 12 n
<< end >>
