magic
tech sky130B
magscale 1 2
timestamp 1735941024
<< nwell >>
rect 16853 -216 17140 -215
rect 18000 -216 18235 -215
rect 14371 -270 14611 -269
rect 14368 -503 14611 -270
rect 14368 -685 14612 -503
rect 16850 -613 17140 -216
rect 17827 -609 18309 -216
rect 13930 -1009 15122 -685
rect 16255 -1080 17140 -613
rect 16255 -1133 17141 -1080
rect 17397 -1133 18309 -609
rect 16255 -1137 17142 -1133
rect 16684 -1422 17142 -1137
rect 17827 -1392 18309 -1133
rect 16684 -1720 17168 -1422
rect 17826 -1716 18310 -1392
rect 14385 -1920 14625 -1919
rect 14382 -2153 14625 -1920
rect 14382 -2335 14626 -2153
rect 13944 -2659 15136 -2335
rect 18096 -2752 18324 -2262
rect 15407 -2952 16730 -2752
rect 17790 -2952 18628 -2752
rect 15407 -3276 19111 -2952
rect 14380 -3524 14620 -3523
rect 14377 -3757 14620 -3524
rect 14377 -3939 14621 -3757
rect 13939 -4263 15131 -3939
rect 15835 -3969 16673 -3276
rect 17733 -3969 18571 -3276
<< nmos >>
rect 14261 -1584 14321 -1184
rect 14379 -1584 14439 -1184
rect 14614 -1384 14674 -1184
rect 16259 -1658 16319 -1458
rect 16377 -1658 16437 -1458
rect 16495 -1658 16555 -1458
rect 17401 -1654 17461 -1454
rect 17519 -1654 17579 -1454
rect 17637 -1654 17697 -1454
rect 14275 -3234 14335 -2834
rect 14393 -3234 14453 -2834
rect 14628 -3034 14688 -2834
rect 14270 -4838 14330 -4438
rect 14388 -4838 14448 -4438
rect 14623 -4638 14683 -4438
rect 15627 -4439 15687 -4239
rect 16047 -4639 16107 -4239
rect 16165 -4639 16225 -4239
rect 16283 -4639 16343 -4239
rect 16401 -4639 16461 -4239
rect 16925 -4439 16985 -4239
rect 17525 -4439 17585 -4239
rect 17945 -4639 18005 -4239
rect 18063 -4639 18123 -4239
rect 18181 -4639 18241 -4239
rect 18299 -4639 18359 -4239
rect 18823 -4439 18883 -4239
<< pmos >>
rect 14024 -947 14084 -747
rect 14142 -947 14202 -747
rect 14260 -947 14320 -747
rect 14378 -947 14438 -747
rect 14496 -947 14556 -747
rect 14614 -947 14674 -747
rect 14732 -947 14792 -747
rect 14850 -947 14910 -747
rect 14968 -947 15028 -747
rect 16349 -1075 16409 -675
rect 16467 -1075 16527 -675
rect 16585 -1075 16645 -675
rect 16703 -1075 16763 -675
rect 16821 -1075 16881 -675
rect 16939 -1075 16999 -675
rect 17491 -1071 17551 -671
rect 17609 -1071 17669 -671
rect 17727 -1071 17787 -671
rect 17845 -1071 17905 -671
rect 17963 -1071 18023 -671
rect 18081 -1071 18141 -671
rect 16778 -1658 16838 -1458
rect 16896 -1658 16956 -1458
rect 17014 -1658 17074 -1458
rect 17920 -1654 17980 -1454
rect 18038 -1654 18098 -1454
rect 18156 -1654 18216 -1454
rect 14038 -2597 14098 -2397
rect 14156 -2597 14216 -2397
rect 14274 -2597 14334 -2397
rect 14392 -2597 14452 -2397
rect 14510 -2597 14570 -2397
rect 14628 -2597 14688 -2397
rect 14746 -2597 14806 -2397
rect 14864 -2597 14924 -2397
rect 14982 -2597 15042 -2397
rect 15502 -3214 15562 -3014
rect 15620 -3214 15680 -3014
rect 15738 -3214 15798 -3014
rect 15986 -3214 16046 -2814
rect 16104 -3214 16164 -2814
rect 16222 -3214 16282 -2814
rect 16340 -3214 16400 -2814
rect 16458 -3214 16518 -2814
rect 16576 -3214 16636 -2814
rect 16823 -3214 16883 -3014
rect 16941 -3214 17001 -3014
rect 17059 -3214 17119 -3014
rect 17400 -3214 17460 -3014
rect 17518 -3214 17578 -3014
rect 17636 -3214 17696 -3014
rect 17884 -3214 17944 -2814
rect 18002 -3214 18062 -2814
rect 18120 -3214 18180 -2814
rect 18238 -3214 18298 -2814
rect 18356 -3214 18416 -2814
rect 18474 -3214 18534 -2814
rect 18721 -3214 18781 -3014
rect 18839 -3214 18899 -3014
rect 18957 -3214 19017 -3014
rect 14033 -4201 14093 -4001
rect 14151 -4201 14211 -4001
rect 14269 -4201 14329 -4001
rect 14387 -4201 14447 -4001
rect 14505 -4201 14565 -4001
rect 14623 -4201 14683 -4001
rect 14741 -4201 14801 -4001
rect 14859 -4201 14919 -4001
rect 14977 -4201 15037 -4001
rect 15929 -3907 15989 -3507
rect 16047 -3907 16107 -3507
rect 16165 -3907 16225 -3507
rect 16283 -3907 16343 -3507
rect 16401 -3907 16461 -3507
rect 16519 -3907 16579 -3507
rect 17827 -3907 17887 -3507
rect 17945 -3907 18005 -3507
rect 18063 -3907 18123 -3507
rect 18181 -3907 18241 -3507
rect 18299 -3907 18359 -3507
rect 18417 -3907 18477 -3507
<< ndiff >>
rect 14203 -1196 14261 -1184
rect 14203 -1572 14215 -1196
rect 14249 -1572 14261 -1196
rect 14203 -1584 14261 -1572
rect 14321 -1196 14379 -1184
rect 14321 -1572 14333 -1196
rect 14367 -1572 14379 -1196
rect 14321 -1584 14379 -1572
rect 14439 -1196 14497 -1184
rect 14439 -1572 14451 -1196
rect 14485 -1572 14497 -1196
rect 14556 -1196 14614 -1184
rect 14556 -1372 14568 -1196
rect 14602 -1372 14614 -1196
rect 14556 -1384 14614 -1372
rect 14674 -1196 14732 -1184
rect 14674 -1372 14686 -1196
rect 14720 -1372 14732 -1196
rect 14674 -1384 14732 -1372
rect 16201 -1470 16259 -1458
rect 14439 -1584 14497 -1572
rect 16201 -1646 16213 -1470
rect 16247 -1646 16259 -1470
rect 16201 -1658 16259 -1646
rect 16319 -1470 16377 -1458
rect 16319 -1646 16331 -1470
rect 16365 -1646 16377 -1470
rect 16319 -1658 16377 -1646
rect 16437 -1470 16495 -1458
rect 16437 -1646 16449 -1470
rect 16483 -1646 16495 -1470
rect 16437 -1658 16495 -1646
rect 16555 -1470 16613 -1458
rect 16555 -1646 16567 -1470
rect 16601 -1646 16613 -1470
rect 16555 -1658 16613 -1646
rect 17343 -1466 17401 -1454
rect 17343 -1642 17355 -1466
rect 17389 -1642 17401 -1466
rect 17343 -1654 17401 -1642
rect 17461 -1466 17519 -1454
rect 17461 -1642 17473 -1466
rect 17507 -1642 17519 -1466
rect 17461 -1654 17519 -1642
rect 17579 -1466 17637 -1454
rect 17579 -1642 17591 -1466
rect 17625 -1642 17637 -1466
rect 17579 -1654 17637 -1642
rect 17697 -1466 17755 -1454
rect 17697 -1642 17709 -1466
rect 17743 -1642 17755 -1466
rect 17697 -1654 17755 -1642
rect 14217 -2846 14275 -2834
rect 14217 -3222 14229 -2846
rect 14263 -3222 14275 -2846
rect 14217 -3234 14275 -3222
rect 14335 -2846 14393 -2834
rect 14335 -3222 14347 -2846
rect 14381 -3222 14393 -2846
rect 14335 -3234 14393 -3222
rect 14453 -2846 14511 -2834
rect 14453 -3222 14465 -2846
rect 14499 -3222 14511 -2846
rect 14570 -2846 14628 -2834
rect 14570 -3022 14582 -2846
rect 14616 -3022 14628 -2846
rect 14570 -3034 14628 -3022
rect 14688 -2846 14746 -2834
rect 14688 -3022 14700 -2846
rect 14734 -3022 14746 -2846
rect 14688 -3034 14746 -3022
rect 14453 -3234 14511 -3222
rect 15569 -4251 15627 -4239
rect 15569 -4427 15581 -4251
rect 15615 -4427 15627 -4251
rect 14212 -4450 14270 -4438
rect 14212 -4826 14224 -4450
rect 14258 -4826 14270 -4450
rect 14212 -4838 14270 -4826
rect 14330 -4450 14388 -4438
rect 14330 -4826 14342 -4450
rect 14376 -4826 14388 -4450
rect 14330 -4838 14388 -4826
rect 14448 -4450 14506 -4438
rect 14448 -4826 14460 -4450
rect 14494 -4826 14506 -4450
rect 14565 -4450 14623 -4438
rect 14565 -4626 14577 -4450
rect 14611 -4626 14623 -4450
rect 14565 -4638 14623 -4626
rect 14683 -4450 14741 -4438
rect 15569 -4439 15627 -4427
rect 15687 -4251 15745 -4239
rect 15687 -4427 15699 -4251
rect 15733 -4427 15745 -4251
rect 15687 -4439 15745 -4427
rect 15989 -4251 16047 -4239
rect 14683 -4626 14695 -4450
rect 14729 -4626 14741 -4450
rect 14683 -4638 14741 -4626
rect 15989 -4627 16001 -4251
rect 16035 -4627 16047 -4251
rect 15989 -4639 16047 -4627
rect 16107 -4251 16165 -4239
rect 16107 -4627 16119 -4251
rect 16153 -4627 16165 -4251
rect 16107 -4639 16165 -4627
rect 16225 -4251 16283 -4239
rect 16225 -4627 16237 -4251
rect 16271 -4627 16283 -4251
rect 16225 -4639 16283 -4627
rect 16343 -4251 16401 -4239
rect 16343 -4627 16355 -4251
rect 16389 -4627 16401 -4251
rect 16343 -4639 16401 -4627
rect 16461 -4251 16519 -4239
rect 16461 -4627 16473 -4251
rect 16507 -4627 16519 -4251
rect 16867 -4251 16925 -4239
rect 16867 -4427 16879 -4251
rect 16913 -4427 16925 -4251
rect 16867 -4439 16925 -4427
rect 16985 -4251 17043 -4239
rect 16985 -4427 16997 -4251
rect 17031 -4427 17043 -4251
rect 16985 -4439 17043 -4427
rect 17467 -4251 17525 -4239
rect 17467 -4427 17479 -4251
rect 17513 -4427 17525 -4251
rect 17467 -4439 17525 -4427
rect 17585 -4251 17643 -4239
rect 17585 -4427 17597 -4251
rect 17631 -4427 17643 -4251
rect 17585 -4439 17643 -4427
rect 17887 -4251 17945 -4239
rect 16461 -4639 16519 -4627
rect 17887 -4627 17899 -4251
rect 17933 -4627 17945 -4251
rect 17887 -4639 17945 -4627
rect 18005 -4251 18063 -4239
rect 18005 -4627 18017 -4251
rect 18051 -4627 18063 -4251
rect 18005 -4639 18063 -4627
rect 18123 -4251 18181 -4239
rect 18123 -4627 18135 -4251
rect 18169 -4627 18181 -4251
rect 18123 -4639 18181 -4627
rect 18241 -4251 18299 -4239
rect 18241 -4627 18253 -4251
rect 18287 -4627 18299 -4251
rect 18241 -4639 18299 -4627
rect 18359 -4251 18417 -4239
rect 18359 -4627 18371 -4251
rect 18405 -4627 18417 -4251
rect 18765 -4251 18823 -4239
rect 18765 -4427 18777 -4251
rect 18811 -4427 18823 -4251
rect 18765 -4439 18823 -4427
rect 18883 -4251 18941 -4239
rect 18883 -4427 18895 -4251
rect 18929 -4427 18941 -4251
rect 18883 -4439 18941 -4427
rect 18359 -4639 18417 -4627
rect 14448 -4838 14506 -4826
<< pdiff >>
rect 16291 -687 16349 -675
rect 13966 -759 14024 -747
rect 13966 -935 13978 -759
rect 14012 -935 14024 -759
rect 13966 -947 14024 -935
rect 14084 -759 14142 -747
rect 14084 -935 14096 -759
rect 14130 -935 14142 -759
rect 14084 -947 14142 -935
rect 14202 -759 14260 -747
rect 14202 -935 14214 -759
rect 14248 -935 14260 -759
rect 14202 -947 14260 -935
rect 14320 -759 14378 -747
rect 14320 -935 14332 -759
rect 14366 -935 14378 -759
rect 14320 -947 14378 -935
rect 14438 -759 14496 -747
rect 14438 -935 14450 -759
rect 14484 -935 14496 -759
rect 14438 -947 14496 -935
rect 14556 -759 14614 -747
rect 14556 -935 14568 -759
rect 14602 -935 14614 -759
rect 14556 -947 14614 -935
rect 14674 -759 14732 -747
rect 14674 -935 14686 -759
rect 14720 -935 14732 -759
rect 14674 -947 14732 -935
rect 14792 -759 14850 -747
rect 14792 -935 14804 -759
rect 14838 -935 14850 -759
rect 14792 -947 14850 -935
rect 14910 -759 14968 -747
rect 14910 -935 14922 -759
rect 14956 -935 14968 -759
rect 14910 -947 14968 -935
rect 15028 -759 15086 -747
rect 15028 -935 15040 -759
rect 15074 -935 15086 -759
rect 15028 -947 15086 -935
rect 16291 -1063 16303 -687
rect 16337 -1063 16349 -687
rect 16291 -1075 16349 -1063
rect 16409 -687 16467 -675
rect 16409 -1063 16421 -687
rect 16455 -1063 16467 -687
rect 16409 -1075 16467 -1063
rect 16527 -687 16585 -675
rect 16527 -1063 16539 -687
rect 16573 -1063 16585 -687
rect 16527 -1075 16585 -1063
rect 16645 -687 16703 -675
rect 16645 -1063 16657 -687
rect 16691 -1063 16703 -687
rect 16645 -1075 16703 -1063
rect 16763 -687 16821 -675
rect 16763 -1063 16775 -687
rect 16809 -1063 16821 -687
rect 16763 -1075 16821 -1063
rect 16881 -687 16939 -675
rect 16881 -1063 16893 -687
rect 16927 -1063 16939 -687
rect 16881 -1075 16939 -1063
rect 16999 -687 17057 -675
rect 16999 -1063 17011 -687
rect 17045 -1063 17057 -687
rect 16999 -1075 17057 -1063
rect 17433 -683 17491 -671
rect 17433 -1059 17445 -683
rect 17479 -1059 17491 -683
rect 17433 -1071 17491 -1059
rect 17551 -683 17609 -671
rect 17551 -1059 17563 -683
rect 17597 -1059 17609 -683
rect 17551 -1071 17609 -1059
rect 17669 -683 17727 -671
rect 17669 -1059 17681 -683
rect 17715 -1059 17727 -683
rect 17669 -1071 17727 -1059
rect 17787 -683 17845 -671
rect 17787 -1059 17799 -683
rect 17833 -1059 17845 -683
rect 17787 -1071 17845 -1059
rect 17905 -683 17963 -671
rect 17905 -1059 17917 -683
rect 17951 -1059 17963 -683
rect 17905 -1071 17963 -1059
rect 18023 -683 18081 -671
rect 18023 -1059 18035 -683
rect 18069 -1059 18081 -683
rect 18023 -1071 18081 -1059
rect 18141 -683 18199 -671
rect 18141 -1059 18153 -683
rect 18187 -1059 18199 -683
rect 18141 -1071 18199 -1059
rect 16720 -1470 16778 -1458
rect 16720 -1646 16732 -1470
rect 16766 -1646 16778 -1470
rect 16720 -1658 16778 -1646
rect 16838 -1470 16896 -1458
rect 16838 -1646 16850 -1470
rect 16884 -1646 16896 -1470
rect 16838 -1658 16896 -1646
rect 16956 -1470 17014 -1458
rect 16956 -1646 16968 -1470
rect 17002 -1646 17014 -1470
rect 16956 -1658 17014 -1646
rect 17074 -1470 17132 -1458
rect 17074 -1646 17086 -1470
rect 17120 -1646 17132 -1470
rect 17074 -1658 17132 -1646
rect 17862 -1466 17920 -1454
rect 17862 -1642 17874 -1466
rect 17908 -1642 17920 -1466
rect 17862 -1654 17920 -1642
rect 17980 -1466 18038 -1454
rect 17980 -1642 17992 -1466
rect 18026 -1642 18038 -1466
rect 17980 -1654 18038 -1642
rect 18098 -1466 18156 -1454
rect 18098 -1642 18110 -1466
rect 18144 -1642 18156 -1466
rect 18098 -1654 18156 -1642
rect 18216 -1466 18274 -1454
rect 18216 -1642 18228 -1466
rect 18262 -1642 18274 -1466
rect 18216 -1654 18274 -1642
rect 13980 -2409 14038 -2397
rect 13980 -2585 13992 -2409
rect 14026 -2585 14038 -2409
rect 13980 -2597 14038 -2585
rect 14098 -2409 14156 -2397
rect 14098 -2585 14110 -2409
rect 14144 -2585 14156 -2409
rect 14098 -2597 14156 -2585
rect 14216 -2409 14274 -2397
rect 14216 -2585 14228 -2409
rect 14262 -2585 14274 -2409
rect 14216 -2597 14274 -2585
rect 14334 -2409 14392 -2397
rect 14334 -2585 14346 -2409
rect 14380 -2585 14392 -2409
rect 14334 -2597 14392 -2585
rect 14452 -2409 14510 -2397
rect 14452 -2585 14464 -2409
rect 14498 -2585 14510 -2409
rect 14452 -2597 14510 -2585
rect 14570 -2409 14628 -2397
rect 14570 -2585 14582 -2409
rect 14616 -2585 14628 -2409
rect 14570 -2597 14628 -2585
rect 14688 -2409 14746 -2397
rect 14688 -2585 14700 -2409
rect 14734 -2585 14746 -2409
rect 14688 -2597 14746 -2585
rect 14806 -2409 14864 -2397
rect 14806 -2585 14818 -2409
rect 14852 -2585 14864 -2409
rect 14806 -2597 14864 -2585
rect 14924 -2409 14982 -2397
rect 14924 -2585 14936 -2409
rect 14970 -2585 14982 -2409
rect 14924 -2597 14982 -2585
rect 15042 -2409 15100 -2397
rect 15042 -2585 15054 -2409
rect 15088 -2585 15100 -2409
rect 15042 -2597 15100 -2585
rect 15928 -2826 15986 -2814
rect 15444 -3026 15502 -3014
rect 15444 -3202 15456 -3026
rect 15490 -3202 15502 -3026
rect 15444 -3214 15502 -3202
rect 15562 -3026 15620 -3014
rect 15562 -3202 15574 -3026
rect 15608 -3202 15620 -3026
rect 15562 -3214 15620 -3202
rect 15680 -3026 15738 -3014
rect 15680 -3202 15692 -3026
rect 15726 -3202 15738 -3026
rect 15680 -3214 15738 -3202
rect 15798 -3026 15856 -3014
rect 15798 -3202 15810 -3026
rect 15844 -3202 15856 -3026
rect 15798 -3214 15856 -3202
rect 15928 -3202 15940 -2826
rect 15974 -3202 15986 -2826
rect 15928 -3214 15986 -3202
rect 16046 -2826 16104 -2814
rect 16046 -3202 16058 -2826
rect 16092 -3202 16104 -2826
rect 16046 -3214 16104 -3202
rect 16164 -2826 16222 -2814
rect 16164 -3202 16176 -2826
rect 16210 -3202 16222 -2826
rect 16164 -3214 16222 -3202
rect 16282 -2826 16340 -2814
rect 16282 -3202 16294 -2826
rect 16328 -3202 16340 -2826
rect 16282 -3214 16340 -3202
rect 16400 -2826 16458 -2814
rect 16400 -3202 16412 -2826
rect 16446 -3202 16458 -2826
rect 16400 -3214 16458 -3202
rect 16518 -2826 16576 -2814
rect 16518 -3202 16530 -2826
rect 16564 -3202 16576 -2826
rect 16518 -3214 16576 -3202
rect 16636 -2826 16694 -2814
rect 16636 -3202 16648 -2826
rect 16682 -3202 16694 -2826
rect 17826 -2826 17884 -2814
rect 16636 -3214 16694 -3202
rect 16765 -3026 16823 -3014
rect 16765 -3202 16777 -3026
rect 16811 -3202 16823 -3026
rect 16765 -3214 16823 -3202
rect 16883 -3026 16941 -3014
rect 16883 -3202 16895 -3026
rect 16929 -3202 16941 -3026
rect 16883 -3214 16941 -3202
rect 17001 -3026 17059 -3014
rect 17001 -3202 17013 -3026
rect 17047 -3202 17059 -3026
rect 17001 -3214 17059 -3202
rect 17119 -3026 17177 -3014
rect 17119 -3202 17131 -3026
rect 17165 -3202 17177 -3026
rect 17119 -3214 17177 -3202
rect 17342 -3026 17400 -3014
rect 17342 -3202 17354 -3026
rect 17388 -3202 17400 -3026
rect 17342 -3214 17400 -3202
rect 17460 -3026 17518 -3014
rect 17460 -3202 17472 -3026
rect 17506 -3202 17518 -3026
rect 17460 -3214 17518 -3202
rect 17578 -3026 17636 -3014
rect 17578 -3202 17590 -3026
rect 17624 -3202 17636 -3026
rect 17578 -3214 17636 -3202
rect 17696 -3026 17754 -3014
rect 17696 -3202 17708 -3026
rect 17742 -3202 17754 -3026
rect 17696 -3214 17754 -3202
rect 17826 -3202 17838 -2826
rect 17872 -3202 17884 -2826
rect 17826 -3214 17884 -3202
rect 17944 -2826 18002 -2814
rect 17944 -3202 17956 -2826
rect 17990 -3202 18002 -2826
rect 17944 -3214 18002 -3202
rect 18062 -2826 18120 -2814
rect 18062 -3202 18074 -2826
rect 18108 -3202 18120 -2826
rect 18062 -3214 18120 -3202
rect 18180 -2826 18238 -2814
rect 18180 -3202 18192 -2826
rect 18226 -3202 18238 -2826
rect 18180 -3214 18238 -3202
rect 18298 -2826 18356 -2814
rect 18298 -3202 18310 -2826
rect 18344 -3202 18356 -2826
rect 18298 -3214 18356 -3202
rect 18416 -2826 18474 -2814
rect 18416 -3202 18428 -2826
rect 18462 -3202 18474 -2826
rect 18416 -3214 18474 -3202
rect 18534 -2826 18592 -2814
rect 18534 -3202 18546 -2826
rect 18580 -3202 18592 -2826
rect 18534 -3214 18592 -3202
rect 18663 -3026 18721 -3014
rect 18663 -3202 18675 -3026
rect 18709 -3202 18721 -3026
rect 18663 -3214 18721 -3202
rect 18781 -3026 18839 -3014
rect 18781 -3202 18793 -3026
rect 18827 -3202 18839 -3026
rect 18781 -3214 18839 -3202
rect 18899 -3026 18957 -3014
rect 18899 -3202 18911 -3026
rect 18945 -3202 18957 -3026
rect 18899 -3214 18957 -3202
rect 19017 -3026 19075 -3014
rect 19017 -3202 19029 -3026
rect 19063 -3202 19075 -3026
rect 19017 -3214 19075 -3202
rect 13975 -4013 14033 -4001
rect 13975 -4189 13987 -4013
rect 14021 -4189 14033 -4013
rect 13975 -4201 14033 -4189
rect 14093 -4013 14151 -4001
rect 14093 -4189 14105 -4013
rect 14139 -4189 14151 -4013
rect 14093 -4201 14151 -4189
rect 14211 -4013 14269 -4001
rect 14211 -4189 14223 -4013
rect 14257 -4189 14269 -4013
rect 14211 -4201 14269 -4189
rect 14329 -4013 14387 -4001
rect 14329 -4189 14341 -4013
rect 14375 -4189 14387 -4013
rect 14329 -4201 14387 -4189
rect 14447 -4013 14505 -4001
rect 14447 -4189 14459 -4013
rect 14493 -4189 14505 -4013
rect 14447 -4201 14505 -4189
rect 14565 -4013 14623 -4001
rect 14565 -4189 14577 -4013
rect 14611 -4189 14623 -4013
rect 14565 -4201 14623 -4189
rect 14683 -4013 14741 -4001
rect 14683 -4189 14695 -4013
rect 14729 -4189 14741 -4013
rect 14683 -4201 14741 -4189
rect 14801 -4013 14859 -4001
rect 14801 -4189 14813 -4013
rect 14847 -4189 14859 -4013
rect 14801 -4201 14859 -4189
rect 14919 -4013 14977 -4001
rect 14919 -4189 14931 -4013
rect 14965 -4189 14977 -4013
rect 14919 -4201 14977 -4189
rect 15037 -4013 15095 -4001
rect 15037 -4189 15049 -4013
rect 15083 -4189 15095 -4013
rect 15037 -4201 15095 -4189
rect 15871 -3519 15929 -3507
rect 15871 -3895 15883 -3519
rect 15917 -3895 15929 -3519
rect 15871 -3907 15929 -3895
rect 15989 -3519 16047 -3507
rect 15989 -3895 16001 -3519
rect 16035 -3895 16047 -3519
rect 15989 -3907 16047 -3895
rect 16107 -3519 16165 -3507
rect 16107 -3895 16119 -3519
rect 16153 -3895 16165 -3519
rect 16107 -3907 16165 -3895
rect 16225 -3519 16283 -3507
rect 16225 -3895 16237 -3519
rect 16271 -3895 16283 -3519
rect 16225 -3907 16283 -3895
rect 16343 -3519 16401 -3507
rect 16343 -3895 16355 -3519
rect 16389 -3895 16401 -3519
rect 16343 -3907 16401 -3895
rect 16461 -3519 16519 -3507
rect 16461 -3895 16473 -3519
rect 16507 -3895 16519 -3519
rect 16461 -3907 16519 -3895
rect 16579 -3519 16637 -3507
rect 16579 -3895 16591 -3519
rect 16625 -3895 16637 -3519
rect 16579 -3907 16637 -3895
rect 17769 -3519 17827 -3507
rect 17769 -3895 17781 -3519
rect 17815 -3895 17827 -3519
rect 17769 -3907 17827 -3895
rect 17887 -3519 17945 -3507
rect 17887 -3895 17899 -3519
rect 17933 -3895 17945 -3519
rect 17887 -3907 17945 -3895
rect 18005 -3519 18063 -3507
rect 18005 -3895 18017 -3519
rect 18051 -3895 18063 -3519
rect 18005 -3907 18063 -3895
rect 18123 -3519 18181 -3507
rect 18123 -3895 18135 -3519
rect 18169 -3895 18181 -3519
rect 18123 -3907 18181 -3895
rect 18241 -3519 18299 -3507
rect 18241 -3895 18253 -3519
rect 18287 -3895 18299 -3519
rect 18241 -3907 18299 -3895
rect 18359 -3519 18417 -3507
rect 18359 -3895 18371 -3519
rect 18405 -3895 18417 -3519
rect 18359 -3907 18417 -3895
rect 18477 -3519 18535 -3507
rect 18477 -3895 18489 -3519
rect 18523 -3895 18535 -3519
rect 18477 -3907 18535 -3895
<< ndiffc >>
rect 14215 -1572 14249 -1196
rect 14333 -1572 14367 -1196
rect 14451 -1572 14485 -1196
rect 14568 -1372 14602 -1196
rect 14686 -1372 14720 -1196
rect 16213 -1646 16247 -1470
rect 16331 -1646 16365 -1470
rect 16449 -1646 16483 -1470
rect 16567 -1646 16601 -1470
rect 17355 -1642 17389 -1466
rect 17473 -1642 17507 -1466
rect 17591 -1642 17625 -1466
rect 17709 -1642 17743 -1466
rect 14229 -3222 14263 -2846
rect 14347 -3222 14381 -2846
rect 14465 -3222 14499 -2846
rect 14582 -3022 14616 -2846
rect 14700 -3022 14734 -2846
rect 15581 -4427 15615 -4251
rect 14224 -4826 14258 -4450
rect 14342 -4826 14376 -4450
rect 14460 -4826 14494 -4450
rect 14577 -4626 14611 -4450
rect 15699 -4427 15733 -4251
rect 14695 -4626 14729 -4450
rect 16001 -4627 16035 -4251
rect 16119 -4627 16153 -4251
rect 16237 -4627 16271 -4251
rect 16355 -4627 16389 -4251
rect 16473 -4627 16507 -4251
rect 16879 -4427 16913 -4251
rect 16997 -4427 17031 -4251
rect 17479 -4427 17513 -4251
rect 17597 -4427 17631 -4251
rect 17899 -4627 17933 -4251
rect 18017 -4627 18051 -4251
rect 18135 -4627 18169 -4251
rect 18253 -4627 18287 -4251
rect 18371 -4627 18405 -4251
rect 18777 -4427 18811 -4251
rect 18895 -4427 18929 -4251
<< pdiffc >>
rect 13978 -935 14012 -759
rect 14096 -935 14130 -759
rect 14214 -935 14248 -759
rect 14332 -935 14366 -759
rect 14450 -935 14484 -759
rect 14568 -935 14602 -759
rect 14686 -935 14720 -759
rect 14804 -935 14838 -759
rect 14922 -935 14956 -759
rect 15040 -935 15074 -759
rect 16303 -1063 16337 -687
rect 16421 -1063 16455 -687
rect 16539 -1063 16573 -687
rect 16657 -1063 16691 -687
rect 16775 -1063 16809 -687
rect 16893 -1063 16927 -687
rect 17011 -1063 17045 -687
rect 17445 -1059 17479 -683
rect 17563 -1059 17597 -683
rect 17681 -1059 17715 -683
rect 17799 -1059 17833 -683
rect 17917 -1059 17951 -683
rect 18035 -1059 18069 -683
rect 18153 -1059 18187 -683
rect 16732 -1646 16766 -1470
rect 16850 -1646 16884 -1470
rect 16968 -1646 17002 -1470
rect 17086 -1646 17120 -1470
rect 17874 -1642 17908 -1466
rect 17992 -1642 18026 -1466
rect 18110 -1642 18144 -1466
rect 18228 -1642 18262 -1466
rect 13992 -2585 14026 -2409
rect 14110 -2585 14144 -2409
rect 14228 -2585 14262 -2409
rect 14346 -2585 14380 -2409
rect 14464 -2585 14498 -2409
rect 14582 -2585 14616 -2409
rect 14700 -2585 14734 -2409
rect 14818 -2585 14852 -2409
rect 14936 -2585 14970 -2409
rect 15054 -2585 15088 -2409
rect 15456 -3202 15490 -3026
rect 15574 -3202 15608 -3026
rect 15692 -3202 15726 -3026
rect 15810 -3202 15844 -3026
rect 15940 -3202 15974 -2826
rect 16058 -3202 16092 -2826
rect 16176 -3202 16210 -2826
rect 16294 -3202 16328 -2826
rect 16412 -3202 16446 -2826
rect 16530 -3202 16564 -2826
rect 16648 -3202 16682 -2826
rect 16777 -3202 16811 -3026
rect 16895 -3202 16929 -3026
rect 17013 -3202 17047 -3026
rect 17131 -3202 17165 -3026
rect 17354 -3202 17388 -3026
rect 17472 -3202 17506 -3026
rect 17590 -3202 17624 -3026
rect 17708 -3202 17742 -3026
rect 17838 -3202 17872 -2826
rect 17956 -3202 17990 -2826
rect 18074 -3202 18108 -2826
rect 18192 -3202 18226 -2826
rect 18310 -3202 18344 -2826
rect 18428 -3202 18462 -2826
rect 18546 -3202 18580 -2826
rect 18675 -3202 18709 -3026
rect 18793 -3202 18827 -3026
rect 18911 -3202 18945 -3026
rect 19029 -3202 19063 -3026
rect 13987 -4189 14021 -4013
rect 14105 -4189 14139 -4013
rect 14223 -4189 14257 -4013
rect 14341 -4189 14375 -4013
rect 14459 -4189 14493 -4013
rect 14577 -4189 14611 -4013
rect 14695 -4189 14729 -4013
rect 14813 -4189 14847 -4013
rect 14931 -4189 14965 -4013
rect 15049 -4189 15083 -4013
rect 15883 -3895 15917 -3519
rect 16001 -3895 16035 -3519
rect 16119 -3895 16153 -3519
rect 16237 -3895 16271 -3519
rect 16355 -3895 16389 -3519
rect 16473 -3895 16507 -3519
rect 16591 -3895 16625 -3519
rect 17781 -3895 17815 -3519
rect 17899 -3895 17933 -3519
rect 18017 -3895 18051 -3519
rect 18135 -3895 18169 -3519
rect 18253 -3895 18287 -3519
rect 18371 -3895 18405 -3519
rect 18489 -3895 18523 -3519
<< psubdiff >>
rect 14739 -1522 14973 -1488
rect 14739 -1612 14785 -1522
rect 14948 -1612 14973 -1522
rect 14739 -1643 14973 -1612
rect 16236 -1893 16391 -1847
rect 16236 -2056 16267 -1893
rect 16357 -2056 16391 -1893
rect 16236 -2081 16391 -2056
rect 17378 -1895 17533 -1849
rect 17378 -2058 17409 -1895
rect 17499 -2058 17533 -1895
rect 17378 -2083 17533 -2058
rect 14753 -3172 14987 -3138
rect 14753 -3262 14799 -3172
rect 14962 -3262 14987 -3172
rect 14753 -3293 14987 -3262
rect 14748 -4776 14982 -4742
rect 14748 -4866 14794 -4776
rect 14957 -4866 14982 -4776
rect 14748 -4897 14982 -4866
rect 16180 -4936 16335 -4890
rect 16180 -5099 16211 -4936
rect 16301 -5099 16335 -4936
rect 16180 -5124 16335 -5099
<< nsubdiff >>
rect 16891 -291 17044 -251
rect 14409 -345 14562 -305
rect 14409 -494 14452 -345
rect 14519 -494 14562 -345
rect 14409 -563 14562 -494
rect 16891 -440 16934 -291
rect 17001 -440 17044 -291
rect 16891 -509 17044 -440
rect 18038 -291 18191 -251
rect 18038 -440 18081 -291
rect 18148 -440 18191 -291
rect 18038 -509 18191 -440
rect 14423 -1995 14576 -1955
rect 14423 -2144 14466 -1995
rect 14533 -2144 14576 -1995
rect 14423 -2213 14576 -2144
rect 18134 -2338 18287 -2298
rect 18134 -2487 18177 -2338
rect 18244 -2487 18287 -2338
rect 18134 -2556 18287 -2487
rect 14418 -3599 14571 -3559
rect 14418 -3748 14461 -3599
rect 14528 -3748 14571 -3599
rect 14418 -3817 14571 -3748
<< psubdiffcont >>
rect 14785 -1612 14948 -1522
rect 16267 -2056 16357 -1893
rect 17409 -2058 17499 -1895
rect 14799 -3262 14962 -3172
rect 14794 -4866 14957 -4776
rect 16211 -5099 16301 -4936
<< nsubdiffcont >>
rect 14452 -494 14519 -345
rect 16934 -440 17001 -291
rect 18081 -440 18148 -291
rect 14466 -2144 14533 -1995
rect 18177 -2487 18244 -2338
rect 14461 -3748 14528 -3599
<< poly >>
rect 16172 -511 16238 -495
rect 17302 -505 17368 -489
rect 16172 -545 16188 -511
rect 16222 -518 16238 -511
rect 16222 -545 16747 -518
rect 16172 -561 16747 -545
rect 17302 -539 17318 -505
rect 17352 -514 17368 -505
rect 17352 -539 17889 -514
rect 17302 -557 17889 -539
rect 16703 -613 16747 -561
rect 17845 -609 17889 -557
rect 16172 -629 16645 -613
rect 16172 -663 16188 -629
rect 16222 -654 16645 -629
rect 16222 -655 16409 -654
rect 16222 -663 16238 -655
rect 16172 -679 16238 -663
rect 16349 -675 16409 -655
rect 16467 -675 16527 -654
rect 16585 -675 16645 -654
rect 16703 -654 16999 -613
rect 16703 -675 16763 -654
rect 16821 -675 16881 -654
rect 16939 -675 16999 -654
rect 17302 -625 17787 -609
rect 17302 -659 17318 -625
rect 17352 -650 17787 -625
rect 17352 -651 17551 -650
rect 17352 -659 17368 -651
rect 17302 -675 17368 -659
rect 17491 -671 17551 -651
rect 17609 -671 17669 -650
rect 17727 -671 17787 -650
rect 17845 -650 18141 -609
rect 17845 -671 17905 -650
rect 17963 -671 18023 -650
rect 18081 -671 18141 -650
rect 14024 -726 14320 -690
rect 14024 -747 14084 -726
rect 14142 -747 14202 -726
rect 14260 -747 14320 -726
rect 14378 -727 14674 -691
rect 14378 -747 14438 -727
rect 14496 -747 14556 -727
rect 14614 -747 14674 -727
rect 14732 -727 15028 -691
rect 14732 -747 14792 -727
rect 14850 -747 14910 -727
rect 14968 -747 15028 -727
rect 14024 -973 14084 -947
rect 14142 -973 14202 -947
rect 14260 -973 14320 -947
rect 14378 -967 14438 -947
rect 14378 -973 14439 -967
rect 14496 -973 14556 -947
rect 14614 -973 14674 -947
rect 14261 -1158 14319 -973
rect 14261 -1184 14321 -1158
rect 14379 -1184 14439 -973
rect 14732 -979 14792 -947
rect 14850 -973 14910 -947
rect 14968 -973 15028 -947
rect 14729 -995 14795 -979
rect 14729 -1029 14745 -995
rect 14779 -1029 14795 -995
rect 14729 -1045 14795 -1029
rect 16349 -1092 16409 -1075
rect 14611 -1112 14677 -1096
rect 14611 -1146 14627 -1112
rect 14661 -1146 14677 -1112
rect 14611 -1162 14677 -1146
rect 14614 -1184 14674 -1162
rect 16349 -1181 16410 -1092
rect 16467 -1101 16527 -1075
rect 16585 -1101 16645 -1075
rect 16259 -1234 16410 -1181
rect 14614 -1410 14674 -1384
rect 16259 -1458 16319 -1234
rect 16703 -1276 16763 -1075
rect 16821 -1101 16881 -1075
rect 16939 -1101 16999 -1075
rect 17491 -1088 17551 -1071
rect 17491 -1177 17552 -1088
rect 17609 -1097 17669 -1071
rect 17727 -1097 17787 -1071
rect 16377 -1327 16763 -1276
rect 17401 -1230 17552 -1177
rect 16377 -1458 16437 -1327
rect 16492 -1385 16558 -1369
rect 16492 -1419 16508 -1385
rect 16542 -1419 16558 -1385
rect 16492 -1435 16558 -1419
rect 16495 -1458 16555 -1435
rect 16778 -1458 16838 -1432
rect 16896 -1458 16956 -1432
rect 17014 -1458 17074 -1432
rect 17401 -1454 17461 -1230
rect 17845 -1272 17905 -1071
rect 17963 -1097 18023 -1071
rect 18081 -1097 18141 -1071
rect 17519 -1323 17905 -1272
rect 17519 -1454 17579 -1323
rect 17634 -1381 17700 -1365
rect 17634 -1415 17650 -1381
rect 17684 -1415 17700 -1381
rect 17634 -1431 17700 -1415
rect 17637 -1454 17697 -1431
rect 17920 -1454 17980 -1428
rect 18038 -1454 18098 -1428
rect 18156 -1454 18216 -1428
rect 14261 -1606 14321 -1584
rect 14379 -1606 14439 -1584
rect 14258 -1622 14324 -1606
rect 14258 -1656 14274 -1622
rect 14308 -1656 14324 -1622
rect 14258 -1672 14324 -1656
rect 14376 -1622 14442 -1606
rect 14376 -1656 14392 -1622
rect 14426 -1656 14442 -1622
rect 14376 -1672 14442 -1656
rect 16259 -1684 16319 -1658
rect 16377 -1684 16437 -1658
rect 16495 -1690 16555 -1658
rect 16778 -1690 16838 -1658
rect 16896 -1690 16956 -1658
rect 17014 -1690 17074 -1658
rect 17401 -1680 17461 -1654
rect 17519 -1680 17579 -1654
rect 16495 -1731 17074 -1690
rect 17637 -1686 17697 -1654
rect 17920 -1686 17980 -1654
rect 18038 -1686 18098 -1654
rect 18156 -1686 18216 -1654
rect 17637 -1727 18216 -1686
rect 14038 -2376 14334 -2340
rect 14038 -2397 14098 -2376
rect 14156 -2397 14216 -2376
rect 14274 -2397 14334 -2376
rect 14392 -2377 14688 -2341
rect 14392 -2397 14452 -2377
rect 14510 -2397 14570 -2377
rect 14628 -2397 14688 -2377
rect 14746 -2377 15042 -2341
rect 14746 -2397 14806 -2377
rect 14864 -2397 14924 -2377
rect 14982 -2397 15042 -2377
rect 14038 -2623 14098 -2597
rect 14156 -2623 14216 -2597
rect 14274 -2623 14334 -2597
rect 14392 -2617 14452 -2597
rect 14392 -2623 14453 -2617
rect 14510 -2623 14570 -2597
rect 14628 -2623 14688 -2597
rect 14275 -2808 14333 -2623
rect 14275 -2834 14335 -2808
rect 14393 -2834 14453 -2623
rect 14746 -2629 14806 -2597
rect 14864 -2623 14924 -2597
rect 14982 -2623 15042 -2597
rect 14743 -2645 14809 -2629
rect 14743 -2679 14759 -2645
rect 14793 -2679 14809 -2645
rect 14743 -2695 14809 -2679
rect 14625 -2762 14691 -2746
rect 14625 -2796 14641 -2762
rect 14675 -2796 14691 -2762
rect 14625 -2812 14691 -2796
rect 15986 -2799 16282 -2748
rect 14628 -2834 14688 -2812
rect 15986 -2814 16046 -2799
rect 16104 -2814 16164 -2799
rect 16222 -2814 16282 -2799
rect 16340 -2814 16400 -2788
rect 16458 -2814 16518 -2788
rect 16576 -2814 16636 -2788
rect 17884 -2799 18180 -2748
rect 17884 -2814 17944 -2799
rect 18002 -2814 18062 -2799
rect 18120 -2814 18180 -2799
rect 18238 -2814 18298 -2788
rect 18356 -2814 18416 -2788
rect 18474 -2814 18534 -2788
rect 15502 -3014 15562 -2988
rect 15620 -3014 15680 -2988
rect 15738 -3014 15798 -2988
rect 14628 -3060 14688 -3034
rect 14275 -3256 14335 -3234
rect 14393 -3250 14453 -3234
rect 14272 -3272 14338 -3256
rect 14272 -3306 14288 -3272
rect 14322 -3306 14338 -3272
rect 14272 -3322 14338 -3306
rect 14387 -3272 14461 -3250
rect 14387 -3306 14406 -3272
rect 14440 -3306 14461 -3272
rect 16823 -2997 17119 -2946
rect 16823 -3014 16883 -2997
rect 16941 -3014 17001 -2997
rect 17059 -3014 17119 -2997
rect 17400 -3014 17460 -2988
rect 17518 -3014 17578 -2988
rect 17636 -3014 17696 -2988
rect 18721 -2997 19017 -2946
rect 18721 -3014 18781 -2997
rect 18839 -3014 18899 -2997
rect 18957 -3014 19017 -2997
rect 15502 -3231 15562 -3214
rect 15620 -3231 15680 -3214
rect 15738 -3231 15798 -3214
rect 15986 -3231 16046 -3214
rect 15502 -3282 16046 -3231
rect 16104 -3240 16164 -3214
rect 16222 -3240 16282 -3214
rect 16340 -3233 16400 -3214
rect 16458 -3233 16518 -3214
rect 16576 -3233 16636 -3214
rect 16823 -3233 16883 -3214
rect 16941 -3233 17001 -3214
rect 14387 -3363 14461 -3306
rect 15627 -3363 15687 -3282
rect 16340 -3284 16883 -3233
rect 16925 -3240 17001 -3233
rect 17059 -3240 17119 -3214
rect 17400 -3231 17460 -3214
rect 17518 -3231 17578 -3214
rect 17636 -3231 17696 -3214
rect 17884 -3231 17944 -3214
rect 16925 -3284 17000 -3240
rect 17400 -3282 17944 -3231
rect 18002 -3240 18062 -3214
rect 18120 -3240 18180 -3214
rect 18238 -3233 18298 -3214
rect 18356 -3233 18416 -3214
rect 18474 -3233 18534 -3214
rect 18721 -3233 18781 -3214
rect 18839 -3233 18899 -3214
rect 14387 -3388 15687 -3363
rect 14386 -3436 15687 -3388
rect 16925 -3404 16985 -3284
rect 14033 -3980 14329 -3944
rect 14033 -4001 14093 -3980
rect 14151 -4001 14211 -3980
rect 14269 -4001 14329 -3980
rect 14387 -3981 14683 -3945
rect 14387 -4001 14447 -3981
rect 14505 -4001 14565 -3981
rect 14623 -4001 14683 -3981
rect 14741 -3981 15037 -3945
rect 14741 -4001 14801 -3981
rect 14859 -4001 14919 -3981
rect 14977 -4001 15037 -3981
rect 15627 -4134 15687 -3436
rect 15929 -3484 16225 -3424
rect 15929 -3507 15989 -3484
rect 16047 -3507 16107 -3484
rect 16165 -3507 16225 -3484
rect 16283 -3483 16579 -3423
rect 16924 -3424 16985 -3404
rect 16283 -3507 16343 -3483
rect 16401 -3507 16461 -3483
rect 16519 -3507 16579 -3483
rect 16905 -3440 16985 -3424
rect 16905 -3474 16920 -3440
rect 16954 -3474 16985 -3440
rect 16905 -3490 16985 -3474
rect 16924 -3513 16985 -3490
rect 16925 -3659 16985 -3513
rect 16924 -3832 16985 -3659
rect 15929 -3933 15989 -3907
rect 15897 -4074 15964 -4067
rect 16047 -4074 16107 -3907
rect 16165 -3933 16225 -3907
rect 16283 -3933 16343 -3907
rect 15897 -4083 16107 -4074
rect 15897 -4117 15913 -4083
rect 15947 -4117 16107 -4083
rect 15897 -4133 16107 -4117
rect 15627 -4150 15778 -4134
rect 15627 -4184 15728 -4150
rect 15762 -4184 15778 -4150
rect 15627 -4200 15778 -4184
rect 14033 -4227 14093 -4201
rect 14151 -4227 14211 -4201
rect 14269 -4227 14329 -4201
rect 14387 -4221 14447 -4201
rect 14387 -4227 14448 -4221
rect 14505 -4227 14565 -4201
rect 14623 -4227 14683 -4201
rect 14270 -4412 14328 -4227
rect 14270 -4438 14330 -4412
rect 14388 -4438 14448 -4227
rect 14741 -4233 14801 -4201
rect 14859 -4227 14919 -4201
rect 14977 -4227 15037 -4201
rect 14738 -4249 14804 -4233
rect 15627 -4239 15687 -4200
rect 16047 -4239 16107 -4133
rect 16401 -4074 16461 -3907
rect 16519 -3933 16579 -3907
rect 16544 -4074 16611 -4067
rect 16401 -4083 16611 -4074
rect 16401 -4117 16561 -4083
rect 16595 -4117 16611 -4083
rect 16401 -4133 16611 -4117
rect 16163 -4167 16229 -4151
rect 16163 -4201 16179 -4167
rect 16213 -4201 16229 -4167
rect 16163 -4217 16229 -4201
rect 16281 -4166 16347 -4151
rect 16281 -4200 16297 -4166
rect 16331 -4200 16347 -4166
rect 16281 -4216 16347 -4200
rect 16165 -4239 16225 -4217
rect 16283 -4239 16343 -4216
rect 16401 -4239 16461 -4133
rect 16925 -4135 16985 -3832
rect 16835 -4151 16985 -4135
rect 16835 -4185 16851 -4151
rect 16885 -4185 16985 -4151
rect 16835 -4201 16985 -4185
rect 16925 -4239 16985 -4201
rect 17525 -3940 17585 -3282
rect 18238 -3284 18781 -3233
rect 18823 -3240 18899 -3233
rect 18957 -3240 19017 -3214
rect 18823 -3284 18898 -3240
rect 17827 -3484 18123 -3424
rect 17827 -3507 17887 -3484
rect 17945 -3507 18005 -3484
rect 18063 -3507 18123 -3484
rect 18181 -3483 18477 -3423
rect 18181 -3507 18241 -3483
rect 18299 -3507 18359 -3483
rect 18417 -3507 18477 -3483
rect 18823 -3437 18883 -3284
rect 18823 -3461 19077 -3437
rect 18823 -3495 19027 -3461
rect 19061 -3495 19077 -3461
rect 18823 -3511 19077 -3495
rect 17827 -3933 17887 -3907
rect 17525 -3956 17592 -3940
rect 17525 -3990 17541 -3956
rect 17575 -3990 17592 -3956
rect 17525 -4006 17592 -3990
rect 17525 -4134 17585 -4006
rect 17795 -4074 17862 -4067
rect 17945 -4074 18005 -3907
rect 18063 -3933 18123 -3907
rect 18181 -3933 18241 -3907
rect 17795 -4083 18005 -4074
rect 17795 -4117 17811 -4083
rect 17845 -4117 18005 -4083
rect 17795 -4133 18005 -4117
rect 17525 -4150 17676 -4134
rect 17525 -4184 17626 -4150
rect 17660 -4184 17676 -4150
rect 17525 -4200 17676 -4184
rect 17525 -4239 17585 -4200
rect 17945 -4239 18005 -4133
rect 18299 -4074 18359 -3907
rect 18417 -3933 18477 -3907
rect 18440 -4073 18507 -4066
rect 18434 -4074 18507 -4073
rect 18299 -4082 18507 -4074
rect 18299 -4116 18457 -4082
rect 18491 -4116 18507 -4082
rect 18299 -4132 18507 -4116
rect 18299 -4133 18496 -4132
rect 18061 -4167 18127 -4151
rect 18061 -4201 18077 -4167
rect 18111 -4201 18127 -4167
rect 18061 -4217 18127 -4201
rect 18179 -4166 18245 -4151
rect 18179 -4200 18195 -4166
rect 18229 -4200 18245 -4166
rect 18179 -4216 18245 -4200
rect 18063 -4239 18123 -4217
rect 18181 -4239 18241 -4216
rect 18299 -4239 18359 -4133
rect 18823 -4135 18883 -3511
rect 18733 -4151 18883 -4135
rect 18733 -4185 18749 -4151
rect 18783 -4185 18883 -4151
rect 18733 -4201 18883 -4185
rect 18823 -4239 18883 -4201
rect 14738 -4283 14754 -4249
rect 14788 -4283 14804 -4249
rect 14738 -4299 14804 -4283
rect 14620 -4366 14686 -4350
rect 14620 -4400 14636 -4366
rect 14670 -4400 14686 -4366
rect 14620 -4416 14686 -4400
rect 14623 -4438 14683 -4416
rect 15627 -4465 15687 -4439
rect 14623 -4664 14683 -4638
rect 16925 -4465 16985 -4439
rect 17525 -4465 17585 -4439
rect 18823 -4465 18883 -4439
rect 16047 -4665 16107 -4639
rect 16165 -4665 16225 -4639
rect 16283 -4665 16343 -4639
rect 16401 -4665 16461 -4639
rect 17945 -4665 18005 -4639
rect 18063 -4665 18123 -4639
rect 18181 -4665 18241 -4639
rect 18299 -4665 18359 -4639
rect 14270 -4860 14330 -4838
rect 14388 -4860 14448 -4838
rect 14267 -4876 14333 -4860
rect 14267 -4910 14283 -4876
rect 14317 -4910 14333 -4876
rect 14267 -4926 14333 -4910
rect 14385 -4876 14451 -4860
rect 14385 -4910 14401 -4876
rect 14435 -4910 14451 -4876
rect 14385 -4926 14451 -4910
<< polycont >>
rect 16188 -545 16222 -511
rect 17318 -539 17352 -505
rect 16188 -663 16222 -629
rect 17318 -659 17352 -625
rect 14745 -1029 14779 -995
rect 14627 -1146 14661 -1112
rect 16508 -1419 16542 -1385
rect 17650 -1415 17684 -1381
rect 14274 -1656 14308 -1622
rect 14392 -1656 14426 -1622
rect 14759 -2679 14793 -2645
rect 14641 -2796 14675 -2762
rect 14288 -3306 14322 -3272
rect 14406 -3306 14440 -3272
rect 16920 -3474 16954 -3440
rect 15913 -4117 15947 -4083
rect 15728 -4184 15762 -4150
rect 16561 -4117 16595 -4083
rect 16179 -4201 16213 -4167
rect 16297 -4200 16331 -4166
rect 16851 -4185 16885 -4151
rect 19027 -3495 19061 -3461
rect 17541 -3990 17575 -3956
rect 17811 -4117 17845 -4083
rect 17626 -4184 17660 -4150
rect 18457 -4116 18491 -4082
rect 18077 -4201 18111 -4167
rect 18195 -4200 18229 -4166
rect 18749 -4185 18783 -4151
rect 14754 -4283 14788 -4249
rect 14636 -4400 14670 -4366
rect 14283 -4910 14317 -4876
rect 14401 -4910 14435 -4876
<< locali >>
rect 14373 -345 14596 -269
rect 14373 -494 14452 -345
rect 14519 -494 14596 -345
rect 14373 -600 14596 -494
rect 16855 -291 17078 -215
rect 16855 -440 16934 -291
rect 17001 -440 17078 -291
rect 16188 -511 16222 -495
rect 16188 -561 16222 -545
rect 16855 -546 17078 -440
rect 18002 -291 18225 -215
rect 18002 -440 18081 -291
rect 18148 -440 18225 -291
rect 17318 -505 17352 -489
rect 17318 -555 17352 -539
rect 18002 -546 18225 -440
rect 16188 -629 16222 -613
rect 14804 -709 15074 -675
rect 16188 -679 16222 -663
rect 17318 -625 17352 -609
rect 13978 -759 14012 -743
rect 13978 -951 14012 -935
rect 14096 -759 14130 -743
rect 14096 -951 14130 -935
rect 14214 -759 14248 -743
rect 14214 -951 14248 -935
rect 14332 -759 14366 -743
rect 14332 -951 14366 -935
rect 14450 -759 14484 -743
rect 14450 -951 14484 -935
rect 14568 -759 14602 -743
rect 14568 -951 14602 -935
rect 14686 -759 14720 -743
rect 14686 -951 14720 -935
rect 14804 -759 14838 -709
rect 14804 -951 14838 -935
rect 14922 -759 14956 -743
rect 14922 -951 14956 -935
rect 15040 -759 15074 -709
rect 15040 -951 15074 -935
rect 16303 -687 16337 -671
rect 14729 -1029 14745 -995
rect 14779 -1029 14795 -995
rect 16303 -1079 16337 -1063
rect 16421 -687 16455 -671
rect 16421 -1079 16455 -1063
rect 16539 -687 16573 -671
rect 16539 -1079 16573 -1063
rect 16657 -687 16691 -671
rect 16657 -1079 16691 -1063
rect 16775 -687 16809 -671
rect 16775 -1079 16809 -1063
rect 16893 -687 16927 -671
rect 16893 -1079 16927 -1063
rect 17011 -687 17045 -671
rect 17318 -675 17352 -659
rect 17011 -1079 17045 -1063
rect 17445 -683 17479 -667
rect 17445 -1075 17479 -1059
rect 17563 -683 17597 -667
rect 17563 -1075 17597 -1059
rect 17681 -683 17715 -667
rect 17681 -1075 17715 -1059
rect 17799 -683 17833 -667
rect 17799 -1075 17833 -1059
rect 17917 -683 17951 -667
rect 17917 -1075 17951 -1059
rect 18035 -683 18069 -667
rect 18035 -1075 18069 -1059
rect 18153 -683 18187 -667
rect 18153 -1075 18187 -1059
rect 14611 -1146 14627 -1112
rect 14661 -1146 14677 -1112
rect 14215 -1196 14249 -1180
rect 14215 -1588 14249 -1572
rect 14333 -1196 14367 -1180
rect 14333 -1588 14367 -1572
rect 14451 -1196 14485 -1180
rect 14568 -1196 14602 -1180
rect 14568 -1388 14602 -1372
rect 14686 -1196 14720 -1180
rect 14686 -1388 14720 -1372
rect 16492 -1419 16508 -1385
rect 16542 -1419 16558 -1385
rect 17634 -1415 17650 -1381
rect 17684 -1415 17700 -1381
rect 16213 -1470 16247 -1454
rect 14451 -1588 14485 -1572
rect 14738 -1522 14987 -1479
rect 14738 -1612 14785 -1522
rect 14948 -1612 14987 -1522
rect 14258 -1656 14274 -1622
rect 14308 -1656 14324 -1622
rect 14376 -1656 14392 -1622
rect 14426 -1656 14442 -1622
rect 14738 -1651 14987 -1612
rect 16213 -1662 16247 -1646
rect 16331 -1470 16365 -1454
rect 16331 -1662 16365 -1646
rect 16449 -1470 16483 -1454
rect 16449 -1662 16483 -1646
rect 16567 -1470 16601 -1454
rect 16567 -1662 16601 -1646
rect 16732 -1470 16766 -1454
rect 16732 -1662 16766 -1646
rect 16850 -1470 16884 -1454
rect 16850 -1662 16884 -1646
rect 16968 -1470 17002 -1454
rect 16968 -1662 17002 -1646
rect 17086 -1470 17120 -1454
rect 17086 -1662 17120 -1646
rect 17355 -1466 17389 -1450
rect 17355 -1658 17389 -1642
rect 17473 -1466 17507 -1450
rect 17473 -1658 17507 -1642
rect 17591 -1466 17625 -1450
rect 17591 -1658 17625 -1642
rect 17709 -1466 17743 -1450
rect 17709 -1658 17743 -1642
rect 17874 -1466 17908 -1450
rect 17874 -1658 17908 -1642
rect 17992 -1466 18026 -1450
rect 17992 -1658 18026 -1642
rect 18110 -1466 18144 -1450
rect 18110 -1658 18144 -1642
rect 18228 -1466 18262 -1450
rect 18228 -1658 18262 -1642
rect 16228 -1893 16400 -1846
rect 14387 -1995 14610 -1919
rect 14387 -2144 14466 -1995
rect 14533 -2144 14610 -1995
rect 16228 -2056 16267 -1893
rect 16357 -2056 16400 -1893
rect 16228 -2095 16400 -2056
rect 17370 -1895 17542 -1848
rect 17370 -2058 17409 -1895
rect 17499 -2058 17542 -1895
rect 17370 -2097 17542 -2058
rect 14387 -2250 14610 -2144
rect 14818 -2359 15088 -2325
rect 13992 -2409 14026 -2393
rect 13992 -2601 14026 -2585
rect 14110 -2409 14144 -2393
rect 14110 -2601 14144 -2585
rect 14228 -2409 14262 -2393
rect 14228 -2601 14262 -2585
rect 14346 -2409 14380 -2393
rect 14346 -2601 14380 -2585
rect 14464 -2409 14498 -2393
rect 14464 -2601 14498 -2585
rect 14582 -2409 14616 -2393
rect 14582 -2601 14616 -2585
rect 14700 -2409 14734 -2393
rect 14700 -2601 14734 -2585
rect 14818 -2409 14852 -2359
rect 14818 -2601 14852 -2585
rect 14936 -2409 14970 -2393
rect 14936 -2601 14970 -2585
rect 15054 -2409 15088 -2359
rect 15054 -2601 15088 -2585
rect 18098 -2338 18323 -2262
rect 18098 -2487 18177 -2338
rect 18244 -2487 18323 -2338
rect 18098 -2593 18323 -2487
rect 14743 -2679 14759 -2645
rect 14793 -2679 14809 -2645
rect 14625 -2796 14641 -2762
rect 14675 -2796 14691 -2762
rect 16294 -2773 16564 -2738
rect 15940 -2826 15974 -2810
rect 14229 -2846 14263 -2830
rect 14229 -3238 14263 -3222
rect 14347 -2846 14381 -2830
rect 14347 -3238 14381 -3222
rect 14465 -2846 14499 -2830
rect 14582 -2846 14616 -2830
rect 14582 -3038 14616 -3022
rect 14700 -2846 14734 -2830
rect 14700 -3038 14734 -3022
rect 15456 -2972 15726 -2937
rect 15456 -3026 15490 -2972
rect 14465 -3238 14499 -3222
rect 14752 -3172 15001 -3129
rect 14752 -3262 14799 -3172
rect 14962 -3262 15001 -3172
rect 15456 -3218 15490 -3202
rect 15574 -3026 15608 -3010
rect 15574 -3218 15608 -3202
rect 15692 -3026 15726 -2972
rect 15692 -3218 15726 -3202
rect 15810 -3026 15844 -3010
rect 15810 -3218 15844 -3202
rect 15940 -3218 15974 -3202
rect 16058 -2826 16092 -2810
rect 16058 -3218 16092 -3202
rect 16176 -2826 16210 -2810
rect 16176 -3218 16210 -3202
rect 16294 -2826 16328 -2773
rect 16294 -3218 16328 -3202
rect 16412 -2826 16446 -2810
rect 16412 -3218 16446 -3202
rect 16530 -2826 16564 -2773
rect 18192 -2773 18462 -2738
rect 16530 -3218 16564 -3202
rect 16648 -2826 16682 -2810
rect 17838 -2826 17872 -2810
rect 17354 -2972 17624 -2937
rect 16648 -3218 16682 -3202
rect 16777 -3026 16811 -3010
rect 16777 -3218 16811 -3202
rect 16895 -3026 16929 -3010
rect 16895 -3218 16929 -3202
rect 17013 -3026 17047 -3010
rect 17013 -3218 17047 -3202
rect 17131 -3026 17165 -3010
rect 17131 -3218 17165 -3202
rect 17354 -3026 17388 -2972
rect 17354 -3218 17388 -3202
rect 17472 -3026 17506 -3010
rect 17472 -3218 17506 -3202
rect 17590 -3026 17624 -2972
rect 17590 -3218 17624 -3202
rect 17708 -3026 17742 -3010
rect 17708 -3218 17742 -3202
rect 17838 -3218 17872 -3202
rect 17956 -2826 17990 -2810
rect 17956 -3218 17990 -3202
rect 18074 -2826 18108 -2810
rect 18074 -3218 18108 -3202
rect 18192 -2826 18226 -2773
rect 18192 -3218 18226 -3202
rect 18310 -2826 18344 -2810
rect 18310 -3218 18344 -3202
rect 18428 -2826 18462 -2773
rect 18428 -3218 18462 -3202
rect 18546 -2826 18580 -2810
rect 18546 -3218 18580 -3202
rect 18675 -3026 18709 -3010
rect 18675 -3218 18709 -3202
rect 18793 -3026 18827 -3010
rect 18793 -3218 18827 -3202
rect 18911 -3026 18945 -3010
rect 18911 -3218 18945 -3202
rect 19029 -3026 19063 -3010
rect 19029 -3218 19063 -3202
rect 14272 -3306 14288 -3272
rect 14322 -3306 14338 -3272
rect 14390 -3306 14406 -3272
rect 14440 -3306 14456 -3272
rect 14752 -3301 15001 -3262
rect 16920 -3440 16954 -3424
rect 16920 -3490 16954 -3474
rect 19010 -3461 19077 -3445
rect 19010 -3495 19027 -3461
rect 19061 -3495 19077 -3461
rect 15883 -3519 15917 -3503
rect 14382 -3599 14605 -3523
rect 14382 -3748 14461 -3599
rect 14528 -3748 14605 -3599
rect 14382 -3854 14605 -3748
rect 16001 -3519 16035 -3503
rect 15883 -3911 15917 -3895
rect 16000 -3895 16001 -3848
rect 16119 -3519 16153 -3503
rect 16035 -3895 16036 -3848
rect 14813 -3963 15083 -3929
rect 13987 -4013 14021 -3997
rect 13987 -4205 14021 -4189
rect 14105 -4013 14139 -3997
rect 14105 -4205 14139 -4189
rect 14223 -4013 14257 -3997
rect 14223 -4205 14257 -4189
rect 14341 -4013 14375 -3997
rect 14341 -4205 14375 -4189
rect 14459 -4013 14493 -3997
rect 14459 -4205 14493 -4189
rect 14577 -4013 14611 -3997
rect 14577 -4205 14611 -4189
rect 14695 -4013 14729 -3997
rect 14695 -4205 14729 -4189
rect 14813 -4013 14847 -3963
rect 14813 -4205 14847 -4189
rect 14931 -4013 14965 -3997
rect 14931 -4205 14965 -4189
rect 15049 -4013 15083 -3963
rect 16000 -3953 16036 -3895
rect 16237 -3519 16271 -3503
rect 16119 -3911 16153 -3895
rect 16235 -3895 16237 -3848
rect 16235 -3953 16271 -3895
rect 16355 -3519 16389 -3503
rect 16355 -3911 16389 -3895
rect 16473 -3519 16507 -3503
rect 16591 -3519 16625 -3503
rect 16507 -3895 16509 -3849
rect 16473 -3953 16509 -3895
rect 16591 -3911 16625 -3895
rect 17781 -3519 17815 -3503
rect 17899 -3519 17933 -3503
rect 17781 -3911 17815 -3895
rect 17898 -3895 17899 -3848
rect 18017 -3519 18051 -3503
rect 17933 -3895 17934 -3848
rect 17096 -3953 17593 -3935
rect 16000 -3956 17593 -3953
rect 16000 -3990 17541 -3956
rect 17575 -3990 17593 -3956
rect 16000 -3993 17593 -3990
rect 17898 -3953 17934 -3895
rect 18135 -3519 18169 -3503
rect 18017 -3911 18051 -3895
rect 18133 -3895 18135 -3848
rect 18133 -3953 18169 -3895
rect 18253 -3519 18287 -3503
rect 18253 -3911 18287 -3895
rect 18371 -3519 18405 -3503
rect 18489 -3519 18523 -3503
rect 19010 -3511 19077 -3495
rect 18405 -3895 18407 -3849
rect 18371 -3953 18407 -3895
rect 18489 -3911 18523 -3895
rect 18994 -3924 19094 -3923
rect 18994 -3953 19150 -3924
rect 17898 -3993 19150 -3953
rect 16019 -3994 17593 -3993
rect 17917 -3994 19150 -3993
rect 15897 -4083 15964 -4067
rect 15897 -4117 15913 -4083
rect 15947 -4117 15964 -4083
rect 15897 -4133 15964 -4117
rect 15049 -4205 15083 -4189
rect 15728 -4150 15762 -4134
rect 15728 -4200 15762 -4184
rect 16074 -4235 16108 -3994
rect 17096 -4011 17593 -3994
rect 16544 -4083 16611 -4067
rect 16544 -4117 16561 -4083
rect 16595 -4117 16611 -4083
rect 16544 -4133 16611 -4117
rect 17795 -4083 17862 -4067
rect 17795 -4117 17811 -4083
rect 17845 -4117 17862 -4083
rect 17795 -4133 17862 -4117
rect 16851 -4151 16885 -4135
rect 16163 -4201 16179 -4167
rect 16213 -4201 16229 -4167
rect 16281 -4200 16297 -4166
rect 16331 -4200 16347 -4166
rect 16851 -4201 16885 -4185
rect 17626 -4150 17660 -4134
rect 17626 -4200 17660 -4184
rect 17972 -4235 18006 -3994
rect 18994 -4022 19150 -3994
rect 18994 -4023 19094 -4022
rect 18440 -4082 18507 -4066
rect 18440 -4116 18457 -4082
rect 18491 -4116 18507 -4082
rect 18440 -4132 18507 -4116
rect 18749 -4151 18783 -4135
rect 18061 -4201 18077 -4167
rect 18111 -4201 18127 -4167
rect 18179 -4200 18195 -4166
rect 18229 -4200 18245 -4166
rect 18749 -4201 18783 -4185
rect 14738 -4283 14754 -4249
rect 14788 -4283 14804 -4249
rect 15581 -4251 15615 -4235
rect 14620 -4400 14636 -4366
rect 14670 -4400 14686 -4366
rect 14224 -4450 14258 -4434
rect 14224 -4842 14258 -4826
rect 14342 -4450 14376 -4434
rect 14342 -4842 14376 -4826
rect 14460 -4450 14494 -4434
rect 14577 -4450 14611 -4434
rect 14577 -4642 14611 -4626
rect 14695 -4450 14729 -4434
rect 15581 -4443 15615 -4427
rect 15699 -4251 15733 -4235
rect 15699 -4443 15733 -4427
rect 16001 -4251 16035 -4235
rect 14695 -4642 14729 -4626
rect 16074 -4251 16153 -4235
rect 16074 -4281 16119 -4251
rect 16001 -4694 16036 -4627
rect 16119 -4643 16153 -4627
rect 16237 -4251 16271 -4235
rect 16237 -4643 16271 -4627
rect 16355 -4251 16389 -4235
rect 16473 -4251 16507 -4235
rect 16879 -4251 16913 -4235
rect 16879 -4443 16913 -4427
rect 16997 -4251 17031 -4235
rect 16997 -4443 17031 -4427
rect 17479 -4251 17513 -4235
rect 17479 -4443 17513 -4427
rect 17597 -4251 17631 -4235
rect 17597 -4443 17631 -4427
rect 17899 -4251 17933 -4235
rect 16355 -4643 16389 -4627
rect 16472 -4694 16507 -4627
rect 16001 -4729 16507 -4694
rect 17972 -4251 18051 -4235
rect 17972 -4281 18017 -4251
rect 17899 -4694 17934 -4627
rect 18017 -4643 18051 -4627
rect 18135 -4251 18169 -4235
rect 18135 -4643 18169 -4627
rect 18253 -4251 18287 -4235
rect 18371 -4251 18405 -4235
rect 18777 -4251 18811 -4235
rect 18777 -4443 18811 -4427
rect 18895 -4251 18929 -4235
rect 18895 -4443 18929 -4427
rect 18253 -4643 18287 -4627
rect 18370 -4694 18405 -4627
rect 17899 -4729 18405 -4694
rect 14460 -4842 14494 -4826
rect 14747 -4776 14996 -4733
rect 14747 -4866 14794 -4776
rect 14957 -4866 14996 -4776
rect 14267 -4910 14283 -4876
rect 14317 -4910 14333 -4876
rect 14385 -4910 14401 -4876
rect 14435 -4910 14451 -4876
rect 14747 -4905 14996 -4866
rect 16172 -4936 16344 -4889
rect 16172 -5099 16211 -4936
rect 16301 -5099 16344 -4936
rect 16172 -5139 16344 -5099
<< viali >>
rect 16188 -545 16222 -511
rect 17318 -539 17352 -505
rect 16188 -663 16222 -629
rect 17318 -659 17352 -625
rect 13978 -935 14012 -759
rect 14096 -935 14130 -759
rect 14214 -935 14248 -759
rect 14332 -935 14366 -759
rect 14450 -935 14484 -759
rect 14568 -935 14602 -759
rect 14686 -935 14720 -759
rect 14804 -935 14838 -759
rect 14922 -935 14956 -759
rect 15040 -935 15074 -759
rect 14745 -1029 14779 -995
rect 16303 -1063 16337 -687
rect 16421 -1063 16455 -687
rect 16539 -1063 16573 -687
rect 16657 -1063 16691 -687
rect 16775 -1063 16809 -687
rect 16893 -1063 16927 -687
rect 17011 -1063 17045 -687
rect 17445 -1059 17479 -683
rect 17563 -1059 17597 -683
rect 17681 -1059 17715 -683
rect 17799 -1059 17833 -683
rect 17917 -1059 17951 -683
rect 18035 -1059 18069 -683
rect 18153 -1059 18187 -683
rect 14627 -1146 14661 -1112
rect 14215 -1572 14249 -1196
rect 14333 -1572 14367 -1196
rect 14451 -1572 14485 -1196
rect 14568 -1372 14602 -1196
rect 14686 -1372 14720 -1196
rect 16508 -1419 16542 -1385
rect 17650 -1415 17684 -1381
rect 14274 -1656 14308 -1622
rect 14392 -1656 14426 -1622
rect 16213 -1646 16247 -1470
rect 16331 -1646 16365 -1470
rect 16449 -1646 16483 -1470
rect 16567 -1646 16601 -1470
rect 16732 -1646 16766 -1470
rect 16850 -1646 16884 -1470
rect 16968 -1646 17002 -1470
rect 17086 -1646 17120 -1470
rect 17355 -1642 17389 -1466
rect 17473 -1642 17507 -1466
rect 17591 -1642 17625 -1466
rect 17709 -1642 17743 -1466
rect 17874 -1642 17908 -1466
rect 17992 -1642 18026 -1466
rect 18110 -1642 18144 -1466
rect 18228 -1642 18262 -1466
rect 13992 -2585 14026 -2409
rect 14110 -2585 14144 -2409
rect 14228 -2585 14262 -2409
rect 14346 -2585 14380 -2409
rect 14464 -2585 14498 -2409
rect 14582 -2585 14616 -2409
rect 14700 -2585 14734 -2409
rect 14818 -2585 14852 -2409
rect 14936 -2585 14970 -2409
rect 15054 -2585 15088 -2409
rect 14759 -2679 14793 -2645
rect 14641 -2796 14675 -2762
rect 14229 -3222 14263 -2846
rect 14347 -3222 14381 -2846
rect 14465 -3222 14499 -2846
rect 14582 -3022 14616 -2846
rect 14700 -3022 14734 -2846
rect 15456 -3202 15490 -3026
rect 15574 -3202 15608 -3026
rect 15692 -3202 15726 -3026
rect 15810 -3202 15844 -3026
rect 15940 -3202 15974 -2826
rect 16058 -3202 16092 -2826
rect 16176 -3202 16210 -2826
rect 16294 -3202 16328 -2826
rect 16412 -3202 16446 -2826
rect 16530 -3202 16564 -2826
rect 16648 -3202 16682 -2826
rect 16777 -3202 16811 -3026
rect 16895 -3202 16929 -3026
rect 17013 -3202 17047 -3026
rect 17131 -3202 17165 -3026
rect 17354 -3202 17388 -3026
rect 17472 -3202 17506 -3026
rect 17590 -3202 17624 -3026
rect 17708 -3202 17742 -3026
rect 17838 -3202 17872 -2826
rect 17956 -3202 17990 -2826
rect 18074 -3202 18108 -2826
rect 18192 -3202 18226 -2826
rect 18310 -3202 18344 -2826
rect 18428 -3202 18462 -2826
rect 18546 -3202 18580 -2826
rect 18675 -3202 18709 -3026
rect 18793 -3202 18827 -3026
rect 18911 -3202 18945 -3026
rect 19029 -3202 19063 -3026
rect 14288 -3306 14322 -3272
rect 14406 -3306 14440 -3272
rect 16920 -3474 16954 -3440
rect 19027 -3495 19061 -3461
rect 15883 -3895 15917 -3519
rect 16001 -3895 16035 -3519
rect 13987 -4189 14021 -4013
rect 14105 -4189 14139 -4013
rect 14223 -4189 14257 -4013
rect 14341 -4189 14375 -4013
rect 14459 -4189 14493 -4013
rect 14577 -4189 14611 -4013
rect 14695 -4189 14729 -4013
rect 14813 -4189 14847 -4013
rect 14931 -4189 14965 -4013
rect 16119 -3895 16153 -3519
rect 16237 -3895 16271 -3519
rect 16355 -3895 16389 -3519
rect 16473 -3895 16507 -3519
rect 16591 -3895 16625 -3519
rect 17781 -3895 17815 -3519
rect 17899 -3895 17933 -3519
rect 18017 -3895 18051 -3519
rect 18135 -3895 18169 -3519
rect 18253 -3895 18287 -3519
rect 18371 -3895 18405 -3519
rect 18489 -3895 18523 -3519
rect 15049 -4189 15083 -4013
rect 15913 -4117 15947 -4083
rect 15728 -4184 15762 -4150
rect 16561 -4117 16595 -4083
rect 17811 -4117 17845 -4083
rect 16179 -4201 16213 -4167
rect 16297 -4200 16331 -4166
rect 16851 -4185 16885 -4151
rect 17626 -4184 17660 -4150
rect 19150 -4022 19282 -3924
rect 18457 -4116 18491 -4082
rect 18077 -4201 18111 -4167
rect 18195 -4200 18229 -4166
rect 18749 -4185 18783 -4151
rect 14754 -4283 14788 -4249
rect 14636 -4400 14670 -4366
rect 15581 -4427 15615 -4251
rect 14224 -4826 14258 -4450
rect 14342 -4826 14376 -4450
rect 14460 -4826 14494 -4450
rect 14577 -4626 14611 -4450
rect 15699 -4427 15733 -4251
rect 14695 -4626 14729 -4450
rect 16001 -4627 16035 -4251
rect 16119 -4627 16153 -4251
rect 16237 -4627 16271 -4251
rect 16355 -4627 16389 -4251
rect 16473 -4627 16507 -4251
rect 16879 -4427 16913 -4251
rect 16997 -4427 17031 -4251
rect 17479 -4427 17513 -4251
rect 17597 -4427 17631 -4251
rect 17899 -4627 17933 -4251
rect 18017 -4627 18051 -4251
rect 18135 -4627 18169 -4251
rect 18253 -4627 18287 -4251
rect 18371 -4627 18405 -4251
rect 18777 -4427 18811 -4251
rect 18895 -4427 18929 -4251
rect 14283 -4910 14317 -4876
rect 14401 -4910 14435 -4876
<< metal1 >>
rect 14375 -461 14595 -441
rect 14375 -569 14419 -461
rect 14551 -569 14595 -461
rect 16172 -503 16228 -495
rect 14375 -611 14595 -569
rect 15246 -511 16228 -503
rect 15246 -545 16188 -511
rect 16222 -545 16228 -511
rect 16891 -515 16901 -407
rect 17033 -470 17043 -407
rect 17033 -481 17045 -470
rect 17033 -515 17046 -481
rect 17302 -491 17358 -489
rect 15246 -561 16228 -545
rect 16901 -553 17046 -515
rect 15246 -562 16225 -561
rect 13979 -641 14956 -611
rect 13979 -747 14011 -641
rect 14215 -747 14247 -641
rect 14451 -747 14483 -641
rect 14687 -747 14719 -641
rect 14922 -747 14956 -641
rect 13972 -759 14018 -747
rect 13972 -935 13978 -759
rect 14012 -935 14018 -759
rect 13972 -947 14018 -935
rect 14090 -759 14136 -747
rect 14090 -935 14096 -759
rect 14130 -935 14136 -759
rect 14090 -947 14136 -935
rect 14208 -759 14254 -747
rect 14208 -935 14214 -759
rect 14248 -935 14254 -759
rect 14208 -947 14254 -935
rect 14326 -759 14372 -747
rect 14326 -935 14332 -759
rect 14366 -935 14372 -759
rect 14326 -947 14372 -935
rect 14444 -759 14490 -747
rect 14444 -935 14450 -759
rect 14484 -935 14490 -759
rect 14444 -947 14490 -935
rect 14562 -759 14608 -747
rect 14562 -935 14568 -759
rect 14602 -935 14608 -759
rect 14562 -947 14608 -935
rect 14680 -759 14726 -747
rect 14680 -935 14686 -759
rect 14720 -935 14726 -759
rect 14680 -947 14726 -935
rect 14798 -759 14844 -747
rect 14798 -935 14804 -759
rect 14838 -935 14844 -759
rect 14798 -947 14844 -935
rect 14916 -759 14962 -747
rect 14916 -935 14922 -759
rect 14956 -935 14962 -759
rect 14916 -947 14962 -935
rect 15034 -759 15080 -747
rect 15034 -935 15040 -759
rect 15074 -935 15080 -759
rect 15034 -947 15080 -935
rect 14095 -1041 14131 -947
rect 14331 -1041 14367 -947
rect 14567 -1040 14603 -947
rect 14729 -995 14795 -988
rect 14729 -1029 14745 -995
rect 14779 -1029 14795 -995
rect 14729 -1040 14795 -1029
rect 14567 -1041 14795 -1040
rect 14095 -1070 14795 -1041
rect 14095 -1071 14677 -1070
rect 14215 -1184 14249 -1071
rect 14611 -1112 14677 -1071
rect 14611 -1146 14627 -1112
rect 14661 -1146 14677 -1112
rect 14611 -1153 14677 -1146
rect 15039 -1152 15074 -947
rect 15246 -1152 15313 -562
rect 17005 -585 17046 -553
rect 17292 -557 17302 -491
rect 17358 -557 17368 -491
rect 18038 -515 18048 -407
rect 18180 -470 18190 -407
rect 18180 -481 18192 -470
rect 18180 -515 18193 -481
rect 18048 -553 18193 -515
rect 18152 -581 18193 -553
rect 16421 -613 16691 -585
rect 16162 -679 16172 -613
rect 16238 -679 16248 -613
rect 16421 -675 16455 -613
rect 16657 -675 16691 -613
rect 16775 -613 17046 -585
rect 17563 -609 17833 -581
rect 16775 -675 16809 -613
rect 17011 -675 17046 -613
rect 17187 -625 17358 -609
rect 17187 -659 17318 -625
rect 17352 -659 17358 -625
rect 17187 -675 17358 -659
rect 17563 -671 17597 -609
rect 17799 -671 17833 -609
rect 17917 -609 18193 -581
rect 17917 -671 17951 -609
rect 18153 -671 18193 -609
rect 16297 -687 16343 -675
rect 16297 -1063 16303 -687
rect 16337 -1063 16343 -687
rect 16297 -1075 16343 -1063
rect 16415 -687 16461 -675
rect 16415 -1063 16421 -687
rect 16455 -1063 16461 -687
rect 16415 -1075 16461 -1063
rect 16533 -687 16579 -675
rect 16533 -1063 16539 -687
rect 16573 -1063 16579 -687
rect 16533 -1075 16579 -1063
rect 16651 -687 16697 -675
rect 16651 -1063 16657 -687
rect 16691 -1063 16697 -687
rect 16651 -1075 16697 -1063
rect 16769 -687 16815 -675
rect 16769 -1063 16775 -687
rect 16809 -1063 16815 -687
rect 16769 -1075 16815 -1063
rect 16887 -687 16933 -675
rect 16887 -1063 16893 -687
rect 16927 -1063 16933 -687
rect 16887 -1075 16933 -1063
rect 17005 -687 17051 -675
rect 17005 -1063 17011 -687
rect 17045 -1063 17051 -687
rect 17005 -1075 17051 -1063
rect 15039 -1180 15313 -1152
rect 14685 -1184 15313 -1180
rect 14209 -1196 14255 -1184
rect 13037 -1589 13326 -1414
rect 14209 -1572 14215 -1196
rect 14249 -1572 14255 -1196
rect 14209 -1584 14255 -1572
rect 14327 -1196 14373 -1184
rect 14327 -1572 14333 -1196
rect 14367 -1572 14373 -1196
rect 14327 -1584 14373 -1572
rect 14445 -1196 14491 -1184
rect 14445 -1572 14451 -1196
rect 14485 -1548 14491 -1196
rect 14562 -1196 14608 -1184
rect 14562 -1372 14568 -1196
rect 14602 -1372 14608 -1196
rect 14562 -1384 14608 -1372
rect 14680 -1196 15313 -1184
rect 14680 -1372 14686 -1196
rect 14720 -1209 15313 -1196
rect 16303 -1117 16337 -1075
rect 16539 -1117 16573 -1075
rect 16303 -1145 16573 -1117
rect 16657 -1116 16691 -1075
rect 16893 -1116 16927 -1075
rect 16657 -1145 16927 -1116
rect 16303 -1193 16337 -1145
rect 14720 -1372 14726 -1209
rect 16303 -1223 16366 -1193
rect 14680 -1384 14726 -1372
rect 16331 -1315 16366 -1223
rect 16331 -1351 16558 -1315
rect 16828 -1326 16838 -1229
rect 16937 -1326 16947 -1229
rect 17011 -1258 17045 -1075
rect 17011 -1312 17120 -1258
rect 14568 -1500 14603 -1384
rect 16331 -1458 16366 -1351
rect 16492 -1385 16558 -1351
rect 16492 -1419 16508 -1385
rect 16542 -1419 16558 -1385
rect 16839 -1327 16936 -1326
rect 16839 -1394 16896 -1327
rect 16492 -1425 16558 -1419
rect 16733 -1430 17002 -1394
rect 16733 -1458 16766 -1430
rect 16969 -1458 17002 -1430
rect 17086 -1458 17120 -1312
rect 16207 -1470 16253 -1458
rect 14699 -1500 14807 -1490
rect 14568 -1548 14699 -1500
rect 14485 -1572 14699 -1548
rect 14445 -1584 14699 -1572
rect 14451 -1588 14699 -1584
rect 13037 -1616 14087 -1589
rect 13037 -1622 14324 -1616
rect 13037 -1656 14274 -1622
rect 14308 -1656 14324 -1622
rect 13037 -1672 14324 -1656
rect 14376 -1622 14442 -1616
rect 14376 -1656 14392 -1622
rect 14426 -1656 14442 -1622
rect 14625 -1632 14699 -1588
rect 14699 -1642 14807 -1632
rect 13037 -1688 14087 -1672
rect 13037 -1689 14024 -1688
rect 13037 -1693 13559 -1689
rect 13037 -1694 13326 -1693
rect 13054 -2104 13343 -1942
rect 13054 -2210 13191 -2104
rect 13303 -2117 13343 -2104
rect 13303 -2210 13345 -2117
rect 13054 -2221 13345 -2210
rect 13054 -2222 13343 -2221
rect 13054 -3216 13342 -3054
rect 13054 -3322 13190 -3216
rect 13302 -3218 13342 -3216
rect 13308 -3229 13342 -3218
rect 13054 -3324 13196 -3322
rect 13308 -3324 13343 -3229
rect 13054 -3333 13343 -3324
rect 13054 -3334 13342 -3333
rect 13054 -3335 13310 -3334
rect 13466 -3587 13559 -1693
rect 13622 -1752 14088 -1730
rect 14376 -1752 14442 -1656
rect 16207 -1646 16213 -1470
rect 16247 -1646 16253 -1470
rect 16207 -1658 16253 -1646
rect 16325 -1470 16371 -1458
rect 16325 -1646 16331 -1470
rect 16365 -1646 16371 -1470
rect 16325 -1658 16371 -1646
rect 16443 -1470 16489 -1458
rect 16443 -1646 16449 -1470
rect 16483 -1646 16489 -1470
rect 16443 -1658 16489 -1646
rect 16561 -1470 16607 -1458
rect 16561 -1646 16567 -1470
rect 16601 -1525 16607 -1470
rect 16726 -1470 16772 -1458
rect 16726 -1525 16732 -1470
rect 16601 -1613 16732 -1525
rect 16601 -1646 16607 -1613
rect 16561 -1658 16607 -1646
rect 16726 -1646 16732 -1613
rect 16766 -1646 16772 -1470
rect 16726 -1658 16772 -1646
rect 16844 -1470 16890 -1458
rect 16844 -1646 16850 -1470
rect 16884 -1646 16890 -1470
rect 16844 -1658 16890 -1646
rect 16962 -1470 17008 -1458
rect 16962 -1646 16968 -1470
rect 17002 -1646 17008 -1470
rect 16962 -1658 17008 -1646
rect 17080 -1470 17126 -1458
rect 17080 -1646 17086 -1470
rect 17120 -1646 17126 -1470
rect 17080 -1658 17126 -1646
rect 16213 -1697 16247 -1658
rect 16449 -1697 16483 -1658
rect 16213 -1732 16483 -1697
rect 16850 -1696 16883 -1658
rect 17086 -1696 17119 -1658
rect 16850 -1732 17119 -1696
rect 13622 -1800 14442 -1752
rect 16247 -1733 16483 -1732
rect 13622 -1831 14088 -1800
rect 16247 -1807 16379 -1733
rect 13622 -2087 13727 -1831
rect 16237 -1915 16247 -1807
rect 16379 -1915 16389 -1807
rect 13622 -2193 13685 -2087
rect 13797 -2193 13807 -2087
rect 14389 -2111 14609 -2091
rect 13622 -2204 13771 -2193
rect 13622 -3381 13727 -2204
rect 14389 -2219 14433 -2111
rect 14565 -2219 14609 -2111
rect 14389 -2261 14609 -2219
rect 17187 -2246 17249 -675
rect 17439 -683 17485 -671
rect 17439 -1059 17445 -683
rect 17479 -1059 17485 -683
rect 17439 -1071 17485 -1059
rect 17557 -683 17603 -671
rect 17557 -1059 17563 -683
rect 17597 -1059 17603 -683
rect 17557 -1071 17603 -1059
rect 17675 -683 17721 -671
rect 17675 -1059 17681 -683
rect 17715 -1059 17721 -683
rect 17675 -1071 17721 -1059
rect 17793 -683 17839 -671
rect 17793 -1059 17799 -683
rect 17833 -1059 17839 -683
rect 17793 -1071 17839 -1059
rect 17911 -683 17957 -671
rect 17911 -1059 17917 -683
rect 17951 -1059 17957 -683
rect 17911 -1071 17957 -1059
rect 18029 -683 18075 -671
rect 18029 -1059 18035 -683
rect 18069 -1059 18075 -683
rect 18029 -1071 18075 -1059
rect 18147 -683 18193 -671
rect 18147 -1059 18153 -683
rect 18187 -1059 18193 -683
rect 18147 -1071 18193 -1059
rect 17445 -1113 17479 -1071
rect 17681 -1113 17715 -1071
rect 17445 -1141 17715 -1113
rect 17799 -1112 17833 -1071
rect 18035 -1112 18069 -1071
rect 17799 -1141 18069 -1112
rect 17445 -1189 17479 -1141
rect 17445 -1219 17508 -1189
rect 17473 -1311 17508 -1219
rect 17980 -1249 18080 -1228
rect 17980 -1303 17994 -1249
rect 18059 -1303 18080 -1249
rect 17980 -1308 18080 -1303
rect 18153 -1254 18187 -1071
rect 18153 -1308 18262 -1254
rect 17473 -1347 17700 -1311
rect 17473 -1454 17508 -1347
rect 17634 -1381 17700 -1347
rect 17634 -1415 17650 -1381
rect 17684 -1415 17700 -1381
rect 17981 -1323 18078 -1308
rect 17981 -1390 18038 -1323
rect 17634 -1421 17700 -1415
rect 17875 -1426 18144 -1390
rect 17875 -1454 17908 -1426
rect 18111 -1454 18144 -1426
rect 18228 -1454 18262 -1308
rect 19079 -1315 19089 -1240
rect 19157 -1315 19257 -1240
rect 19106 -1316 19257 -1315
rect 17349 -1466 17395 -1454
rect 17349 -1642 17355 -1466
rect 17389 -1642 17395 -1466
rect 17349 -1654 17395 -1642
rect 17467 -1466 17513 -1454
rect 17467 -1642 17473 -1466
rect 17507 -1642 17513 -1466
rect 17467 -1654 17513 -1642
rect 17585 -1466 17631 -1454
rect 17585 -1642 17591 -1466
rect 17625 -1642 17631 -1466
rect 17585 -1654 17631 -1642
rect 17703 -1466 17749 -1454
rect 17703 -1642 17709 -1466
rect 17743 -1521 17749 -1466
rect 17868 -1466 17914 -1454
rect 17868 -1521 17874 -1466
rect 17743 -1609 17874 -1521
rect 17743 -1642 17749 -1609
rect 17703 -1654 17749 -1642
rect 17868 -1642 17874 -1609
rect 17908 -1642 17914 -1466
rect 17868 -1654 17914 -1642
rect 17986 -1466 18032 -1454
rect 17986 -1642 17992 -1466
rect 18026 -1642 18032 -1466
rect 17986 -1654 18032 -1642
rect 18104 -1466 18150 -1454
rect 18104 -1642 18110 -1466
rect 18144 -1642 18150 -1466
rect 18104 -1654 18150 -1642
rect 18222 -1466 18268 -1454
rect 18222 -1642 18228 -1466
rect 18262 -1642 18268 -1466
rect 18222 -1654 18268 -1642
rect 17355 -1693 17389 -1654
rect 17591 -1693 17625 -1654
rect 17355 -1729 17625 -1693
rect 17992 -1692 18025 -1654
rect 18228 -1692 18261 -1654
rect 17992 -1728 18261 -1692
rect 17355 -1730 17521 -1729
rect 17389 -1809 17521 -1730
rect 17379 -1917 17389 -1809
rect 17521 -1917 17531 -1809
rect 13993 -2291 14970 -2261
rect 17187 -2263 17250 -2246
rect 17112 -2267 17250 -2263
rect 13993 -2397 14025 -2291
rect 14229 -2397 14261 -2291
rect 14465 -2397 14497 -2291
rect 14701 -2397 14733 -2291
rect 14936 -2397 14970 -2291
rect 15280 -2301 17250 -2267
rect 15278 -2330 17250 -2301
rect 15278 -2346 15324 -2330
rect 17112 -2332 17250 -2330
rect 13986 -2409 14032 -2397
rect 13986 -2585 13992 -2409
rect 14026 -2585 14032 -2409
rect 13986 -2597 14032 -2585
rect 14104 -2409 14150 -2397
rect 14104 -2585 14110 -2409
rect 14144 -2585 14150 -2409
rect 14104 -2597 14150 -2585
rect 14222 -2409 14268 -2397
rect 14222 -2585 14228 -2409
rect 14262 -2585 14268 -2409
rect 14222 -2597 14268 -2585
rect 14340 -2409 14386 -2397
rect 14340 -2585 14346 -2409
rect 14380 -2585 14386 -2409
rect 14340 -2597 14386 -2585
rect 14458 -2409 14504 -2397
rect 14458 -2585 14464 -2409
rect 14498 -2585 14504 -2409
rect 14458 -2597 14504 -2585
rect 14576 -2409 14622 -2397
rect 14576 -2585 14582 -2409
rect 14616 -2585 14622 -2409
rect 14576 -2597 14622 -2585
rect 14694 -2409 14740 -2397
rect 14694 -2585 14700 -2409
rect 14734 -2585 14740 -2409
rect 14694 -2597 14740 -2585
rect 14812 -2409 14858 -2397
rect 14812 -2585 14818 -2409
rect 14852 -2585 14858 -2409
rect 14812 -2597 14858 -2585
rect 14930 -2409 14976 -2397
rect 14930 -2585 14936 -2409
rect 14970 -2585 14976 -2409
rect 14930 -2597 14976 -2585
rect 15048 -2409 15094 -2397
rect 15048 -2585 15054 -2409
rect 15088 -2585 15094 -2409
rect 15048 -2597 15094 -2585
rect 14109 -2691 14145 -2597
rect 14345 -2691 14381 -2597
rect 14581 -2690 14617 -2597
rect 14743 -2645 14809 -2638
rect 14743 -2679 14759 -2645
rect 14793 -2679 14809 -2645
rect 14743 -2690 14809 -2679
rect 14581 -2691 14809 -2690
rect 14109 -2720 14809 -2691
rect 14109 -2721 14691 -2720
rect 14229 -2834 14263 -2721
rect 14625 -2762 14691 -2721
rect 14625 -2796 14641 -2762
rect 14675 -2796 14691 -2762
rect 14625 -2803 14691 -2796
rect 15053 -2815 15088 -2597
rect 15277 -2798 15324 -2346
rect 16236 -2562 16246 -2454
rect 16378 -2562 16388 -2454
rect 18134 -2562 18144 -2454
rect 18276 -2562 18286 -2454
rect 16246 -2602 16378 -2562
rect 18144 -2602 18276 -2562
rect 16245 -2668 16378 -2602
rect 18143 -2668 18276 -2602
rect 15574 -2711 17047 -2668
rect 15277 -2814 15323 -2798
rect 15242 -2815 15323 -2814
rect 15053 -2830 15323 -2815
rect 14699 -2834 15323 -2830
rect 14223 -2846 14269 -2834
rect 13958 -3324 13968 -3206
rect 14086 -3238 14096 -3206
rect 14223 -3222 14229 -2846
rect 14263 -3222 14269 -2846
rect 14223 -3234 14269 -3222
rect 14341 -2846 14387 -2834
rect 14341 -3222 14347 -2846
rect 14381 -3222 14387 -2846
rect 14341 -3234 14387 -3222
rect 14459 -2846 14505 -2834
rect 14459 -3222 14465 -2846
rect 14499 -3198 14505 -2846
rect 14576 -2846 14622 -2834
rect 14576 -3022 14582 -2846
rect 14616 -3022 14622 -2846
rect 14576 -3034 14622 -3022
rect 14694 -2846 15323 -2834
rect 14694 -3022 14700 -2846
rect 14734 -2858 15323 -2846
rect 14734 -2859 14976 -2858
rect 14734 -3022 14740 -2859
rect 15242 -2860 15323 -2858
rect 15574 -3014 15608 -2711
rect 15940 -2814 15974 -2711
rect 16176 -2814 16210 -2711
rect 16412 -2814 16446 -2711
rect 16648 -2814 16682 -2711
rect 15934 -2826 15980 -2814
rect 14694 -3034 14740 -3022
rect 15450 -3026 15496 -3014
rect 14582 -3150 14617 -3034
rect 14713 -3150 14821 -3140
rect 14582 -3198 14713 -3150
rect 14499 -3222 14713 -3198
rect 14459 -3234 14713 -3222
rect 14465 -3238 14713 -3234
rect 14086 -3266 14101 -3238
rect 14086 -3272 14338 -3266
rect 14086 -3306 14288 -3272
rect 14322 -3306 14338 -3272
rect 14086 -3322 14338 -3306
rect 14390 -3272 14456 -3266
rect 14390 -3306 14406 -3272
rect 14440 -3306 14456 -3272
rect 14639 -3282 14713 -3238
rect 15450 -3202 15456 -3026
rect 15490 -3202 15496 -3026
rect 15450 -3214 15496 -3202
rect 15568 -3026 15614 -3014
rect 15568 -3202 15574 -3026
rect 15608 -3202 15614 -3026
rect 15568 -3214 15614 -3202
rect 15686 -3026 15732 -3014
rect 15686 -3202 15692 -3026
rect 15726 -3202 15732 -3026
rect 15686 -3214 15732 -3202
rect 15804 -3026 15850 -3014
rect 15934 -3026 15940 -2826
rect 15804 -3202 15810 -3026
rect 15844 -3202 15940 -3026
rect 15974 -3202 15980 -2826
rect 15804 -3214 15850 -3202
rect 15934 -3214 15980 -3202
rect 16052 -2826 16098 -2814
rect 16052 -3202 16058 -2826
rect 16092 -3202 16098 -2826
rect 16052 -3214 16098 -3202
rect 16170 -2826 16216 -2814
rect 16170 -3202 16176 -2826
rect 16210 -3202 16216 -2826
rect 16170 -3214 16216 -3202
rect 16288 -2826 16334 -2814
rect 16288 -3202 16294 -2826
rect 16328 -3202 16334 -2826
rect 16288 -3214 16334 -3202
rect 16406 -2826 16452 -2814
rect 16406 -3202 16412 -2826
rect 16446 -3202 16452 -2826
rect 16406 -3214 16452 -3202
rect 16524 -2826 16570 -2814
rect 16524 -3202 16530 -2826
rect 16564 -3202 16570 -2826
rect 16524 -3214 16570 -3202
rect 16642 -2826 16688 -2814
rect 16642 -3202 16648 -2826
rect 16682 -3026 16688 -2826
rect 17013 -3014 17047 -2711
rect 17472 -2711 18945 -2668
rect 17472 -3014 17506 -2711
rect 17838 -2814 17872 -2711
rect 18074 -2814 18108 -2711
rect 18310 -2814 18344 -2711
rect 18546 -2814 18580 -2711
rect 17832 -2826 17878 -2814
rect 16771 -3026 16817 -3014
rect 16682 -3202 16777 -3026
rect 16811 -3202 16817 -3026
rect 16642 -3214 16688 -3202
rect 16771 -3214 16817 -3202
rect 16889 -3026 16935 -3014
rect 16889 -3202 16895 -3026
rect 16929 -3202 16935 -3026
rect 16889 -3214 16935 -3202
rect 17007 -3026 17053 -3014
rect 17007 -3202 17013 -3026
rect 17047 -3202 17053 -3026
rect 17007 -3214 17053 -3202
rect 17125 -3026 17171 -3014
rect 17125 -3202 17131 -3026
rect 17165 -3202 17171 -3026
rect 17125 -3214 17171 -3202
rect 17348 -3026 17394 -3014
rect 17348 -3202 17354 -3026
rect 17388 -3202 17394 -3026
rect 17348 -3214 17394 -3202
rect 17466 -3026 17512 -3014
rect 17466 -3202 17472 -3026
rect 17506 -3202 17512 -3026
rect 17466 -3214 17512 -3202
rect 17584 -3026 17630 -3014
rect 17584 -3202 17590 -3026
rect 17624 -3202 17630 -3026
rect 17584 -3214 17630 -3202
rect 17702 -3026 17748 -3014
rect 17832 -3026 17838 -2826
rect 17702 -3202 17708 -3026
rect 17742 -3202 17838 -3026
rect 17872 -3202 17878 -2826
rect 17702 -3214 17748 -3202
rect 17832 -3214 17878 -3202
rect 17950 -2826 17996 -2814
rect 17950 -3202 17956 -2826
rect 17990 -3202 17996 -2826
rect 17950 -3214 17996 -3202
rect 18068 -2826 18114 -2814
rect 18068 -3202 18074 -2826
rect 18108 -3202 18114 -2826
rect 18068 -3214 18114 -3202
rect 18186 -2826 18232 -2814
rect 18186 -3202 18192 -2826
rect 18226 -3202 18232 -2826
rect 18186 -3214 18232 -3202
rect 18304 -2826 18350 -2814
rect 18304 -3202 18310 -2826
rect 18344 -3202 18350 -2826
rect 18304 -3214 18350 -3202
rect 18422 -2826 18468 -2814
rect 18422 -3202 18428 -2826
rect 18462 -3202 18468 -2826
rect 18422 -3214 18468 -3202
rect 18540 -2826 18586 -2814
rect 18540 -3202 18546 -2826
rect 18580 -3026 18586 -2826
rect 18911 -3014 18945 -2711
rect 18669 -3026 18715 -3014
rect 18580 -3202 18675 -3026
rect 18709 -3202 18715 -3026
rect 18540 -3214 18586 -3202
rect 18669 -3214 18715 -3202
rect 18787 -3026 18833 -3014
rect 18787 -3202 18793 -3026
rect 18827 -3202 18833 -3026
rect 18787 -3214 18833 -3202
rect 18905 -3026 18951 -3014
rect 18905 -3202 18911 -3026
rect 18945 -3202 18951 -3026
rect 18905 -3214 18951 -3202
rect 19023 -3026 19069 -3014
rect 19023 -3202 19029 -3026
rect 19063 -3202 19069 -3026
rect 19023 -3214 19069 -3202
rect 14713 -3292 14821 -3282
rect 15456 -3248 15490 -3214
rect 16058 -3248 16092 -3214
rect 16294 -3248 16328 -3214
rect 15456 -3283 15615 -3248
rect 16058 -3283 16328 -3248
rect 16895 -3248 16929 -3214
rect 17131 -3248 17165 -3214
rect 16895 -3283 17165 -3248
rect 17354 -3248 17388 -3214
rect 17956 -3248 17990 -3214
rect 18192 -3248 18226 -3214
rect 17354 -3283 17513 -3248
rect 17956 -3283 18226 -3248
rect 18793 -3248 18827 -3214
rect 19029 -3248 19063 -3214
rect 18793 -3283 19063 -3248
rect 14086 -3324 14101 -3322
rect 14001 -3338 14101 -3324
rect 14001 -3381 14101 -3380
rect 13622 -3402 14101 -3381
rect 14390 -3402 14456 -3306
rect 13622 -3450 14456 -3402
rect 13622 -3479 14101 -3450
rect 13622 -3481 13727 -3479
rect 14001 -3480 14101 -3479
rect 13455 -3666 13465 -3587
rect 13558 -3666 13568 -3587
rect 13466 -4840 13559 -3666
rect 14384 -3715 14604 -3695
rect 14384 -3823 14428 -3715
rect 14560 -3823 14604 -3715
rect 14384 -3865 14604 -3823
rect 13988 -3895 14965 -3865
rect 13988 -4001 14020 -3895
rect 14224 -4001 14256 -3895
rect 14460 -4001 14492 -3895
rect 14696 -4001 14728 -3895
rect 14931 -4001 14965 -3895
rect 13981 -4013 14027 -4001
rect 13981 -4189 13987 -4013
rect 14021 -4189 14027 -4013
rect 13981 -4201 14027 -4189
rect 14099 -4013 14145 -4001
rect 14099 -4189 14105 -4013
rect 14139 -4189 14145 -4013
rect 14099 -4201 14145 -4189
rect 14217 -4013 14263 -4001
rect 14217 -4189 14223 -4013
rect 14257 -4189 14263 -4013
rect 14217 -4201 14263 -4189
rect 14335 -4013 14381 -4001
rect 14335 -4189 14341 -4013
rect 14375 -4189 14381 -4013
rect 14335 -4201 14381 -4189
rect 14453 -4013 14499 -4001
rect 14453 -4189 14459 -4013
rect 14493 -4189 14499 -4013
rect 14453 -4201 14499 -4189
rect 14571 -4013 14617 -4001
rect 14571 -4189 14577 -4013
rect 14611 -4189 14617 -4013
rect 14571 -4201 14617 -4189
rect 14689 -4013 14735 -4001
rect 14689 -4189 14695 -4013
rect 14729 -4189 14735 -4013
rect 14689 -4201 14735 -4189
rect 14807 -4013 14853 -4001
rect 14807 -4189 14813 -4013
rect 14847 -4189 14853 -4013
rect 14807 -4201 14853 -4189
rect 14925 -4013 14971 -4001
rect 14925 -4189 14931 -4013
rect 14965 -4189 14971 -4013
rect 14925 -4201 14971 -4189
rect 15043 -4013 15089 -4001
rect 15043 -4189 15049 -4013
rect 15083 -4189 15089 -4013
rect 15043 -4201 15089 -4189
rect 15581 -4067 15615 -3283
rect 16294 -3345 16328 -3283
rect 15883 -3383 16625 -3345
rect 15883 -3507 15917 -3383
rect 16119 -3507 16153 -3383
rect 16355 -3507 16389 -3383
rect 16591 -3507 16625 -3383
rect 16881 -3490 16891 -3424
rect 16954 -3490 16964 -3424
rect 15877 -3519 15923 -3507
rect 15877 -3895 15883 -3519
rect 15917 -3895 15923 -3519
rect 15877 -3907 15923 -3895
rect 15995 -3519 16041 -3507
rect 15995 -3895 16001 -3519
rect 16035 -3895 16041 -3519
rect 15995 -3907 16041 -3895
rect 16113 -3519 16159 -3507
rect 16113 -3895 16119 -3519
rect 16153 -3895 16159 -3519
rect 16113 -3907 16159 -3895
rect 16231 -3519 16277 -3507
rect 16231 -3895 16237 -3519
rect 16271 -3895 16277 -3519
rect 16231 -3907 16277 -3895
rect 16349 -3519 16395 -3507
rect 16349 -3895 16355 -3519
rect 16389 -3895 16395 -3519
rect 16349 -3907 16395 -3895
rect 16467 -3519 16513 -3507
rect 16467 -3895 16473 -3519
rect 16507 -3895 16513 -3519
rect 16467 -3907 16513 -3895
rect 16585 -3519 16631 -3507
rect 16585 -3895 16591 -3519
rect 16625 -3895 16631 -3519
rect 16585 -3907 16631 -3895
rect 16997 -4066 17031 -3283
rect 16724 -4067 17031 -4066
rect 15581 -4072 15897 -4067
rect 16611 -4072 17031 -4067
rect 15581 -4083 15964 -4072
rect 15581 -4110 15913 -4083
rect 14104 -4295 14140 -4201
rect 14340 -4295 14376 -4201
rect 14576 -4294 14612 -4201
rect 14738 -4249 14804 -4242
rect 14738 -4283 14754 -4249
rect 14788 -4283 14804 -4249
rect 14738 -4294 14804 -4283
rect 14576 -4295 14804 -4294
rect 14104 -4324 14804 -4295
rect 14104 -4325 14686 -4324
rect 14224 -4438 14258 -4325
rect 14620 -4366 14686 -4325
rect 14620 -4400 14636 -4366
rect 14670 -4400 14686 -4366
rect 14620 -4407 14686 -4400
rect 15048 -4434 15083 -4201
rect 15581 -4239 15615 -4110
rect 15897 -4117 15913 -4110
rect 15947 -4117 15964 -4083
rect 15897 -4123 15964 -4117
rect 16544 -4083 17031 -4072
rect 16544 -4117 16561 -4083
rect 16595 -4110 17031 -4083
rect 16595 -4117 16611 -4110
rect 16724 -4111 17031 -4110
rect 16544 -4123 16611 -4117
rect 15722 -4150 15778 -4138
rect 15722 -4184 15728 -4150
rect 15762 -4151 15778 -4150
rect 16835 -4151 16891 -4139
rect 15762 -4167 16229 -4151
rect 15762 -4184 16179 -4167
rect 15722 -4200 16179 -4184
rect 16163 -4201 16179 -4200
rect 16213 -4201 16229 -4167
rect 16163 -4208 16229 -4201
rect 16281 -4166 16851 -4151
rect 16281 -4200 16297 -4166
rect 16331 -4185 16851 -4166
rect 16885 -4185 16891 -4151
rect 16331 -4200 16891 -4185
rect 16281 -4210 16348 -4200
rect 16835 -4201 16891 -4200
rect 16997 -4239 17031 -4111
rect 17479 -4067 17513 -3283
rect 18192 -3345 18226 -3283
rect 17781 -3383 18523 -3345
rect 17781 -3507 17815 -3383
rect 18017 -3507 18051 -3383
rect 18253 -3507 18287 -3383
rect 18489 -3507 18523 -3383
rect 17775 -3519 17821 -3507
rect 17775 -3895 17781 -3519
rect 17815 -3895 17821 -3519
rect 17775 -3907 17821 -3895
rect 17893 -3519 17939 -3507
rect 17893 -3895 17899 -3519
rect 17933 -3895 17939 -3519
rect 17893 -3907 17939 -3895
rect 18011 -3519 18057 -3507
rect 18011 -3895 18017 -3519
rect 18051 -3895 18057 -3519
rect 18011 -3907 18057 -3895
rect 18129 -3519 18175 -3507
rect 18129 -3895 18135 -3519
rect 18169 -3895 18175 -3519
rect 18129 -3907 18175 -3895
rect 18247 -3519 18293 -3507
rect 18247 -3895 18253 -3519
rect 18287 -3895 18293 -3519
rect 18247 -3907 18293 -3895
rect 18365 -3519 18411 -3507
rect 18365 -3895 18371 -3519
rect 18405 -3895 18411 -3519
rect 18365 -3907 18411 -3895
rect 18483 -3519 18529 -3507
rect 18483 -3895 18489 -3519
rect 18523 -3895 18529 -3519
rect 18483 -3907 18529 -3895
rect 18895 -4066 18929 -3283
rect 18507 -4067 18576 -4066
rect 18622 -4067 18929 -4066
rect 17479 -4072 17795 -4067
rect 18507 -4071 18929 -4067
rect 17479 -4083 17862 -4072
rect 17479 -4110 17811 -4083
rect 17479 -4239 17513 -4110
rect 17795 -4117 17811 -4110
rect 17845 -4117 17862 -4083
rect 17795 -4123 17862 -4117
rect 18440 -4082 18929 -4071
rect 18440 -4116 18457 -4082
rect 18491 -4110 18929 -4082
rect 18491 -4116 18507 -4110
rect 18622 -4111 18929 -4110
rect 18440 -4122 18507 -4116
rect 17620 -4150 17676 -4138
rect 17620 -4184 17626 -4150
rect 17660 -4151 17676 -4150
rect 18733 -4151 18789 -4139
rect 17660 -4167 18127 -4151
rect 17660 -4184 18077 -4167
rect 17620 -4200 18077 -4184
rect 18061 -4201 18077 -4200
rect 18111 -4201 18127 -4167
rect 18061 -4208 18127 -4201
rect 18179 -4166 18749 -4151
rect 18179 -4200 18195 -4166
rect 18229 -4185 18749 -4166
rect 18783 -4185 18789 -4151
rect 18229 -4200 18789 -4185
rect 18179 -4210 18246 -4200
rect 18733 -4201 18789 -4200
rect 18895 -4239 18929 -4111
rect 19010 -3461 19077 -3437
rect 19010 -3495 19027 -3461
rect 19061 -3495 19077 -3461
rect 14694 -4438 15083 -4434
rect 14218 -4450 14264 -4438
rect 14218 -4826 14224 -4450
rect 14258 -4826 14264 -4450
rect 14218 -4838 14264 -4826
rect 14336 -4450 14382 -4438
rect 14336 -4826 14342 -4450
rect 14376 -4826 14382 -4450
rect 14336 -4838 14382 -4826
rect 14454 -4450 14500 -4438
rect 14454 -4826 14460 -4450
rect 14494 -4802 14500 -4450
rect 14571 -4450 14617 -4438
rect 14571 -4626 14577 -4450
rect 14611 -4626 14617 -4450
rect 14571 -4638 14617 -4626
rect 14689 -4450 15083 -4438
rect 15575 -4251 15621 -4239
rect 15575 -4427 15581 -4251
rect 15615 -4427 15621 -4251
rect 15575 -4439 15621 -4427
rect 15693 -4251 15739 -4239
rect 15693 -4427 15699 -4251
rect 15733 -4427 15739 -4251
rect 15693 -4439 15739 -4427
rect 15995 -4251 16041 -4239
rect 14689 -4626 14695 -4450
rect 14729 -4463 15083 -4450
rect 14729 -4626 14735 -4463
rect 15005 -4466 15083 -4463
rect 15005 -4518 15015 -4466
rect 15078 -4518 15088 -4466
rect 15010 -4524 15083 -4518
rect 14689 -4638 14735 -4626
rect 14577 -4754 14612 -4638
rect 15698 -4733 15732 -4439
rect 15995 -4627 16001 -4251
rect 16035 -4627 16041 -4251
rect 15995 -4639 16041 -4627
rect 16113 -4251 16159 -4239
rect 16113 -4627 16119 -4251
rect 16153 -4627 16159 -4251
rect 16113 -4639 16159 -4627
rect 16231 -4251 16277 -4239
rect 16231 -4627 16237 -4251
rect 16271 -4627 16277 -4251
rect 16231 -4639 16277 -4627
rect 16349 -4251 16395 -4239
rect 16349 -4627 16355 -4251
rect 16389 -4627 16395 -4251
rect 16349 -4639 16395 -4627
rect 16467 -4251 16513 -4239
rect 16467 -4627 16473 -4251
rect 16507 -4627 16513 -4251
rect 16873 -4251 16919 -4239
rect 16873 -4427 16879 -4251
rect 16913 -4427 16919 -4251
rect 16873 -4439 16919 -4427
rect 16991 -4251 17037 -4239
rect 16991 -4427 16997 -4251
rect 17031 -4427 17037 -4251
rect 16991 -4439 17037 -4427
rect 17473 -4251 17519 -4239
rect 17473 -4427 17479 -4251
rect 17513 -4427 17519 -4251
rect 17473 -4439 17519 -4427
rect 17591 -4251 17637 -4239
rect 17591 -4427 17597 -4251
rect 17631 -4427 17637 -4251
rect 17591 -4439 17637 -4427
rect 17893 -4251 17939 -4239
rect 16467 -4639 16513 -4627
rect 16355 -4733 16389 -4639
rect 16879 -4733 16912 -4439
rect 14708 -4754 14816 -4744
rect 14577 -4802 14708 -4754
rect 14494 -4826 14708 -4802
rect 14454 -4838 14708 -4826
rect 13466 -4842 14051 -4840
rect 14460 -4842 14708 -4838
rect 13466 -4870 14096 -4842
rect 13466 -4876 14333 -4870
rect 13466 -4910 14283 -4876
rect 14317 -4910 14333 -4876
rect 13466 -4926 14333 -4910
rect 14385 -4876 14451 -4870
rect 14385 -4910 14401 -4876
rect 14435 -4910 14451 -4876
rect 14634 -4886 14708 -4842
rect 15698 -4765 16912 -4733
rect 17596 -4733 17630 -4439
rect 17893 -4627 17899 -4251
rect 17933 -4627 17939 -4251
rect 17893 -4639 17939 -4627
rect 18011 -4251 18057 -4239
rect 18011 -4627 18017 -4251
rect 18051 -4627 18057 -4251
rect 18011 -4639 18057 -4627
rect 18129 -4251 18175 -4239
rect 18129 -4627 18135 -4251
rect 18169 -4627 18175 -4251
rect 18129 -4639 18175 -4627
rect 18247 -4251 18293 -4239
rect 18247 -4627 18253 -4251
rect 18287 -4627 18293 -4251
rect 18247 -4639 18293 -4627
rect 18365 -4251 18411 -4239
rect 18365 -4627 18371 -4251
rect 18405 -4627 18411 -4251
rect 18771 -4251 18817 -4239
rect 18771 -4427 18777 -4251
rect 18811 -4427 18817 -4251
rect 18771 -4439 18817 -4427
rect 18889 -4251 18935 -4239
rect 18889 -4427 18895 -4251
rect 18929 -4427 18935 -4251
rect 18889 -4439 18935 -4427
rect 18365 -4639 18411 -4627
rect 18253 -4733 18287 -4639
rect 18777 -4733 18810 -4439
rect 17596 -4765 18810 -4733
rect 16191 -4850 16323 -4765
rect 18089 -4850 18221 -4765
rect 14708 -4896 14816 -4886
rect 13466 -4942 14096 -4926
rect 13466 -4946 14051 -4942
rect 13466 -4947 13567 -4946
rect 13996 -4995 14096 -4984
rect 13960 -5101 13970 -4995
rect 14082 -5006 14096 -4995
rect 14385 -5006 14451 -4910
rect 16181 -4958 16191 -4850
rect 16323 -4958 16333 -4850
rect 18079 -4958 18089 -4850
rect 18221 -4958 18231 -4850
rect 19010 -4878 19077 -3495
rect 19138 -3924 19294 -3918
rect 19138 -4022 19150 -3924
rect 19282 -4022 19294 -3924
rect 19138 -4028 19294 -4022
rect 14082 -5054 14451 -5006
rect 14082 -5084 14096 -5054
rect 14082 -5101 14092 -5084
rect 14384 -5157 14450 -5054
rect 19010 -5157 19076 -4878
rect 14382 -5237 19076 -5157
<< via1 >>
rect 14419 -569 14551 -461
rect 16901 -515 17033 -407
rect 17302 -505 17358 -491
rect 17302 -539 17318 -505
rect 17318 -539 17352 -505
rect 17352 -539 17358 -505
rect 17302 -557 17358 -539
rect 18048 -515 18180 -407
rect 16172 -629 16238 -613
rect 16172 -663 16188 -629
rect 16188 -663 16222 -629
rect 16222 -663 16238 -629
rect 16172 -679 16238 -663
rect 16838 -1326 16937 -1229
rect 14699 -1632 14807 -1500
rect 13191 -2210 13303 -2104
rect 13190 -3218 13302 -3216
rect 13190 -3322 13308 -3218
rect 13196 -3324 13308 -3322
rect 16247 -1915 16379 -1807
rect 13685 -2193 13797 -2087
rect 14433 -2219 14565 -2111
rect 17994 -1303 18059 -1249
rect 19089 -1315 19157 -1240
rect 17389 -1917 17521 -1809
rect 16246 -2562 16378 -2454
rect 18144 -2562 18276 -2454
rect 13968 -3324 14086 -3206
rect 14713 -3282 14821 -3150
rect 13465 -3666 13558 -3587
rect 14428 -3823 14560 -3715
rect 16891 -3440 16954 -3424
rect 16891 -3474 16920 -3440
rect 16920 -3474 16954 -3440
rect 16891 -3490 16954 -3474
rect 15015 -4518 15078 -4466
rect 14708 -4886 14816 -4754
rect 13970 -5101 14082 -4995
rect 16191 -4958 16323 -4850
rect 18089 -4958 18221 -4850
<< metal2 >>
rect 16890 -396 17043 -386
rect 14408 -450 14561 -440
rect 18037 -396 18190 -386
rect 17302 -491 17358 -481
rect 16890 -535 17043 -525
rect 14408 -589 14561 -579
rect 17177 -557 17302 -495
rect 17358 -557 17359 -495
rect 18037 -535 18190 -525
rect 16172 -606 16238 -603
rect 15246 -613 16238 -606
rect 15246 -679 16172 -613
rect 14679 -1642 14689 -1489
rect 14818 -1642 14828 -1489
rect 13179 -2077 13346 -2076
rect 13686 -2077 13802 -2076
rect 13179 -2087 13802 -2077
rect 13179 -2104 13685 -2087
rect 13179 -2210 13191 -2104
rect 13303 -2193 13685 -2104
rect 13797 -2193 13802 -2087
rect 13303 -2210 13802 -2193
rect 13179 -2219 13802 -2210
rect 14422 -2100 14575 -2090
rect 14422 -2239 14575 -2229
rect 13178 -3198 13343 -3188
rect 13178 -3199 13346 -3198
rect 13968 -3199 14086 -3196
rect 13178 -3206 14086 -3199
rect 13178 -3216 13968 -3206
rect 13178 -3322 13190 -3216
rect 13302 -3218 13968 -3216
rect 13178 -3324 13196 -3322
rect 13308 -3324 13968 -3218
rect 14693 -3292 14703 -3139
rect 14832 -3292 14842 -3139
rect 13178 -3331 14086 -3324
rect 13184 -3333 14086 -3331
rect 13221 -3334 14086 -3333
rect 13455 -3578 13570 -3568
rect 13455 -3685 13570 -3675
rect 13965 -4985 14081 -3334
rect 14417 -3704 14570 -3694
rect 14417 -3843 14570 -3833
rect 15015 -4462 15078 -4456
rect 15246 -4462 15314 -679
rect 16172 -689 16238 -679
rect 17177 -1218 17237 -557
rect 17302 -567 17358 -557
rect 17099 -1219 17237 -1218
rect 16837 -1229 17237 -1219
rect 16837 -1326 16838 -1229
rect 16937 -1326 17237 -1229
rect 17994 -1240 18059 -1239
rect 19089 -1240 19157 -1230
rect 17993 -1249 19089 -1240
rect 17993 -1303 17994 -1249
rect 18059 -1303 19089 -1249
rect 17993 -1314 19089 -1303
rect 19089 -1325 19157 -1315
rect 16837 -1334 17237 -1326
rect 16837 -1338 17146 -1334
rect 16237 -1797 16390 -1787
rect 16237 -1936 16390 -1926
rect 17379 -1799 17532 -1789
rect 17379 -1938 17532 -1928
rect 16235 -2443 16388 -2433
rect 16235 -2582 16388 -2572
rect 18133 -2443 18286 -2433
rect 18133 -2582 18286 -2572
rect 16876 -3414 16954 -3404
rect 16876 -3510 16954 -3500
rect 15010 -4466 15314 -4462
rect 15010 -4518 15015 -4466
rect 15078 -4518 15314 -4466
rect 15010 -4524 15314 -4518
rect 15015 -4528 15078 -4524
rect 14688 -4896 14698 -4743
rect 14827 -4896 14837 -4743
rect 16181 -4840 16334 -4830
rect 16181 -4979 16334 -4969
rect 18079 -4840 18232 -4830
rect 18079 -4979 18232 -4969
rect 13965 -4995 14082 -4985
rect 13965 -5101 13970 -4995
rect 13965 -5111 14082 -5101
rect 13965 -5112 14081 -5111
<< via2 >>
rect 16890 -407 17043 -396
rect 14408 -461 14561 -450
rect 14408 -569 14419 -461
rect 14419 -569 14551 -461
rect 14551 -569 14561 -461
rect 16890 -515 16901 -407
rect 16901 -515 17033 -407
rect 17033 -515 17043 -407
rect 18037 -407 18190 -396
rect 16890 -525 17043 -515
rect 14408 -579 14561 -569
rect 18037 -515 18048 -407
rect 18048 -515 18180 -407
rect 18180 -515 18190 -407
rect 18037 -525 18190 -515
rect 14689 -1500 14818 -1489
rect 14689 -1632 14699 -1500
rect 14699 -1632 14807 -1500
rect 14807 -1632 14818 -1500
rect 14689 -1642 14818 -1632
rect 14422 -2111 14575 -2100
rect 14422 -2219 14433 -2111
rect 14433 -2219 14565 -2111
rect 14565 -2219 14575 -2111
rect 14422 -2229 14575 -2219
rect 14703 -3150 14832 -3139
rect 14703 -3282 14713 -3150
rect 14713 -3282 14821 -3150
rect 14821 -3282 14832 -3150
rect 14703 -3292 14832 -3282
rect 13455 -3587 13570 -3578
rect 13455 -3666 13465 -3587
rect 13465 -3666 13558 -3587
rect 13558 -3666 13570 -3587
rect 13455 -3675 13570 -3666
rect 14417 -3715 14570 -3704
rect 14417 -3823 14428 -3715
rect 14428 -3823 14560 -3715
rect 14560 -3823 14570 -3715
rect 14417 -3833 14570 -3823
rect 16237 -1807 16390 -1797
rect 16237 -1915 16247 -1807
rect 16247 -1915 16379 -1807
rect 16379 -1915 16390 -1807
rect 16237 -1926 16390 -1915
rect 17379 -1809 17532 -1799
rect 17379 -1917 17389 -1809
rect 17389 -1917 17521 -1809
rect 17521 -1917 17532 -1809
rect 17379 -1928 17532 -1917
rect 16235 -2454 16388 -2443
rect 16235 -2562 16246 -2454
rect 16246 -2562 16378 -2454
rect 16378 -2562 16388 -2454
rect 16235 -2572 16388 -2562
rect 18133 -2454 18286 -2443
rect 18133 -2562 18144 -2454
rect 18144 -2562 18276 -2454
rect 18276 -2562 18286 -2454
rect 18133 -2572 18286 -2562
rect 16876 -3424 16954 -3414
rect 16876 -3490 16891 -3424
rect 16891 -3490 16954 -3424
rect 16876 -3500 16954 -3490
rect 14698 -4754 14827 -4743
rect 14698 -4886 14708 -4754
rect 14708 -4886 14816 -4754
rect 14816 -4886 14827 -4754
rect 14698 -4896 14827 -4886
rect 16181 -4850 16334 -4840
rect 16181 -4958 16191 -4850
rect 16191 -4958 16323 -4850
rect 16323 -4958 16334 -4850
rect 16181 -4969 16334 -4958
rect 18079 -4850 18232 -4840
rect 18079 -4958 18089 -4850
rect 18089 -4958 18221 -4850
rect 18221 -4958 18232 -4850
rect 18079 -4969 18232 -4958
<< metal3 >>
rect 14376 -598 14386 -419
rect 14585 -598 14595 -419
rect 16858 -544 16868 -365
rect 17067 -544 17077 -365
rect 18005 -544 18015 -365
rect 18214 -544 18224 -365
rect 14670 -1467 14849 -1457
rect 14670 -1675 14849 -1666
rect 16204 -1957 16213 -1778
rect 16412 -1957 16422 -1778
rect 17346 -1959 17355 -1780
rect 17554 -1959 17564 -1780
rect 14390 -2248 14400 -2069
rect 14599 -2248 14609 -2069
rect 16203 -2591 16213 -2412
rect 16412 -2591 16422 -2412
rect 18101 -2591 18111 -2412
rect 18310 -2591 18320 -2412
rect 14684 -3117 14863 -3107
rect 14684 -3325 14863 -3316
rect 13466 -3410 13558 -3409
rect 16864 -3410 16968 -3408
rect 13466 -3414 16968 -3410
rect 13466 -3500 16876 -3414
rect 16954 -3500 16968 -3414
rect 13466 -3513 16968 -3500
rect 13466 -3573 13558 -3513
rect 13445 -3578 13580 -3573
rect 13445 -3675 13455 -3578
rect 13570 -3675 13580 -3578
rect 13445 -3680 13580 -3675
rect 14385 -3852 14395 -3673
rect 14594 -3852 14604 -3673
rect 14679 -4721 14858 -4711
rect 14679 -4929 14858 -4920
rect 16147 -5000 16157 -4821
rect 16356 -5000 16366 -4821
rect 18045 -5000 18055 -4821
rect 18254 -5000 18264 -4821
<< via3 >>
rect 14386 -450 14585 -419
rect 14386 -579 14408 -450
rect 14408 -579 14561 -450
rect 14561 -579 14585 -450
rect 14386 -598 14585 -579
rect 16868 -396 17067 -365
rect 16868 -525 16890 -396
rect 16890 -525 17043 -396
rect 17043 -525 17067 -396
rect 16868 -544 17067 -525
rect 18015 -396 18214 -365
rect 18015 -525 18037 -396
rect 18037 -525 18190 -396
rect 18190 -525 18214 -396
rect 18015 -544 18214 -525
rect 14670 -1489 14849 -1467
rect 14670 -1642 14689 -1489
rect 14689 -1642 14818 -1489
rect 14818 -1642 14849 -1489
rect 14670 -1666 14849 -1642
rect 16213 -1797 16412 -1778
rect 16213 -1926 16237 -1797
rect 16237 -1926 16390 -1797
rect 16390 -1926 16412 -1797
rect 16213 -1957 16412 -1926
rect 17355 -1799 17554 -1780
rect 17355 -1928 17379 -1799
rect 17379 -1928 17532 -1799
rect 17532 -1928 17554 -1799
rect 17355 -1959 17554 -1928
rect 14400 -2100 14599 -2069
rect 14400 -2229 14422 -2100
rect 14422 -2229 14575 -2100
rect 14575 -2229 14599 -2100
rect 14400 -2248 14599 -2229
rect 16213 -2443 16412 -2412
rect 16213 -2572 16235 -2443
rect 16235 -2572 16388 -2443
rect 16388 -2572 16412 -2443
rect 16213 -2591 16412 -2572
rect 18111 -2443 18310 -2412
rect 18111 -2572 18133 -2443
rect 18133 -2572 18286 -2443
rect 18286 -2572 18310 -2443
rect 18111 -2591 18310 -2572
rect 14684 -3139 14863 -3117
rect 14684 -3292 14703 -3139
rect 14703 -3292 14832 -3139
rect 14832 -3292 14863 -3139
rect 14684 -3316 14863 -3292
rect 14395 -3704 14594 -3673
rect 14395 -3833 14417 -3704
rect 14417 -3833 14570 -3704
rect 14570 -3833 14594 -3704
rect 14395 -3852 14594 -3833
rect 14679 -4743 14858 -4721
rect 14679 -4896 14698 -4743
rect 14698 -4896 14827 -4743
rect 14827 -4896 14858 -4743
rect 14679 -4920 14858 -4896
rect 16157 -4840 16356 -4821
rect 16157 -4969 16181 -4840
rect 16181 -4969 16334 -4840
rect 16334 -4969 16356 -4840
rect 16157 -5000 16356 -4969
rect 18055 -4840 18254 -4821
rect 18055 -4969 18079 -4840
rect 18079 -4969 18232 -4840
rect 18232 -4969 18254 -4840
rect 18055 -5000 18254 -4969
<< metal4 >>
rect 14364 -259 18797 -94
rect 14365 -365 18793 -259
rect 14365 -419 16868 -365
rect 14365 -598 14386 -419
rect 14585 -544 16868 -419
rect 17067 -544 18015 -365
rect 18214 -544 18793 -365
rect 14585 -598 18793 -544
rect 14365 -804 18793 -598
rect 13845 -2069 14740 -1855
rect 13845 -2248 14400 -2069
rect 14599 -2237 14740 -2069
rect 14599 -2242 15085 -2237
rect 16963 -2242 17310 -2239
rect 18177 -2242 18793 -804
rect 14599 -2248 18793 -2242
rect 13845 -2412 18793 -2248
rect 13845 -2591 16213 -2412
rect 16412 -2591 18111 -2412
rect 18310 -2591 18793 -2412
rect 13845 -2747 18793 -2591
rect 13845 -3477 14015 -2747
rect 18177 -2752 18793 -2747
rect 13845 -3673 15113 -3477
rect 13845 -3852 14395 -3673
rect 14594 -3852 15113 -3673
rect 13845 -4121 15113 -3852
rect 16133 -4821 16378 -4818
rect 16133 -4839 16157 -4821
rect 16356 -4839 16378 -4821
rect 18031 -4821 18276 -4818
rect 18031 -4839 18055 -4821
rect 18254 -4839 18276 -4821
rect 16029 -5143 16053 -4906
rect 16563 -5143 17899 -4957
rect 16029 -5148 18396 -5143
rect 16417 -5150 18088 -5148
<< via4 >>
rect 14611 -1467 15121 -1389
rect 14611 -1666 14670 -1467
rect 14670 -1666 14849 -1467
rect 14849 -1666 15121 -1467
rect 14611 -1693 15121 -1666
rect 16179 -1778 16483 -1627
rect 16179 -1957 16213 -1778
rect 16213 -1957 16412 -1778
rect 16412 -1957 16483 -1778
rect 16179 -2137 16483 -1957
rect 17313 -1780 17617 -1617
rect 17313 -1959 17355 -1780
rect 17355 -1959 17554 -1780
rect 17554 -1959 17617 -1780
rect 17313 -2127 17617 -1959
rect 14605 -3117 15115 -3049
rect 14605 -3316 14684 -3117
rect 14684 -3316 14863 -3117
rect 14863 -3316 15115 -3117
rect 14605 -3353 15115 -3316
rect 14604 -4721 15114 -4654
rect 14604 -4920 14679 -4721
rect 14679 -4920 14858 -4721
rect 14858 -4920 15114 -4721
rect 14604 -4958 15114 -4920
rect 16053 -5000 16157 -4839
rect 16157 -5000 16356 -4839
rect 16356 -5000 16563 -4839
rect 16053 -5143 16563 -5000
rect 17899 -5000 18055 -4839
rect 18055 -5000 18254 -4839
rect 18254 -5000 18409 -4839
rect 17899 -5143 18409 -5000
<< metal5 >>
rect 14460 -1389 18434 -1225
rect 14460 -1693 14611 -1389
rect 15121 -1617 18434 -1389
rect 15121 -1627 17313 -1617
rect 15121 -1693 16179 -1627
rect 14460 -2137 16179 -1693
rect 16483 -2127 17313 -1627
rect 17617 -2127 18434 -1617
rect 16483 -2137 18434 -2127
rect 14460 -3049 18434 -2137
rect 14460 -3353 14605 -3049
rect 15115 -3353 18434 -3049
rect 14460 -4654 18434 -3353
rect 14460 -4958 14604 -4654
rect 15114 -4839 18434 -4654
rect 15114 -4958 16053 -4839
rect 14460 -5143 16053 -4958
rect 16563 -5143 17899 -4839
rect 18409 -5143 18434 -4839
rect 14460 -5604 18434 -5143
use fulladder  fulladder_0 ~/Desktop/design4/mag/Full_Adder
timestamp 1735941024
transform 1 0 21956 0 1 -5144
box -2361 -464 3896 5054
use fulladder  fulladder_1
timestamp 1735941024
transform 1 0 2351 0 1 -5140
box -2361 -464 3896 5054
use fulladder  fulladder_2
timestamp 1735941024
transform 1 0 8864 0 1 -5143
box -2361 -464 3896 5054
use fulladder  fulladder_3
timestamp 1735941024
transform 1 0 15398 0 1 456
box -2361 -464 3896 5054
use fulladder  fulladder_4
timestamp 1735941024
transform 1 0 21956 0 1 460
box -2361 -464 3896 5054
use fulladder  fulladder_5
timestamp 1735941024
transform 1 0 8864 0 1 461
box -2361 -464 3896 5054
use fulladder  fulladder_6
timestamp 1735941024
transform 1 0 2351 0 1 464
box -2361 -464 3896 5054
<< end >>
