* NGSPICE file created from fulladder_pex.ext - technology: sky130B

.subckt fulladder A B carry_in VDD VSS carry_out Y
X0 a_n710_2114.t3 a_n1300_2551.t7 VDD.t35 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 VDD.t32 carry_in.t0 a_2783_1215.t2 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 VDD.t7 a_591_1241.t8 a_1944_1934.t2 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 a_827_509.t1 B.t0 a_591_1241.t1 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 VDD.t49 a_1157_3490.t4 a_2153_4077.t5 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X5 a_591_509.t0 a_885_1215.t4 VSS.t10 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X6 VDD.t10 a_591_1241.t9 a_2371_1241.t8 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 VDD.t26 a_n724_3764.t4 a_1011_4073.t2 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 a_n724_3764.t0 a_n1314_4201.t7 VDD.t31 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 a_n1063_1914.t1 carry_in.t1 a_n1300_2551.t2 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 VDD.t39 B.t1 a_n1314_4201.t3 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X11 VSS.t9 a_591_1241.t10 a_1944_1934.t3 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X12 VDD.t2 a_591_1241.t11 a_1944_1934.t1 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 a_n1068_310.t0 A.t0 a_n1305_947.t3 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 a_885_1215.t0 A.t1 VDD.t3 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 a_885_1215.t2 A.t2 VSS.t4 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 a_n715_510.t2 a_n1305_947.t7 VDD.t58 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X17 VDD.t45 B.t2 a_46_1934.t2 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X18 a_2371_1241.t0 a_1944_1934.t4 Y.t3 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 VDD.t19 A.t3 a_473_1241.t5 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 a_1157_3490.t1 a_893_4073.t5 VDD.t20 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X21 a_591_1241.t5 a_46_1934.t4 a_591_509.t1 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 VDD.t25 A.t4 a_473_1241.t4 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 a_1011_4073.t5 a_n715_510.t4 a_893_4073.t4 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 VDD.t33 carry_in.t2 a_n1300_2551.t4 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 VSS.t18 a_1157_3490.t5 a_2035_4077.t4 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VSS.t13 carry_in.t3 a_n1068_310.t1 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X27 a_1011_4073.t4 a_n715_510.t5 a_893_4073.t3 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X28 VSS.t7 B.t3 a_46_1934.t3 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 a_473_1241.t8 a_885_1215.t5 a_591_1241.t6 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X30 VDD.t47 A.t5 a_n1314_4201.t5 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 VDD.t57 a_n1305_947.t8 a_n715_510.t1 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X32 a_2783_1215.t1 carry_in.t4 VDD.t8 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X33 a_n710_2114.t2 a_n1300_2551.t8 VDD.t34 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 a_473_1241.t7 a_885_1215.t6 a_591_1241.t7 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X35 a_n1305_947.t2 A.t6 VDD.t1 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X36 a_2153_4077.t2 a_n710_2114.t4 a_2035_4077.t3 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X37 a_n1077_3564.t1 A.t7 a_n1314_4201.t6 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 VDD.t13 a_1157_3490.t6 a_2153_4077.t4 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 a_1011_4073.t1 a_n724_3764.t5 VDD.t0 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X40 VDD.t16 carry_in.t5 a_2371_1241.t11 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X41 VSS.t6 B.t4 a_n1063_1914.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X42 a_n724_3764.t3 a_n1314_4201.t8 VDD.t61 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 a_2783_1215.t0 carry_in.t6 VDD.t62 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X44 a_473_1241.t2 B.t5 VDD.t15 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X45 a_n710_2114.t0 a_n1300_2551.t9 VSS.t15 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 a_n1300_2551.t5 B.t6 VDD.t46 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X47 a_n715_510.t0 a_n1305_947.t9 VDD.t56 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X48 VDD.t43 A.t8 a_885_1215.t3 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X49 a_46_1934.t1 B.t7 VDD.t37 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X50 a_n1314_4201.t2 B.t8 VDD.t24 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 Y.t2 a_1944_1934.t5 a_2371_1241.t2 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 a_2371_1241.t3 a_2783_1215.t4 Y.t6 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 a_473_1241.t1 B.t9 VDD.t29 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 carry_out.t2 a_2035_4077.t5 VDD.t21 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X55 VDD.t22 A.t9 a_n1305_947.t1 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 a_2153_4077.t1 a_n710_2114.t5 a_2035_4077.t2 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X57 a_591_1241.t2 a_46_1934.t5 a_473_1241.t11 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X58 a_893_4073.t1 a_n715_510.t6 VSS.t19 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X59 a_n1300_2551.t3 carry_in.t7 VDD.t23 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X60 a_2783_1215.t3 carry_in.t8 VSS.t11 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 a_2035_4077.t0 a_n710_2114.t6 VSS.t2 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 VDD.t28 a_893_4073.t6 a_1157_3490.t2 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_1157_3490.t0 a_893_4073.t7 VSS.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X64 a_893_4073.t2 a_n715_510.t7 a_1011_4073.t3 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X65 a_591_1241.t4 a_46_1934.t6 a_473_1241.t10 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X66 a_2371_1241.t7 a_591_1241.t12 VDD.t44 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X67 a_n1314_4201.t4 A.t10 VDD.t27 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X68 a_n1300_2551.t6 carry_in.t9 VDD.t60 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 VSS.t12 carry_in.t10 a_2725_509.t1 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X70 carry_out.t3 a_2035_4077.t6 VSS.t14 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 a_2371_1241.t4 a_2783_1215.t5 Y.t5 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X72 VDD.t36 a_n1300_2551.t10 a_n710_2114.t1 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 a_591_1241.t0 a_885_1215.t7 a_473_1241.t6 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 a_1944_1934.t0 a_591_1241.t13 VDD.t5 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 a_n1305_947.t0 A.t11 VDD.t52 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 VSS.t5 B.t10 a_n1077_3564.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X77 a_2153_4077.t3 a_1157_3490.t7 VDD.t9 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X78 a_2371_1241.t6 a_591_1241.t14 VDD.t40 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X79 VDD.t50 a_n724_3764.t6 a_1011_4073.t0 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X80 VDD.t59 a_n1314_4201.t9 a_n724_3764.t2 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X81 a_2489_509.t1 a_2783_1215.t6 VSS.t8 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X82 VDD.t14 B.t11 a_n1300_2551.t1 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X83 a_885_1215.t1 A.t12 VDD.t17 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 VDD.t53 a_893_4073.t8 a_1157_3490.t3 w_857_4011# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 a_2371_1241.t10 carry_in.t11 VDD.t48 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X86 a_n1305_947.t6 carry_in.t12 VDD.t6 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X87 VDD.t42 carry_in.t13 a_2371_1241.t9 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 VDD.t30 B.t12 a_46_1934.t0 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 a_2725_509.t0 a_591_1241.t15 Y.t7 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 Y.t1 a_1944_1934.t6 a_2371_1241.t1 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X91 VDD.t41 carry_in.t14 a_n1305_947.t5 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X92 a_473_1241.t3 A.t13 VDD.t51 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 VDD.t38 a_2035_4077.t7 carry_out.t1 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X94 VDD.t55 B.t13 a_473_1241.t0 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X95 VSS.t3 A.t14 a_827_509.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X96 VDD.t12 B.t14 a_n1300_2551.t0 w_n1454_2489# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X97 VDD.t54 a_2035_4077.t8 carry_out.t0 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X98 Y.t4 a_2783_1215.t7 a_2371_1241.t5 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X99 a_n724_3764.t1 a_n1314_4201.t10 VSS.t16 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X100 a_n715_510.t3 a_n1305_947.t10 VSS.t17 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X101 a_473_1241.t9 a_46_1934.t7 a_591_1241.t3 w_9_1872# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X102 a_2035_4077.t1 a_n710_2114.t7 a_2153_4077.t0 w_1999_4015# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X103 VDD.t11 B.t15 a_n1314_4201.t1 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X104 VSS.t1 a_n724_3764.t7 a_893_4073.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X105 a_n1314_4201.t0 A.t15 VDD.t18 w_n1468_4139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X106 VDD.t4 carry_in.t15 a_n1305_947.t4 w_n1459_885# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X107 Y.t0 a_1944_1934.t7 a_2489_509.t0 a_n659_3505# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
R0 a_n1300_2551.n2 a_n1300_2551.t7 214.335
R1 a_n1300_2551.t8 a_n1300_2551.n2 214.335
R2 a_n1300_2551.n3 a_n1300_2551.t8 143.851
R3 a_n1300_2551.n3 a_n1300_2551.t9 135.658
R4 a_n1300_2551.n2 a_n1300_2551.t10 80.333
R5 a_n1300_2551.n4 a_n1300_2551.t1 28.565
R6 a_n1300_2551.n4 a_n1300_2551.t5 28.565
R7 a_n1300_2551.n0 a_n1300_2551.t4 28.565
R8 a_n1300_2551.n0 a_n1300_2551.t6 28.565
R9 a_n1300_2551.t0 a_n1300_2551.n7 28.565
R10 a_n1300_2551.n7 a_n1300_2551.t3 28.565
R11 a_n1300_2551.n1 a_n1300_2551.t2 9.714
R12 a_n1300_2551.n1 a_n1300_2551.n0 1.003
R13 a_n1300_2551.n6 a_n1300_2551.n5 0.833
R14 a_n1300_2551.n5 a_n1300_2551.n4 0.653
R15 a_n1300_2551.n7 a_n1300_2551.n6 0.653
R16 a_n1300_2551.n6 a_n1300_2551.n1 0.341
R17 a_n1300_2551.n5 a_n1300_2551.n3 0.032
R18 VDD.n58 VDD.t18 30.163
R19 VDD.n20 VDD.t60 30.163
R20 VDD.n12 VDD.t1 30.163
R21 VDD.n40 VDD.t2 28.664
R22 VDD.n45 VDD.t8 28.664
R23 VDD.n28 VDD.t45 28.664
R24 VDD.n33 VDD.t17 28.664
R25 VDD.n2 VDD.t28 28.57
R26 VDD.n7 VDD.t54 28.57
R27 VDD.n1 VDD.t20 28.565
R28 VDD.n1 VDD.t53 28.565
R29 VDD.n6 VDD.t21 28.565
R30 VDD.n6 VDD.t38 28.565
R31 VDD.n57 VDD.t27 28.565
R32 VDD.n57 VDD.t47 28.565
R33 VDD.n53 VDD.t31 28.565
R34 VDD.n53 VDD.t59 28.565
R35 VDD.n54 VDD.t61 28.565
R36 VDD.n54 VDD.t39 28.565
R37 VDD.n56 VDD.t24 28.565
R38 VDD.n56 VDD.t11 28.565
R39 VDD.n41 VDD.t5 28.565
R40 VDD.n41 VDD.t7 28.565
R41 VDD.n46 VDD.t62 28.565
R42 VDD.n46 VDD.t32 28.565
R43 VDD.n29 VDD.t37 28.565
R44 VDD.n29 VDD.t30 28.565
R45 VDD.n34 VDD.t3 28.565
R46 VDD.n34 VDD.t43 28.565
R47 VDD.n19 VDD.t23 28.565
R48 VDD.n19 VDD.t33 28.565
R49 VDD.n22 VDD.t35 28.565
R50 VDD.n22 VDD.t36 28.565
R51 VDD.n23 VDD.t34 28.565
R52 VDD.n23 VDD.t14 28.565
R53 VDD.n18 VDD.t46 28.565
R54 VDD.n18 VDD.t12 28.565
R55 VDD.n11 VDD.t52 28.565
R56 VDD.n11 VDD.t22 28.565
R57 VDD.n14 VDD.t56 28.565
R58 VDD.n14 VDD.t57 28.565
R59 VDD.n15 VDD.t58 28.565
R60 VDD.n15 VDD.t4 28.565
R61 VDD.n10 VDD.t6 28.565
R62 VDD.n10 VDD.t41 28.565
R63 VDD.n3 VDD.t26 14.284
R64 VDD.n8 VDD.t13 14.284
R65 VDD.n40 VDD.t44 14.284
R66 VDD.n45 VDD.t42 14.284
R67 VDD.n28 VDD.t15 14.284
R68 VDD.n33 VDD.t25 14.284
R69 VDD.n0 VDD.t0 14.282
R70 VDD.n0 VDD.t50 14.282
R71 VDD.n5 VDD.t9 14.282
R72 VDD.n5 VDD.t49 14.282
R73 VDD.n39 VDD.t40 14.282
R74 VDD.n39 VDD.t10 14.282
R75 VDD.n44 VDD.t48 14.282
R76 VDD.n44 VDD.t16 14.282
R77 VDD.n27 VDD.t29 14.282
R78 VDD.n27 VDD.t55 14.282
R79 VDD.n32 VDD.t51 14.282
R80 VDD.n32 VDD.t19 14.282
R81 VDD.n49 VDD.n43 4.276
R82 VDD.n37 VDD.n31 4.276
R83 VDD.n42 VDD.n41 2.451
R84 VDD.n30 VDD.n29 2.451
R85 VDD.n47 VDD.n46 2.449
R86 VDD.n35 VDD.n34 2.449
R87 VDD.n3 VDD.n2 2.195
R88 VDD.n8 VDD.n7 2.195
R89 VDD.n9 VDD.n5 1.72
R90 VDD.n4 VDD.n0 1.698
R91 VDD.n2 VDD.n1 1.651
R92 VDD.n7 VDD.n6 1.651
R93 VDD.n55 VDD.n53 1.564
R94 VDD.n24 VDD.n22 1.564
R95 VDD.n16 VDD.n14 1.564
R96 VDD.n43 VDD.n39 0.922
R97 VDD.n48 VDD.n44 0.922
R98 VDD.n31 VDD.n27 0.922
R99 VDD.n36 VDD.n32 0.922
R100 VDD.n42 VDD.n40 0.921
R101 VDD.n47 VDD.n45 0.921
R102 VDD.n30 VDD.n28 0.921
R103 VDD.n35 VDD.n33 0.921
R104 VDD.n4 VDD.n3 0.806
R105 VDD.n9 VDD.n8 0.778
R106 VDD.n58 VDD.n57 0.747
R107 VDD.n55 VDD.n54 0.747
R108 VDD.n20 VDD.n19 0.747
R109 VDD.n24 VDD.n23 0.747
R110 VDD.n12 VDD.n11 0.747
R111 VDD.n16 VDD.n15 0.747
R112 VDD.n59 VDD.n56 0.689
R113 VDD.n21 VDD.n18 0.689
R114 VDD.n13 VDD.n10 0.689
R115 VDD.n43 VDD.n42 0.686
R116 VDD.n48 VDD.n47 0.686
R117 VDD.n31 VDD.n30 0.686
R118 VDD.n36 VDD.n35 0.686
R119 VDD.n59 VDD.n58 0.59
R120 VDD.n21 VDD.n20 0.59
R121 VDD.n13 VDD.n12 0.59
R122 VDD.n60 VDD.n55 0.451
R123 VDD.n25 VDD.n24 0.451
R124 VDD.n17 VDD.n16 0.451
R125 VDD.n26 VDD.n17 0.276
R126 VDD.n52 VDD.n4 0.253
R127 VDD.n51 VDD.n9 0.241
R128 VDD.n49 VDD.n48 0.179
R129 VDD.n37 VDD.n36 0.179
R130 VDD.n50 VDD.n38 0.174
R131 VDD.n38 VDD.n26 0.161
R132 VDD.n51 VDD.n50 0.153
R133 VDD.n38 VDD.n37 0.142
R134 VDD.n50 VDD.n49 0.141
R135 VDD VDD.n52 0.081
R136 VDD.n52 VDD.n51 0.078
R137 VDD VDD.n60 0.04
R138 VDD.n60 VDD.n59 0.011
R139 VDD.n25 VDD.n21 0.011
R140 VDD.n17 VDD.n13 0.011
R141 VDD.n26 VDD.n25 0.001
R142 a_n710_2114.t5 a_n710_2114.t6 574.43
R143 a_n710_2114.n1 a_n710_2114.t4 285.109
R144 a_n710_2114.n3 a_n710_2114.n2 211.136
R145 a_n710_2114.n4 a_n710_2114.n0 192.754
R146 a_n710_2114.n1 a_n710_2114.t7 160.666
R147 a_n710_2114.n2 a_n710_2114.t5 160.666
R148 a_n710_2114.n2 a_n710_2114.n1 114.829
R149 a_n710_2114.t3 a_n710_2114.n4 28.568
R150 a_n710_2114.n0 a_n710_2114.t1 28.565
R151 a_n710_2114.n0 a_n710_2114.t2 28.565
R152 a_n710_2114.n3 a_n710_2114.t0 19.084
R153 a_n710_2114.n4 a_n710_2114.n3 1.051
R154 carry_in.n5 carry_in.n4 501.28
R155 carry_in.t1 carry_in.t7 437.233
R156 carry_in.t3 carry_in.t14 415.315
R157 carry_in.t4 carry_in.n2 313.873
R158 carry_in.n4 carry_in.t10 294.986
R159 carry_in.n1 carry_in.t5 272.288
R160 carry_in.n5 carry_in.t0 236.01
R161 carry_in.n8 carry_in.t1 216.627
R162 carry_in.n6 carry_in.t3 216.111
R163 carry_in.n7 carry_in.t9 214.686
R164 carry_in.t7 carry_in.n7 214.686
R165 carry_in.n0 carry_in.t15 214.335
R166 carry_in.t14 carry_in.n0 214.335
R167 carry_in.n3 carry_in.t4 190.152
R168 carry_in.n3 carry_in.t6 190.152
R169 carry_in.n1 carry_in.t11 160.666
R170 carry_in.n2 carry_in.t13 160.666
R171 carry_in.n6 carry_in.n5 148.428
R172 carry_in.n4 carry_in.t8 110.859
R173 carry_in.n2 carry_in.n1 96.129
R174 carry_in.n7 carry_in.t2 80.333
R175 carry_in.n0 carry_in.t12 80.333
R176 carry_in.t0 carry_in.n3 80.333
R177 carry_in.n8 carry_in.n6 2.923
R178 carry_in carry_in.n8 0.732
R179 a_2783_1215.n1 a_2783_1215.t7 318.922
R180 a_2783_1215.n0 a_2783_1215.t4 274.739
R181 a_2783_1215.n0 a_2783_1215.t5 274.739
R182 a_2783_1215.n1 a_2783_1215.t6 269.116
R183 a_2783_1215.t7 a_2783_1215.n0 179.946
R184 a_2783_1215.n2 a_2783_1215.n1 105.178
R185 a_2783_1215.n3 a_2783_1215.t0 29.444
R186 a_2783_1215.t2 a_2783_1215.n4 28.565
R187 a_2783_1215.n4 a_2783_1215.t1 28.565
R188 a_2783_1215.n2 a_2783_1215.t3 18.145
R189 a_2783_1215.n3 a_2783_1215.n2 2.878
R190 a_2783_1215.n4 a_2783_1215.n3 0.764
R191 a_591_1241.t0 a_591_1241.n0 14.282
R192 a_591_1241.n0 a_591_1241.t7 14.282
R193 a_591_1241.n0 a_591_1241.n12 90.436
R194 a_591_1241.n8 a_591_1241.n11 50.575
R195 a_591_1241.n12 a_591_1241.n8 74.302
R196 a_591_1241.n11 a_591_1241.n10 157.665
R197 a_591_1241.n10 a_591_1241.t5 8.7
R198 a_591_1241.n10 a_591_1241.t1 8.7
R199 a_591_1241.n11 a_591_1241.n9 122.999
R200 a_591_1241.n9 a_591_1241.t2 14.282
R201 a_591_1241.n9 a_591_1241.t3 14.282
R202 a_591_1241.n8 a_591_1241.n7 90.416
R203 a_591_1241.n7 a_591_1241.t4 14.282
R204 a_591_1241.n7 a_591_1241.t6 14.282
R205 a_591_1241.n12 a_591_1241.n1 342.688
R206 a_591_1241.n1 a_591_1241.n6 126.566
R207 a_591_1241.n6 a_591_1241.t15 294.653
R208 a_591_1241.n6 a_591_1241.t10 111.663
R209 a_591_1241.n1 a_591_1241.n5 552.333
R210 a_591_1241.n5 a_591_1241.n4 6.615
R211 a_591_1241.n4 a_591_1241.t13 93.989
R212 a_591_1241.n5 a_591_1241.n3 97.816
R213 a_591_1241.n3 a_591_1241.t11 80.333
R214 a_591_1241.n3 a_591_1241.t12 394.151
R215 a_591_1241.t12 a_591_1241.n2 269.523
R216 a_591_1241.n2 a_591_1241.t9 160.666
R217 a_591_1241.n2 a_591_1241.t14 269.523
R218 a_591_1241.n4 a_591_1241.t8 198.043
R219 a_1944_1934.n2 a_1944_1934.t4 318.922
R220 a_1944_1934.n1 a_1944_1934.t5 273.935
R221 a_1944_1934.n1 a_1944_1934.t6 273.935
R222 a_1944_1934.n2 a_1944_1934.t7 269.116
R223 a_1944_1934.n4 a_1944_1934.n0 193.227
R224 a_1944_1934.t4 a_1944_1934.n1 179.142
R225 a_1944_1934.n3 a_1944_1934.n2 106.999
R226 a_1944_1934.t2 a_1944_1934.n4 28.568
R227 a_1944_1934.n0 a_1944_1934.t1 28.565
R228 a_1944_1934.n0 a_1944_1934.t0 28.565
R229 a_1944_1934.n3 a_1944_1934.t3 18.149
R230 a_1944_1934.n4 a_1944_1934.n3 3.726
R231 B.n7 B.n6 861.987
R232 B.n6 B.n5 560.726
R233 B.t10 B.t15 415.315
R234 B.t4 B.t14 415.315
R235 B.n2 B.t5 394.151
R236 B.n5 B.t0 294.653
R237 B.n1 B.t9 269.523
R238 B.t5 B.n1 269.523
R239 B.n9 B.t10 217.716
R240 B.n8 B.t1 214.335
R241 B.t15 B.n8 214.335
R242 B.n0 B.t11 214.335
R243 B.t14 B.n0 214.335
R244 B.n7 B.t4 198.921
R245 B.n3 B.t12 198.043
R246 B.n1 B.t13 160.666
R247 B.n5 B.t3 111.663
R248 B.n4 B.n2 97.816
R249 B.n3 B.t7 93.989
R250 B.n8 B.t8 80.333
R251 B.n2 B.t2 80.333
R252 B.n0 B.t6 80.333
R253 B.n6 B.n4 65.07
R254 B.n9 B.n7 16.411
R255 B.n4 B.n3 6.615
R256 B B.n9 0.455
R257 a_827_509.t0 a_827_509.t1 17.4
R258 a_1157_3490.t4 a_1157_3490.t5 800.071
R259 a_1157_3490.n3 a_1157_3490.n2 672.951
R260 a_1157_3490.n1 a_1157_3490.t6 285.109
R261 a_1157_3490.n2 a_1157_3490.t4 193.602
R262 a_1157_3490.n1 a_1157_3490.t7 160.666
R263 a_1157_3490.n2 a_1157_3490.n1 91.507
R264 a_1157_3490.n0 a_1157_3490.t3 28.57
R265 a_1157_3490.n4 a_1157_3490.t2 28.565
R266 a_1157_3490.t1 a_1157_3490.n4 28.565
R267 a_1157_3490.n0 a_1157_3490.t0 17.638
R268 a_1157_3490.n4 a_1157_3490.n3 0.69
R269 a_1157_3490.n3 a_1157_3490.n0 0.6
R270 a_2153_4077.n0 a_2153_4077.t5 14.282
R271 a_2153_4077.n0 a_2153_4077.t2 14.282
R272 a_2153_4077.n1 a_2153_4077.t4 14.282
R273 a_2153_4077.n1 a_2153_4077.t3 14.282
R274 a_2153_4077.t0 a_2153_4077.n3 14.282
R275 a_2153_4077.n3 a_2153_4077.t1 14.282
R276 a_2153_4077.n3 a_2153_4077.n2 2.546
R277 a_2153_4077.n2 a_2153_4077.n1 2.367
R278 a_2153_4077.n2 a_2153_4077.n0 0.001
R279 a_885_1215.n1 a_885_1215.t7 318.922
R280 a_885_1215.n0 a_885_1215.t5 274.739
R281 a_885_1215.n0 a_885_1215.t6 274.739
R282 a_885_1215.n1 a_885_1215.t4 269.116
R283 a_885_1215.t7 a_885_1215.n0 179.946
R284 a_885_1215.n2 a_885_1215.n1 107.263
R285 a_885_1215.t0 a_885_1215.n4 29.444
R286 a_885_1215.n3 a_885_1215.t3 28.565
R287 a_885_1215.n3 a_885_1215.t1 28.565
R288 a_885_1215.n2 a_885_1215.t2 18.145
R289 a_885_1215.n4 a_885_1215.n2 2.878
R290 a_885_1215.n4 a_885_1215.n3 0.764
R291 VSS.n13 VSS.t11 20.763
R292 VSS.n1 VSS.t4 20.763
R293 VSS.n14 VSS.t9 20.606
R294 VSS.n2 VSS.t7 20.606
R295 VSS.n11 VSS.t17 18.185
R296 VSS.n9 VSS.t15 18.185
R297 VSS.n7 VSS.t16 18.185
R298 VSS.n4 VSS.t2 17.929
R299 VSS.n6 VSS.t19 17.925
R300 VSS.n5 VSS.t0 17.4
R301 VSS.n5 VSS.t1 17.4
R302 VSS.n3 VSS.t14 17.4
R303 VSS.n3 VSS.t18 17.4
R304 VSS.n11 VSS.t13 9.487
R305 VSS.n9 VSS.t6 9.487
R306 VSS.n7 VSS.t5 9.487
R307 VSS.n12 VSS.t8 8.7
R308 VSS.n12 VSS.t12 8.7
R309 VSS.n0 VSS.t10 8.7
R310 VSS.n0 VSS.t3 8.7
R311 VSS.n13 VSS.n12 0.948
R312 VSS.n1 VSS.n0 0.948
R313 VSS.n6 VSS.n5 0.72
R314 VSS.n4 VSS.n3 0.72
R315 VSS.n15 VSS.n14 0.146
R316 VSS.n15 VSS.n2 0.146
R317 VSS.n8 VSS.n4 0.142
R318 VSS.n8 VSS.n6 0.138
R319 VSS.n14 VSS.n13 0.125
R320 VSS.n2 VSS.n1 0.125
R321 VSS.n8 VSS.n7 0.019
R322 VSS.n15 VSS.n11 0.015
R323 VSS.n10 VSS.n9 0.015
R324 VSS.n15 VSS.n10 0.009
R325 VSS.n10 VSS.n8 0.009
R326 VSS VSS.n15 0.001
R327 a_591_509.t0 a_591_509.t1 380.209
R328 a_2371_1241.t0 a_2371_1241.n0 14.282
R329 a_2371_1241.n0 a_2371_1241.t1 14.282
R330 a_2371_1241.n0 a_2371_1241.n9 0.999
R331 a_2371_1241.n9 a_2371_1241.n6 0.575
R332 a_2371_1241.n6 a_2371_1241.n8 0.2
R333 a_2371_1241.n8 a_2371_1241.t4 16.058
R334 a_2371_1241.n8 a_2371_1241.n7 0.999
R335 a_2371_1241.n7 a_2371_1241.t3 14.282
R336 a_2371_1241.n7 a_2371_1241.t5 14.282
R337 a_2371_1241.n9 a_2371_1241.t2 16.058
R338 a_2371_1241.n6 a_2371_1241.n4 0.227
R339 a_2371_1241.n4 a_2371_1241.n5 1.511
R340 a_2371_1241.n5 a_2371_1241.t7 14.282
R341 a_2371_1241.n5 a_2371_1241.t8 14.282
R342 a_2371_1241.n4 a_2371_1241.n1 0.669
R343 a_2371_1241.n1 a_2371_1241.n2 0.001
R344 a_2371_1241.n1 a_2371_1241.n3 267.767
R345 a_2371_1241.n3 a_2371_1241.t10 14.282
R346 a_2371_1241.n3 a_2371_1241.t9 14.282
R347 a_2371_1241.n2 a_2371_1241.t6 14.282
R348 a_2371_1241.n2 a_2371_1241.t11 14.282
R349 a_n724_3764.t6 a_n724_3764.t7 800.071
R350 a_n724_3764.n3 a_n724_3764.n2 659.097
R351 a_n724_3764.n1 a_n724_3764.t4 285.109
R352 a_n724_3764.n2 a_n724_3764.t6 193.602
R353 a_n724_3764.n4 a_n724_3764.n0 192.754
R354 a_n724_3764.n1 a_n724_3764.t5 160.666
R355 a_n724_3764.n2 a_n724_3764.n1 91.507
R356 a_n724_3764.t0 a_n724_3764.n4 28.568
R357 a_n724_3764.n0 a_n724_3764.t2 28.565
R358 a_n724_3764.n0 a_n724_3764.t3 28.565
R359 a_n724_3764.n3 a_n724_3764.t1 19.061
R360 a_n724_3764.n4 a_n724_3764.n3 1.005
R361 a_1011_4073.n0 a_1011_4073.t0 14.282
R362 a_1011_4073.n0 a_1011_4073.t4 14.282
R363 a_1011_4073.n1 a_1011_4073.t2 14.282
R364 a_1011_4073.n1 a_1011_4073.t1 14.282
R365 a_1011_4073.t3 a_1011_4073.n3 14.282
R366 a_1011_4073.n3 a_1011_4073.t5 14.282
R367 a_1011_4073.n3 a_1011_4073.n2 2.546
R368 a_1011_4073.n2 a_1011_4073.n1 2.367
R369 a_1011_4073.n2 a_1011_4073.n0 0.001
R370 a_n1314_4201.n0 a_n1314_4201.t7 214.335
R371 a_n1314_4201.t8 a_n1314_4201.n0 214.335
R372 a_n1314_4201.n1 a_n1314_4201.t8 143.851
R373 a_n1314_4201.n1 a_n1314_4201.t10 135.658
R374 a_n1314_4201.n0 a_n1314_4201.t9 80.333
R375 a_n1314_4201.n2 a_n1314_4201.t3 28.565
R376 a_n1314_4201.n2 a_n1314_4201.t2 28.565
R377 a_n1314_4201.n4 a_n1314_4201.t1 28.565
R378 a_n1314_4201.n4 a_n1314_4201.t4 28.565
R379 a_n1314_4201.n7 a_n1314_4201.t5 28.565
R380 a_n1314_4201.t0 a_n1314_4201.n7 28.565
R381 a_n1314_4201.n6 a_n1314_4201.t6 9.714
R382 a_n1314_4201.n7 a_n1314_4201.n6 1.003
R383 a_n1314_4201.n5 a_n1314_4201.n3 0.833
R384 a_n1314_4201.n3 a_n1314_4201.n2 0.653
R385 a_n1314_4201.n5 a_n1314_4201.n4 0.653
R386 a_n1314_4201.n6 a_n1314_4201.n5 0.341
R387 a_n1314_4201.n3 a_n1314_4201.n1 0.032
R388 a_n1063_1914.t0 a_n1063_1914.t1 17.4
R389 A.n4 A.n3 535.449
R390 A.t7 A.t10 437.233
R391 A.t0 A.t11 437.233
R392 A.t12 A.n1 313.873
R393 A.n3 A.t14 294.986
R394 A.n0 A.t3 272.288
R395 A.n4 A.t8 245.184
R396 A.n6 A.t0 218.628
R397 A.n8 A.t7 217.024
R398 A.n7 A.t15 214.686
R399 A.t10 A.n7 214.686
R400 A.n5 A.t6 214.686
R401 A.t11 A.n5 214.686
R402 A.n2 A.t12 190.152
R403 A.n2 A.t1 190.152
R404 A.n0 A.t13 160.666
R405 A.n1 A.t4 160.666
R406 A.n3 A.t2 110.859
R407 A.n1 A.n0 96.129
R408 A.n7 A.t5 80.333
R409 A.t8 A.n2 80.333
R410 A.n5 A.t9 80.333
R411 A.n6 A.n4 14.9
R412 A.n8 A.n6 2.599
R413 A A.n8 0.289
R414 a_n1305_947.n0 a_n1305_947.t9 214.335
R415 a_n1305_947.t7 a_n1305_947.n0 214.335
R416 a_n1305_947.n1 a_n1305_947.t7 143.851
R417 a_n1305_947.n1 a_n1305_947.t10 135.658
R418 a_n1305_947.n0 a_n1305_947.t8 80.333
R419 a_n1305_947.n2 a_n1305_947.t4 28.565
R420 a_n1305_947.n2 a_n1305_947.t6 28.565
R421 a_n1305_947.n4 a_n1305_947.t5 28.565
R422 a_n1305_947.n4 a_n1305_947.t0 28.565
R423 a_n1305_947.n7 a_n1305_947.t1 28.565
R424 a_n1305_947.t2 a_n1305_947.n7 28.565
R425 a_n1305_947.n6 a_n1305_947.t3 9.714
R426 a_n1305_947.n7 a_n1305_947.n6 1.003
R427 a_n1305_947.n5 a_n1305_947.n3 0.833
R428 a_n1305_947.n3 a_n1305_947.n2 0.653
R429 a_n1305_947.n5 a_n1305_947.n4 0.653
R430 a_n1305_947.n6 a_n1305_947.n5 0.341
R431 a_n1305_947.n3 a_n1305_947.n1 0.032
R432 a_n1068_310.t0 a_n1068_310.t1 17.4
R433 a_n715_510.t4 a_n715_510.t6 574.43
R434 a_n715_510.n0 a_n715_510.t5 285.109
R435 a_n715_510.n2 a_n715_510.n1 197.217
R436 a_n715_510.n4 a_n715_510.n3 192.754
R437 a_n715_510.n0 a_n715_510.t7 160.666
R438 a_n715_510.n1 a_n715_510.t4 160.666
R439 a_n715_510.n1 a_n715_510.n0 114.829
R440 a_n715_510.n3 a_n715_510.t0 28.568
R441 a_n715_510.n4 a_n715_510.t1 28.565
R442 a_n715_510.t2 a_n715_510.n4 28.565
R443 a_n715_510.n2 a_n715_510.t3 18.838
R444 a_n715_510.n3 a_n715_510.n2 1.129
R445 a_46_1934.n1 a_46_1934.t7 318.922
R446 a_46_1934.n0 a_46_1934.t5 273.935
R447 a_46_1934.n0 a_46_1934.t6 273.935
R448 a_46_1934.n1 a_46_1934.t4 269.116
R449 a_46_1934.n4 a_46_1934.n3 193.227
R450 a_46_1934.t7 a_46_1934.n0 179.142
R451 a_46_1934.n2 a_46_1934.n1 106.999
R452 a_46_1934.n3 a_46_1934.t0 28.568
R453 a_46_1934.t2 a_46_1934.n4 28.565
R454 a_46_1934.n4 a_46_1934.t1 28.565
R455 a_46_1934.n2 a_46_1934.t3 18.149
R456 a_46_1934.n3 a_46_1934.n2 3.726
R457 Y.n7 Y.n6 208.992
R458 Y.n4 Y.n2 157.665
R459 Y.n4 Y.n3 122.999
R460 Y.n6 Y.n0 90.436
R461 Y.n5 Y.n1 90.416
R462 Y.n6 Y.n5 74.302
R463 Y.n5 Y.n4 50.575
R464 Y.n0 Y.t5 14.282
R465 Y.n0 Y.t4 14.282
R466 Y.n1 Y.t6 14.282
R467 Y.n1 Y.t1 14.282
R468 Y.n3 Y.t3 14.282
R469 Y.n3 Y.t2 14.282
R470 Y.n2 Y.t7 8.7
R471 Y.n2 Y.t0 8.7
R472 Y.n8 Y.n7 8.62
R473 Y Y.n8 0.039
R474 Y.n8 Y 0.039
R475 a_473_1241.n2 a_473_1241.n0 267.767
R476 a_473_1241.n6 a_473_1241.t11 16.058
R477 a_473_1241.n4 a_473_1241.t7 16.058
R478 a_473_1241.n5 a_473_1241.t10 14.282
R479 a_473_1241.n5 a_473_1241.t9 14.282
R480 a_473_1241.n3 a_473_1241.t6 14.282
R481 a_473_1241.n3 a_473_1241.t8 14.282
R482 a_473_1241.n1 a_473_1241.t5 14.282
R483 a_473_1241.n1 a_473_1241.t1 14.282
R484 a_473_1241.n0 a_473_1241.t4 14.282
R485 a_473_1241.n0 a_473_1241.t3 14.282
R486 a_473_1241.n9 a_473_1241.t0 14.282
R487 a_473_1241.t2 a_473_1241.n9 14.282
R488 a_473_1241.n9 a_473_1241.n8 1.511
R489 a_473_1241.n6 a_473_1241.n5 0.999
R490 a_473_1241.n4 a_473_1241.n3 0.999
R491 a_473_1241.n8 a_473_1241.n2 0.669
R492 a_473_1241.n7 a_473_1241.n6 0.575
R493 a_473_1241.n8 a_473_1241.n7 0.227
R494 a_473_1241.n7 a_473_1241.n4 0.2
R495 a_473_1241.n2 a_473_1241.n1 0.001
R496 a_893_4073.t7 a_893_4073.n3 404.877
R497 a_893_4073.n2 a_893_4073.t6 210.902
R498 a_893_4073.n4 a_893_4073.t7 136.943
R499 a_893_4073.n3 a_893_4073.n2 107.801
R500 a_893_4073.n2 a_893_4073.t5 80.333
R501 a_893_4073.n3 a_893_4073.t8 80.333
R502 a_893_4073.n1 a_893_4073.t0 17.4
R503 a_893_4073.n1 a_893_4073.t1 17.4
R504 a_893_4073.t4 a_893_4073.n5 15.032
R505 a_893_4073.n0 a_893_4073.t3 14.282
R506 a_893_4073.n0 a_893_4073.t2 14.282
R507 a_893_4073.n5 a_893_4073.n0 1.65
R508 a_893_4073.n4 a_893_4073.n1 0.672
R509 a_893_4073.n5 a_893_4073.n4 0.665
R510 a_2035_4077.t6 a_2035_4077.n2 404.877
R511 a_2035_4077.n1 a_2035_4077.t8 210.902
R512 a_2035_4077.n3 a_2035_4077.t6 136.943
R513 a_2035_4077.n2 a_2035_4077.n1 107.801
R514 a_2035_4077.n1 a_2035_4077.t5 80.333
R515 a_2035_4077.n2 a_2035_4077.t7 80.333
R516 a_2035_4077.n0 a_2035_4077.t4 17.4
R517 a_2035_4077.n0 a_2035_4077.t0 17.4
R518 a_2035_4077.n4 a_2035_4077.t2 15.032
R519 a_2035_4077.t3 a_2035_4077.n5 14.282
R520 a_2035_4077.n5 a_2035_4077.t1 14.282
R521 a_2035_4077.n5 a_2035_4077.n4 1.65
R522 a_2035_4077.n3 a_2035_4077.n0 0.672
R523 a_2035_4077.n4 a_2035_4077.n3 0.665
R524 a_n1077_3564.t0 a_n1077_3564.t1 17.4
R525 carry_out.n0 carry_out.t1 28.57
R526 carry_out.n1 carry_out.t0 28.565
R527 carry_out.n1 carry_out.t2 28.565
R528 carry_out.n0 carry_out.t3 17.638
R529 carry_out.n3 carry_out.n2 2.061
R530 carry_out.n2 carry_out.n1 0.69
R531 carry_out.n2 carry_out.n0 0.6
R532 carry_out carry_out.n3 0.097
R533 carry_out.n3 carry_out 0.004
R534 a_2725_509.t0 a_2725_509.t1 17.4
R535 a_2489_509.t0 a_2489_509.t1 380.209
C0 VDD w_9_1872# 0.92fF
C1 Y VSS 0.19fF
C2 A w_9_1872# 0.60fF
C3 VDD w_1999_4015# 0.66fF
C4 B w_n1459_885# 0.17fF
C5 carry_in w_n1459_885# 0.20fF
C6 B VSS 0.62fF
C7 carry_in VSS 1.49fF
C8 VDD carry_out 1.13fF
C9 B w_n1468_4139# 0.14fF
C10 carry_in w_n1468_4139# 0.00fF
C11 w_n1459_885# w_9_1872# 0.00fF
C12 VSS w_9_1872# 0.29fF
C13 Y carry_in 0.23fF
C14 VSS w_1999_4015# 0.14fF
C15 B carry_in 0.63fF
C16 VSS carry_out 0.27fF
C17 VDD w_857_4011# 0.53fF
C18 Y w_9_1872# 0.15fF
C19 A w_857_4011# 0.01fF
C20 B w_9_1872# 0.43fF
C21 carry_in w_9_1872# 0.39fF
C22 carry_in w_1999_4015# 0.00fF
C23 carry_in carry_out 0.00fF
C24 VSS w_857_4011# 0.15fF
C25 VDD A 1.32fF
C26 VDD w_n1454_2489# 0.37fF
C27 A w_n1454_2489# 0.07fF
C28 w_9_1872# w_1999_4015# 0.01fF
C29 carry_out w_9_1872# 0.02fF
C30 VDD w_n1459_885# 0.32fF
C31 VDD VSS 11.68fF
C32 carry_out w_1999_4015# 0.16fF
C33 A w_n1459_885# 0.19fF
C34 B w_857_4011# 0.00fF
C35 w_n1459_885# w_n1454_2489# 0.02fF
C36 VSS A 1.71fF
C37 VSS w_n1454_2489# 0.16fF
C38 VDD w_n1468_4139# 0.37fF
C39 VDD Y 0.07fF
C40 A w_n1468_4139# 0.06fF
C41 w_n1454_2489# w_n1468_4139# 0.01fF
C42 Y A 0.01fF
C43 VSS w_n1459_885# 0.17fF
C44 B VDD 0.87fF
C45 VDD carry_in 0.63fF
C46 w_1999_4015# w_857_4011# 0.03fF
C47 B A 2.23fF
C48 carry_in A 0.88fF
C49 B w_n1454_2489# 0.29fF
C50 carry_in w_n1454_2489# 0.07fF
C51 carry_out w_857_4011# 0.01fF
C52 VSS w_n1468_4139# 0.09fF
C53 Y a_n659_3505# 0.46fF
C54 carry_in a_n659_3505# 5.72fF
C55 carry_out a_n659_3505# 0.43fF
C56 VSS a_n659_3505# 7.97fF
C57 VDD a_n659_3505# 8.39fF
C58 B a_n659_3505# 3.79fF
C59 A a_n659_3505# 4.31fF
C60 w_n1459_885# a_n659_3505# 1.62fF
C61 w_9_1872# a_n659_3505# 8.86fF
C62 w_n1454_2489# a_n659_3505# 1.62fF
C63 w_n1468_4139# a_n659_3505# 1.65fF
C64 w_1999_4015# a_n659_3505# 2.98fF
C65 w_857_4011# a_n659_3505# 2.70fF
C66 a_473_1241.t0 a_n659_3505# 0.06fF
C67 a_473_1241.t4 a_n659_3505# 0.06fF
C68 a_473_1241.t3 a_n659_3505# 0.06fF
C69 a_473_1241.n0 a_n659_3505# 0.53fF $ **FLOATING
C70 a_473_1241.t5 a_n659_3505# 0.06fF
C71 a_473_1241.t1 a_n659_3505# 0.06fF
C72 a_473_1241.n1 a_n659_3505# 0.12fF $ **FLOATING
C73 a_473_1241.n2 a_n659_3505# 0.37fF $ **FLOATING
C74 a_473_1241.t6 a_n659_3505# 0.06fF
C75 a_473_1241.t8 a_n659_3505# 0.06fF
C76 a_473_1241.n3 a_n659_3505# 0.45fF $ **FLOATING
C77 a_473_1241.t7 a_n659_3505# 0.12fF
C78 a_473_1241.n4 a_n659_3505# 0.69fF $ **FLOATING
C79 a_473_1241.t10 a_n659_3505# 0.06fF
C80 a_473_1241.t9 a_n659_3505# 0.06fF
C81 a_473_1241.n5 a_n659_3505# 0.45fF $ **FLOATING
C82 a_473_1241.t11 a_n659_3505# 0.12fF
C83 a_473_1241.n6 a_n659_3505# 0.71fF $ **FLOATING
C84 a_473_1241.n7 a_n659_3505# 0.06fF $ **FLOATING
C85 a_473_1241.n8 a_n659_3505# 0.16fF $ **FLOATING
C86 a_473_1241.n9 a_n659_3505# 0.48fF $ **FLOATING
C87 a_473_1241.t2 a_n659_3505# 0.06fF
C88 Y.t5 a_n659_3505# 0.04fF
C89 Y.t4 a_n659_3505# 0.04fF
C90 Y.n0 a_n659_3505# 0.29fF $ **FLOATING
C91 Y.t6 a_n659_3505# 0.04fF
C92 Y.t1 a_n659_3505# 0.04fF
C93 Y.n1 a_n659_3505# 0.29fF $ **FLOATING
C94 Y.t7 a_n659_3505# 0.04fF
C95 Y.t0 a_n659_3505# 0.04fF
C96 Y.n2 a_n659_3505# 0.33fF $ **FLOATING
C97 Y.t3 a_n659_3505# 0.04fF
C98 Y.t2 a_n659_3505# 0.04fF
C99 Y.n3 a_n659_3505# 0.30fF $ **FLOATING
C100 Y.n4 a_n659_3505# 0.14fF $ **FLOATING
C101 Y.n5 a_n659_3505# 0.09fF $ **FLOATING
C102 Y.n6 a_n659_3505# 0.17fF $ **FLOATING
C103 Y.n7 a_n659_3505# 0.21fF $ **FLOATING
C104 Y.n8 a_n659_3505# 0.12fF $ **FLOATING
C105 A.t1 a_n659_3505# 0.05fF
C106 A.t4 a_n659_3505# 0.07fF
C107 A.t13 a_n659_3505# 0.07fF
C108 A.t3 a_n659_3505# 0.09fF
C109 A.n0 a_n659_3505# 0.09fF $ **FLOATING
C110 A.n1 a_n659_3505# 0.09fF $ **FLOATING
C111 A.t12 a_n659_3505# 0.08fF
C112 A.n2 a_n659_3505# 0.08fF $ **FLOATING
C113 A.t8 a_n659_3505# 0.06fF
C114 A.t2 a_n659_3505# 0.04fF
C115 A.t14 a_n659_3505# 0.14fF
C116 A.n3 a_n659_3505# 0.29fF $ **FLOATING
C117 A.n4 a_n659_3505# 0.23fF $ **FLOATING
C118 A.t9 a_n659_3505# 0.03fF
C119 A.t6 a_n659_3505# 0.05fF
C120 A.n5 a_n659_3505# 0.06fF $ **FLOATING
C121 A.t11 a_n659_3505# 0.10fF
C122 A.t0 a_n659_3505# 0.11fF
C123 A.n6 a_n659_3505# 2.93fF $ **FLOATING
C124 A.t5 a_n659_3505# 0.03fF
C125 A.t15 a_n659_3505# 0.05fF
C126 A.n7 a_n659_3505# 0.06fF $ **FLOATING
C127 A.t10 a_n659_3505# 0.10fF
C128 A.t7 a_n659_3505# 0.11fF
C129 A.n8 a_n659_3505# 0.81fF $ **FLOATING
C130 a_2371_1241.t0 a_n659_3505# 0.06fF
C131 a_2371_1241.n0 a_n659_3505# 0.45fF $ **FLOATING
C132 a_2371_1241.n1 a_n659_3505# 0.37fF $ **FLOATING
C133 a_2371_1241.n2 a_n659_3505# 0.12fF $ **FLOATING
C134 a_2371_1241.t6 a_n659_3505# 0.06fF
C135 a_2371_1241.t11 a_n659_3505# 0.06fF
C136 a_2371_1241.n3 a_n659_3505# 0.53fF $ **FLOATING
C137 a_2371_1241.t10 a_n659_3505# 0.06fF
C138 a_2371_1241.t9 a_n659_3505# 0.06fF
C139 a_2371_1241.n4 a_n659_3505# 0.16fF $ **FLOATING
C140 a_2371_1241.n5 a_n659_3505# 0.48fF $ **FLOATING
C141 a_2371_1241.t7 a_n659_3505# 0.06fF
C142 a_2371_1241.t8 a_n659_3505# 0.06fF
C143 a_2371_1241.n6 a_n659_3505# 0.06fF $ **FLOATING
C144 a_2371_1241.t2 a_n659_3505# 0.12fF
C145 a_2371_1241.n7 a_n659_3505# 0.45fF $ **FLOATING
C146 a_2371_1241.t3 a_n659_3505# 0.06fF
C147 a_2371_1241.t5 a_n659_3505# 0.06fF
C148 a_2371_1241.n8 a_n659_3505# 0.69fF $ **FLOATING
C149 a_2371_1241.t4 a_n659_3505# 0.12fF
C150 a_2371_1241.n9 a_n659_3505# 0.71fF $ **FLOATING
C151 a_2371_1241.t1 a_n659_3505# 0.06fF
C152 VSS.t7 a_n659_3505# 0.01fF
C153 VSS.t4 a_n659_3505# 0.01fF
C154 VSS.t10 a_n659_3505# 0.01fF
C155 VSS.t3 a_n659_3505# 0.01fF
C156 VSS.n0 a_n659_3505# 0.04fF $ **FLOATING
C157 VSS.n1 a_n659_3505# 0.05fF $ **FLOATING
C158 VSS.n2 a_n659_3505# 0.05fF $ **FLOATING
C159 VSS.t2 a_n659_3505# 0.00fF
C160 VSS.t14 a_n659_3505# 0.00fF
C161 VSS.t18 a_n659_3505# 0.00fF
C162 VSS.n3 a_n659_3505# 0.02fF $ **FLOATING
C163 VSS.n4 a_n659_3505# 0.04fF $ **FLOATING
C164 VSS.t19 a_n659_3505# 0.00fF
C165 VSS.t0 a_n659_3505# 0.00fF
C166 VSS.t1 a_n659_3505# 0.00fF
C167 VSS.n5 a_n659_3505# 0.02fF $ **FLOATING
C168 VSS.n6 a_n659_3505# 0.04fF $ **FLOATING
C169 VSS.t16 a_n659_3505# 0.00fF
C170 VSS.t5 a_n659_3505# 0.01fF
C171 VSS.n7 a_n659_3505# 0.21fF $ **FLOATING
C172 VSS.n8 a_n659_3505# 4.80fF $ **FLOATING
C173 VSS.t15 a_n659_3505# 0.00fF
C174 VSS.t6 a_n659_3505# 0.01fF
C175 VSS.n9 a_n659_3505# 0.08fF $ **FLOATING
C176 VSS.n10 a_n659_3505# 5.87fF $ **FLOATING
C177 VSS.t17 a_n659_3505# 0.00fF
C178 VSS.t13 a_n659_3505# 0.01fF
C179 VSS.n11 a_n659_3505# 0.08fF $ **FLOATING
C180 VSS.t9 a_n659_3505# 0.01fF
C181 VSS.t11 a_n659_3505# 0.01fF
C182 VSS.t8 a_n659_3505# 0.01fF
C183 VSS.t12 a_n659_3505# 0.01fF
C184 VSS.n12 a_n659_3505# 0.04fF $ **FLOATING
C185 VSS.n13 a_n659_3505# 0.05fF $ **FLOATING
C186 VSS.n14 a_n659_3505# 0.05fF $ **FLOATING
C187 VSS.n15 a_n659_3505# 5.06fF $ **FLOATING
C188 B.t6 a_n659_3505# 0.04fF
C189 B.t11 a_n659_3505# 0.06fF
C190 B.n0 a_n659_3505# 0.07fF $ **FLOATING
C191 B.t14 a_n659_3505# 0.12fF
C192 B.t4 a_n659_3505# 0.12fF
C193 B.t2 a_n659_3505# 0.04fF
C194 B.t13 a_n659_3505# 0.08fF
C195 B.t9 a_n659_3505# 0.11fF
C196 B.n1 a_n659_3505# 0.14fF $ **FLOATING
C197 B.t5 a_n659_3505# 0.13fF
C198 B.n2 a_n659_3505# 0.10fF $ **FLOATING
C199 B.t7 a_n659_3505# 0.04fF
C200 B.t12 a_n659_3505# 0.06fF
C201 B.n3 a_n659_3505# 0.05fF $ **FLOATING
C202 B.n4 a_n659_3505# 0.03fF $ **FLOATING
C203 B.t3 a_n659_3505# 0.04fF
C204 B.t0 a_n659_3505# 0.16fF
C205 B.n5 a_n659_3505# 0.33fF $ **FLOATING
C206 B.n6 a_n659_3505# 0.38fF $ **FLOATING
C207 B.n7 a_n659_3505# 0.38fF $ **FLOATING
C208 B.t8 a_n659_3505# 0.04fF
C209 B.t1 a_n659_3505# 0.06fF
C210 B.n8 a_n659_3505# 0.07fF $ **FLOATING
C211 B.t15 a_n659_3505# 0.12fF
C212 B.t10 a_n659_3505# 0.13fF
C213 B.n9 a_n659_3505# 1.84fF $ **FLOATING
C214 a_591_1241.t0 a_n659_3505# 0.02fF
C215 a_591_1241.n0 a_n659_3505# 0.16fF $ **FLOATING
C216 a_591_1241.n1 a_n659_3505# 0.23fF $ **FLOATING
C217 a_591_1241.t8 a_n659_3505# 0.05fF
C218 a_591_1241.t12 a_n659_3505# 0.10fF
C219 a_591_1241.t14 a_n659_3505# 0.08fF
C220 a_591_1241.t9 a_n659_3505# 0.06fF
C221 a_591_1241.n2 a_n659_3505# 0.11fF $ **FLOATING
C222 a_591_1241.t11 a_n659_3505# 0.03fF
C223 a_591_1241.n3 a_n659_3505# 0.08fF $ **FLOATING
C224 a_591_1241.t13 a_n659_3505# 0.03fF
C225 a_591_1241.n4 a_n659_3505# 0.04fF $ **FLOATING
C226 a_591_1241.n5 a_n659_3505# 0.09fF $ **FLOATING
C227 a_591_1241.t10 a_n659_3505# 0.03fF
C228 a_591_1241.n6 a_n659_3505# 0.18fF $ **FLOATING
C229 a_591_1241.t15 a_n659_3505# 0.12fF
C230 a_591_1241.n7 a_n659_3505# 0.16fF $ **FLOATING
C231 a_591_1241.t4 a_n659_3505# 0.02fF
C232 a_591_1241.t6 a_n659_3505# 0.02fF
C233 a_591_1241.n8 a_n659_3505# 0.05fF $ **FLOATING
C234 a_591_1241.n9 a_n659_3505# 0.16fF $ **FLOATING
C235 a_591_1241.t2 a_n659_3505# 0.02fF
C236 a_591_1241.t3 a_n659_3505# 0.02fF
C237 a_591_1241.n10 a_n659_3505# 0.18fF $ **FLOATING
C238 a_591_1241.t5 a_n659_3505# 0.02fF
C239 a_591_1241.t1 a_n659_3505# 0.02fF
C240 a_591_1241.n11 a_n659_3505# 0.07fF $ **FLOATING
C241 a_591_1241.n12 a_n659_3505# 0.15fF $ **FLOATING
C242 a_591_1241.t7 a_n659_3505# 0.02fF
C243 carry_in.t12 a_n659_3505# 0.03fF
C244 carry_in.t15 a_n659_3505# 0.04fF
C245 carry_in.n0 a_n659_3505# 0.05fF $ **FLOATING
C246 carry_in.t14 a_n659_3505# 0.08fF
C247 carry_in.t3 a_n659_3505# 0.08fF
C248 carry_in.t6 a_n659_3505# 0.04fF
C249 carry_in.t13 a_n659_3505# 0.06fF
C250 carry_in.t11 a_n659_3505# 0.06fF
C251 carry_in.t5 a_n659_3505# 0.07fF
C252 carry_in.n1 a_n659_3505# 0.07fF $ **FLOATING
C253 carry_in.n2 a_n659_3505# 0.07fF $ **FLOATING
C254 carry_in.t4 a_n659_3505# 0.07fF
C255 carry_in.n3 a_n659_3505# 0.06fF $ **FLOATING
C256 carry_in.t0 a_n659_3505# 0.05fF
C257 carry_in.t8 a_n659_3505# 0.03fF
C258 carry_in.t10 a_n659_3505# 0.11fF
C259 carry_in.n4 a_n659_3505# 0.23fF $ **FLOATING
C260 carry_in.n5 a_n659_3505# 0.20fF $ **FLOATING
C261 carry_in.n6 a_n659_3505# 2.14fF $ **FLOATING
C262 carry_in.t2 a_n659_3505# 0.03fF
C263 carry_in.t9 a_n659_3505# 0.04fF
C264 carry_in.n7 a_n659_3505# 0.05fF $ **FLOATING
C265 carry_in.t7 a_n659_3505# 0.08fF
C266 carry_in.t1 a_n659_3505# 0.09fF
C267 carry_in.n8 a_n659_3505# 0.89fF $ **FLOATING
C268 VDD.t0 a_n659_3505# 0.01fF
C269 VDD.t50 a_n659_3505# 0.01fF
C270 VDD.n0 a_n659_3505# 0.10fF $ **FLOATING
C271 VDD.t26 a_n659_3505# 0.01fF
C272 VDD.t28 a_n659_3505# 0.01fF
C273 VDD.t20 a_n659_3505# 0.01fF
C274 VDD.t53 a_n659_3505# 0.01fF
C275 VDD.n1 a_n659_3505# 0.06fF $ **FLOATING
C276 VDD.n2 a_n659_3505# 0.09fF $ **FLOATING
C277 VDD.n3 a_n659_3505# 0.12fF $ **FLOATING
C278 VDD.n4 a_n659_3505# 0.04fF $ **FLOATING
C279 VDD.t9 a_n659_3505# 0.01fF
C280 VDD.t49 a_n659_3505# 0.01fF
C281 VDD.n5 a_n659_3505# 0.10fF $ **FLOATING
C282 VDD.t13 a_n659_3505# 0.01fF
C283 VDD.t54 a_n659_3505# 0.01fF
C284 VDD.t21 a_n659_3505# 0.01fF
C285 VDD.t38 a_n659_3505# 0.01fF
C286 VDD.n6 a_n659_3505# 0.06fF $ **FLOATING
C287 VDD.n7 a_n659_3505# 0.09fF $ **FLOATING
C288 VDD.n8 a_n659_3505# 0.12fF $ **FLOATING
C289 VDD.n9 a_n659_3505# 0.04fF $ **FLOATING
C290 VDD.t6 a_n659_3505# 0.01fF
C291 VDD.t41 a_n659_3505# 0.01fF
C292 VDD.n10 a_n659_3505# 0.05fF $ **FLOATING
C293 VDD.t1 a_n659_3505# 0.01fF
C294 VDD.t52 a_n659_3505# 0.01fF
C295 VDD.t22 a_n659_3505# 0.01fF
C296 VDD.n11 a_n659_3505# 0.05fF $ **FLOATING
C297 VDD.n12 a_n659_3505# 0.09fF $ **FLOATING
C298 VDD.n13 a_n659_3505# 0.05fF $ **FLOATING
C299 VDD.t56 a_n659_3505# 0.01fF
C300 VDD.t57 a_n659_3505# 0.01fF
C301 VDD.n14 a_n659_3505# 0.06fF $ **FLOATING
C302 VDD.t58 a_n659_3505# 0.01fF
C303 VDD.t4 a_n659_3505# 0.01fF
C304 VDD.n15 a_n659_3505# 0.05fF $ **FLOATING
C305 VDD.n16 a_n659_3505# 0.03fF $ **FLOATING
C306 VDD.n17 a_n659_3505# 2.10fF $ **FLOATING
C307 VDD.t46 a_n659_3505# 0.01fF
C308 VDD.t12 a_n659_3505# 0.01fF
C309 VDD.n18 a_n659_3505# 0.05fF $ **FLOATING
C310 VDD.t60 a_n659_3505# 0.01fF
C311 VDD.t23 a_n659_3505# 0.01fF
C312 VDD.t33 a_n659_3505# 0.01fF
C313 VDD.n19 a_n659_3505# 0.05fF $ **FLOATING
C314 VDD.n20 a_n659_3505# 0.09fF $ **FLOATING
C315 VDD.n21 a_n659_3505# 0.05fF $ **FLOATING
C316 VDD.t35 a_n659_3505# 0.01fF
C317 VDD.t36 a_n659_3505# 0.01fF
C318 VDD.n22 a_n659_3505# 0.06fF $ **FLOATING
C319 VDD.t34 a_n659_3505# 0.01fF
C320 VDD.t14 a_n659_3505# 0.01fF
C321 VDD.n23 a_n659_3505# 0.05fF $ **FLOATING
C322 VDD.n24 a_n659_3505# 0.03fF $ **FLOATING
C323 VDD.n25 a_n659_3505# 0.19fF $ **FLOATING
C324 VDD.n26 a_n659_3505# 2.69fF $ **FLOATING
C325 VDD.t29 a_n659_3505# 0.01fF
C326 VDD.t55 a_n659_3505# 0.01fF
C327 VDD.n27 a_n659_3505# 0.09fF $ **FLOATING
C328 VDD.t15 a_n659_3505# 0.01fF
C329 VDD.t45 a_n659_3505# 0.01fF
C330 VDD.n28 a_n659_3505# 0.18fF $ **FLOATING
C331 VDD.t37 a_n659_3505# 0.01fF
C332 VDD.t30 a_n659_3505# 0.01fF
C333 VDD.n29 a_n659_3505# 0.07fF $ **FLOATING
C334 VDD.n30 a_n659_3505# 0.06fF $ **FLOATING
C335 VDD.n31 a_n659_3505# 0.03fF $ **FLOATING
C336 VDD.t51 a_n659_3505# 0.01fF
C337 VDD.t19 a_n659_3505# 0.01fF
C338 VDD.n32 a_n659_3505# 0.09fF $ **FLOATING
C339 VDD.t25 a_n659_3505# 0.01fF
C340 VDD.t17 a_n659_3505# 0.01fF
C341 VDD.n33 a_n659_3505# 0.18fF $ **FLOATING
C342 VDD.t3 a_n659_3505# 0.01fF
C343 VDD.t43 a_n659_3505# 0.01fF
C344 VDD.n34 a_n659_3505# 0.07fF $ **FLOATING
C345 VDD.n35 a_n659_3505# 0.06fF $ **FLOATING
C346 VDD.n36 a_n659_3505# 0.03fF $ **FLOATING
C347 VDD.n37 a_n659_3505# 0.04fF $ **FLOATING
C348 VDD.n38 a_n659_3505# 2.14fF $ **FLOATING
C349 VDD.t40 a_n659_3505# 0.01fF
C350 VDD.t10 a_n659_3505# 0.01fF
C351 VDD.n39 a_n659_3505# 0.09fF $ **FLOATING
C352 VDD.t44 a_n659_3505# 0.01fF
C353 VDD.t2 a_n659_3505# 0.01fF
C354 VDD.n40 a_n659_3505# 0.18fF $ **FLOATING
C355 VDD.t5 a_n659_3505# 0.01fF
C356 VDD.t7 a_n659_3505# 0.01fF
C357 VDD.n41 a_n659_3505# 0.07fF $ **FLOATING
C358 VDD.n42 a_n659_3505# 0.06fF $ **FLOATING
C359 VDD.n43 a_n659_3505# 0.03fF $ **FLOATING
C360 VDD.t48 a_n659_3505# 0.01fF
C361 VDD.t16 a_n659_3505# 0.01fF
C362 VDD.n44 a_n659_3505# 0.09fF $ **FLOATING
C363 VDD.t42 a_n659_3505# 0.01fF
C364 VDD.t8 a_n659_3505# 0.01fF
C365 VDD.n45 a_n659_3505# 0.18fF $ **FLOATING
C366 VDD.t62 a_n659_3505# 0.01fF
C367 VDD.t32 a_n659_3505# 0.01fF
C368 VDD.n46 a_n659_3505# 0.07fF $ **FLOATING
C369 VDD.n47 a_n659_3505# 0.06fF $ **FLOATING
C370 VDD.n48 a_n659_3505# 0.03fF $ **FLOATING
C371 VDD.n49 a_n659_3505# 0.04fF $ **FLOATING
C372 VDD.n50 a_n659_3505# 2.98fF $ **FLOATING
C373 VDD.n51 a_n659_3505# 2.95fF $ **FLOATING
C374 VDD.n52 a_n659_3505# 1.99fF $ **FLOATING
C375 VDD.t31 a_n659_3505# 0.01fF
C376 VDD.t59 a_n659_3505# 0.01fF
C377 VDD.n53 a_n659_3505# 0.06fF $ **FLOATING
C378 VDD.t61 a_n659_3505# 0.01fF
C379 VDD.t39 a_n659_3505# 0.01fF
C380 VDD.n54 a_n659_3505# 0.05fF $ **FLOATING
C381 VDD.n55 a_n659_3505# 0.03fF $ **FLOATING
C382 VDD.t24 a_n659_3505# 0.01fF
C383 VDD.t11 a_n659_3505# 0.01fF
C384 VDD.n56 a_n659_3505# 0.05fF $ **FLOATING
C385 VDD.t18 a_n659_3505# 0.01fF
C386 VDD.t27 a_n659_3505# 0.01fF
C387 VDD.t47 a_n659_3505# 0.01fF
C388 VDD.n57 a_n659_3505# 0.05fF $ **FLOATING
C389 VDD.n58 a_n659_3505# 0.09fF $ **FLOATING
C390 VDD.n59 a_n659_3505# 0.05fF $ **FLOATING
C391 VDD.n60 a_n659_3505# 0.82fF $ **FLOATING
.ends

