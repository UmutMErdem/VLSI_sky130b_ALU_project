magic
tech sky130B
magscale 1 2
timestamp 1735468497
<< error_p >>
rect -29 141 29 147
rect -29 107 -17 141
rect -29 101 29 107
<< nmos >>
rect -30 -131 30 69
<< ndiff >>
rect -88 57 -30 69
rect -88 -119 -76 57
rect -42 -119 -30 57
rect -88 -131 -30 -119
rect 30 57 88 69
rect 30 -119 42 57
rect 76 -119 88 57
rect 30 -131 88 -119
<< ndiffc >>
rect -76 -119 -42 57
rect 42 -119 76 57
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -30 69 30 91
rect -30 -157 30 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -33 107 -17 141
rect 17 107 33 141
rect -76 57 -42 73
rect -76 -135 -42 -119
rect 42 57 76 73
rect 42 -135 76 -119
<< viali >>
rect -17 107 17 141
rect -76 -119 -42 57
rect 42 -119 76 57
<< metal1 >>
rect -29 141 29 147
rect -29 107 -17 141
rect 17 107 29 141
rect -29 101 29 107
rect -82 57 -36 69
rect -82 -119 -76 57
rect -42 -119 -36 57
rect -82 -131 -36 -119
rect 36 57 82 69
rect 36 -119 42 57
rect 76 -119 82 57
rect 36 -131 82 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
