magic
tech sky130B
magscale 1 2
timestamp 1736524681
<< nwell >>
rect 458 726 1372 1504
rect 1626 726 2540 1504
rect 888 136 1372 726
rect 2056 466 2540 726
rect 2794 724 3708 1504
rect 3962 726 4876 1504
rect 5136 728 6050 1506
rect 3224 466 3708 724
rect 2055 418 2540 466
rect 3223 418 3708 466
rect 2055 142 2539 418
rect 3223 142 3707 418
rect 4392 142 4876 726
rect 5566 462 6050 728
rect 6304 726 7218 1506
rect 7472 728 8386 1506
rect 5564 420 6050 462
rect 6734 461 7218 726
rect 7902 461 8386 728
rect 8640 726 9554 1506
rect 9070 462 9554 726
rect 6733 420 7218 461
rect 7901 420 8386 461
rect 9069 420 9554 462
rect 5564 138 6048 420
rect 6733 137 7217 420
rect 7901 137 8385 420
rect 9069 138 9553 420
<< nmos >>
rect 462 202 522 402
rect 580 202 640 402
rect 698 202 758 402
rect 1630 204 1690 404
rect 1748 204 1808 404
rect 1866 204 1926 404
rect 2798 204 2858 404
rect 2916 204 2976 404
rect 3034 204 3094 404
rect 3966 204 4026 404
rect 4084 204 4144 404
rect 4202 204 4262 404
rect 5140 204 5200 404
rect 5258 204 5318 404
rect 5376 204 5436 404
rect 6308 204 6368 404
rect 6426 204 6486 404
rect 6544 204 6604 404
rect 7476 206 7536 406
rect 7594 206 7654 406
rect 7712 206 7772 406
rect 8644 206 8704 406
rect 8762 206 8822 406
rect 8880 206 8940 406
<< pmos >>
rect 552 788 612 1188
rect 670 788 730 1188
rect 788 788 848 1188
rect 906 788 966 1188
rect 1024 788 1084 1188
rect 1142 788 1202 1188
rect 1720 788 1780 1188
rect 1838 788 1898 1188
rect 1956 788 2016 1188
rect 2074 788 2134 1188
rect 2192 788 2252 1188
rect 2310 788 2370 1188
rect 2888 786 2948 1186
rect 3006 786 3066 1186
rect 3124 786 3184 1186
rect 3242 786 3302 1186
rect 3360 786 3420 1186
rect 3478 786 3538 1186
rect 4056 788 4116 1188
rect 4174 788 4234 1188
rect 4292 788 4352 1188
rect 4410 788 4470 1188
rect 4528 788 4588 1188
rect 4646 788 4706 1188
rect 5230 790 5290 1190
rect 5348 790 5408 1190
rect 5466 790 5526 1190
rect 5584 790 5644 1190
rect 5702 790 5762 1190
rect 5820 790 5880 1190
rect 6398 788 6458 1188
rect 6516 788 6576 1188
rect 6634 788 6694 1188
rect 6752 788 6812 1188
rect 6870 788 6930 1188
rect 6988 788 7048 1188
rect 7566 790 7626 1190
rect 7684 790 7744 1190
rect 7802 790 7862 1190
rect 7920 790 7980 1190
rect 8038 790 8098 1190
rect 8156 790 8216 1190
rect 982 198 1042 398
rect 1100 198 1160 398
rect 1218 198 1278 398
rect 2149 204 2209 404
rect 2267 204 2327 404
rect 2385 204 2445 404
rect 3317 204 3377 404
rect 3435 204 3495 404
rect 3553 204 3613 404
rect 4486 204 4546 404
rect 4604 204 4664 404
rect 4722 204 4782 404
rect 5658 200 5718 400
rect 5776 200 5836 400
rect 5894 200 5954 400
rect 8734 788 8794 1188
rect 8852 788 8912 1188
rect 8970 788 9030 1188
rect 9088 788 9148 1188
rect 9206 788 9266 1188
rect 9324 788 9384 1188
rect 6827 199 6887 399
rect 6945 199 7005 399
rect 7063 199 7123 399
rect 7995 199 8055 399
rect 8113 199 8173 399
rect 8231 199 8291 399
rect 9163 200 9223 400
rect 9281 200 9341 400
rect 9399 200 9459 400
<< ndiff >>
rect 404 390 462 402
rect 404 214 416 390
rect 450 214 462 390
rect 404 202 462 214
rect 522 390 580 402
rect 522 214 534 390
rect 568 214 580 390
rect 522 202 580 214
rect 640 390 698 402
rect 640 214 652 390
rect 686 214 698 390
rect 640 202 698 214
rect 758 390 816 402
rect 758 214 770 390
rect 804 214 816 390
rect 758 202 816 214
rect 1572 392 1630 404
rect 1572 216 1584 392
rect 1618 216 1630 392
rect 1572 204 1630 216
rect 1690 392 1748 404
rect 1690 216 1702 392
rect 1736 216 1748 392
rect 1690 204 1748 216
rect 1808 392 1866 404
rect 1808 216 1820 392
rect 1854 216 1866 392
rect 1808 204 1866 216
rect 1926 392 1984 404
rect 1926 216 1938 392
rect 1972 216 1984 392
rect 1926 204 1984 216
rect 2740 392 2798 404
rect 2740 216 2752 392
rect 2786 216 2798 392
rect 2740 204 2798 216
rect 2858 392 2916 404
rect 2858 216 2870 392
rect 2904 216 2916 392
rect 2858 204 2916 216
rect 2976 392 3034 404
rect 2976 216 2988 392
rect 3022 216 3034 392
rect 2976 204 3034 216
rect 3094 392 3152 404
rect 3094 216 3106 392
rect 3140 216 3152 392
rect 3094 204 3152 216
rect 3908 392 3966 404
rect 3908 216 3920 392
rect 3954 216 3966 392
rect 3908 204 3966 216
rect 4026 392 4084 404
rect 4026 216 4038 392
rect 4072 216 4084 392
rect 4026 204 4084 216
rect 4144 392 4202 404
rect 4144 216 4156 392
rect 4190 216 4202 392
rect 4144 204 4202 216
rect 4262 392 4320 404
rect 4262 216 4274 392
rect 4308 216 4320 392
rect 4262 204 4320 216
rect 5082 392 5140 404
rect 5082 216 5094 392
rect 5128 216 5140 392
rect 5082 204 5140 216
rect 5200 392 5258 404
rect 5200 216 5212 392
rect 5246 216 5258 392
rect 5200 204 5258 216
rect 5318 392 5376 404
rect 5318 216 5330 392
rect 5364 216 5376 392
rect 5318 204 5376 216
rect 5436 392 5494 404
rect 5436 216 5448 392
rect 5482 216 5494 392
rect 5436 204 5494 216
rect 6250 392 6308 404
rect 6250 216 6262 392
rect 6296 216 6308 392
rect 6250 204 6308 216
rect 6368 392 6426 404
rect 6368 216 6380 392
rect 6414 216 6426 392
rect 6368 204 6426 216
rect 6486 392 6544 404
rect 6486 216 6498 392
rect 6532 216 6544 392
rect 6486 204 6544 216
rect 6604 392 6662 404
rect 6604 216 6616 392
rect 6650 216 6662 392
rect 6604 204 6662 216
rect 7418 394 7476 406
rect 7418 218 7430 394
rect 7464 218 7476 394
rect 7418 206 7476 218
rect 7536 394 7594 406
rect 7536 218 7548 394
rect 7582 218 7594 394
rect 7536 206 7594 218
rect 7654 394 7712 406
rect 7654 218 7666 394
rect 7700 218 7712 394
rect 7654 206 7712 218
rect 7772 394 7830 406
rect 7772 218 7784 394
rect 7818 218 7830 394
rect 7772 206 7830 218
rect 8586 394 8644 406
rect 8586 218 8598 394
rect 8632 218 8644 394
rect 8586 206 8644 218
rect 8704 394 8762 406
rect 8704 218 8716 394
rect 8750 218 8762 394
rect 8704 206 8762 218
rect 8822 394 8880 406
rect 8822 218 8834 394
rect 8868 218 8880 394
rect 8822 206 8880 218
rect 8940 394 8998 406
rect 8940 218 8952 394
rect 8986 218 8998 394
rect 8940 206 8998 218
<< pdiff >>
rect 494 1176 552 1188
rect 494 800 506 1176
rect 540 800 552 1176
rect 494 788 552 800
rect 612 1176 670 1188
rect 612 800 624 1176
rect 658 800 670 1176
rect 612 788 670 800
rect 730 1176 788 1188
rect 730 800 742 1176
rect 776 800 788 1176
rect 730 788 788 800
rect 848 1176 906 1188
rect 848 800 860 1176
rect 894 800 906 1176
rect 848 788 906 800
rect 966 1176 1024 1188
rect 966 800 978 1176
rect 1012 800 1024 1176
rect 966 788 1024 800
rect 1084 1176 1142 1188
rect 1084 800 1096 1176
rect 1130 800 1142 1176
rect 1084 788 1142 800
rect 1202 1176 1260 1188
rect 1202 800 1214 1176
rect 1248 800 1260 1176
rect 1202 788 1260 800
rect 1662 1176 1720 1188
rect 1662 800 1674 1176
rect 1708 800 1720 1176
rect 1662 788 1720 800
rect 1780 1176 1838 1188
rect 1780 800 1792 1176
rect 1826 800 1838 1176
rect 1780 788 1838 800
rect 1898 1176 1956 1188
rect 1898 800 1910 1176
rect 1944 800 1956 1176
rect 1898 788 1956 800
rect 2016 1176 2074 1188
rect 2016 800 2028 1176
rect 2062 800 2074 1176
rect 2016 788 2074 800
rect 2134 1176 2192 1188
rect 2134 800 2146 1176
rect 2180 800 2192 1176
rect 2134 788 2192 800
rect 2252 1176 2310 1188
rect 2252 800 2264 1176
rect 2298 800 2310 1176
rect 2252 788 2310 800
rect 2370 1176 2428 1188
rect 2370 800 2382 1176
rect 2416 800 2428 1176
rect 2370 788 2428 800
rect 2830 1174 2888 1186
rect 2830 798 2842 1174
rect 2876 798 2888 1174
rect 2830 786 2888 798
rect 2948 1174 3006 1186
rect 2948 798 2960 1174
rect 2994 798 3006 1174
rect 2948 786 3006 798
rect 3066 1174 3124 1186
rect 3066 798 3078 1174
rect 3112 798 3124 1174
rect 3066 786 3124 798
rect 3184 1174 3242 1186
rect 3184 798 3196 1174
rect 3230 798 3242 1174
rect 3184 786 3242 798
rect 3302 1174 3360 1186
rect 3302 798 3314 1174
rect 3348 798 3360 1174
rect 3302 786 3360 798
rect 3420 1174 3478 1186
rect 3420 798 3432 1174
rect 3466 798 3478 1174
rect 3420 786 3478 798
rect 3538 1174 3596 1186
rect 3538 798 3550 1174
rect 3584 798 3596 1174
rect 3538 786 3596 798
rect 3998 1176 4056 1188
rect 3998 800 4010 1176
rect 4044 800 4056 1176
rect 3998 788 4056 800
rect 4116 1176 4174 1188
rect 4116 800 4128 1176
rect 4162 800 4174 1176
rect 4116 788 4174 800
rect 4234 1176 4292 1188
rect 4234 800 4246 1176
rect 4280 800 4292 1176
rect 4234 788 4292 800
rect 4352 1176 4410 1188
rect 4352 800 4364 1176
rect 4398 800 4410 1176
rect 4352 788 4410 800
rect 4470 1176 4528 1188
rect 4470 800 4482 1176
rect 4516 800 4528 1176
rect 4470 788 4528 800
rect 4588 1176 4646 1188
rect 4588 800 4600 1176
rect 4634 800 4646 1176
rect 4588 788 4646 800
rect 4706 1176 4764 1188
rect 4706 800 4718 1176
rect 4752 800 4764 1176
rect 4706 788 4764 800
rect 5172 1178 5230 1190
rect 5172 802 5184 1178
rect 5218 802 5230 1178
rect 5172 790 5230 802
rect 5290 1178 5348 1190
rect 5290 802 5302 1178
rect 5336 802 5348 1178
rect 5290 790 5348 802
rect 5408 1178 5466 1190
rect 5408 802 5420 1178
rect 5454 802 5466 1178
rect 5408 790 5466 802
rect 5526 1178 5584 1190
rect 5526 802 5538 1178
rect 5572 802 5584 1178
rect 5526 790 5584 802
rect 5644 1178 5702 1190
rect 5644 802 5656 1178
rect 5690 802 5702 1178
rect 5644 790 5702 802
rect 5762 1178 5820 1190
rect 5762 802 5774 1178
rect 5808 802 5820 1178
rect 5762 790 5820 802
rect 5880 1178 5938 1190
rect 5880 802 5892 1178
rect 5926 802 5938 1178
rect 5880 790 5938 802
rect 6340 1176 6398 1188
rect 6340 800 6352 1176
rect 6386 800 6398 1176
rect 6340 788 6398 800
rect 6458 1176 6516 1188
rect 6458 800 6470 1176
rect 6504 800 6516 1176
rect 6458 788 6516 800
rect 6576 1176 6634 1188
rect 6576 800 6588 1176
rect 6622 800 6634 1176
rect 6576 788 6634 800
rect 6694 1176 6752 1188
rect 6694 800 6706 1176
rect 6740 800 6752 1176
rect 6694 788 6752 800
rect 6812 1176 6870 1188
rect 6812 800 6824 1176
rect 6858 800 6870 1176
rect 6812 788 6870 800
rect 6930 1176 6988 1188
rect 6930 800 6942 1176
rect 6976 800 6988 1176
rect 6930 788 6988 800
rect 7048 1176 7106 1188
rect 7048 800 7060 1176
rect 7094 800 7106 1176
rect 7048 788 7106 800
rect 7508 1178 7566 1190
rect 7508 802 7520 1178
rect 7554 802 7566 1178
rect 7508 790 7566 802
rect 7626 1178 7684 1190
rect 7626 802 7638 1178
rect 7672 802 7684 1178
rect 7626 790 7684 802
rect 7744 1178 7802 1190
rect 7744 802 7756 1178
rect 7790 802 7802 1178
rect 7744 790 7802 802
rect 7862 1178 7920 1190
rect 7862 802 7874 1178
rect 7908 802 7920 1178
rect 7862 790 7920 802
rect 7980 1178 8038 1190
rect 7980 802 7992 1178
rect 8026 802 8038 1178
rect 7980 790 8038 802
rect 8098 1178 8156 1190
rect 8098 802 8110 1178
rect 8144 802 8156 1178
rect 8098 790 8156 802
rect 8216 1178 8274 1190
rect 8216 802 8228 1178
rect 8262 802 8274 1178
rect 8216 790 8274 802
rect 8676 1176 8734 1188
rect 8676 800 8688 1176
rect 8722 800 8734 1176
rect 924 386 982 398
rect 924 210 936 386
rect 970 210 982 386
rect 924 198 982 210
rect 1042 386 1100 398
rect 1042 210 1054 386
rect 1088 210 1100 386
rect 1042 198 1100 210
rect 1160 386 1218 398
rect 1160 210 1172 386
rect 1206 210 1218 386
rect 1160 198 1218 210
rect 1278 386 1336 398
rect 1278 210 1290 386
rect 1324 210 1336 386
rect 1278 198 1336 210
rect 2091 392 2149 404
rect 2091 216 2103 392
rect 2137 216 2149 392
rect 2091 204 2149 216
rect 2209 392 2267 404
rect 2209 216 2221 392
rect 2255 216 2267 392
rect 2209 204 2267 216
rect 2327 392 2385 404
rect 2327 216 2339 392
rect 2373 216 2385 392
rect 2327 204 2385 216
rect 2445 392 2503 404
rect 2445 216 2457 392
rect 2491 216 2503 392
rect 2445 204 2503 216
rect 3259 392 3317 404
rect 3259 216 3271 392
rect 3305 216 3317 392
rect 3259 204 3317 216
rect 3377 392 3435 404
rect 3377 216 3389 392
rect 3423 216 3435 392
rect 3377 204 3435 216
rect 3495 392 3553 404
rect 3495 216 3507 392
rect 3541 216 3553 392
rect 3495 204 3553 216
rect 3613 392 3671 404
rect 3613 216 3625 392
rect 3659 216 3671 392
rect 3613 204 3671 216
rect 4428 392 4486 404
rect 4428 216 4440 392
rect 4474 216 4486 392
rect 4428 204 4486 216
rect 4546 392 4604 404
rect 4546 216 4558 392
rect 4592 216 4604 392
rect 4546 204 4604 216
rect 4664 392 4722 404
rect 4664 216 4676 392
rect 4710 216 4722 392
rect 4664 204 4722 216
rect 4782 392 4840 404
rect 4782 216 4794 392
rect 4828 216 4840 392
rect 4782 204 4840 216
rect 5600 388 5658 400
rect 5600 212 5612 388
rect 5646 212 5658 388
rect 5600 200 5658 212
rect 5718 388 5776 400
rect 5718 212 5730 388
rect 5764 212 5776 388
rect 5718 200 5776 212
rect 5836 388 5894 400
rect 5836 212 5848 388
rect 5882 212 5894 388
rect 5836 200 5894 212
rect 5954 388 6012 400
rect 5954 212 5966 388
rect 6000 212 6012 388
rect 5954 200 6012 212
rect 8676 788 8734 800
rect 8794 1176 8852 1188
rect 8794 800 8806 1176
rect 8840 800 8852 1176
rect 8794 788 8852 800
rect 8912 1176 8970 1188
rect 8912 800 8924 1176
rect 8958 800 8970 1176
rect 8912 788 8970 800
rect 9030 1176 9088 1188
rect 9030 800 9042 1176
rect 9076 800 9088 1176
rect 9030 788 9088 800
rect 9148 1176 9206 1188
rect 9148 800 9160 1176
rect 9194 800 9206 1176
rect 9148 788 9206 800
rect 9266 1176 9324 1188
rect 9266 800 9278 1176
rect 9312 800 9324 1176
rect 9266 788 9324 800
rect 9384 1176 9442 1188
rect 9384 800 9396 1176
rect 9430 800 9442 1176
rect 9384 788 9442 800
rect 6769 387 6827 399
rect 6769 211 6781 387
rect 6815 211 6827 387
rect 6769 199 6827 211
rect 6887 387 6945 399
rect 6887 211 6899 387
rect 6933 211 6945 387
rect 6887 199 6945 211
rect 7005 387 7063 399
rect 7005 211 7017 387
rect 7051 211 7063 387
rect 7005 199 7063 211
rect 7123 387 7181 399
rect 7123 211 7135 387
rect 7169 211 7181 387
rect 7123 199 7181 211
rect 7937 387 7995 399
rect 7937 211 7949 387
rect 7983 211 7995 387
rect 7937 199 7995 211
rect 8055 387 8113 399
rect 8055 211 8067 387
rect 8101 211 8113 387
rect 8055 199 8113 211
rect 8173 387 8231 399
rect 8173 211 8185 387
rect 8219 211 8231 387
rect 8173 199 8231 211
rect 8291 387 8349 399
rect 8291 211 8303 387
rect 8337 211 8349 387
rect 8291 199 8349 211
rect 9105 388 9163 400
rect 9105 212 9117 388
rect 9151 212 9163 388
rect 9105 200 9163 212
rect 9223 388 9281 400
rect 9223 212 9235 388
rect 9269 212 9281 388
rect 9223 200 9281 212
rect 9341 388 9399 400
rect 9341 212 9353 388
rect 9387 212 9399 388
rect 9341 200 9399 212
rect 9459 388 9517 400
rect 9459 212 9471 388
rect 9505 212 9517 388
rect 9459 200 9517 212
<< ndiffc >>
rect 416 214 450 390
rect 534 214 568 390
rect 652 214 686 390
rect 770 214 804 390
rect 1584 216 1618 392
rect 1702 216 1736 392
rect 1820 216 1854 392
rect 1938 216 1972 392
rect 2752 216 2786 392
rect 2870 216 2904 392
rect 2988 216 3022 392
rect 3106 216 3140 392
rect 3920 216 3954 392
rect 4038 216 4072 392
rect 4156 216 4190 392
rect 4274 216 4308 392
rect 5094 216 5128 392
rect 5212 216 5246 392
rect 5330 216 5364 392
rect 5448 216 5482 392
rect 6262 216 6296 392
rect 6380 216 6414 392
rect 6498 216 6532 392
rect 6616 216 6650 392
rect 7430 218 7464 394
rect 7548 218 7582 394
rect 7666 218 7700 394
rect 7784 218 7818 394
rect 8598 218 8632 394
rect 8716 218 8750 394
rect 8834 218 8868 394
rect 8952 218 8986 394
<< pdiffc >>
rect 506 800 540 1176
rect 624 800 658 1176
rect 742 800 776 1176
rect 860 800 894 1176
rect 978 800 1012 1176
rect 1096 800 1130 1176
rect 1214 800 1248 1176
rect 1674 800 1708 1176
rect 1792 800 1826 1176
rect 1910 800 1944 1176
rect 2028 800 2062 1176
rect 2146 800 2180 1176
rect 2264 800 2298 1176
rect 2382 800 2416 1176
rect 2842 798 2876 1174
rect 2960 798 2994 1174
rect 3078 798 3112 1174
rect 3196 798 3230 1174
rect 3314 798 3348 1174
rect 3432 798 3466 1174
rect 3550 798 3584 1174
rect 4010 800 4044 1176
rect 4128 800 4162 1176
rect 4246 800 4280 1176
rect 4364 800 4398 1176
rect 4482 800 4516 1176
rect 4600 800 4634 1176
rect 4718 800 4752 1176
rect 5184 802 5218 1178
rect 5302 802 5336 1178
rect 5420 802 5454 1178
rect 5538 802 5572 1178
rect 5656 802 5690 1178
rect 5774 802 5808 1178
rect 5892 802 5926 1178
rect 6352 800 6386 1176
rect 6470 800 6504 1176
rect 6588 800 6622 1176
rect 6706 800 6740 1176
rect 6824 800 6858 1176
rect 6942 800 6976 1176
rect 7060 800 7094 1176
rect 7520 802 7554 1178
rect 7638 802 7672 1178
rect 7756 802 7790 1178
rect 7874 802 7908 1178
rect 7992 802 8026 1178
rect 8110 802 8144 1178
rect 8228 802 8262 1178
rect 8688 800 8722 1176
rect 936 210 970 386
rect 1054 210 1088 386
rect 1172 210 1206 386
rect 1290 210 1324 386
rect 2103 216 2137 392
rect 2221 216 2255 392
rect 2339 216 2373 392
rect 2457 216 2491 392
rect 3271 216 3305 392
rect 3389 216 3423 392
rect 3507 216 3541 392
rect 3625 216 3659 392
rect 4440 216 4474 392
rect 4558 216 4592 392
rect 4676 216 4710 392
rect 4794 216 4828 392
rect 5612 212 5646 388
rect 5730 212 5764 388
rect 5848 212 5882 388
rect 5966 212 6000 388
rect 8806 800 8840 1176
rect 8924 800 8958 1176
rect 9042 800 9076 1176
rect 9160 800 9194 1176
rect 9278 800 9312 1176
rect 9396 800 9430 1176
rect 6781 211 6815 387
rect 6899 211 6933 387
rect 7017 211 7051 387
rect 7135 211 7169 387
rect 7949 211 7983 387
rect 8067 211 8101 387
rect 8185 211 8219 387
rect 8303 211 8337 387
rect 9117 212 9151 388
rect 9235 212 9269 388
rect 9353 212 9387 388
rect 9471 212 9505 388
<< psubdiff >>
rect 538 82 734 112
rect 538 16 578 82
rect 696 16 734 82
rect 538 -32 734 16
rect 1706 82 1902 112
rect 1706 16 1746 82
rect 1864 16 1902 82
rect 1706 -32 1902 16
rect 2874 82 3070 112
rect 2874 16 2914 82
rect 3032 16 3070 82
rect 2874 -32 3070 16
rect 4042 82 4238 112
rect 4042 16 4082 82
rect 4200 16 4238 82
rect 4042 -32 4238 16
rect 5216 84 5412 114
rect 5216 18 5256 84
rect 5374 18 5412 84
rect 5216 -30 5412 18
rect 6384 84 6580 114
rect 6384 18 6424 84
rect 6542 18 6580 84
rect 6384 -30 6580 18
rect 7552 84 7748 114
rect 7552 18 7592 84
rect 7710 18 7748 84
rect 7552 -30 7748 18
rect 8720 84 8916 114
rect 8720 18 8760 84
rect 8878 18 8916 84
rect 8720 -30 8916 18
<< nsubdiff >>
rect 978 1426 1244 1464
rect 978 1354 1034 1426
rect 1178 1354 1244 1426
rect 2146 1426 2412 1464
rect 978 1324 1244 1354
rect 2146 1354 2202 1426
rect 2346 1354 2412 1426
rect 3314 1426 3580 1464
rect 2146 1324 2412 1354
rect 3314 1354 3370 1426
rect 3514 1354 3580 1426
rect 4482 1426 4748 1464
rect 3314 1324 3580 1354
rect 4482 1354 4538 1426
rect 4682 1354 4748 1426
rect 5656 1428 5922 1466
rect 4482 1324 4748 1354
rect 5656 1356 5712 1428
rect 5856 1356 5922 1428
rect 6824 1428 7090 1466
rect 5656 1326 5922 1356
rect 6824 1356 6880 1428
rect 7024 1356 7090 1428
rect 7992 1428 8258 1466
rect 6824 1326 7090 1356
rect 7992 1356 8048 1428
rect 8192 1356 8258 1428
rect 9160 1428 9426 1466
rect 7992 1326 8258 1356
rect 9160 1356 9216 1428
rect 9360 1356 9426 1428
rect 9160 1326 9426 1356
<< psubdiffcont >>
rect 578 16 696 82
rect 1746 16 1864 82
rect 2914 16 3032 82
rect 4082 16 4200 82
rect 5256 18 5374 84
rect 6424 18 6542 84
rect 7592 18 7710 84
rect 8760 18 8878 84
<< nsubdiffcont >>
rect 1034 1354 1178 1426
rect 2202 1354 2346 1426
rect 3370 1354 3514 1426
rect 4538 1354 4682 1426
rect 5712 1356 5856 1428
rect 6880 1356 7024 1428
rect 8048 1356 8192 1428
rect 9216 1356 9360 1428
<< poly >>
rect 400 1348 466 1364
rect 400 1314 416 1348
rect 450 1344 466 1348
rect 450 1314 950 1344
rect 1568 1348 1634 1364
rect 400 1301 950 1314
rect 400 1298 466 1301
rect 400 1249 466 1256
rect 906 1249 950 1301
rect 1568 1314 1584 1348
rect 1618 1344 1634 1348
rect 1618 1314 2118 1344
rect 2736 1348 2802 1364
rect 1568 1301 2118 1314
rect 1568 1298 1634 1301
rect 1568 1249 1634 1256
rect 2074 1249 2118 1301
rect 2736 1314 2752 1348
rect 2786 1344 2802 1348
rect 2786 1314 3286 1344
rect 3904 1348 3970 1364
rect 2736 1301 3286 1314
rect 2736 1298 2802 1301
rect 2736 1249 2802 1256
rect 3242 1249 3286 1301
rect 3904 1314 3920 1348
rect 3954 1344 3970 1348
rect 3954 1314 4454 1344
rect 5078 1350 5144 1366
rect 3904 1301 4454 1314
rect 3904 1298 3970 1301
rect 3904 1249 3970 1256
rect 4410 1249 4454 1301
rect 5078 1316 5094 1350
rect 5128 1346 5144 1350
rect 5128 1316 5628 1346
rect 6246 1350 6312 1366
rect 5078 1303 5628 1316
rect 5078 1300 5144 1303
rect 5078 1251 5144 1258
rect 5584 1251 5628 1303
rect 6246 1316 6262 1350
rect 6296 1346 6312 1350
rect 6296 1316 6796 1346
rect 7414 1350 7480 1366
rect 6246 1303 6796 1316
rect 6246 1300 6312 1303
rect 6246 1251 6312 1258
rect 6752 1251 6796 1303
rect 7414 1316 7430 1350
rect 7464 1346 7480 1350
rect 7464 1316 7964 1346
rect 8582 1350 8648 1366
rect 7414 1303 7964 1316
rect 7414 1300 7480 1303
rect 7414 1251 7480 1258
rect 7920 1251 7964 1303
rect 8582 1316 8598 1350
rect 8632 1346 8648 1350
rect 8632 1316 9132 1346
rect 8582 1303 9132 1316
rect 8582 1300 8648 1303
rect 8582 1251 8648 1258
rect 9088 1251 9132 1303
rect 400 1240 848 1249
rect 400 1206 416 1240
rect 450 1208 848 1240
rect 450 1207 612 1208
rect 450 1206 466 1207
rect 400 1190 466 1206
rect 552 1188 612 1207
rect 670 1188 730 1208
rect 788 1188 848 1208
rect 906 1208 1202 1249
rect 906 1188 966 1208
rect 1024 1188 1084 1208
rect 1142 1188 1202 1208
rect 1568 1240 2016 1249
rect 1568 1206 1584 1240
rect 1618 1208 2016 1240
rect 1618 1207 1780 1208
rect 1618 1206 1634 1207
rect 1568 1190 1634 1206
rect 1720 1188 1780 1207
rect 1838 1188 1898 1208
rect 1956 1188 2016 1208
rect 2074 1208 2370 1249
rect 2074 1188 2134 1208
rect 2192 1188 2252 1208
rect 2310 1188 2370 1208
rect 2736 1240 3184 1249
rect 2736 1206 2752 1240
rect 2786 1208 3184 1240
rect 2786 1207 2948 1208
rect 2786 1206 2802 1207
rect 2736 1190 2802 1206
rect 2888 1186 2948 1207
rect 3006 1186 3066 1208
rect 3124 1186 3184 1208
rect 3242 1208 3538 1249
rect 3242 1186 3302 1208
rect 3360 1186 3420 1208
rect 3478 1186 3538 1208
rect 3904 1240 4352 1249
rect 3904 1206 3920 1240
rect 3954 1208 4352 1240
rect 3954 1207 4116 1208
rect 3954 1206 3970 1207
rect 3904 1190 3970 1206
rect 4056 1188 4116 1207
rect 4174 1188 4234 1208
rect 4292 1188 4352 1208
rect 4410 1208 4706 1249
rect 4410 1188 4470 1208
rect 4528 1188 4588 1208
rect 4646 1188 4706 1208
rect 5078 1242 5526 1251
rect 5078 1208 5094 1242
rect 5128 1210 5526 1242
rect 5128 1209 5290 1210
rect 5128 1208 5144 1209
rect 5078 1192 5144 1208
rect 5230 1190 5290 1209
rect 5348 1190 5408 1210
rect 5466 1190 5526 1210
rect 5584 1210 5880 1251
rect 5584 1190 5644 1210
rect 5702 1190 5762 1210
rect 5820 1190 5880 1210
rect 6246 1242 6694 1251
rect 6246 1208 6262 1242
rect 6296 1210 6694 1242
rect 6296 1209 6458 1210
rect 6296 1208 6312 1209
rect 6246 1192 6312 1208
rect 552 770 612 788
rect 552 681 613 770
rect 670 762 730 788
rect 788 762 848 788
rect 462 628 613 681
rect 462 402 522 628
rect 906 586 966 788
rect 1024 762 1084 788
rect 1142 762 1202 788
rect 1720 770 1780 788
rect 1720 681 1781 770
rect 1838 762 1898 788
rect 1956 762 2016 788
rect 580 535 966 586
rect 1630 628 1781 681
rect 580 402 640 535
rect 695 477 761 493
rect 695 443 711 477
rect 745 443 761 477
rect 695 427 761 443
rect 698 402 758 427
rect 982 398 1042 424
rect 1100 398 1160 424
rect 1218 398 1278 424
rect 1630 404 1690 628
rect 2074 586 2134 788
rect 2192 762 2252 788
rect 2310 762 2370 788
rect 6398 1188 6458 1209
rect 6516 1188 6576 1210
rect 6634 1188 6694 1210
rect 6752 1210 7048 1251
rect 6752 1188 6812 1210
rect 6870 1188 6930 1210
rect 6988 1188 7048 1210
rect 7414 1242 7862 1251
rect 7414 1208 7430 1242
rect 7464 1210 7862 1242
rect 7464 1209 7626 1210
rect 7464 1208 7480 1209
rect 7414 1192 7480 1208
rect 7566 1190 7626 1209
rect 7684 1190 7744 1210
rect 7802 1190 7862 1210
rect 7920 1210 8216 1251
rect 7920 1190 7980 1210
rect 8038 1190 8098 1210
rect 8156 1190 8216 1210
rect 8582 1242 9030 1251
rect 8582 1208 8598 1242
rect 8632 1210 9030 1242
rect 8632 1209 8794 1210
rect 8632 1208 8648 1209
rect 8582 1192 8648 1208
rect 2888 770 2948 786
rect 2888 681 2949 770
rect 3006 760 3066 786
rect 3124 760 3184 786
rect 1748 535 2134 586
rect 2798 628 2949 681
rect 1748 404 1808 535
rect 1863 477 1929 493
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 1863 427 1929 443
rect 1866 404 1926 427
rect 2149 404 2209 430
rect 2267 404 2327 430
rect 2385 404 2445 430
rect 2798 404 2858 628
rect 3242 586 3302 786
rect 3360 760 3420 786
rect 3478 760 3538 786
rect 4056 770 4116 788
rect 4056 681 4117 770
rect 4174 762 4234 788
rect 4292 762 4352 788
rect 2916 535 3302 586
rect 3966 628 4117 681
rect 2916 404 2976 535
rect 3031 477 3097 493
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 3031 427 3097 443
rect 3034 404 3094 427
rect 3317 404 3377 430
rect 3435 404 3495 430
rect 3553 404 3613 430
rect 3966 404 4026 628
rect 4410 586 4470 788
rect 4528 762 4588 788
rect 4646 762 4706 788
rect 5230 772 5290 790
rect 5230 683 5291 772
rect 5348 764 5408 790
rect 5466 764 5526 790
rect 4084 535 4470 586
rect 5140 630 5291 683
rect 4084 404 4144 535
rect 4199 477 4265 493
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 4199 427 4265 443
rect 4202 404 4262 427
rect 4486 404 4546 430
rect 4604 404 4664 430
rect 4722 404 4782 430
rect 5140 404 5200 630
rect 5584 588 5644 790
rect 5702 764 5762 790
rect 5820 764 5880 790
rect 8734 1188 8794 1209
rect 8852 1188 8912 1210
rect 8970 1188 9030 1210
rect 9088 1210 9384 1251
rect 9088 1188 9148 1210
rect 9206 1188 9266 1210
rect 9324 1188 9384 1210
rect 6398 772 6458 788
rect 6398 683 6459 772
rect 6516 762 6576 788
rect 6634 762 6694 788
rect 5258 537 5644 588
rect 6308 630 6459 683
rect 5258 404 5318 537
rect 5373 479 5439 495
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 5373 429 5439 445
rect 5376 404 5436 429
rect 462 176 522 202
rect 580 176 640 202
rect 698 172 758 202
rect 5658 400 5718 426
rect 5776 400 5836 426
rect 5894 400 5954 426
rect 6308 404 6368 630
rect 6752 588 6812 788
rect 6870 762 6930 788
rect 6988 762 7048 788
rect 7566 772 7626 790
rect 7566 683 7627 772
rect 7684 764 7744 790
rect 7802 764 7862 790
rect 6426 537 6812 588
rect 7476 630 7627 683
rect 6426 404 6486 537
rect 6541 479 6607 495
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 6541 429 6607 445
rect 6544 404 6604 429
rect 982 172 1042 198
rect 1100 172 1160 198
rect 1218 172 1278 198
rect 1630 178 1690 204
rect 1748 178 1808 204
rect 1866 172 1926 204
rect 2149 172 2209 204
rect 2267 172 2327 204
rect 2385 172 2445 204
rect 2798 178 2858 204
rect 2916 178 2976 204
rect 698 131 1277 172
rect 1866 131 2445 172
rect 3034 172 3094 204
rect 3317 172 3377 204
rect 3435 172 3495 204
rect 3553 172 3613 204
rect 3966 178 4026 204
rect 4084 178 4144 204
rect 3034 131 3613 172
rect 4202 172 4262 204
rect 4486 172 4546 204
rect 4604 172 4664 204
rect 4722 178 4782 204
rect 5140 178 5200 204
rect 5258 178 5318 204
rect 4722 172 4781 178
rect 4202 131 4781 172
rect 5376 174 5436 204
rect 6827 399 6887 425
rect 6945 399 7005 425
rect 7063 399 7123 425
rect 7476 406 7536 630
rect 7920 588 7980 790
rect 8038 764 8098 790
rect 8156 764 8216 790
rect 8734 772 8794 788
rect 8734 683 8795 772
rect 8852 762 8912 788
rect 8970 762 9030 788
rect 7594 537 7980 588
rect 8644 630 8795 683
rect 7594 406 7654 537
rect 7709 479 7775 495
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 7709 429 7775 445
rect 7712 406 7772 429
rect 5658 174 5718 200
rect 5776 174 5836 200
rect 5894 174 5954 200
rect 6308 178 6368 204
rect 6426 178 6486 204
rect 5376 168 5954 174
rect 6544 174 6604 204
rect 7995 399 8055 425
rect 8113 399 8173 425
rect 8231 399 8291 425
rect 8644 406 8704 630
rect 9088 588 9148 788
rect 9206 762 9266 788
rect 9324 762 9384 788
rect 8762 537 9148 588
rect 8762 406 8822 537
rect 8877 479 8943 495
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 8877 429 8943 445
rect 8880 406 8940 429
rect 6827 174 6887 199
rect 6945 174 7005 199
rect 7063 174 7123 199
rect 7476 180 7536 206
rect 7594 180 7654 206
rect 5376 133 5955 168
rect 6544 133 7123 174
rect 7712 174 7772 206
rect 9163 400 9223 426
rect 9281 400 9341 426
rect 9399 400 9459 426
rect 7995 174 8055 199
rect 8113 174 8173 199
rect 8231 174 8291 199
rect 8644 180 8704 206
rect 8762 180 8822 206
rect 7712 133 8291 174
rect 8880 174 8940 206
rect 9163 174 9223 200
rect 9281 174 9341 200
rect 9399 174 9459 200
rect 8880 133 9459 174
<< polycont >>
rect 416 1314 450 1348
rect 1584 1314 1618 1348
rect 2752 1314 2786 1348
rect 3920 1314 3954 1348
rect 5094 1316 5128 1350
rect 6262 1316 6296 1350
rect 7430 1316 7464 1350
rect 8598 1316 8632 1350
rect 416 1206 450 1240
rect 1584 1206 1618 1240
rect 2752 1206 2786 1240
rect 3920 1206 3954 1240
rect 5094 1208 5128 1242
rect 6262 1208 6296 1242
rect 711 443 745 477
rect 7430 1208 7464 1242
rect 8598 1208 8632 1242
rect 1879 443 1913 477
rect 3047 443 3081 477
rect 4215 443 4249 477
rect 5389 445 5423 479
rect 6557 445 6591 479
rect 7725 445 7759 479
rect 8893 445 8927 479
<< locali >>
rect 1002 1426 1206 1438
rect 1002 1354 1034 1426
rect 1178 1354 1206 1426
rect 1002 1352 1064 1354
rect 1144 1352 1206 1354
rect 400 1314 416 1348
rect 450 1314 466 1348
rect 1002 1336 1206 1352
rect 2170 1426 2374 1438
rect 2170 1354 2202 1426
rect 2346 1354 2374 1426
rect 2170 1352 2232 1354
rect 2312 1352 2374 1354
rect 1568 1314 1584 1348
rect 1618 1314 1634 1348
rect 2170 1336 2374 1352
rect 3338 1426 3542 1438
rect 3338 1354 3370 1426
rect 3514 1354 3542 1426
rect 3338 1352 3400 1354
rect 3480 1352 3542 1354
rect 2736 1314 2752 1348
rect 2786 1314 2802 1348
rect 3338 1336 3542 1352
rect 4506 1426 4710 1438
rect 4506 1354 4538 1426
rect 4682 1354 4710 1426
rect 4506 1352 4568 1354
rect 4648 1352 4710 1354
rect 3904 1314 3920 1348
rect 3954 1314 3970 1348
rect 4506 1336 4710 1352
rect 5680 1428 5884 1440
rect 5680 1356 5712 1428
rect 5856 1356 5884 1428
rect 5680 1354 5742 1356
rect 5822 1354 5884 1356
rect 5078 1316 5094 1350
rect 5128 1316 5144 1350
rect 5680 1338 5884 1354
rect 6848 1428 7052 1440
rect 6848 1356 6880 1428
rect 7024 1356 7052 1428
rect 6848 1354 6910 1356
rect 6990 1354 7052 1356
rect 6246 1316 6262 1350
rect 6296 1316 6312 1350
rect 6848 1338 7052 1354
rect 8016 1428 8220 1440
rect 8016 1356 8048 1428
rect 8192 1356 8220 1428
rect 8016 1354 8078 1356
rect 8158 1354 8220 1356
rect 7414 1316 7430 1350
rect 7464 1316 7480 1350
rect 8016 1338 8220 1354
rect 9184 1428 9388 1440
rect 9184 1356 9216 1428
rect 9360 1356 9388 1428
rect 9184 1354 9246 1356
rect 9326 1354 9388 1356
rect 8582 1316 8598 1350
rect 8632 1316 8648 1350
rect 9184 1338 9388 1354
rect 400 1206 416 1240
rect 450 1206 466 1240
rect 1568 1206 1584 1240
rect 1618 1206 1634 1240
rect 2736 1206 2752 1240
rect 2786 1206 2802 1240
rect 3904 1206 3920 1240
rect 3954 1206 3970 1240
rect 5078 1208 5094 1242
rect 5128 1208 5144 1242
rect 6246 1208 6262 1242
rect 6296 1208 6312 1242
rect 7414 1208 7430 1242
rect 7464 1208 7480 1242
rect 8582 1208 8598 1242
rect 8632 1208 8648 1242
rect 506 1176 540 1192
rect 506 784 540 800
rect 624 1176 658 1192
rect 624 784 658 800
rect 742 1176 776 1192
rect 742 784 776 800
rect 860 1176 894 1192
rect 860 784 894 800
rect 978 1176 1012 1192
rect 978 784 1012 800
rect 1096 1176 1130 1192
rect 1096 784 1130 800
rect 1214 1176 1248 1192
rect 1214 784 1248 800
rect 1674 1176 1708 1192
rect 1674 784 1708 800
rect 1792 1176 1826 1192
rect 1792 784 1826 800
rect 1910 1176 1944 1192
rect 1910 784 1944 800
rect 2028 1176 2062 1192
rect 2028 784 2062 800
rect 2146 1176 2180 1192
rect 2146 784 2180 800
rect 2264 1176 2298 1192
rect 2264 784 2298 800
rect 2382 1176 2416 1192
rect 2382 784 2416 800
rect 2842 1174 2876 1190
rect 2842 782 2876 798
rect 2960 1174 2994 1190
rect 2960 782 2994 798
rect 3078 1174 3112 1190
rect 3078 782 3112 798
rect 3196 1174 3230 1190
rect 3196 782 3230 798
rect 3314 1174 3348 1190
rect 3314 782 3348 798
rect 3432 1174 3466 1190
rect 3432 782 3466 798
rect 3550 1174 3584 1190
rect 3550 782 3584 798
rect 4010 1176 4044 1192
rect 4010 784 4044 800
rect 4128 1176 4162 1192
rect 4128 784 4162 800
rect 4246 1176 4280 1192
rect 4246 784 4280 800
rect 4364 1176 4398 1192
rect 4364 784 4398 800
rect 4482 1176 4516 1192
rect 4482 784 4516 800
rect 4600 1176 4634 1192
rect 4600 784 4634 800
rect 4718 1176 4752 1192
rect 4718 784 4752 800
rect 5184 1178 5218 1194
rect 5184 786 5218 802
rect 5302 1178 5336 1194
rect 5302 786 5336 802
rect 5420 1178 5454 1194
rect 5420 786 5454 802
rect 5538 1178 5572 1194
rect 5538 786 5572 802
rect 5656 1178 5690 1194
rect 5656 786 5690 802
rect 5774 1178 5808 1194
rect 5774 786 5808 802
rect 5892 1178 5926 1194
rect 5892 786 5926 802
rect 6352 1176 6386 1192
rect 6352 784 6386 800
rect 6470 1176 6504 1192
rect 6470 784 6504 800
rect 6588 1176 6622 1192
rect 6588 784 6622 800
rect 6706 1176 6740 1192
rect 6706 784 6740 800
rect 6824 1176 6858 1192
rect 6824 784 6858 800
rect 6942 1176 6976 1192
rect 6942 784 6976 800
rect 7060 1176 7094 1192
rect 7060 784 7094 800
rect 7520 1178 7554 1194
rect 7520 786 7554 802
rect 7638 1178 7672 1194
rect 7638 786 7672 802
rect 7756 1178 7790 1194
rect 7756 786 7790 802
rect 7874 1178 7908 1194
rect 7874 786 7908 802
rect 7992 1178 8026 1194
rect 7992 786 8026 802
rect 8110 1178 8144 1194
rect 8110 786 8144 802
rect 8228 1178 8262 1194
rect 8228 786 8262 802
rect 8688 1176 8722 1192
rect 8688 784 8722 800
rect 8806 1176 8840 1192
rect 8806 784 8840 800
rect 8924 1176 8958 1192
rect 8924 784 8958 800
rect 9042 1176 9076 1192
rect 9042 784 9076 800
rect 9160 1176 9194 1192
rect 9160 784 9194 800
rect 9278 1176 9312 1192
rect 9278 784 9312 800
rect 9396 1176 9430 1192
rect 9396 784 9430 800
rect 695 443 711 477
rect 745 443 761 477
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 416 390 450 406
rect 416 198 450 214
rect 534 390 568 406
rect 534 198 568 214
rect 652 390 686 406
rect 652 198 686 214
rect 770 390 804 406
rect 770 198 804 214
rect 936 386 970 402
rect 936 194 970 210
rect 1054 386 1088 402
rect 1054 194 1088 210
rect 1172 386 1206 402
rect 1172 194 1206 210
rect 1290 386 1324 402
rect 1290 194 1324 210
rect 1584 392 1618 408
rect 1584 200 1618 216
rect 1702 392 1736 408
rect 1702 200 1736 216
rect 1820 392 1854 408
rect 1820 200 1854 216
rect 1938 392 1972 408
rect 1938 200 1972 216
rect 2103 392 2137 408
rect 2103 200 2137 216
rect 2221 392 2255 408
rect 2221 200 2255 216
rect 2339 392 2373 408
rect 2339 200 2373 216
rect 2457 392 2491 408
rect 2457 200 2491 216
rect 2752 392 2786 408
rect 2752 200 2786 216
rect 2870 392 2904 408
rect 2870 200 2904 216
rect 2988 392 3022 408
rect 2988 200 3022 216
rect 3106 392 3140 408
rect 3106 200 3140 216
rect 3271 392 3305 408
rect 3271 200 3305 216
rect 3389 392 3423 408
rect 3389 200 3423 216
rect 3507 392 3541 408
rect 3507 200 3541 216
rect 3625 392 3659 408
rect 3625 200 3659 216
rect 3920 392 3954 408
rect 3920 200 3954 216
rect 4038 392 4072 408
rect 4038 200 4072 216
rect 4156 392 4190 408
rect 4156 200 4190 216
rect 4274 392 4308 408
rect 4274 200 4308 216
rect 4440 392 4474 408
rect 4440 200 4474 216
rect 4558 392 4592 408
rect 4558 200 4592 216
rect 4676 392 4710 408
rect 4676 200 4710 216
rect 4794 392 4828 408
rect 4794 200 4828 216
rect 5094 392 5128 408
rect 5094 200 5128 216
rect 5212 392 5246 408
rect 5212 200 5246 216
rect 5330 392 5364 408
rect 5330 200 5364 216
rect 5448 392 5482 408
rect 5448 200 5482 216
rect 5612 388 5646 404
rect 5612 196 5646 212
rect 5730 388 5764 404
rect 5730 196 5764 212
rect 5848 388 5882 404
rect 5848 196 5882 212
rect 5966 388 6000 404
rect 5966 196 6000 212
rect 6262 392 6296 408
rect 6262 200 6296 216
rect 6380 392 6414 408
rect 6380 200 6414 216
rect 6498 392 6532 408
rect 6498 200 6532 216
rect 6616 392 6650 408
rect 6616 200 6650 216
rect 6781 387 6815 403
rect 6781 195 6815 211
rect 6899 387 6933 403
rect 6899 195 6933 211
rect 7017 387 7051 403
rect 7017 195 7051 211
rect 7135 387 7169 403
rect 7135 195 7169 211
rect 7430 394 7464 410
rect 7430 202 7464 218
rect 7548 394 7582 410
rect 7548 202 7582 218
rect 7666 394 7700 410
rect 7666 202 7700 218
rect 7784 394 7818 410
rect 7784 202 7818 218
rect 7949 387 7983 403
rect 7949 195 7983 211
rect 8067 387 8101 403
rect 8067 195 8101 211
rect 8185 387 8219 403
rect 8185 195 8219 211
rect 8303 387 8337 403
rect 8303 195 8337 211
rect 8598 394 8632 410
rect 8598 202 8632 218
rect 8716 394 8750 410
rect 8716 202 8750 218
rect 8834 394 8868 410
rect 8834 202 8868 218
rect 8952 394 8986 410
rect 8952 202 8986 218
rect 9117 388 9151 404
rect 9117 196 9151 212
rect 9235 388 9269 404
rect 9235 196 9269 212
rect 9353 388 9387 404
rect 9353 196 9387 212
rect 9471 388 9505 404
rect 9471 196 9505 212
rect 560 86 702 98
rect 560 82 600 86
rect 666 82 702 86
rect 560 16 578 82
rect 696 16 702 82
rect 560 -10 702 16
rect 1728 86 1870 98
rect 1728 82 1768 86
rect 1834 82 1870 86
rect 1728 16 1746 82
rect 1864 16 1870 82
rect 1728 -10 1870 16
rect 2896 86 3038 98
rect 2896 82 2936 86
rect 3002 82 3038 86
rect 2896 16 2914 82
rect 3032 16 3038 82
rect 2896 -10 3038 16
rect 4064 86 4206 98
rect 4064 82 4104 86
rect 4170 82 4206 86
rect 4064 16 4082 82
rect 4200 16 4206 82
rect 4064 -10 4206 16
rect 5238 88 5380 100
rect 5238 84 5278 88
rect 5344 84 5380 88
rect 5238 18 5256 84
rect 5374 18 5380 84
rect 5238 -8 5380 18
rect 6406 88 6548 100
rect 6406 84 6446 88
rect 6512 84 6548 88
rect 6406 18 6424 84
rect 6542 18 6548 84
rect 6406 -8 6548 18
rect 7574 88 7716 100
rect 7574 84 7614 88
rect 7680 84 7716 88
rect 7574 18 7592 84
rect 7710 18 7716 84
rect 7574 -8 7716 18
rect 8742 88 8884 100
rect 8742 84 8782 88
rect 8848 84 8884 88
rect 8742 18 8760 84
rect 8878 18 8884 84
rect 8742 -8 8884 18
<< viali >>
rect 1064 1354 1144 1424
rect 1064 1352 1144 1354
rect 416 1314 450 1348
rect 2232 1354 2312 1424
rect 2232 1352 2312 1354
rect 1584 1314 1618 1348
rect 3400 1354 3480 1424
rect 3400 1352 3480 1354
rect 2752 1314 2786 1348
rect 4568 1354 4648 1424
rect 4568 1352 4648 1354
rect 3920 1314 3954 1348
rect 5742 1356 5822 1426
rect 5742 1354 5822 1356
rect 5094 1316 5128 1350
rect 6910 1356 6990 1426
rect 6910 1354 6990 1356
rect 6262 1316 6296 1350
rect 8078 1356 8158 1426
rect 8078 1354 8158 1356
rect 7430 1316 7464 1350
rect 9246 1356 9326 1426
rect 9246 1354 9326 1356
rect 8598 1316 8632 1350
rect 416 1206 450 1240
rect 1584 1206 1618 1240
rect 2752 1206 2786 1240
rect 3920 1206 3954 1240
rect 5094 1208 5128 1242
rect 6262 1208 6296 1242
rect 7430 1208 7464 1242
rect 8598 1208 8632 1242
rect 506 800 540 1176
rect 624 800 658 1176
rect 742 800 776 1176
rect 860 800 894 1176
rect 978 800 1012 1176
rect 1096 800 1130 1176
rect 1214 800 1248 1176
rect 1674 800 1708 1176
rect 1792 800 1826 1176
rect 1910 800 1944 1176
rect 2028 800 2062 1176
rect 2146 800 2180 1176
rect 2264 800 2298 1176
rect 2382 800 2416 1176
rect 2842 798 2876 1174
rect 2960 798 2994 1174
rect 3078 798 3112 1174
rect 3196 798 3230 1174
rect 3314 798 3348 1174
rect 3432 798 3466 1174
rect 3550 798 3584 1174
rect 4010 800 4044 1176
rect 4128 800 4162 1176
rect 4246 800 4280 1176
rect 4364 800 4398 1176
rect 4482 800 4516 1176
rect 4600 800 4634 1176
rect 4718 800 4752 1176
rect 5184 802 5218 1178
rect 5302 802 5336 1178
rect 5420 802 5454 1178
rect 5538 802 5572 1178
rect 5656 802 5690 1178
rect 5774 802 5808 1178
rect 5892 802 5926 1178
rect 6352 800 6386 1176
rect 6470 800 6504 1176
rect 6588 800 6622 1176
rect 6706 800 6740 1176
rect 6824 800 6858 1176
rect 6942 800 6976 1176
rect 7060 800 7094 1176
rect 7520 802 7554 1178
rect 7638 802 7672 1178
rect 7756 802 7790 1178
rect 7874 802 7908 1178
rect 7992 802 8026 1178
rect 8110 802 8144 1178
rect 8228 802 8262 1178
rect 8688 800 8722 1176
rect 8806 800 8840 1176
rect 8924 800 8958 1176
rect 9042 800 9076 1176
rect 9160 800 9194 1176
rect 9278 800 9312 1176
rect 9396 800 9430 1176
rect 711 443 745 477
rect 1879 443 1913 477
rect 3047 443 3081 477
rect 4215 443 4249 477
rect 5389 445 5423 479
rect 6557 445 6591 479
rect 7725 445 7759 479
rect 8893 445 8927 479
rect 416 214 450 390
rect 534 214 568 390
rect 652 214 686 390
rect 770 214 804 390
rect 936 210 970 386
rect 1054 210 1088 386
rect 1172 210 1206 386
rect 1290 210 1324 386
rect 1584 216 1618 392
rect 1702 216 1736 392
rect 1820 216 1854 392
rect 1938 216 1972 392
rect 2103 216 2137 392
rect 2221 216 2255 392
rect 2339 216 2373 392
rect 2457 216 2491 392
rect 2752 216 2786 392
rect 2870 216 2904 392
rect 2988 216 3022 392
rect 3106 216 3140 392
rect 3271 216 3305 392
rect 3389 216 3423 392
rect 3507 216 3541 392
rect 3625 216 3659 392
rect 3920 216 3954 392
rect 4038 216 4072 392
rect 4156 216 4190 392
rect 4274 216 4308 392
rect 4440 216 4474 392
rect 4558 216 4592 392
rect 4676 216 4710 392
rect 4794 216 4828 392
rect 5094 216 5128 392
rect 5212 216 5246 392
rect 5330 216 5364 392
rect 5448 216 5482 392
rect 5612 212 5646 388
rect 5730 212 5764 388
rect 5848 212 5882 388
rect 5966 212 6000 388
rect 6262 216 6296 392
rect 6380 216 6414 392
rect 6498 216 6532 392
rect 6616 216 6650 392
rect 6781 211 6815 387
rect 6899 211 6933 387
rect 7017 211 7051 387
rect 7135 211 7169 387
rect 7430 218 7464 394
rect 7548 218 7582 394
rect 7666 218 7700 394
rect 7784 218 7818 394
rect 7949 211 7983 387
rect 8067 211 8101 387
rect 8185 211 8219 387
rect 8303 211 8337 387
rect 8598 218 8632 394
rect 8716 218 8750 394
rect 8834 218 8868 394
rect 8952 218 8986 394
rect 9117 212 9151 388
rect 9235 212 9269 388
rect 9353 212 9387 388
rect 9471 212 9505 388
rect 600 82 666 86
rect 600 16 666 82
rect 1768 82 1834 86
rect 1768 16 1834 82
rect 2936 82 3002 86
rect 2936 16 3002 82
rect 4104 82 4170 86
rect 4104 16 4170 82
rect 5278 84 5344 88
rect 5278 18 5344 84
rect 6446 84 6512 88
rect 6446 18 6512 84
rect 7614 84 7680 88
rect 7614 18 7680 84
rect 8782 84 8848 88
rect 8782 18 8848 84
<< metal1 >>
rect 366 1348 466 1450
rect 366 1314 416 1348
rect 450 1314 466 1348
rect 1052 1424 1156 1430
rect 1052 1352 1064 1424
rect 1144 1352 1156 1424
rect 1052 1346 1156 1352
rect 1534 1348 1634 1450
rect 366 1288 466 1314
rect 1087 1290 1122 1346
rect 1534 1314 1584 1348
rect 1618 1314 1634 1348
rect 2220 1424 2324 1430
rect 2220 1352 2232 1424
rect 2312 1352 2324 1424
rect 2220 1346 2324 1352
rect 2702 1348 2802 1450
rect 366 1240 466 1260
rect 366 1206 416 1240
rect 450 1206 466 1240
rect 366 1108 466 1206
rect 624 1249 894 1277
rect 624 1188 658 1249
rect 860 1188 894 1249
rect 978 1249 1248 1290
rect 1534 1288 1634 1314
rect 2255 1290 2290 1346
rect 2702 1314 2752 1348
rect 2786 1314 2802 1348
rect 3388 1424 3492 1430
rect 3388 1352 3400 1424
rect 3480 1352 3492 1424
rect 3388 1346 3492 1352
rect 3870 1348 3970 1450
rect 978 1188 1012 1249
rect 1214 1188 1248 1249
rect 1534 1240 1634 1260
rect 1534 1206 1584 1240
rect 1618 1206 1634 1240
rect 500 1176 546 1188
rect 500 800 506 1176
rect 540 800 546 1176
rect 500 788 546 800
rect 618 1176 664 1188
rect 618 800 624 1176
rect 658 800 664 1176
rect 618 788 664 800
rect 736 1176 782 1188
rect 736 800 742 1176
rect 776 800 782 1176
rect 736 788 782 800
rect 854 1176 900 1188
rect 854 800 860 1176
rect 894 800 900 1176
rect 854 788 900 800
rect 972 1176 1018 1188
rect 972 800 978 1176
rect 1012 800 1018 1176
rect 972 788 1018 800
rect 1090 1176 1136 1188
rect 1090 800 1096 1176
rect 1130 800 1136 1176
rect 1090 788 1136 800
rect 1208 1176 1254 1188
rect 1208 800 1214 1176
rect 1248 800 1254 1176
rect 1534 1108 1634 1206
rect 1792 1249 2062 1277
rect 1792 1188 1826 1249
rect 2028 1188 2062 1249
rect 2146 1249 2416 1290
rect 2702 1288 2802 1314
rect 3423 1290 3458 1346
rect 3870 1314 3920 1348
rect 3954 1314 3970 1348
rect 4556 1424 4660 1430
rect 4556 1352 4568 1424
rect 4648 1352 4660 1424
rect 4556 1346 4660 1352
rect 5044 1350 5144 1452
rect 2146 1188 2180 1249
rect 2382 1188 2416 1249
rect 2702 1240 2802 1260
rect 2702 1206 2752 1240
rect 2786 1206 2802 1240
rect 1668 1176 1714 1188
rect 1208 788 1254 800
rect 1668 800 1674 1176
rect 1708 800 1714 1176
rect 1668 788 1714 800
rect 1786 1176 1832 1188
rect 1786 800 1792 1176
rect 1826 800 1832 1176
rect 1786 788 1832 800
rect 1904 1176 1950 1188
rect 1904 800 1910 1176
rect 1944 800 1950 1176
rect 1904 788 1950 800
rect 2022 1176 2068 1188
rect 2022 800 2028 1176
rect 2062 800 2068 1176
rect 2022 788 2068 800
rect 2140 1176 2186 1188
rect 2140 800 2146 1176
rect 2180 800 2186 1176
rect 2140 788 2186 800
rect 2258 1176 2304 1188
rect 2258 800 2264 1176
rect 2298 800 2304 1176
rect 2258 788 2304 800
rect 2376 1176 2422 1188
rect 2376 800 2382 1176
rect 2416 800 2422 1176
rect 2702 1108 2802 1206
rect 2960 1249 3230 1277
rect 2960 1186 2994 1249
rect 3196 1186 3230 1249
rect 3314 1249 3584 1290
rect 3870 1288 3970 1314
rect 4591 1290 4626 1346
rect 5044 1316 5094 1350
rect 5128 1316 5144 1350
rect 5730 1426 5834 1432
rect 5730 1354 5742 1426
rect 5822 1354 5834 1426
rect 5730 1348 5834 1354
rect 6212 1350 6312 1452
rect 5044 1290 5144 1316
rect 5765 1292 5800 1348
rect 6212 1316 6262 1350
rect 6296 1316 6312 1350
rect 6898 1426 7002 1432
rect 6898 1354 6910 1426
rect 6990 1354 7002 1426
rect 6898 1348 7002 1354
rect 7380 1350 7480 1452
rect 3314 1186 3348 1249
rect 3550 1186 3584 1249
rect 3870 1240 3970 1260
rect 3870 1206 3920 1240
rect 3954 1206 3970 1240
rect 2836 1174 2882 1186
rect 2376 788 2422 800
rect 2836 798 2842 1174
rect 2876 798 2882 1174
rect 506 745 540 788
rect 742 745 776 788
rect 506 717 776 745
rect 860 746 894 788
rect 1096 746 1130 788
rect 860 717 1130 746
rect 506 669 540 717
rect 506 639 569 669
rect 534 547 569 639
rect 1214 604 1248 788
rect 1674 745 1708 788
rect 1910 745 1944 788
rect 1674 717 1944 745
rect 2028 746 2062 788
rect 2264 746 2298 788
rect 2028 717 2298 746
rect 1674 669 1708 717
rect 1674 639 1737 669
rect 534 511 761 547
rect 534 402 569 511
rect 695 477 761 511
rect 695 443 711 477
rect 745 443 761 477
rect 1042 535 1139 586
rect 1214 550 1323 604
rect 1042 468 1099 535
rect 695 437 761 443
rect 936 432 1205 468
rect 410 390 456 402
rect 410 214 416 390
rect 450 214 456 390
rect 410 202 456 214
rect 528 390 574 402
rect 528 214 534 390
rect 568 214 574 390
rect 528 202 574 214
rect 646 390 692 402
rect 646 214 652 390
rect 686 214 692 390
rect 646 202 692 214
rect 764 390 810 402
rect 936 398 969 432
rect 1172 398 1205 432
rect 1289 398 1323 550
rect 1702 547 1737 639
rect 2382 604 2416 788
rect 2836 786 2882 798
rect 2954 1174 3000 1186
rect 2954 798 2960 1174
rect 2994 798 3000 1174
rect 2954 786 3000 798
rect 3072 1174 3118 1186
rect 3072 798 3078 1174
rect 3112 798 3118 1174
rect 3072 786 3118 798
rect 3190 1174 3236 1186
rect 3190 798 3196 1174
rect 3230 798 3236 1174
rect 3190 786 3236 798
rect 3308 1174 3354 1186
rect 3308 798 3314 1174
rect 3348 798 3354 1174
rect 3308 786 3354 798
rect 3426 1174 3472 1186
rect 3426 798 3432 1174
rect 3466 798 3472 1174
rect 3426 786 3472 798
rect 3544 1174 3590 1186
rect 3544 798 3550 1174
rect 3584 798 3590 1174
rect 3870 1108 3970 1206
rect 4128 1249 4398 1277
rect 4128 1188 4162 1249
rect 4364 1188 4398 1249
rect 4482 1249 4752 1290
rect 4482 1188 4516 1249
rect 4718 1188 4752 1249
rect 5044 1242 5144 1262
rect 5044 1208 5094 1242
rect 5128 1208 5144 1242
rect 4004 1176 4050 1188
rect 3544 786 3590 798
rect 4004 800 4010 1176
rect 4044 800 4050 1176
rect 4004 788 4050 800
rect 4122 1176 4168 1188
rect 4122 800 4128 1176
rect 4162 800 4168 1176
rect 4122 788 4168 800
rect 4240 1176 4286 1188
rect 4240 800 4246 1176
rect 4280 800 4286 1176
rect 4240 788 4286 800
rect 4358 1176 4404 1188
rect 4358 800 4364 1176
rect 4398 800 4404 1176
rect 4358 788 4404 800
rect 4476 1176 4522 1188
rect 4476 800 4482 1176
rect 4516 800 4522 1176
rect 4476 788 4522 800
rect 4594 1176 4640 1188
rect 4594 800 4600 1176
rect 4634 800 4640 1176
rect 4594 788 4640 800
rect 4712 1176 4758 1188
rect 4712 800 4718 1176
rect 4752 800 4758 1176
rect 5044 1110 5144 1208
rect 5302 1251 5572 1279
rect 5302 1190 5336 1251
rect 5538 1190 5572 1251
rect 5656 1251 5926 1292
rect 6212 1290 6312 1316
rect 6933 1292 6968 1348
rect 7380 1316 7430 1350
rect 7464 1316 7480 1350
rect 8066 1426 8170 1432
rect 8066 1354 8078 1426
rect 8158 1354 8170 1426
rect 8066 1348 8170 1354
rect 8548 1350 8648 1452
rect 5656 1190 5690 1251
rect 5892 1190 5926 1251
rect 6212 1242 6312 1262
rect 6212 1208 6262 1242
rect 6296 1208 6312 1242
rect 5178 1178 5224 1190
rect 4712 788 4758 800
rect 5178 802 5184 1178
rect 5218 802 5224 1178
rect 5178 790 5224 802
rect 5296 1178 5342 1190
rect 5296 802 5302 1178
rect 5336 802 5342 1178
rect 5296 790 5342 802
rect 5414 1178 5460 1190
rect 5414 802 5420 1178
rect 5454 802 5460 1178
rect 5414 790 5460 802
rect 5532 1178 5578 1190
rect 5532 802 5538 1178
rect 5572 802 5578 1178
rect 5532 790 5578 802
rect 5650 1178 5696 1190
rect 5650 802 5656 1178
rect 5690 802 5696 1178
rect 5650 790 5696 802
rect 5768 1178 5814 1190
rect 5768 802 5774 1178
rect 5808 802 5814 1178
rect 5768 790 5814 802
rect 5886 1178 5932 1190
rect 5886 802 5892 1178
rect 5926 802 5932 1178
rect 6212 1110 6312 1208
rect 6470 1251 6740 1279
rect 6470 1188 6504 1251
rect 6706 1188 6740 1251
rect 6824 1251 7094 1292
rect 7380 1290 7480 1316
rect 8101 1292 8136 1348
rect 8548 1316 8598 1350
rect 8632 1316 8648 1350
rect 9234 1426 9338 1432
rect 9234 1354 9246 1426
rect 9326 1354 9338 1426
rect 9234 1348 9338 1354
rect 6824 1188 6858 1251
rect 7060 1188 7094 1251
rect 7380 1242 7480 1262
rect 7380 1208 7430 1242
rect 7464 1208 7480 1242
rect 6346 1176 6392 1188
rect 5886 790 5932 802
rect 6346 800 6352 1176
rect 6386 800 6392 1176
rect 2842 745 2876 786
rect 3078 745 3112 786
rect 2842 717 3112 745
rect 3196 746 3230 786
rect 3432 746 3466 786
rect 3196 717 3466 746
rect 2842 669 2876 717
rect 2842 639 2905 669
rect 1702 511 1929 547
rect 1702 404 1737 511
rect 1863 477 1929 511
rect 1863 443 1879 477
rect 1913 443 1929 477
rect 2210 535 2307 586
rect 2382 550 2491 604
rect 2210 468 2267 535
rect 1863 437 1929 443
rect 2104 432 2373 468
rect 2104 404 2137 432
rect 2340 404 2373 432
rect 2457 404 2491 550
rect 2870 547 2905 639
rect 3550 604 3584 786
rect 4010 745 4044 788
rect 4246 745 4280 788
rect 4010 717 4280 745
rect 4364 746 4398 788
rect 4600 746 4634 788
rect 4364 717 4634 746
rect 4010 669 4044 717
rect 4010 639 4073 669
rect 2870 511 3097 547
rect 2870 404 2905 511
rect 3031 477 3097 511
rect 3031 443 3047 477
rect 3081 443 3097 477
rect 3378 535 3475 586
rect 3550 550 3659 604
rect 3378 468 3435 535
rect 3031 437 3097 443
rect 3272 432 3541 468
rect 3272 404 3305 432
rect 3508 404 3541 432
rect 3625 404 3659 550
rect 4038 547 4073 639
rect 4718 604 4752 788
rect 5184 747 5218 790
rect 5420 747 5454 790
rect 5184 719 5454 747
rect 5538 748 5572 790
rect 5774 748 5808 790
rect 5538 719 5808 748
rect 5184 671 5218 719
rect 5184 641 5247 671
rect 4038 511 4265 547
rect 4038 404 4073 511
rect 4199 477 4265 511
rect 4199 443 4215 477
rect 4249 443 4265 477
rect 4546 535 4643 586
rect 4718 550 4827 604
rect 4546 468 4603 535
rect 4199 437 4265 443
rect 4440 432 4709 468
rect 4440 404 4473 432
rect 4676 404 4709 432
rect 4793 404 4827 550
rect 5212 549 5247 641
rect 5892 606 5926 790
rect 6346 788 6392 800
rect 6464 1176 6510 1188
rect 6464 800 6470 1176
rect 6504 800 6510 1176
rect 6464 788 6510 800
rect 6582 1176 6628 1188
rect 6582 800 6588 1176
rect 6622 800 6628 1176
rect 6582 788 6628 800
rect 6700 1176 6746 1188
rect 6700 800 6706 1176
rect 6740 800 6746 1176
rect 6700 788 6746 800
rect 6818 1176 6864 1188
rect 6818 800 6824 1176
rect 6858 800 6864 1176
rect 6818 788 6864 800
rect 6936 1176 6982 1188
rect 6936 800 6942 1176
rect 6976 800 6982 1176
rect 6936 788 6982 800
rect 7054 1176 7100 1188
rect 7054 800 7060 1176
rect 7094 800 7100 1176
rect 7380 1110 7480 1208
rect 7638 1251 7908 1279
rect 7638 1190 7672 1251
rect 7874 1190 7908 1251
rect 7992 1251 8262 1292
rect 8548 1290 8648 1316
rect 9269 1292 9304 1348
rect 7992 1190 8026 1251
rect 8228 1190 8262 1251
rect 8548 1242 8648 1262
rect 8548 1208 8598 1242
rect 8632 1208 8648 1242
rect 7514 1178 7560 1190
rect 7054 788 7100 800
rect 7514 802 7520 1178
rect 7554 802 7560 1178
rect 7514 790 7560 802
rect 7632 1178 7678 1190
rect 7632 802 7638 1178
rect 7672 802 7678 1178
rect 7632 790 7678 802
rect 7750 1178 7796 1190
rect 7750 802 7756 1178
rect 7790 802 7796 1178
rect 7750 790 7796 802
rect 7868 1178 7914 1190
rect 7868 802 7874 1178
rect 7908 802 7914 1178
rect 7868 790 7914 802
rect 7986 1178 8032 1190
rect 7986 802 7992 1178
rect 8026 802 8032 1178
rect 7986 790 8032 802
rect 8104 1178 8150 1190
rect 8104 802 8110 1178
rect 8144 802 8150 1178
rect 8104 790 8150 802
rect 8222 1178 8268 1190
rect 8222 802 8228 1178
rect 8262 802 8268 1178
rect 8548 1110 8648 1208
rect 8806 1251 9076 1279
rect 8806 1188 8840 1251
rect 9042 1188 9076 1251
rect 9160 1251 9430 1292
rect 9160 1188 9194 1251
rect 9396 1188 9430 1251
rect 8682 1176 8728 1188
rect 8222 790 8268 802
rect 8682 800 8688 1176
rect 8722 800 8728 1176
rect 6352 747 6386 788
rect 6588 747 6622 788
rect 6352 719 6622 747
rect 6706 748 6740 788
rect 6942 748 6976 788
rect 6706 719 6976 748
rect 6352 671 6386 719
rect 6352 641 6415 671
rect 5212 513 5439 549
rect 5212 404 5247 513
rect 5373 479 5439 513
rect 5373 445 5389 479
rect 5423 445 5439 479
rect 5720 537 5817 588
rect 5892 552 6001 606
rect 5720 470 5777 537
rect 5373 439 5439 445
rect 5614 434 5883 470
rect 764 214 770 390
rect 804 337 810 390
rect 930 386 976 398
rect 930 337 936 386
rect 804 249 936 337
rect 804 214 810 249
rect 764 202 810 214
rect 930 210 936 249
rect 970 210 976 386
rect 416 165 450 202
rect 652 165 686 202
rect 930 198 976 210
rect 1048 386 1094 398
rect 1048 210 1054 386
rect 1088 210 1094 386
rect 1048 198 1094 210
rect 1166 386 1212 398
rect 1166 210 1172 386
rect 1206 210 1212 386
rect 1166 198 1212 210
rect 1284 386 1330 398
rect 1284 210 1290 386
rect 1324 210 1330 386
rect 1284 198 1330 210
rect 1578 392 1624 404
rect 1578 216 1584 392
rect 1618 216 1624 392
rect 1578 204 1624 216
rect 1696 392 1742 404
rect 1696 216 1702 392
rect 1736 216 1742 392
rect 1696 204 1742 216
rect 1814 392 1860 404
rect 1814 216 1820 392
rect 1854 216 1860 392
rect 1814 204 1860 216
rect 1932 392 1978 404
rect 1932 216 1938 392
rect 1972 337 1978 392
rect 2097 392 2143 404
rect 2097 337 2103 392
rect 1972 249 2103 337
rect 1972 216 1978 249
rect 1932 204 1978 216
rect 2097 216 2103 249
rect 2137 216 2143 392
rect 2097 204 2143 216
rect 2215 392 2261 404
rect 2215 216 2221 392
rect 2255 216 2261 392
rect 2215 204 2261 216
rect 2333 392 2379 404
rect 2333 216 2339 392
rect 2373 216 2379 392
rect 2333 204 2379 216
rect 2451 392 2497 404
rect 2451 216 2457 392
rect 2491 216 2497 392
rect 2451 204 2497 216
rect 2746 392 2792 404
rect 2746 216 2752 392
rect 2786 216 2792 392
rect 2746 204 2792 216
rect 2864 392 2910 404
rect 2864 216 2870 392
rect 2904 216 2910 392
rect 2864 204 2910 216
rect 2982 392 3028 404
rect 2982 216 2988 392
rect 3022 216 3028 392
rect 2982 204 3028 216
rect 3100 392 3146 404
rect 3100 216 3106 392
rect 3140 337 3146 392
rect 3265 392 3311 404
rect 3265 337 3271 392
rect 3140 249 3271 337
rect 3140 216 3146 249
rect 3100 204 3146 216
rect 3265 216 3271 249
rect 3305 216 3311 392
rect 3265 204 3311 216
rect 3383 392 3429 404
rect 3383 216 3389 392
rect 3423 216 3429 392
rect 3383 204 3429 216
rect 3501 392 3547 404
rect 3501 216 3507 392
rect 3541 216 3547 392
rect 3501 204 3547 216
rect 3619 392 3665 404
rect 3619 216 3625 392
rect 3659 216 3665 392
rect 3619 204 3665 216
rect 3914 392 3960 404
rect 3914 216 3920 392
rect 3954 216 3960 392
rect 3914 204 3960 216
rect 4032 392 4078 404
rect 4032 216 4038 392
rect 4072 216 4078 392
rect 4032 204 4078 216
rect 4150 392 4196 404
rect 4150 216 4156 392
rect 4190 216 4196 392
rect 4150 204 4196 216
rect 4268 392 4314 404
rect 4268 216 4274 392
rect 4308 337 4314 392
rect 4434 392 4480 404
rect 4434 337 4440 392
rect 4308 249 4440 337
rect 4308 216 4314 249
rect 4268 204 4314 216
rect 4434 216 4440 249
rect 4474 216 4480 392
rect 4434 204 4480 216
rect 4552 392 4598 404
rect 4552 216 4558 392
rect 4592 216 4598 392
rect 4552 204 4598 216
rect 4670 392 4716 404
rect 4670 216 4676 392
rect 4710 216 4716 392
rect 4670 204 4716 216
rect 4788 392 4834 404
rect 4788 216 4794 392
rect 4828 216 4834 392
rect 4788 204 4834 216
rect 5088 392 5134 404
rect 5088 216 5094 392
rect 5128 216 5134 392
rect 5088 204 5134 216
rect 5206 392 5252 404
rect 5206 216 5212 392
rect 5246 216 5252 392
rect 5206 204 5252 216
rect 5324 392 5370 404
rect 5324 216 5330 392
rect 5364 216 5370 392
rect 5324 204 5370 216
rect 5442 392 5488 404
rect 5614 400 5647 434
rect 5850 400 5883 434
rect 5967 400 6001 552
rect 6380 549 6415 641
rect 7060 606 7094 788
rect 7520 747 7554 790
rect 7756 747 7790 790
rect 7520 719 7790 747
rect 7874 748 7908 790
rect 8110 748 8144 790
rect 7874 719 8144 748
rect 7520 671 7554 719
rect 7520 641 7583 671
rect 6380 513 6607 549
rect 6380 404 6415 513
rect 6541 479 6607 513
rect 6541 445 6557 479
rect 6591 445 6607 479
rect 6888 537 6985 588
rect 7060 552 7169 606
rect 6888 470 6945 537
rect 6541 439 6607 445
rect 6782 434 7051 470
rect 5442 216 5448 392
rect 5482 339 5488 392
rect 5606 388 5652 400
rect 5606 339 5612 388
rect 5482 251 5612 339
rect 5482 216 5488 251
rect 5442 204 5488 216
rect 5606 212 5612 251
rect 5646 212 5652 388
rect 416 126 686 165
rect 1053 166 1086 198
rect 1289 166 1322 198
rect 1053 130 1322 166
rect 1584 165 1618 204
rect 1820 165 1854 204
rect 1584 126 1854 165
rect 2221 166 2254 204
rect 2457 166 2490 204
rect 2221 130 2490 166
rect 2752 165 2786 204
rect 2988 165 3022 204
rect 2752 126 3022 165
rect 3389 166 3422 204
rect 3625 166 3658 204
rect 3389 130 3658 166
rect 3920 165 3954 204
rect 4156 165 4190 204
rect 3920 126 4190 165
rect 4557 166 4590 204
rect 4793 166 4826 204
rect 4557 130 4826 166
rect 5094 167 5128 204
rect 5330 167 5364 204
rect 5606 200 5652 212
rect 5724 388 5770 400
rect 5724 212 5730 388
rect 5764 212 5770 388
rect 5724 200 5770 212
rect 5842 388 5888 400
rect 5842 212 5848 388
rect 5882 212 5888 388
rect 5842 200 5888 212
rect 5960 388 6006 400
rect 5960 212 5966 388
rect 6000 212 6006 388
rect 5960 200 6006 212
rect 6256 392 6302 404
rect 6256 216 6262 392
rect 6296 216 6302 392
rect 6256 204 6302 216
rect 6374 392 6420 404
rect 6374 216 6380 392
rect 6414 216 6420 392
rect 6374 204 6420 216
rect 6492 392 6538 404
rect 6492 216 6498 392
rect 6532 216 6538 392
rect 6492 204 6538 216
rect 6610 392 6656 404
rect 6782 399 6815 434
rect 7018 399 7051 434
rect 7135 399 7169 552
rect 7548 549 7583 641
rect 8228 606 8262 790
rect 8682 788 8728 800
rect 8800 1176 8846 1188
rect 8800 800 8806 1176
rect 8840 800 8846 1176
rect 8800 788 8846 800
rect 8918 1176 8964 1188
rect 8918 800 8924 1176
rect 8958 800 8964 1176
rect 8918 788 8964 800
rect 9036 1176 9082 1188
rect 9036 800 9042 1176
rect 9076 800 9082 1176
rect 9036 788 9082 800
rect 9154 1176 9200 1188
rect 9154 800 9160 1176
rect 9194 800 9200 1176
rect 9154 788 9200 800
rect 9272 1176 9318 1188
rect 9272 800 9278 1176
rect 9312 800 9318 1176
rect 9272 788 9318 800
rect 9390 1176 9436 1188
rect 9390 800 9396 1176
rect 9430 800 9436 1176
rect 9390 788 9436 800
rect 8688 747 8722 788
rect 8924 747 8958 788
rect 8688 719 8958 747
rect 9042 748 9076 788
rect 9278 748 9312 788
rect 9042 719 9312 748
rect 8688 671 8722 719
rect 8688 641 8751 671
rect 7548 513 7775 549
rect 7548 406 7583 513
rect 7709 479 7775 513
rect 7709 445 7725 479
rect 7759 445 7775 479
rect 8056 537 8153 588
rect 8228 552 8337 606
rect 8056 470 8113 537
rect 7709 439 7775 445
rect 7950 434 8219 470
rect 6610 216 6616 392
rect 6650 339 6656 392
rect 6775 387 6821 399
rect 6775 339 6781 387
rect 6650 251 6781 339
rect 6650 216 6656 251
rect 6610 204 6656 216
rect 6775 211 6781 251
rect 6815 211 6821 387
rect 5094 128 5364 167
rect 5731 168 5764 200
rect 5967 168 6000 200
rect 5731 132 6000 168
rect 6262 167 6296 204
rect 6498 167 6532 204
rect 6775 199 6821 211
rect 6893 387 6939 399
rect 6893 211 6899 387
rect 6933 211 6939 387
rect 6893 199 6939 211
rect 7011 387 7057 399
rect 7011 211 7017 387
rect 7051 211 7057 387
rect 7011 199 7057 211
rect 7129 387 7175 399
rect 7129 211 7135 387
rect 7169 211 7175 387
rect 7129 199 7175 211
rect 7424 394 7470 406
rect 7424 218 7430 394
rect 7464 218 7470 394
rect 7424 206 7470 218
rect 7542 394 7588 406
rect 7542 218 7548 394
rect 7582 218 7588 394
rect 7542 206 7588 218
rect 7660 394 7706 406
rect 7660 218 7666 394
rect 7700 218 7706 394
rect 7660 206 7706 218
rect 7778 394 7824 406
rect 7950 399 7983 434
rect 8186 399 8219 434
rect 8303 399 8337 552
rect 8716 549 8751 641
rect 9396 606 9430 788
rect 8716 513 8943 549
rect 8716 406 8751 513
rect 8877 479 8943 513
rect 8877 445 8893 479
rect 8927 445 8943 479
rect 9224 537 9321 588
rect 9396 552 9505 606
rect 9224 470 9281 537
rect 8877 439 8943 445
rect 9118 434 9387 470
rect 7778 218 7784 394
rect 7818 339 7824 394
rect 7943 387 7989 399
rect 7943 339 7949 387
rect 7818 251 7949 339
rect 7818 218 7824 251
rect 7778 206 7824 218
rect 7943 211 7949 251
rect 7983 211 7989 387
rect 6262 128 6532 167
rect 6899 168 6932 199
rect 7135 168 7168 199
rect 6899 132 7168 168
rect 7430 167 7464 206
rect 7666 167 7700 206
rect 7943 199 7989 211
rect 8061 387 8107 399
rect 8061 211 8067 387
rect 8101 211 8107 387
rect 8061 199 8107 211
rect 8179 387 8225 399
rect 8179 211 8185 387
rect 8219 211 8225 387
rect 8179 199 8225 211
rect 8297 387 8343 399
rect 8297 211 8303 387
rect 8337 211 8343 387
rect 8297 199 8343 211
rect 8592 394 8638 406
rect 8592 218 8598 394
rect 8632 218 8638 394
rect 8592 206 8638 218
rect 8710 394 8756 406
rect 8710 218 8716 394
rect 8750 218 8756 394
rect 8710 206 8756 218
rect 8828 394 8874 406
rect 8828 218 8834 394
rect 8868 218 8874 394
rect 8828 206 8874 218
rect 8946 394 8992 406
rect 9118 400 9151 434
rect 9354 400 9387 434
rect 9471 400 9505 552
rect 8946 218 8952 394
rect 8986 339 8992 394
rect 9111 388 9157 400
rect 9111 339 9117 388
rect 8986 251 9117 339
rect 8986 218 8992 251
rect 8946 206 8992 218
rect 9111 212 9117 251
rect 9151 212 9157 388
rect 7430 128 7700 167
rect 8067 168 8100 199
rect 8303 168 8336 199
rect 8067 132 8336 168
rect 8598 167 8632 206
rect 8834 167 8868 206
rect 9111 200 9157 212
rect 9229 388 9275 400
rect 9229 212 9235 388
rect 9269 212 9275 388
rect 9229 200 9275 212
rect 9347 388 9393 400
rect 9347 212 9353 388
rect 9387 212 9393 388
rect 9347 200 9393 212
rect 9465 388 9511 400
rect 9465 212 9471 388
rect 9505 212 9511 388
rect 9465 200 9511 212
rect 8598 128 8868 167
rect 9235 168 9268 200
rect 9471 168 9504 200
rect 9235 132 9504 168
rect 616 98 650 126
rect 1784 98 1818 126
rect 2952 98 2986 126
rect 4120 98 4154 126
rect 5294 100 5328 128
rect 6462 100 6496 128
rect 7630 100 7664 128
rect 8798 100 8832 128
rect 594 86 672 98
rect 594 16 600 86
rect 666 16 672 86
rect 594 4 672 16
rect 1762 86 1840 98
rect 1762 16 1768 86
rect 1834 16 1840 86
rect 1762 4 1840 16
rect 2930 86 3008 98
rect 2930 16 2936 86
rect 3002 16 3008 86
rect 2930 4 3008 16
rect 4098 86 4176 98
rect 4098 16 4104 86
rect 4170 16 4176 86
rect 4098 4 4176 16
rect 5272 88 5350 100
rect 5272 18 5278 88
rect 5344 18 5350 88
rect 5272 6 5350 18
rect 6440 88 6518 100
rect 6440 18 6446 88
rect 6512 18 6518 88
rect 6440 6 6518 18
rect 7608 88 7686 100
rect 7608 18 7614 88
rect 7680 18 7686 88
rect 7608 6 7686 18
rect 8776 88 8854 100
rect 8776 18 8782 88
rect 8848 18 8854 88
rect 8776 6 8854 18
<< via1 >>
rect 1078 1353 1130 1405
rect 2246 1353 2298 1405
rect 3414 1353 3466 1405
rect 4582 1353 4634 1405
rect 5756 1355 5808 1407
rect 6924 1355 6976 1407
rect 8092 1355 8144 1407
rect 9260 1355 9312 1407
rect 607 29 659 81
rect 1775 29 1827 81
rect 2943 29 2995 81
rect 4111 29 4163 81
rect 5285 31 5337 83
rect 6453 31 6505 83
rect 7621 31 7673 83
rect 8789 31 8841 83
<< metal2 >>
rect 1056 1426 1146 1436
rect 1056 1325 1146 1335
rect 2224 1426 2314 1436
rect 2224 1325 2314 1335
rect 3392 1426 3482 1436
rect 3392 1325 3482 1335
rect 4560 1426 4650 1436
rect 4560 1325 4650 1335
rect 5734 1428 5824 1438
rect 5734 1327 5824 1337
rect 6902 1428 6992 1438
rect 6902 1327 6992 1337
rect 8070 1428 8160 1438
rect 8070 1327 8160 1337
rect 9238 1428 9328 1438
rect 9238 1327 9328 1337
rect 591 99 681 109
rect 591 -2 681 8
rect 1759 99 1849 109
rect 1759 -2 1849 8
rect 2927 99 3017 109
rect 2927 -2 3017 8
rect 4095 99 4185 109
rect 4095 -2 4185 8
rect 5269 101 5359 111
rect 5269 0 5359 10
rect 6437 101 6527 111
rect 6437 0 6527 10
rect 7605 101 7695 111
rect 7605 0 7695 10
rect 8773 101 8863 111
rect 8773 0 8863 10
<< via2 >>
rect 1056 1405 1146 1426
rect 1056 1353 1078 1405
rect 1078 1353 1130 1405
rect 1130 1353 1146 1405
rect 1056 1335 1146 1353
rect 2224 1405 2314 1426
rect 2224 1353 2246 1405
rect 2246 1353 2298 1405
rect 2298 1353 2314 1405
rect 2224 1335 2314 1353
rect 3392 1405 3482 1426
rect 3392 1353 3414 1405
rect 3414 1353 3466 1405
rect 3466 1353 3482 1405
rect 3392 1335 3482 1353
rect 4560 1405 4650 1426
rect 4560 1353 4582 1405
rect 4582 1353 4634 1405
rect 4634 1353 4650 1405
rect 4560 1335 4650 1353
rect 5734 1407 5824 1428
rect 5734 1355 5756 1407
rect 5756 1355 5808 1407
rect 5808 1355 5824 1407
rect 5734 1337 5824 1355
rect 6902 1407 6992 1428
rect 6902 1355 6924 1407
rect 6924 1355 6976 1407
rect 6976 1355 6992 1407
rect 6902 1337 6992 1355
rect 8070 1407 8160 1428
rect 8070 1355 8092 1407
rect 8092 1355 8144 1407
rect 8144 1355 8160 1407
rect 8070 1337 8160 1355
rect 9238 1407 9328 1428
rect 9238 1355 9260 1407
rect 9260 1355 9312 1407
rect 9312 1355 9328 1407
rect 9238 1337 9328 1355
rect 591 81 681 99
rect 591 29 607 81
rect 607 29 659 81
rect 659 29 681 81
rect 591 8 681 29
rect 1759 81 1849 99
rect 1759 29 1775 81
rect 1775 29 1827 81
rect 1827 29 1849 81
rect 1759 8 1849 29
rect 2927 81 3017 99
rect 2927 29 2943 81
rect 2943 29 2995 81
rect 2995 29 3017 81
rect 2927 8 3017 29
rect 4095 81 4185 99
rect 4095 29 4111 81
rect 4111 29 4163 81
rect 4163 29 4185 81
rect 4095 8 4185 29
rect 5269 83 5359 101
rect 5269 31 5285 83
rect 5285 31 5337 83
rect 5337 31 5359 83
rect 5269 10 5359 31
rect 6437 83 6527 101
rect 6437 31 6453 83
rect 6453 31 6505 83
rect 6505 31 6527 83
rect 6437 10 6527 31
rect 7605 83 7695 101
rect 7605 31 7621 83
rect 7621 31 7673 83
rect 7673 31 7695 83
rect 7605 10 7695 31
rect 8773 83 8863 101
rect 8773 31 8789 83
rect 8789 31 8841 83
rect 8841 31 8863 83
rect 8773 10 8863 31
<< metal3 >>
rect 1028 1320 1038 1440
rect 1160 1320 1170 1440
rect 2196 1426 2338 1440
rect 2196 1335 2224 1426
rect 2314 1335 2338 1426
rect 2196 1320 2338 1335
rect 3364 1426 3506 1440
rect 3364 1335 3392 1426
rect 3482 1335 3506 1426
rect 3364 1320 3506 1335
rect 4532 1426 4674 1440
rect 4532 1335 4560 1426
rect 4650 1335 4674 1426
rect 4532 1320 4674 1335
rect 5706 1428 5848 1442
rect 5706 1337 5734 1428
rect 5824 1337 5848 1428
rect 5706 1322 5848 1337
rect 6874 1428 7016 1442
rect 6874 1337 6902 1428
rect 6992 1337 7016 1428
rect 6874 1322 7016 1337
rect 8042 1428 8184 1442
rect 8042 1337 8070 1428
rect 8160 1337 8184 1428
rect 8042 1322 8184 1337
rect 9210 1428 9352 1442
rect 9210 1337 9238 1428
rect 9328 1337 9352 1428
rect 9210 1322 9352 1337
rect 571 -2 581 109
rect 691 -2 701 109
rect 1739 -2 1749 109
rect 1859 -2 1869 109
rect 2907 -2 2917 109
rect 3027 -2 3037 109
rect 4075 -2 4085 109
rect 4195 -2 4205 109
rect 5249 0 5259 111
rect 5369 0 5379 111
rect 6417 0 6427 111
rect 6537 0 6547 111
rect 7585 0 7595 111
rect 7705 0 7715 111
rect 8753 0 8763 111
rect 8873 0 8883 111
<< via3 >>
rect 1038 1426 1160 1440
rect 1038 1335 1056 1426
rect 1056 1335 1146 1426
rect 1146 1335 1160 1426
rect 1038 1320 1160 1335
rect 2240 1348 2304 1412
rect 3408 1348 3472 1412
rect 4578 1350 4642 1414
rect 5750 1350 5814 1414
rect 6918 1348 6982 1412
rect 8086 1350 8150 1414
rect 9254 1350 9318 1414
rect 581 99 691 109
rect 581 8 591 99
rect 591 8 681 99
rect 681 8 691 99
rect 581 -2 691 8
rect 1749 99 1859 109
rect 1749 8 1759 99
rect 1759 8 1849 99
rect 1849 8 1859 99
rect 1749 -2 1859 8
rect 2917 99 3027 109
rect 2917 8 2927 99
rect 2927 8 3017 99
rect 3017 8 3027 99
rect 2917 -2 3027 8
rect 4085 99 4195 109
rect 4085 8 4095 99
rect 4095 8 4185 99
rect 4185 8 4195 99
rect 4085 -2 4195 8
rect 5259 101 5369 111
rect 5259 10 5269 101
rect 5269 10 5359 101
rect 5359 10 5369 101
rect 5259 0 5369 10
rect 6427 101 6537 111
rect 6427 10 6437 101
rect 6437 10 6527 101
rect 6527 10 6537 101
rect 6427 0 6537 10
rect 7595 101 7705 111
rect 7595 10 7605 101
rect 7605 10 7695 101
rect 7695 10 7705 101
rect 7595 0 7705 10
rect 8763 101 8873 111
rect 8763 10 8773 101
rect 8773 10 8863 101
rect 8863 10 8873 101
rect 8763 0 8873 10
<< metal4 >>
rect 458 1440 9450 1506
rect 458 1320 1038 1440
rect 1160 1414 9450 1440
rect 1160 1412 4578 1414
rect 1160 1348 2240 1412
rect 2304 1348 3408 1412
rect 3472 1350 4578 1412
rect 4642 1350 5750 1414
rect 5814 1412 8086 1414
rect 5814 1350 6918 1412
rect 3472 1348 6918 1350
rect 6982 1350 8086 1412
rect 8150 1350 9254 1414
rect 9318 1350 9450 1414
rect 6982 1348 9450 1350
rect 1160 1320 9450 1348
rect 458 1310 9450 1320
rect 5258 111 5370 112
rect 5258 110 5259 111
rect 458 109 5259 110
rect 458 -2 581 109
rect 691 -2 1749 109
rect 1859 -2 2917 109
rect 3027 -2 4085 109
rect 4195 0 5259 109
rect 5369 110 5370 111
rect 6426 111 6538 112
rect 6426 110 6427 111
rect 5369 0 6427 110
rect 6537 110 6538 111
rect 7594 111 7706 112
rect 7594 110 7595 111
rect 6537 0 7595 110
rect 7705 110 7706 111
rect 8762 111 8874 112
rect 8762 110 8763 111
rect 7705 0 8763 110
rect 8873 110 8874 111
rect 8873 0 9556 110
rect 4195 -2 9556 0
rect 458 -86 9556 -2
<< labels >>
flabel metal4 4764 -86 5044 110 1 FreeSerif 800 0 0 0 VSS
port 2 n
flabel metal1 366 1368 466 1450 1 FreeSerif 480 0 0 0 B[0]
port 3 n
flabel metal1 366 1108 458 1190 1 FreeSerif 480 0 0 0 A[0]
port 4 n
flabel metal1 1534 1108 1626 1190 1 FreeSerif 480 0 0 0 A[1]
port 5 n
flabel metal1 2702 1108 2794 1190 1 FreeSerif 480 0 0 0 A[2]
port 6 n
flabel metal1 3870 1108 3962 1190 1 FreeSerif 480 0 0 0 A[3]
port 7 n
flabel metal1 5044 1110 5136 1192 1 FreeSerif 480 0 0 0 A[4]
port 8 n
flabel metal1 6212 1110 6304 1192 1 FreeSerif 480 0 0 0 A[5]
port 9 n
flabel metal1 7380 1110 7472 1192 1 FreeSerif 480 0 0 0 A[6]
port 10 n
flabel metal1 8548 1110 8640 1192 1 FreeSerif 480 0 0 0 A[7]
port 11 n
flabel metal1 9224 538 9320 588 1 FreeSerif 480 0 0 0 Y[7]
port 12 n
flabel metal1 8056 538 8152 588 1 FreeSerif 480 0 0 0 Y[6]
port 13 n
flabel metal1 6888 538 6984 588 1 FreeSerif 480 0 0 0 Y[5]
port 14 n
flabel metal1 5720 538 5816 588 1 FreeSerif 480 0 0 0 Y[4]
port 15 n
flabel metal1 4546 536 4642 586 1 FreeSerif 480 0 0 0 Y[3]
port 16 n
flabel metal1 3378 536 3474 586 1 FreeSerif 480 0 0 0 Y[2]
port 17 n
flabel metal1 2210 536 2306 586 1 FreeSerif 480 0 0 0 Y[1]
port 18 n
flabel metal1 1042 536 1138 586 1 FreeSerif 480 0 0 0 Y[0]
port 19 n
flabel metal1 1534 1368 1634 1450 1 FreeSerif 480 0 0 0 B[1]
port 20 n
flabel metal1 2702 1368 2802 1450 1 FreeSerif 480 0 0 0 B[2]
port 21 n
flabel metal1 3870 1368 3970 1450 1 FreeSerif 480 0 0 0 B[3]
port 22 n
flabel metal1 5044 1370 5144 1452 1 FreeSerif 480 0 0 0 B[4]
port 23 n
flabel metal1 6212 1370 6312 1452 1 FreeSerif 480 0 0 0 B[5]
port 24 n
flabel metal1 7380 1370 7480 1452 1 FreeSerif 480 0 0 0 B[6]
port 25 n
flabel metal1 8548 1370 8648 1452 1 FreeSerif 480 0 0 0 B[7]
port 26 n
flabel metal4 4786 1366 4910 1454 1 FreeSerif 800 0 0 0 VDD
port 27 n
<< end >>
