* NGSPICE file created from inverter_pex.ext - technology: sky130B

.subckt inverter IN VDD OUT VSS
X0 OUT.t3 IN.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 OUT.t2 IN.t1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 VDD.t1 IN.t2 OUT.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 OUT.t0 IN.t3 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 IN.n0 IN.t1 188.514
R1 IN.n0 IN.t0 188.514
R2 IN.n1 IN.t3 137.369
R3 IN.n0 IN.t2 110.859
R4 IN.n1 IN.n0 61.856
R5 IN IN.n1 13.908
R6 VDD.n2 VDD.t2 173.615
R7 VDD.n3 VDD.t4 170.169
R8 VDD.n1 VDD.t5 29.197
R9 VDD.n0 VDD.t3 28.565
R10 VDD.n0 VDD.t1 28.565
R11 VDD.n1 VDD.n0 0.375
R12 VDD.n3 VDD.t0 0.244
R13 VDD.n4 VDD.n1 0.078
R14 VDD.n4 VDD 0.034
R15 VDD.t0 VDD.n2 0.021
R16 VDD.n4 VDD.n3 0.002
R17 VDD VDD.n4 0.001
R18 OUT.n1 OUT.n0 194.26
R19 OUT.n1 OUT.t2 28.568
R20 OUT.n0 OUT.t1 28.565
R21 OUT.n0 OUT.t3 28.565
R22 OUT OUT.t0 18.129
R23 OUT OUT.n2 0.593
R24 OUT.n2 OUT 0.593
R25 OUT OUT.n1 0.5
R26 OUT.n2 OUT 0.078
R27 OUT.n2 OUT 0.049
R28 OUT.n2 OUT 0.049
R29 VSS.n0 VSS.t0 17.972
R30 VSS.n0 VSS 0.023
R31 VSS VSS.n0 0.001
C0 VDD IN 0.19fF
C1 OUT IN 0.06fF
C2 OUT VDD 0.90fF
.ends

