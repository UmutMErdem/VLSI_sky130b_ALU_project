magic
tech sky130B
magscale 1 2
timestamp 1736110968
<< nwell >>
rect 458 725 1372 1504
rect 888 466 1372 725
rect 887 418 1372 466
rect 887 142 1371 418
<< nmos >>
rect 462 204 522 404
rect 580 204 640 404
rect 698 204 758 404
<< pmos >>
rect 552 787 612 1187
rect 670 787 730 1187
rect 788 787 848 1187
rect 906 787 966 1187
rect 1024 787 1084 1187
rect 1142 787 1202 1187
rect 981 204 1041 404
rect 1099 204 1159 404
rect 1217 204 1277 404
<< ndiff >>
rect 404 392 462 404
rect 404 216 416 392
rect 450 216 462 392
rect 404 204 462 216
rect 522 392 580 404
rect 522 216 534 392
rect 568 216 580 392
rect 522 204 580 216
rect 640 392 698 404
rect 640 216 652 392
rect 686 216 698 392
rect 640 204 698 216
rect 758 392 816 404
rect 758 216 770 392
rect 804 216 816 392
rect 758 204 816 216
<< pdiff >>
rect 494 1175 552 1187
rect 494 799 506 1175
rect 540 799 552 1175
rect 494 787 552 799
rect 612 1175 670 1187
rect 612 799 624 1175
rect 658 799 670 1175
rect 612 787 670 799
rect 730 1175 788 1187
rect 730 799 742 1175
rect 776 799 788 1175
rect 730 787 788 799
rect 848 1175 906 1187
rect 848 799 860 1175
rect 894 799 906 1175
rect 848 787 906 799
rect 966 1175 1024 1187
rect 966 799 978 1175
rect 1012 799 1024 1175
rect 966 787 1024 799
rect 1084 1175 1142 1187
rect 1084 799 1096 1175
rect 1130 799 1142 1175
rect 1084 787 1142 799
rect 1202 1175 1260 1187
rect 1202 799 1214 1175
rect 1248 799 1260 1175
rect 1202 787 1260 799
rect 923 392 981 404
rect 923 216 935 392
rect 969 216 981 392
rect 923 204 981 216
rect 1041 392 1099 404
rect 1041 216 1053 392
rect 1087 216 1099 392
rect 1041 204 1099 216
rect 1159 392 1217 404
rect 1159 216 1171 392
rect 1205 216 1217 392
rect 1159 204 1217 216
rect 1277 392 1335 404
rect 1277 216 1289 392
rect 1323 216 1335 392
rect 1277 204 1335 216
<< ndiffc >>
rect 416 216 450 392
rect 534 216 568 392
rect 652 216 686 392
rect 770 216 804 392
<< pdiffc >>
rect 506 799 540 1175
rect 624 799 658 1175
rect 742 799 776 1175
rect 860 799 894 1175
rect 978 799 1012 1175
rect 1096 799 1130 1175
rect 1214 799 1248 1175
rect 935 216 969 392
rect 1053 216 1087 392
rect 1171 216 1205 392
rect 1289 216 1323 392
<< psubdiff >>
rect 538 82 734 112
rect 538 16 578 82
rect 696 16 734 82
rect 538 -32 734 16
<< nsubdiff >>
rect 978 1426 1244 1464
rect 978 1354 1034 1426
rect 1178 1354 1244 1426
rect 978 1324 1244 1354
<< psubdiffcont >>
rect 578 16 696 82
<< nsubdiffcont >>
rect 1034 1354 1178 1426
<< poly >>
rect 400 1348 466 1364
rect 400 1314 416 1348
rect 450 1344 466 1348
rect 450 1314 950 1344
rect 400 1301 950 1314
rect 400 1298 466 1301
rect 400 1249 466 1256
rect 906 1249 950 1301
rect 400 1240 848 1249
rect 400 1206 416 1240
rect 450 1208 848 1240
rect 450 1207 612 1208
rect 450 1206 466 1207
rect 400 1190 466 1206
rect 552 1187 612 1207
rect 670 1187 730 1208
rect 788 1187 848 1208
rect 906 1208 1202 1249
rect 906 1187 966 1208
rect 1024 1187 1084 1208
rect 1142 1187 1202 1208
rect 552 770 612 787
rect 552 681 613 770
rect 670 761 730 787
rect 788 761 848 787
rect 462 628 613 681
rect 462 404 522 628
rect 906 586 966 787
rect 1024 761 1084 787
rect 1142 761 1202 787
rect 580 535 966 586
rect 580 404 640 535
rect 695 477 761 493
rect 695 443 711 477
rect 745 443 761 477
rect 695 427 761 443
rect 698 404 758 427
rect 981 404 1041 430
rect 1099 404 1159 430
rect 1217 404 1277 430
rect 462 178 522 204
rect 580 178 640 204
rect 698 172 758 204
rect 981 172 1041 204
rect 1099 172 1159 204
rect 1217 172 1277 204
rect 698 131 1277 172
<< polycont >>
rect 416 1314 450 1348
rect 416 1206 450 1240
rect 711 443 745 477
<< locali >>
rect 1002 1426 1206 1438
rect 1002 1354 1034 1426
rect 1178 1354 1206 1426
rect 1002 1352 1064 1354
rect 1144 1352 1206 1354
rect 400 1314 416 1348
rect 450 1314 466 1348
rect 1002 1336 1206 1352
rect 400 1206 416 1240
rect 450 1206 466 1240
rect 506 1175 540 1191
rect 506 783 540 799
rect 624 1175 658 1191
rect 624 783 658 799
rect 742 1175 776 1191
rect 742 783 776 799
rect 860 1175 894 1191
rect 860 783 894 799
rect 978 1175 1012 1191
rect 978 783 1012 799
rect 1096 1175 1130 1191
rect 1096 783 1130 799
rect 1214 1175 1248 1191
rect 1214 783 1248 799
rect 695 443 711 477
rect 745 443 761 477
rect 416 392 450 408
rect 416 200 450 216
rect 534 392 568 408
rect 534 200 568 216
rect 652 392 686 408
rect 652 200 686 216
rect 770 392 804 408
rect 770 200 804 216
rect 935 392 969 408
rect 935 200 969 216
rect 1053 392 1087 408
rect 1053 200 1087 216
rect 1171 392 1205 408
rect 1171 200 1205 216
rect 1289 392 1323 408
rect 1289 200 1323 216
rect 560 86 702 98
rect 560 82 600 86
rect 666 82 702 86
rect 560 16 578 82
rect 696 16 702 82
rect 560 -10 702 16
<< viali >>
rect 1064 1354 1144 1424
rect 1064 1352 1144 1354
rect 416 1314 450 1348
rect 416 1206 450 1240
rect 506 799 540 1175
rect 624 799 658 1175
rect 742 799 776 1175
rect 860 799 894 1175
rect 978 799 1012 1175
rect 1096 799 1130 1175
rect 1214 799 1248 1175
rect 711 443 745 477
rect 416 216 450 392
rect 534 216 568 392
rect 652 216 686 392
rect 770 216 804 392
rect 935 216 969 392
rect 1053 216 1087 392
rect 1171 216 1205 392
rect 1289 216 1323 392
rect 600 82 666 86
rect 600 16 666 82
<< metal1 >>
rect 366 1348 466 1450
rect 366 1314 416 1348
rect 450 1314 466 1348
rect 1052 1424 1156 1430
rect 1052 1352 1064 1424
rect 1144 1352 1156 1424
rect 1052 1346 1156 1352
rect 366 1288 466 1314
rect 1087 1290 1122 1346
rect 366 1240 466 1260
rect 366 1206 416 1240
rect 450 1206 466 1240
rect 366 1108 466 1206
rect 624 1249 894 1277
rect 624 1187 658 1249
rect 860 1187 894 1249
rect 978 1249 1248 1290
rect 978 1187 1012 1249
rect 1214 1187 1248 1249
rect 500 1175 546 1187
rect 500 799 506 1175
rect 540 799 546 1175
rect 500 787 546 799
rect 618 1175 664 1187
rect 618 799 624 1175
rect 658 799 664 1175
rect 618 787 664 799
rect 736 1175 782 1187
rect 736 799 742 1175
rect 776 799 782 1175
rect 736 787 782 799
rect 854 1175 900 1187
rect 854 799 860 1175
rect 894 799 900 1175
rect 854 787 900 799
rect 972 1175 1018 1187
rect 972 799 978 1175
rect 1012 799 1018 1175
rect 972 787 1018 799
rect 1090 1175 1136 1187
rect 1090 799 1096 1175
rect 1130 799 1136 1175
rect 1090 787 1136 799
rect 1208 1175 1254 1187
rect 1208 799 1214 1175
rect 1248 799 1254 1175
rect 1208 787 1254 799
rect 506 745 540 787
rect 742 745 776 787
rect 506 717 776 745
rect 860 746 894 787
rect 1096 746 1130 787
rect 860 717 1130 746
rect 506 669 540 717
rect 506 639 569 669
rect 534 547 569 639
rect 1214 604 1248 787
rect 534 511 761 547
rect 534 404 569 511
rect 695 477 761 511
rect 695 443 711 477
rect 745 443 761 477
rect 1042 535 1139 586
rect 1214 550 1323 604
rect 1042 468 1099 535
rect 695 437 761 443
rect 936 432 1205 468
rect 936 404 969 432
rect 1172 404 1205 432
rect 1289 404 1323 550
rect 410 392 456 404
rect 410 216 416 392
rect 450 216 456 392
rect 410 204 456 216
rect 528 392 574 404
rect 528 216 534 392
rect 568 216 574 392
rect 528 204 574 216
rect 646 392 692 404
rect 646 216 652 392
rect 686 216 692 392
rect 646 204 692 216
rect 764 392 810 404
rect 764 216 770 392
rect 804 337 810 392
rect 929 392 975 404
rect 929 337 935 392
rect 804 249 935 337
rect 804 216 810 249
rect 764 204 810 216
rect 929 216 935 249
rect 969 216 975 392
rect 929 204 975 216
rect 1047 392 1093 404
rect 1047 216 1053 392
rect 1087 216 1093 392
rect 1047 204 1093 216
rect 1165 392 1211 404
rect 1165 216 1171 392
rect 1205 216 1211 392
rect 1165 204 1211 216
rect 1283 392 1329 404
rect 1283 216 1289 392
rect 1323 216 1329 392
rect 1283 204 1329 216
rect 416 165 450 204
rect 652 165 686 204
rect 416 126 686 165
rect 1053 166 1086 204
rect 1289 166 1322 204
rect 1053 130 1322 166
rect 616 98 650 126
rect 594 86 672 98
rect 594 16 600 86
rect 666 16 672 86
rect 594 4 672 16
<< via1 >>
rect 1078 1353 1130 1405
rect 607 29 659 81
<< metal2 >>
rect 1056 1426 1146 1436
rect 1056 1325 1146 1335
rect 591 99 681 109
rect 591 -2 681 8
<< via2 >>
rect 1056 1405 1146 1426
rect 1056 1353 1078 1405
rect 1078 1353 1130 1405
rect 1130 1353 1146 1405
rect 1056 1335 1146 1353
rect 591 81 681 99
rect 591 29 607 81
rect 607 29 659 81
rect 659 29 681 81
rect 591 8 681 29
<< metal3 >>
rect 1028 1320 1038 1440
rect 1160 1320 1170 1440
rect 571 -2 581 109
rect 691 -2 701 109
<< via3 >>
rect 1038 1426 1160 1440
rect 1038 1335 1056 1426
rect 1056 1335 1146 1426
rect 1146 1335 1160 1426
rect 1038 1320 1160 1335
rect 581 99 691 109
rect 581 8 591 99
rect 591 8 681 99
rect 681 8 691 99
rect 581 -2 691 8
<< metal4 >>
rect 954 1440 1258 1504
rect 954 1320 1038 1440
rect 1160 1320 1258 1440
rect 954 1310 1258 1320
rect 580 109 692 110
rect 580 98 581 109
rect 522 -2 581 98
rect 691 98 692 109
rect 691 -2 752 98
rect 522 -64 752 -2
<< labels >>
flabel metal1 1049 541 1132 580 1 FreeSans 240 0 0 0 OUT
port 6 n
flabel metal4 1024 1320 1188 1432 1 FreeSerif 560 0 0 0 VDD
port 9 n
flabel metal4 548 -22 720 88 1 FreeSerif 560 0 0 0 VSS
port 10 n
flabel metal1 366 1110 464 1208 1 FreeSerif 480 0 0 0 A
port 14 n
flabel metal1 368 1378 466 1446 1 FreeSerif 480 0 0 0 B
port 15 n
<< end >>
