* NGSPICE file created from control_unit_pex.ext - technology: sky130B

.subckt control_unit B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7] A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7] Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7] VDD VSS opcode[0],opcode[1],opcode[2],opcode[3] Cout
X0 VDD.t3602 a_48690_23619.t4 a_49686_24206.t5 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 VDD.t1053 a_3642_11724.t4 a_3951_1740.t5 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2 a_39263_15765.t3 a_38721_16161.t4 VDD.t3539 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3 VDD.t1090 a_13130_8992.t4 a_13711_11724.t5 VDD.t1089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 VDD.t1325 A[3].t0 a_19763_16387.t2 VDD.t1324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 a_59280_15743.t3 a_59223_16436.t8 VSS.t319 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 VSS.t645 a_42301_n1318.t4 a_44682_3363.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 VDD.t1273 a_63527_6198.t7 a_64117_5761.t2 VDD.t1272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 VSS.t300 a_70513_4160.t8 a_7957_1259.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 a_46175_15029.t0 a_45279_16157.t4 VSS.t526 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 a_52710_16433.t2 a_54665_15740.t4 a_54253_15766.t3 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_54914_n1762.t2 B[6].t0 VDD.t1378 VDD.t1377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X12 VDD.t231 a_44405_8194.t4 a_48548_6884.t2 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 VDD.t4607 VSS.t714 a_3591_21596.t5 VDD.t4606 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 VDD.t3008 A[6].t0 a_9867_21592.t2 VDD.t3007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 VSS.t42 a_48124_21370.t8 a_49477_22063.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X16 a_52999_20434.t1 A[2].t0 a_52762_21071.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_31377_10037.t1 a_30152_10818.t4 a_30645_10037.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 VDD.t262 A[4].t0 a_5331_6357.t2 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X19 VDD.t2973 a_53343_23888.t4 a_55078_24197.t2 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 a_56502_14835.t1 a_51813_16162.t4 VSS.t480 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X21 VDD.t3232 a_61518_24201.t5 a_61782_23618.t2 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X22 VDD.t3740 A[7].t0 a_42770_18699.t3 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 VDD.t263 A[4].t1 a_62375_18703.t5 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X24 a_44405_8194.t0 a_47794_3876.t5 VDD.t2884 VDD.t2883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X25 VDD.t884 a_59635_6910.t8 a_61415_6910.t2 VDD.t883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X26 VDD.t233 a_44405_8194.t5 a_44460_6616.t6 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 VDD.t2740 a_53816_17942.t5 a_52749_18576.t2 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 a_31379_12341.t0 B[0].t0 VSS.t352 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X29 a_4332_n2152.t4 a_4857_n2637.t4 a_3983_n2152.t6 VDD.t2737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X30 a_47794_3876.t2 a_45049_1913.t4 VSS.t667 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X31 a_556_13728.t3 a_1735_13585.t4 a_1680_13125.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X32 VDD.t2914 opcode[2].t0 a_3392_1740.t2 VDD.t2913 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X33 a_4243_8992.t6 a_4183_8966.t8 a_3710_8262.t2 VDD.t4514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X34 VDD.t2890 a_70513_7304.t8 a_11101_1259.t2 VDD.t2889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X35 a_566_8262.t6 a_1745_8119.t4 a_1099_8992.t8 VDD.t1774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X36 a_55469_11532.t2 a_54879_11969.t7 VDD.t2098 VDD.t2097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X37 a_23777_10847.t3 opcode[1].t0 VSS.t136 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X38 a_37916_8132.t6 a_35594_7027.t4 VDD.t3701 VDD.t3700 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X39 a_48130_1040.t11 a_48542_1014.t4 a_48248_1040.t7 VDD.t2575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X40 a_67135_3808.t4 a_54908_6842.t8 VDD.t4567 VDD.t4566 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 VDD.t254 a_30645_10037.t8 a_48006_21370.t10 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X42 VSS.t279 a_1974_8339.t4 a_1926_7659.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X43 a_41948_n1318.t0 B[5].t0 a_41711_n1755.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X44 VDD.t1489 a_30647_12105.t8 a_39706_24333.t6 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X45 VDD.t1761 a_70513_19926.t8 a_23723_1259.t2 VDD.t1760 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 VDD.t992 a_49832_23623.t4 a_52762_21071.t0 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X47 a_48124_21370.t7 a_47579_22063.t4 a_48124_20638.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 VDD.t3684 a_16274_8992.t4 a_16855_11724.t11 VDD.t3683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X49 a_1916_10391.t1 opcode[1].t1 a_556_10994.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X50 a_17456_7659.t0 a_16805_8966.t8 VSS.t209 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X51 VDD.t1007 a_7464_n2148.t8 Y[5].t2 VDD.t1006 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X52 a_16865_8992.t10 a_17511_8119.t4 a_16332_8262.t5 VDD.t1798 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 a_29950_n2431.t11 a_30150_n1593.t4 a_30643_n2374.t4 VDD.t1750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 a_54785_1041.t11 a_53005_1041.t8 VDD.t1502 VDD.t1501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 a_20643_8115.t2 opcode[0].t0 VDD.t3690 VDD.t3689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 VDD.t1545 B[7].t0 a_13849_16387.t2 VDD.t1544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 VDD.t1323 A[3].t1 a_63532_11802.t2 VDD.t1322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X58 a_53430_9674.t5 a_51695_9365.t4 VDD.t580 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X59 VDD.t585 a_498_11724.t4 a_807_1740.t11 VDD.t584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X60 a_10519_8988.t2 opcode[0].t1 VDD.t4012 VDD.t4011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X61 a_58329_6179.t2 a_57739_6616.t7 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X62 a_45811_7603.t2 a_41507_3295.t4 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 a_13661_8966.t4 a_18447_5326.t4 a_18035_5352.t3 VDD.t1623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X64 a_7381_20723.t2 opcode[0].t2 VDD.t4535 VDD.t4534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X65 VDD.t1490 a_30647_12105.t9 a_41066_22066.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X66 a_6842_8258.t6 a_7315_8962.t8 a_7375_8988.t8 VDD.t3288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X67 a_44445_4000.t6 a_41697_1042.t8 VDD.t1666 VDD.t1665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X68 a_70513_20044.t11 a_64122_11365.t4 VDD.t2846 VDD.t2845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X69 a_839_n2152.t8 a_1713_n2637.t4 a_1188_n2152.t5 VDD.t2357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X70 VDD.t84 a_51054_2325.t4 a_51109_747.t5 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 a_56850_21339.t2 a_49832_23623.t5 VDD.t993 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X72 a_35602_9612.t2 a_35012_10049.t7 VDD.t4352 VDD.t4351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 VDD.t4137 B[1].t0 a_11640_16408.t2 VDD.t4136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 VDD.t4504 a_46176_16428.t8 a_46233_15735.t2 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X75 a_60193_3291.t3 a_59929_3874.t5 VSS.t334 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X76 VDD.t1573 a_62660_24205.t5 a_58326_16165.t2 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X77 a_1424_n3485.t0 a_779_n2178.t4 VSS.t437 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X78 a_45821_15761.t11 a_46233_15735.t4 a_45939_15761.t6 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X79 VSS.t155 a_6832_13724.t8 a_6774_14454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_15966_5352.t2 B[4].t0 VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X81 VDD.t792 opcode[1].t2 a_70513_4278.t11 VDD.t791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X82 VDD.t895 A[0].t0 a_39706_24333.t0 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X83 VDD.t2902 a_37916_8132.t7 a_38506_7695.t2 VDD.t2901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 VDD.t754 a_30645_5900.t8 a_59311_24329.t2 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 a_52473_15766.t4 a_51815_16459.t4 a_52355_15766.t5 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X86 a_43173_24209.t5 a_42177_23622.t4 VDD.t2799 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 a_54540_21365.t5 a_54113_22058.t4 a_54658_21365.t4 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 VSS.t543 a_6827_15753.t5 a_6887_15819.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 VDD.t3538 a_38721_16161.t5 a_39263_15765.t2 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 a_8021_8115.t3 opcode[0].t3 VSS.t469 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X91 a_7083_1744.t2 a_6774_11720.t4 VDD.t2058 VDD.t2057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X92 a_70513_4278.t0 a_52473_15766.t8 a_70513_4160.t0 VDD.t662 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X93 a_55202_6816.t2 a_51059_8126.t4 VDD.t4285 VDD.t4284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X94 a_11565_15824.t2 a_11505_15751.t5 VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X95 VDD.t4335 a_35602_9612.t4 a_40101_6796.t2 VDD.t4334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X96 a_70455_n1231.t3 opcode[1].t3 VSS.t137 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X97 a_45939_15761.t3 a_46176_16428.t9 a_46175_15029.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X98 a_70455_1913.t3 opcode[1].t4 VSS.t138 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X99 VDD.t86 a_51054_2325.t5 a_54785_1041.t1 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X100 a_51114_6548.t6 a_48815_11511.t4 VDD.t2261 VDD.t2260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X101 a_3591_21596.t4 VSS.t715 VDD.t4605 VDD.t4604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X102 a_63598_4278.t6 A[3].t2 VDD.t1321 VDD.t1320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X103 a_61769_6178.t0 a_59635_6910.t9 a_61533_6910.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X104 a_55853_15446.t6 A[5].t0 a_56502_14835.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X105 a_3424_n2152.t2 opcode[3].t0 VDD.t4551 VDD.t4550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X106 a_61782_23618.t1 a_61518_24201.t6 VDD.t3233 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X107 a_38484_3565.t3 a_37894_4002.t7 VSS.t707 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X108 a_9976_13724.t7 a_11155_13581.t4 a_10509_14454.t8 VDD.t3564 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 a_23787_8115.t2 opcode[0].t4 VDD.t1353 VDD.t1352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X110 VDD.t325 a_60201_9159.t4 a_61197_9746.t5 VDD.t324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X111 VDD.t371 a_3700_13728.t8 a_3642_14458.t2 VDD.t370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X112 VDD.t897 A[0].t1 a_8289_6359.t2 VDD.t896 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X113 a_67372_6666.t1 a_64117_5761.t4 a_67135_7303.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X114 a_3983_n2152.t5 a_4857_n2637.t5 a_4332_n2152.t3 VDD.t2738 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 VDD.t3952 a_16795_16385.t7 a_7305_14428.t2 VDD.t3951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X116 a_1916_13125.t1 opcode[0].t5 a_556_13728.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X117 a_35591_989.t2 a_35001_1426.t7 VDD.t2736 VDD.t2735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X118 VDD.t923 B[4].t1 a_15966_5352.t1 VDD.t922 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X119 a_70509_n1998.t2 a_39381_15765.t8 a_70509_n2116.t1 VDD.t576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X120 a_48248_308.t1 a_48542_1014.t5 VSS.t471 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X121 VDD.t680 a_48855_n1313.t4 a_52887_1041.t8 VDD.t679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X122 a_48254_6910.t2 a_47709_7603.t4 a_48136_6910.t2 VDD.t2159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X123 a_51709_7715.t3 a_51119_8152.t7 VSS.t205 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X124 VDD.t1380 B[6].t1 a_63595_1208.t2 VDD.t1379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X125 VDD.t2195 B[0].t1 a_23700_6043.t2 VDD.t2194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X126 VSS.t26 a_41507_3295.t5 a_44702_7583.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X127 a_20611_n2633.t2 a_20054_1744.t8 VDD.t3044 VDD.t3043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X128 VDD.t379 a_1964_13805.t4 a_1089_14458.t11 VDD.t378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X129 VDD.t4569 a_54908_6842.t9 a_65651_3118.t8 VDD.t4568 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X130 a_55202_6816.t3 a_51059_8126.t5 VSS.t674 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X131 a_53576_9091.t3 a_53312_9674.t5 VSS.t265 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X132 a_4568_n3485.t1 a_3923_n2178.t4 VSS.t50 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X133 a_3951_1740.t7 a_3392_1740.t4 a_4300_1740.t3 VDD.t2290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X134 a_22489_21592.t11 A[0].t2 a_21956_20862.t7 VDD.t898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X135 a_48006_21370.t9 a_30645_10037.t9 VDD.t255 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X136 VDD.t4026 A[2].t1 a_20103_5350.t7 VDD.t4025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X137 a_40296_23896.t2 a_39706_24333.t7 VDD.t1543 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X138 VSS.t523 a_42756_17049.t7 a_40011_18575.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X139 a_1156_1740.t6 a_1681_1255.t4 a_807_1740.t3 VDD.t557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X140 VDD.t794 opcode[1].t5 a_70513_7422.t11 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X141 VDD.t668 A[5].t1 a_55862_18700.t5 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X142 a_1745_8119.t1 opcode[0].t6 VSS.t610 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X143 VSS.t396 a_508_8992.t4 a_1916_10391.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X144 a_44399_2324.t2 a_67133_11394.t7 VDD.t535 VDD.t534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X145 a_41587_6822.t5 a_41999_6796.t4 a_41705_6822.t2 VDD.t972 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X146 a_63010_16442.t0 a_30645_3831.t8 VSS.t94 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X147 a_46215_18571.t2 a_47282_17937.t5 VDD.t3632 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X148 a_16213_21596.t11 a_16859_20723.t4 a_15680_20866.t4 VDD.t3384 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X149 a_63532_11802.t1 A[3].t3 VDD.t1319 VDD.t1318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X150 a_19464_8258.t4 a_20643_8115.t4 a_20588_7655.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X151 VDD.t1317 A[3].t4 a_19357_21596.t8 VDD.t1316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X152 a_41991_1016.t2 a_37848_2326.t4 VDD.t1936 VDD.t1935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X153 a_57722_4002.t6 a_54903_1041.t8 VDD.t1017 VDD.t1016 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 a_41066_22066.t1 a_30647_12105.t10 VDD.t1491 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X155 VDD.t3878 opcode[0].t7 a_29954_7911.t4 VDD.t3877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X156 a_16805_8966.t5 a_19563_6043.t4 a_20103_5350.t8 VDD.t3385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X157 VDD.t542 a_57730_9870.t7 a_58320_9433.t2 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X158 a_13011_21592.t5 A[3].t5 a_12478_20862.t3 VDD.t3282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X159 a_40799_18571.t2 a_42770_18699.t7 VDD.t960 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X160 a_30647_7968.t5 a_30154_7310.t4 a_29954_7911.t7 VDD.t1424 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X161 a_29952_3774.t5 a_30152_3173.t4 a_30645_3831.t1 VDD.t1132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X162 a_37908_2352.t2 a_35591_989.t4 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X163 a_70455_1913.t2 opcode[1].t6 VDD.t796 VDD.t795 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X164 a_1099_8992.t3 a_1974_8339.t5 VDD.t1715 VDD.t1714 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 a_46233_15735.t1 a_46176_16428.t10 VDD.t4505 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X166 a_1188_n2152.t7 opcode[3].t1 a_1424_n3485.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X167 a_41152_1735.t2 a_39799_1042.t8 VDD.t1752 VDD.t1751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X168 a_13657_20719.t2 opcode[0].t8 VDD.t3678 VDD.t3677 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X169 VDD.t4109 B[5].t1 a_30150_1105.t2 VDD.t4108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X170 a_39706_24333.t1 A[0].t3 VDD.t899 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X171 a_59311_24329.t1 a_30645_5900.t9 VDD.t755 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X172 a_52355_15766.t4 a_51815_16459.t5 a_52473_15766.t3 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X173 a_9668_1744.t2 opcode[2].t1 VDD.t2916 VDD.t2915 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X174 a_54658_21365.t3 a_54113_22058.t5 a_54540_21365.t4 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X175 a_6827_15753.t0 B[5].t2 VSS.t648 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X176 VDD.t1260 a_9334_20862.t8 a_7055_n2174.t2 VDD.t1259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X177 a_6813_6359.t2 A[2].t2 VDD.t4028 VDD.t4027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X178 a_3642_11724.t2 a_3700_10994.t8 VDD.t2691 VDD.t2690 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X179 VDD.t642 a_11505_15751.t6 a_11565_15824.t1 VDD.t641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X180 a_58868_15769.t8 a_58326_16165.t4 VDD.t977 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X181 a_70509_1028.t2 a_45939_15761.t8 a_70509_1146.t2 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X182 a_30645_3831.t4 a_30152_4612.t4 a_29952_3774.t9 VDD.t1431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X183 a_61407_1042.t11 a_59627_1042.t8 VDD.t564 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X184 VDD.t756 a_30645_5900.t10 a_60671_22062.t2 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X185 a_45939_15029.t1 a_46233_15735.t5 a_45939_15761.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 VDD.t3880 opcode[3].t2 a_19178_n2148.t2 VDD.t3879 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X187 VDD.t959 a_61518_24201.t7 a_61782_23618.t0 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X188 a_48136_6910.t11 a_44405_8194.t6 VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X189 a_70509_1028.t6 a_70455_1913.t4 a_71842_1737.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X190 a_70509_10624.t2 a_65769_n1230.t8 VDD.t3860 VDD.t3859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 a_40859_18597.t2 a_40799_18571.t4 VDD.t1351 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X192 a_11165_8115.t2 opcode[0].t9 VDD.t3868 VDD.t3867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X193 a_4332_n2152.t2 a_4857_n2637.t6 a_3983_n2152.t4 VDD.t2739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X194 VSS.t65 a_1964_13805.t5 a_1916_13125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X195 a_30645_n306.t2 a_30152_n964.t4 a_29952_n363.t5 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X196 VSS.t646 a_42301_n1318.t5 a_44696_1713.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X197 VDD.t2068 a_63527_9231.t7 a_64117_8794.t2 VDD.t2067 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X198 a_66063_6587.t2 a_64117_5761.t5 VDD.t1139 VDD.t1138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X199 a_1089_14458.t10 a_1964_13805.t6 VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X200 a_59627_1042.t6 a_59082_1735.t4 a_59627_310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X201 a_62375_18703.t0 a_30645_3831.t9 VDD.t536 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X202 a_4332_n2152.t5 opcode[3].t3 a_4568_n3485.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X203 VDD.t2702 a_35575_3749.t4 a_40093_1016.t2 VDD.t2701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X204 a_21956_20862.t6 A[0].t4 a_22489_21592.t10 VDD.t2314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X205 VDD.t147 A[1].t0 a_48006_21370.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 VSS.t283 a_59187_17949.t5 a_51813_16162.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X207 VDD.t3679 a_39706_24333.t8 a_40296_23896.t1 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X208 VDD.t2397 a_54713_3294.t4 a_57744_8220.t2 VDD.t2396 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X209 a_39807_6090.t1 a_40101_6796.t4 VSS.t673 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X210 a_8021_8115.t2 opcode[0].t10 VDD.t3810 VDD.t3809 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X211 a_54790_6842.t11 a_53010_6842.t8 VDD.t2592 VDD.t2591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X212 VDD.t257 a_53891_18572.t4 a_53951_18598.t5 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X213 a_10227_1744.t8 opcode[2].t2 VDD.t2918 VDD.t2917 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X214 VDD.t1492 a_30647_12105.t11 a_41066_22066.t0 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X215 VSS.t353 B[0].t2 a_30154_11447.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X216 a_56102_24201.t3 a_53357_22238.t4 a_56220_24201.t5 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X217 VDD.t798 opcode[1].t7 a_4879_10851.t2 VDD.t797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X218 a_70459_8189.t3 opcode[1].t8 VSS.t139 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X219 a_35594_7027.t0 a_35004_7464.t7 VDD.t2794 VDD.t2793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X220 VDD.t2721 a_43055_24209.t5 a_43319_23626.t2 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X221 a_5794_16410.t5 A[6].t1 a_5659_15753.t4 VDD.t3009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X222 VDD.t612 a_55853_15446.t7 a_54245_18572.t2 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X223 VSS.t46 A[4].t2 a_5331_6357.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X224 a_52762_21071.t5 A[2].t3 VDD.t4029 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X225 a_70513_16900.t11 opcode[1].t9 VDD.t800 VDD.t799 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X226 a_10509_11720.t2 a_9918_14454.t4 a_9976_10990.t2 VDD.t2819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X227 a_49904_21370.t5 a_48124_21370.t9 VDD.t4077 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X228 VSS.t374 a_55848_17050.t7 a_53103_18576.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X229 VDD.t3145 a_46652_3872.t5 a_46916_3289.t2 VDD.t3144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X230 VSS.t222 a_30154_7310.t5 a_31379_7968.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X231 a_70509_13650.t6 a_70455_14535.t4 a_70509_13768.t8 VDD.t2248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X232 a_14357_10851.t3 opcode[1].t10 VSS.t140 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X233 VDD.t4139 B[1].t1 a_29952_9980.t2 VDD.t4138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X234 a_35594_7027.t1 a_35004_7464.t8 VSS.t452 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X235 a_57676_2326.t3 a_67135_3808.t7 VSS.t642 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X236 a_51690_3564.t2 a_51100_4001.t7 VDD.t2188 VDD.t2187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X237 VDD.t757 a_30645_5900.t11 a_59311_24329.t0 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X238 a_70459_17667.t2 opcode[1].t11 VDD.t802 VDD.t801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X239 a_19997_8988.t8 a_19937_8962.t8 a_19464_8258.t1 VDD.t2127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X240 VDD.t3053 a_7432_1744.t8 a_7989_n2633.t2 VDD.t3052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X241 a_54540_21365.t9 a_54952_21339.t4 a_54658_21365.t5 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X242 VSS.t120 A[5].t2 a_6827_15753.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X243 VDD.t4085 a_42301_n1318.t6 a_44459_2350.t6 VDD.t4084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X244 a_7055_n2174.t1 a_9334_20862.t9 VDD.t1262 VDD.t1261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X245 a_15946_15776.t0 B[6].t2 VSS.t215 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X246 VSS.t123 a_42761_15445.t7 a_41153_18571.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X247 a_13721_8992.t6 a_13661_8966.t8 a_13188_8262.t4 VDD.t4235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X248 a_70509_n1998.t3 a_61343_9163.t4 VDD.t357 VDD.t356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X249 VSS.t249 a_38721_16161.t6 a_38723_16458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X250 VDD.t2693 a_3700_10994.t9 a_3642_11724.t3 VDD.t2692 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X251 VDD.t2762 a_9976_10990.t8 a_9918_11720.t2 VDD.t2761 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X252 a_70455_n1231.t2 opcode[1].t12 VDD.t804 VDD.t803 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X253 VDD.t3682 opcode[0].t11 a_22489_21592.t2 VDD.t3681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X254 a_11565_15824.t0 a_11505_15751.t7 VDD.t644 VDD.t643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X255 VDD.t978 a_58326_16165.t5 a_58868_15769.t7 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X256 VDD.t2167 a_48254_6910.t8 a_51105_9802.t2 VDD.t2166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X257 VDD.t2594 a_53010_6842.t9 a_54790_6842.t10 VDD.t2593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X258 a_60671_22062.t1 a_30645_5900.t12 VDD.t758 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X259 a_43509_21373.t4 a_42964_22066.t4 a_43509_20641.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X260 a_14498_15776.t0 B[7].t1 VSS.t243 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X261 VDD.t806 opcode[1].t13 a_70459_5045.t2 VDD.t805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X262 VDD.t2500 a_508_8992.t5 a_1089_11724.t5 VDD.t2499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X263 a_19178_n2148.t1 opcode[3].t4 VDD.t3882 VDD.t3881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X264 a_61189_3878.t5 a_60193_3291.t4 VDD.t1894 VDD.t1893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X265 a_65769_6613.t7 a_65224_7306.t4 a_65651_6613.t11 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X266 VSS.t311 a_56366_23618.t4 a_63350_20637.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X267 a_30645_3831.t0 opcode[0].t12 a_31377_4067.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X268 a_11155_13581.t2 opcode[0].t13 VDD.t3830 VDD.t3829 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X269 VDD.t1110 a_64192_n2074.t4 a_67135_n540.t6 VDD.t1109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X270 a_45279_16157.t0 a_52674_17946.t5 VDD.t395 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X271 a_6832_13724.t4 a_8011_13581.t4 a_7365_14454.t8 VDD.t1328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X272 a_40724_17941.t3 a_41153_18571.t4 a_40859_18597.t3 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X273 VDD.t3884 opcode[3].t5 a_839_n2152.t9 VDD.t3883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X274 VDD.t390 a_37903_748.t7 a_38493_311.t2 VDD.t389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X275 a_47912_3876.t5 a_45049_1913.t5 a_47794_3876.t3 VDD.t4245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X276 VDD.t1092 a_13130_8992.t5 a_13711_11724.t4 VDD.t1091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X277 a_13188_8262.t0 a_14367_8119.t4 a_13721_8992.t0 VDD.t963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X278 VSS.t453 a_60758_18575.t4 a_60329_17945.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X279 a_20515_5324.t2 A[2].t4 VDD.t4031 VDD.t4030 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X280 a_52460_1734.t2 a_48855_n1313.t5 VDD.t1229 VDD.t1228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X281 a_22526_4620.t0 B[1].t2 VSS.t651 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X282 VDD.t4337 a_35602_9612.t5 a_37902_9782.t3 VDD.t4336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X283 VDD.t149 A[1].t1 a_7551_6363.t2 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X284 a_9986_8258.t3 a_11165_8115.t4 a_11110_7655.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X285 a_54914_n1762.t1 B[6].t3 VDD.t1382 VDD.t1381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X286 VDD.t205 a_35591_989.t5 a_37894_4002.t3 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X287 a_70513_19926.t4 a_43509_21373.t8 a_70513_20044.t3 VDD.t2694 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X288 a_4233_11724.t11 opcode[1].t14 VDD.t808 VDD.t807 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X289 a_41161_15765.t10 A[7].t1 VDD.t3741 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X290 a_7989_n2633.t1 a_7432_1744.t9 VDD.t3055 VDD.t3054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X291 a_70459_20811.t2 opcode[1].t15 VDD.t810 VDD.t809 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X292 a_61178_15743.t3 a_30645_3831.t10 VSS.t95 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X293 a_65651_n1230.t11 a_64192_n2074.t5 VDD.t1112 VDD.t1111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X294 VDD.t537 a_30645_3831.t11 a_62375_18703.t1 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X295 VSS.t9 a_30152_n964.t5 a_31377_n306.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X296 a_11080_n3481.t1 a_9700_n2148.t4 a_10608_n2148.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X297 a_4804_n3485.t0 a_3424_n2152.t4 a_4332_n2152.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X298 a_22489_21592.t9 A[0].t5 a_21956_20862.t5 VDD.t2315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X299 a_48006_21370.t1 A[1].t2 VDD.t150 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X300 a_59187_17949.t1 a_59262_18579.t4 VSS.t163 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X301 VDD.t967 a_47800_9746.t5 a_48064_9163.t2 VDD.t966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X302 a_38498_1915.t3 a_37908_2352.t7 VSS.t266 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X303 a_40296_23896.t0 a_39706_24333.t9 VDD.t3680 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X304 VSS.t152 a_3058_20866.t8 a_779_n2178.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X305 a_51709_7715.t2 a_51119_8152.t8 VDD.t1286 VDD.t1285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X306 a_57739_6616.t2 a_55469_11532.t4 VDD.t3500 VDD.t3499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X307 a_54903_309.t0 a_55197_1015.t4 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X308 a_46350_1040.t3 a_45805_1733.t4 a_46350_308.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X309 a_46356_6178.t1 a_46650_6884.t4 VSS.t57 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X310 VSS.t444 a_62361_17053.t7 a_59616_18579.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X311 a_23141_8988.t11 a_23081_8962.t8 a_22608_8258.t7 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X312 VDD.t2718 a_55848_17050.t8 a_53103_18576.t2 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X313 a_38721_16161.t0 a_46140_17941.t5 VDD.t1106 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X314 a_19464_8258.t7 a_20643_8115.t5 a_19997_8988.t5 VDD.t583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X315 VDD.t4339 a_35602_9612.t6 a_39689_6822.t2 VDD.t4338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X316 a_53951_18598.t4 a_53891_18572.t5 VDD.t258 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X317 VDD.t3291 a_45279_16157.t5 a_45281_16454.t2 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X318 a_16865_8992.t2 a_16805_8966.t9 a_16332_8262.t1 VDD.t1334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X319 a_24594_4618.t0 B[0].t3 VSS.t354 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X320 a_14357_13585.t3 opcode[0].t14 VSS.t607 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X321 a_70509_1146.t11 opcode[1].t16 VDD.t812 VDD.t811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X322 a_51059_8126.t0 a_67135_n540.t7 VDD.t2996 VDD.t2995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X323 a_46176_16428.t0 a_47179_16454.t4 a_47719_15761.t8 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X324 VSS.t15 a_51054_2325.t6 a_51346_110.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X325 VDD.t1938 a_37848_2326.t5 a_41579_1042.t8 VDD.t1937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X326 VSS.t52 a_15426_6045.t4 a_16084_4620.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X327 a_56220_24201.t4 a_53357_22238.t5 a_56102_24201.t2 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X328 a_19454_13724.t7 a_19927_14428.t4 a_19987_14454.t11 VDD.t384 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X329 a_4879_10851.t1 opcode[1].t17 VDD.t814 VDD.t813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X330 a_29954_7911.t9 B[2].t0 VDD.t3725 VDD.t3724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X331 a_43319_23626.t1 a_43055_24209.t6 VDD.t345 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X332 a_5659_15753.t3 A[6].t2 a_5794_16410.t4 VDD.t3010 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X333 a_9976_10990.t1 a_9918_14454.t5 a_10509_11720.t1 VDD.t368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X334 a_58312_3565.t3 a_57722_4002.t7 VSS.t223 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X335 VDD.t669 A[5].t3 a_53713_16459.t2 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X336 a_61636_24201.t5 a_59910_20638.t4 a_61518_24201.t0 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X337 a_13602_20259.t0 A[3].t6 VSS.t259 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X338 VDD.t4078 a_48124_21370.t10 a_49904_21370.t4 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X339 a_3652_8992.t2 a_3710_8262.t8 VDD.t2541 VDD.t2540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X340 a_17501_10851.t2 opcode[1].t18 VDD.t816 VDD.t815 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X341 a_43391_21373.t11 a_43803_21347.t4 a_43509_21373.t5 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X342 a_50022_21370.t4 a_49477_22063.t4 a_50022_20638.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X343 a_71842_14595.t1 opcode[1].t19 a_70509_13650.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X344 VDD.t1031 opcode[0].t15 a_30154_12886.t2 VDD.t1030 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X345 VDD.t2102 a_5108_13805.t4 a_4233_14458.t11 VDD.t2101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X346 a_29950_n2431.t0 B[7].t2 VDD.t1547 VDD.t1546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X347 a_65651_3118.t1 a_65224_3811.t4 a_65769_3118.t5 VDD.t376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X348 VDD.t2317 A[0].t6 a_24240_5350.t8 VDD.t2316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X349 VDD.t1264 a_9334_20862.t10 a_7055_n2174.t0 VDD.t1263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X350 a_25633_21592.t11 VSS.t716 a_25100_20862.t7 VDD.t4603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X351 VDD.t3554 a_556_10994.t8 a_498_11724.t2 VDD.t3553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 VSS.t561 a_556_10994.t9 a_498_11724.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X353 a_16014_1740.t2 opcode[2].t3 VDD.t2920 VDD.t2919 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X354 a_29952_5843.t6 a_30152_6681.t4 a_30645_5900.t6 VDD.t3286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X355 a_37848_2326.t0 a_41251_9658.t5 VDD.t2140 VDD.t2139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X356 a_29952_3774.t8 opcode[0].t16 VDD.t4006 VDD.t4005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X357 VDD.t3742 A[7].t2 a_42761_15445.t6 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X358 a_18035_5352.t10 B[3].t0 VDD.t2652 VDD.t2651 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X359 a_44405_8194.t1 a_47794_3876.t6 VSS.t465 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X360 a_65769_6613.t2 a_66063_6587.t4 a_65651_6613.t4 VDD.t2053 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X361 VDD.t759 a_30645_5900.t13 a_60671_22062.t0 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X362 VDD.t264 A[4].t3 a_62366_15449.t3 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X363 a_14310_5328.t3 A[5].t4 VSS.t121 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X364 a_43745_20641.t1 a_41611_21373.t8 a_43509_21373.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X365 a_13849_16387.t6 A[7].t3 a_14498_15776.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X366 VDD.t309 a_53576_9091.t4 a_54572_9678.t2 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X367 a_3983_n2152.t3 a_3424_n2152.t5 a_4332_n2152.t1 VDD.t575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X368 VDD.t3886 opcode[3].t6 a_19178_n2148.t0 VDD.t3885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 a_63114_20637.t0 a_63408_21343.t4 VSS.t324 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X370 VDD.t1900 a_70513_4160.t9 a_7957_1259.t2 VDD.t1899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X371 VDD.t2922 opcode[2].t4 a_22290_1744.t2 VDD.t2921 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X372 a_9986_8258.t5 a_10459_8962.t8 a_10519_8988.t3 VDD.t1976 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X373 a_48130_1040.t10 a_48542_1014.t6 a_48248_1040.t6 VDD.t2907 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X374 a_40859_18597.t4 a_41153_18571.t5 a_40724_17941.t2 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X375 VDD.t1504 a_6842_8258.t8 a_6784_8988.t2 VDD.t1503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X376 VSS.t635 A[2].t5 a_6813_6359.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X377 a_61819_1016.t2 a_57676_2326.t4 VDD.t1639 VDD.t1638 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X378 VDD.t2654 B[3].t1 a_30152_5242.t2 VDD.t2653 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X379 a_30647_12105.t4 a_30154_11447.t4 a_29954_12048.t11 VDD.t3907 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X380 a_4243_8992.t3 opcode[0].t17 VDD.t1338 VDD.t1337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X381 VSS.t239 a_6842_8258.t9 a_6784_8988.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X382 a_29950_1706.t11 a_30150_2544.t4 a_30643_1763.t7 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X383 a_54113_22058.t1 a_30647_7968.t8 VDD.t1915 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X384 VSS.t47 A[4].t4 a_17040_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X385 a_49319_15441.t3 A[6].t3 a_49968_14830.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X386 VDD.t1384 B[6].t4 a_54914_n1762.t0 VDD.t1383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X387 VDD.t818 opcode[1].t20 a_4233_11724.t10 VDD.t817 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X388 a_11100_10387.t0 a_9918_14454.t6 VSS.t63 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X389 VDD.t3743 A[7].t4 a_41161_15765.t9 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X390 VSS.t614 a_55853_15446.t8 a_54245_18572.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X391 VDD.t820 opcode[1].t21 a_10509_11720.t8 VDD.t819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X392 a_46770_3872.t5 a_45035_3563.t4 VDD.t2632 VDD.t2631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 a_59627_1042.t0 a_59921_1016.t4 a_59509_1042.t7 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X394 VDD.t2318 A[0].t7 a_41493_21373.t11 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X395 VDD.t151 A[1].t3 a_48418_21344.t2 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X396 a_62375_18703.t2 a_30645_3831.t12 VDD.t538 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X397 VSS.t440 a_4857_n2637.t7 a_4804_n3485.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X398 a_60980_1735.t2 a_59627_1042.t9 VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X399 VSS.t483 a_59616_18579.t4 a_59187_17949.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X400 a_39681_1042.t2 a_35591_989.t6 VDD.t207 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X401 a_46232_1040.t2 a_45805_1733.t5 a_46350_1040.t2 VDD.t1979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X402 a_35001_1426.t5 B[3].t2 VDD.t2656 VDD.t2655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X403 a_21860_15776.t0 B[2].t1 VSS.t594 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X404 a_21956_20862.t1 a_23135_20719.t4 a_23080_20259.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X405 a_11165_8115.t3 opcode[0].t18 VSS.t536 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X406 a_10227_1744.t0 a_9918_11720.t4 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X407 VDD.t879 a_54658_21365.t8 a_56011_22058.t2 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X408 VDD.t4376 A[3].t7 a_18035_5352.t6 VDD.t4375 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X409 VDD.t2924 opcode[2].t5 a_13429_1740.t5 VDD.t2923 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X410 a_53816_17942.t1 a_54245_18572.t4 a_53951_18598.t0 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X411 a_45281_16454.t1 a_45279_16157.t6 VDD.t3292 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X412 a_70455_n1231.t1 opcode[1].t22 VDD.t822 VDD.t821 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X413 a_51114_2351.t2 a_51054_2325.t7 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X414 a_67135_3808.t3 a_54908_6842.t10 VDD.t4571 VDD.t4570 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X415 a_46650_6884.t0 a_42266_11512.t4 VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X416 VDD.t4032 A[2].t6 a_54952_21339.t2 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X417 a_41697_310.t1 a_41991_1016.t4 VSS.t56 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X418 a_47719_15761.t7 a_47179_16454.t5 a_46176_16428.t1 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X419 VSS.t693 a_55504_n1325.t4 a_57959_3365.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X420 a_54253_15766.t1 A[5].t5 VDD.t670 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X421 a_19987_14454.t10 a_19927_14428.t5 a_19454_13724.t6 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X422 a_17692_7659.t0 opcode[0].t19 a_16332_8262.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X423 a_41697_1042.t5 a_41152_1735.t4 a_41579_1042.t5 VDD.t2149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X424 a_48542_1014.t0 a_44399_2324.t4 VDD.t2064 VDD.t2063 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X425 VSS.t156 a_556_13728.t8 a_498_14458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X426 a_10509_11720.t0 a_9918_14454.t7 a_9976_10990.t0 VDD.t369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X427 VDD.t4374 A[3].t8 a_6071_6357.t2 VDD.t4373 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X428 a_61415_6910.t11 a_57684_8194.t4 VDD.t3580 VDD.t3579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X429 VDD.t496 a_59901_23892.t4 a_61636_24201.t0 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X430 a_12478_20862.t4 a_13657_20719.t4 a_13602_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X431 a_49904_21370.t3 a_48124_21370.t11 VDD.t4079 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X432 VSS.t74 a_566_8262.t8 a_508_8992.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X433 a_40109_9654.t1 a_38501_6091.t4 VSS.t182 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X434 a_7083_1744.t1 a_6774_11720.t5 VDD.t2060 VDD.t2059 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X435 a_55202_6816.t1 a_51059_8126.t6 VDD.t4287 VDD.t4286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X436 VSS.t145 a_54658_21365.t9 a_56011_22058.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X437 a_10519_8988.t10 a_11165_8115.t5 a_9986_8258.t2 VDD.t2716 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X438 VDD.t3537 a_38721_16161.t7 a_42756_17049.t5 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X439 a_44445_4000.t5 a_41697_1042.t9 VDD.t1668 VDD.t1667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X440 VDD.t511 a_42266_11512.t5 a_44451_9870.t2 VDD.t510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_64188_3841.t2 a_63598_4278.t7 VDD.t2801 VDD.t2800 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X442 a_30647_12105.t7 opcode[0].t20 a_31379_12341.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X443 a_46350_1040.t7 a_46644_1014.t4 a_46232_1040.t8 VDD.t3327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X444 a_70513_20044.t8 opcode[1].t23 VDD.t824 VDD.t823 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X445 a_498_11724.t1 a_556_10994.t10 VDD.t3556 VDD.t3555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X446 VSS.t567 a_17447_1255.t4 a_17394_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X447 a_807_1740.t0 a_248_1740.t4 a_1156_1740.t0 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 a_54363_7535.t2 a_53010_6842.t10 VDD.t2596 VDD.t2595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X449 VSS.t432 a_47711_18567.t4 a_47282_17937.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X450 VDD.t1117 a_13778_1740.t8 a_14335_n2637.t2 VDD.t1116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X451 a_19357_21596.t9 A[1].t4 a_18824_20866.t7 VDD.t1921 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X452 VDD.t3329 a_6832_10990.t8 a_6774_11720.t3 VDD.t3328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X453 a_50022_21370.t7 a_49477_22063.t5 a_49904_21370.t11 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X454 a_62366_15449.t2 A[4].t5 VDD.t265 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X455 a_22172_5352.t6 A[1].t5 VDD.t1923 VDD.t1922 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X456 VDD.t2926 opcode[2].t6 a_248_1740.t2 VDD.t2925 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X457 a_49314_17045.t3 a_45279_16157.t7 a_49963_16434.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X458 VDD.t3334 a_8056_15820.t4 a_10509_14454.t9 VDD.t3333 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X459 a_11289_6045.t2 B[6].t5 VDD.t1386 VDD.t1385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X460 VDD.t974 a_48064_9163.t4 a_52887_1041.t2 VDD.t973 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X461 a_48254_6910.t6 a_48548_6884.t4 a_48136_6910.t5 VDD.t4023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X462 a_31377_6136.t1 B[3].t3 VSS.t425 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X463 VDD.t4491 a_19454_10990.t8 a_19396_11720.t2 VDD.t4490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X464 a_4857_n2637.t0 a_4300_1740.t8 VSS.t344 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X465 a_20611_n2633.t1 a_20054_1744.t9 VDD.t3046 VDD.t3045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X466 VSS.t135 a_11101_1259.t4 a_11048_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X467 a_41579_1042.t11 a_41991_1016.t5 a_41697_1042.t6 VDD.t2988 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X468 a_1156_1740.t5 a_1681_1255.t5 a_807_1740.t4 VDD.t558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X469 VDD.t2154 a_18824_20866.t8 a_16545_n2178.t2 VDD.t2153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X470 a_23131_14454.t6 a_23071_14428.t4 a_22598_13724.t5 VDD.t1135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X471 a_22849_1744.t11 a_22290_1744.t4 a_23198_1744.t6 VDD.t3114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X472 a_7115_n2148.t8 a_7055_n2174.t4 VDD.t2772 VDD.t2771 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X473 VDD.t1348 a_56102_24201.t5 a_56366_23618.t2 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X474 a_4233_11724.t9 opcode[1].t24 VDD.t826 VDD.t825 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X475 a_9761_5354.t8 a_9221_6047.t4 a_1039_8966.t4 VDD.t3362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X476 a_10608_n2148.t0 a_11133_n2633.t4 a_10259_n2148.t8 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X477 a_48418_21344.t1 A[1].t6 VDD.t1924 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X478 a_60766_15769.t8 A[4].t6 VDD.t266 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X479 a_44451_9870.t6 a_41507_3295.t6 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X480 VSS.t24 a_11289_6045.t4 a_11947_4620.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X481 a_44399_2324.t3 a_67133_11394.t8 VSS.t93 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X482 a_31375_1763.t1 a_30150_2544.t5 a_30643_1763.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X483 VDD.t3284 a_42756_17049.t8 a_40011_18575.t2 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X484 a_51337_3364.t1 a_48064_9163.t5 a_51100_4001.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X485 a_57722_4002.t5 a_54903_1041.t9 VDD.t1019 VDD.t1018 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X486 a_16805_8966.t6 a_19563_6043.t5 a_20103_5350.t9 VDD.t3386 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 a_46233_22680.t2 a_43319_23626.t4 VDD.t2566 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X488 a_29954_12048.t5 B[0].t4 VDD.t2197 VDD.t2196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X489 VDD.t3940 opcode[0].t21 a_17511_8119.t2 VDD.t3939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X490 a_23316_20259.t0 opcode[0].t22 a_21956_20862.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X491 VDD.t268 A[4].t7 a_15966_5352.t7 VDD.t267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X492 a_12808_16408.t2 B[0].t5 VDD.t2199 VDD.t2198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X493 a_67370_10757.t0 a_64117_8794.t4 a_67133_11394.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X494 a_54908_6842.t0 a_54363_7535.t4 a_54790_6842.t3 VDD.t458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X495 VDD.t2263 a_48815_11511.t5 a_53304_6816.t2 VDD.t2262 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X496 a_25100_20862.t1 a_26279_20719.t4 a_25633_21592.t6 VDD.t2182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X497 a_38498_1915.t2 a_37908_2352.t8 VDD.t1633 VDD.t1632 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X498 a_53425_3873.t5 a_51699_310.t4 a_53307_3873.t4 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X499 a_53951_18598.t1 a_54245_18572.t5 a_53816_17942.t2 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X500 VDD.t3293 a_45279_16157.t8 a_45281_16454.t0 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X501 a_41153_18571.t2 a_42761_15445.t8 VDD.t677 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X502 VDD.t3117 a_40101_3874.t5 a_40365_3291.t2 VDD.t3116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X503 a_51059_8126.t1 a_67135_n540.t8 VSS.t485 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X504 VDD.t2074 A[5].t6 a_54253_15766.t5 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X505 VDD.t1693 a_6813_6359.t4 a_16865_8992.t4 VDD.t1692 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X506 VDD.t2169 a_48254_6910.t9 a_52465_7535.t2 VDD.t2168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X507 VDD.t3923 opcode[0].t23 a_29954_12048.t2 VDD.t3922 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X508 VDD.t2567 a_43319_23626.t5 a_49904_21370.t8 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X509 a_48124_21370.t3 a_47579_22063.t5 a_48006_21370.t5 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X510 a_61407_1042.t10 a_59627_1042.t10 VDD.t568 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X511 VDD.t943 a_3058_20866.t9 a_779_n2178.t1 VDD.t942 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X512 a_54903_1041.t4 a_54358_1734.t4 a_54785_1041.t7 VDD.t1552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X513 a_46809_23893.t3 a_46219_24330.t7 VSS.t423 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X514 a_46238_6910.t8 a_46650_6884.t5 a_46356_6910.t6 VDD.t330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X515 a_59322_18605.t5 a_59262_18579.t5 VDD.t989 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X516 a_20290_411.t1 a_19396_11720.t4 VSS.t202 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X517 a_20003_20723.t3 opcode[0].t24 VSS.t281 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X518 VSS.t71 a_52674_17946.t6 a_45279_16157.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X519 a_35591_989.t3 a_35001_1426.t8 VSS.t317 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X520 a_70513_4160.t4 a_70459_5045.t4 a_71846_4869.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X521 VSS.t467 a_22709_16385.t7 a_19927_14428.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X522 a_64185_771.t2 a_63595_1208.t7 VDD.t1791 VDD.t1790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X523 VDD.t4372 A[3].t9 a_18447_5326.t2 VDD.t4371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X524 Y[4].t2 a_10608_n2148.t8 VDD.t746 VDD.t745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X525 VSS.t185 a_64192_n2074.t6 a_65224_n537.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X526 a_58986_15037.t0 a_59280_15743.t4 a_58986_15769.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X527 VDD.t1595 a_556_10994.t11 a_498_11724.t0 VDD.t1594 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X528 a_53304_6816.t1 a_48815_11511.t6 VDD.t2265 VDD.t2264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X529 a_58326_1915.t3 a_57736_2352.t7 VSS.t493 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X530 a_18243_16385.t5 A[4].t8 VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X531 a_47918_9746.t2 a_45055_7783.t4 a_47800_9746.t1 VDD.t4536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X532 a_30643_n2374.t0 opcode[0].t25 a_31375_n2138.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X533 a_13657_20719.t3 opcode[0].t26 VSS.t562 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X534 a_46922_9159.t2 a_46658_9742.t5 VDD.t1756 VDD.t1755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X535 a_59635_6178.t0 a_59929_6884.t4 VSS.t39 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X536 VSS.t43 a_30645_10037.t10 a_46470_22043.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X537 a_49328_18695.t6 a_30645_n306.t8 VDD.t3364 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X538 a_62375_18703.t6 A[4].t9 a_63024_18092.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X539 a_19396_11720.t1 a_19454_10990.t9 VDD.t4493 VDD.t4492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X540 VDD.t2658 B[3].t4 a_17495_6045.t2 VDD.t2657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X541 VSS.t36 a_9168_15798.t5 a_9228_15824.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X542 a_65224_n537.t2 a_64192_n2074.t7 VDD.t3480 VDD.t3479 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X543 a_53005_1041.t1 a_52460_1734.t4 a_52887_1041.t3 VDD.t2136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X544 a_52355_15766.t2 a_52710_16433.t8 VDD.t1130 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 a_44465_8220.t6 a_44405_8194.t7 VDD.t237 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X546 a_59517_6910.t2 a_54713_3294.t5 VDD.t2399 VDD.t2398 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X547 VDD.t1096 a_5331_6357.t4 a_10519_8988.t9 VDD.t1095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X548 VSS.t129 a_30645_5900.t14 a_60671_22062.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X549 VDD.t2774 a_7055_n2174.t5 a_7115_n2148.t7 VDD.t2773 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 a_70455_11391.t3 opcode[1].t25 VSS.t141 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X551 a_48130_1040.t6 a_46350_1040.t8 VDD.t4425 VDD.t4424 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 VSS.t596 A[7].t5 a_40621_16458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X553 a_20579_1259.t2 a_70513_16782.t8 VDD.t3322 VDD.t3321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X554 VDD.t271 A[4].t10 a_60766_15769.t7 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X555 a_44454_746.t2 a_44399_2324.t5 VDD.t2066 VDD.t2065 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X556 VDD.t925 B[4].t2 a_29952_3774.t2 VDD.t924 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X557 a_30645_5900.t0 a_30152_5242.t4 a_29952_5843.t0 VDD.t441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X558 a_40011_18575.t1 a_42756_17049.t9 VDD.t3285 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X559 a_1735_10851.t2 opcode[1].t26 VDD.t828 VDD.t827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X560 VDD.t2279 a_13120_11724.t4 a_13429_1740.t6 VDD.t2278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X561 a_11165_8115.t1 opcode[0].t27 VDD.t1604 VDD.t1603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X562 VDD.t256 a_30645_10037.t11 a_46233_22680.t6 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X563 VDD.t4196 a_40799_18571.t5 a_40859_18597.t1 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X564 a_70513_7304.t4 a_70459_8189.t4 a_70513_7422.t6 VDD.t3242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X565 VDD.t830 opcode[1].t27 a_70455_1913.t1 VDD.t829 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X566 a_59548_23692.t1 A[3].t10 a_59311_24329.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X567 VSS.t626 A[2].t7 a_23316_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X568 VDD.t57 a_37856_8106.t4 a_37911_6528.t6 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X569 VSS.t172 a_60329_17945.t5 a_59262_18579.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X570 VDD.t2201 B[0].t6 a_12808_16408.t1 VDD.t2200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X571 a_35594_7027.t2 a_35004_7464.t9 VDD.t2796 VDD.t2795 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X572 a_45821_15761.t5 a_45279_16157.t9 VDD.t3294 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X573 a_41676_11949.t6 A[6].t4 VDD.t3012 VDD.t3011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X574 VDD.t2110 a_4593_6357.t4 a_7375_8988.t5 VDD.t2109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X575 a_30152_475.t2 opcode[0].t28 VDD.t3494 VDD.t3493 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X576 a_53816_17942.t3 a_54245_18572.t6 a_53951_18598.t2 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 a_52887_1041.t4 a_52460_1734.t5 a_53005_1041.t2 VDD.t2137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X578 VDD.t678 a_42761_15445.t9 a_41153_18571.t1 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X579 a_1681_1255.t2 a_70509_n2116.t8 VDD.t3038 VDD.t3037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X580 a_13898_5354.t2 B[5].t3 VDD.t4111 VDD.t4110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X581 VSS.t694 a_55504_n1325.t5 a_59082_1735.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X582 a_30645_10037.t0 a_30152_9379.t4 a_29952_9980.t6 VDD.t2150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X583 VDD.t2361 a_57744_8220.t7 a_58334_7783.t2 VDD.t2360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X584 a_21632_6045.t2 B[1].t3 VDD.t4141 VDD.t4140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X585 a_59863_310.t1 a_55504_n1325.t6 a_59627_1042.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X586 VSS.t3 a_7995_15753.t5 a_8056_15820.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X587 VDD.t1597 opcode[0].t29 a_30150_n1593.t0 VDD.t1596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X588 a_51109_747.t4 a_51054_2325.t8 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X589 VDD.t513 a_42266_11512.t6 a_46238_6910.t5 VDD.t512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X590 a_54253_15766.t6 A[5].t7 VDD.t2075 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X591 a_53571_3290.t2 a_53307_3873.t5 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X592 VDD.t4087 a_42301_n1318.t7 a_44459_2350.t5 VDD.t4086 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X593 a_13721_8992.t5 a_13661_8966.t9 a_13188_8262.t3 VDD.t4236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X594 a_49568_24206.t3 a_46823_22243.t4 VSS.t492 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X595 a_49904_21370.t7 a_43319_23626.t6 VDD.t2568 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X596 VDD.t2719 a_55848_17050.t9 a_53103_18576.t1 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X597 VDD.t3858 a_61533_6910.t8 a_70509_1146.t5 VDD.t3857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X598 VDD.t4289 a_51059_8126.t7 a_54790_6842.t8 VDD.t4288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X599 a_779_n2178.t2 a_3058_20866.t10 VDD.t945 VDD.t944 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X600 VSS.t426 a_51690_3564.t4 a_53307_3873.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X601 a_30647_12105.t0 a_30154_12886.t4 a_29954_12048.t8 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X602 a_7083_1744.t8 a_7957_1259.t4 a_7432_1744.t3 VDD.t2898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X603 VDD.t273 A[4].t11 a_16378_5326.t2 VDD.t272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X604 a_41991_1016.t3 a_37848_2326.t6 VSS.t308 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X605 VSS.t413 a_30645_10037.t12 a_46456_23693.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X606 a_4879_10851.t0 opcode[1].t28 VDD.t832 VDD.t831 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X607 VDD.t275 A[4].t12 a_63527_6198.t0 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X608 VDD.t277 A[4].t13 a_18243_16385.t4 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X609 VSS.t305 A[1].t7 a_7551_6363.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X610 a_1039_8966.t7 A[7].t6 a_10115_4622.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X611 a_55139_309.t1 a_53005_1041.t9 a_54903_1041.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X612 a_53010_6842.t4 a_52465_7535.t4 a_53010_6110.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X613 a_41369_9658.t5 a_38506_7695.t4 a_41251_9658.t3 VDD.t767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X614 a_22550_8988.t2 a_22608_8258.t8 VDD.t2768 VDD.t2767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X615 VDD.t2453 a_13401_n2178.t4 a_13461_n2152.t2 VDD.t2452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X616 VSS.t306 A[1].t8 a_26460_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X617 a_62361_17053.t2 a_30645_3831.t13 VDD.t539 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X618 VDD.t4222 a_19454_10990.t10 a_19396_11720.t0 VDD.t4221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X619 a_30152_10818.t2 opcode[0].t30 VSS.t633 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X620 VDD.t3162 a_53307_3873.t6 a_53571_3290.t1 VDD.t3161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X621 VDD.t1131 a_52710_16433.t9 a_52355_15766.t1 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X622 a_46776_9742.t5 a_45050_6179.t4 a_46658_9742.t0 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X623 a_10259_n2148.t5 a_9700_n2148.t5 a_10608_n2148.t6 VDD.t3574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X624 a_30152_4612.t2 opcode[0].t31 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X625 a_13178_13728.t4 a_14357_13585.t4 a_13711_14458.t8 VDD.t387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 a_37903_748.t6 a_35575_3749.t5 VDD.t2704 VDD.t2703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X627 a_22489_21592.t1 opcode[0].t32 VDD.t3812 VDD.t3811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X628 VSS.t549 a_46922_9159.t4 a_47800_9746.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X629 a_61525_1042.t5 a_60980_1735.t4 a_61407_1042.t6 VDD.t2840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X630 a_7115_n2148.t6 a_7055_n2174.t6 VDD.t2118 VDD.t2117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X631 VSS.t472 opcode[2].t7 a_22290_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X632 a_61415_6910.t9 a_61827_6884.t4 a_61533_6910.t6 VDD.t3140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X633 VDD.t979 a_58326_16165.t6 a_62366_15449.t6 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X634 a_16378_5326.t1 A[4].t14 VDD.t279 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X635 VSS.t647 a_42301_n1318.t8 a_45805_1733.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X636 a_70513_4278.t10 opcode[1].t29 VDD.t834 VDD.t833 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X637 VSS.t312 a_56366_23618.t5 a_59557_20438.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X638 a_47912_3876.t2 a_46916_3289.t4 VDD.t2776 VDD.t2775 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X639 a_62996_21369.t2 a_61216_21369.t8 VDD.t527 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X640 VDD.t1660 a_42756_17049.t10 a_40011_18575.t0 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X641 VDD.t836 opcode[1].t30 a_1735_10851.t1 VDD.t835 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 a_13188_8262.t5 a_14367_8119.t5 a_13721_8992.t7 VDD.t3471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X643 VDD.t2569 a_43319_23626.t7 a_46228_21076.t6 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X644 a_22290_4620.t0 a_22584_5326.t4 a_19937_8962.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X645 a_24240_5350.t11 a_23700_6043.t4 a_23081_8962.t7 VDD.t1478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X646 a_46233_22680.t5 a_30645_10037.t13 VDD.t2585 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X647 a_51813_16162.t1 a_59187_17949.t6 VDD.t1747 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X648 a_23141_8988.t2 opcode[0].t33 VDD.t3876 VDD.t3875 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X649 VDD.t209 a_35591_989.t7 a_37894_4002.t4 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X650 VSS.t181 a_5331_6357.t5 a_11346_7655.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X651 a_10459_8962.t0 A[4].t15 a_16320_4620.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X652 a_60329_17945.t4 a_60404_18575.t4 VSS.t525 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X653 a_12808_16408.t0 B[0].t7 VDD.t2203 VDD.t2202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X654 VDD.t4506 a_46176_16428.t11 a_45821_15761.t8 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X655 VDD.t3874 a_16332_8262.t8 a_16274_8992.t3 VDD.t3873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X656 a_39807_6822.t2 a_39262_7515.t4 a_39689_6822.t3 VDD.t2882 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X657 a_52892_6842.t2 a_48254_6910.t10 VDD.t901 VDD.t900 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X658 a_70513_16900.t0 a_50022_21370.t8 a_70513_16782.t2 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X659 VSS.t91 a_22550_8988.t4 a_23958_10387.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X660 VDD.t969 a_47800_9746.t6 a_48064_9163.t1 VDD.t968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X661 a_23131_11720.t8 a_23777_10847.t4 a_22598_10990.t4 VDD.t2362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X662 VDD.t658 a_45041_9433.t4 a_46776_9742.t0 VDD.t657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X663 a_55197_1015.t3 a_51054_2325.t9 VSS.t16 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X664 a_57739_6616.t1 a_55469_11532.t5 VDD.t3498 VDD.t3497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X665 a_23135_20719.t2 opcode[0].t34 VDD.t3832 VDD.t3831 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X666 VDD.t2785 a_65769_6613.t8 a_70513_16900.t3 VDD.t2784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X667 VSS.t197 a_48855_n1313.t6 a_52460_1734.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X668 a_7995_15753.t0 B[4].t3 VSS.t150 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X669 a_65649_10704.t10 a_41705_6822.t8 VDD.t3617 VDD.t3616 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X670 VDD.t1388 B[6].t6 a_30152_n964.t2 VDD.t1387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X671 a_10608_n2148.t7 opcode[3].t7 a_10844_n3481.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 VSS.t328 A[5].t8 a_53713_16459.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X673 a_35238_789.t1 B[3].t5 a_35001_1426.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X674 a_41611_21373.t4 a_41905_21347.t4 a_41493_21373.t3 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X675 VSS.t350 a_9986_8258.t8 a_9928_8988.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X676 a_70459_5045.t1 opcode[1].t31 VDD.t682 VDD.t681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X677 VSS.t572 a_48690_23619.t5 a_49568_24206.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X678 a_53103_18576.t0 a_55848_17050.t10 VDD.t2720 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X679 a_70455_14535.t2 opcode[1].t32 VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X680 a_22322_n2148.t2 opcode[3].t8 VDD.t3888 VDD.t3887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X681 a_41251_9658.t2 a_38506_7695.t5 VSS.t132 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X682 VSS.t584 a_30150_1105.t4 a_31375_1763.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X683 VDD.t947 a_3058_20866.t11 a_779_n2178.t3 VDD.t946 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X684 a_59280_15743.t2 a_59223_16436.t9 VDD.t4560 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 VDD.t211 a_35591_989.t8 a_39254_1735.t2 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X686 a_39582_17945.t3 a_40011_18575.t4 a_39717_18601.t3 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X687 a_58329_6179.t3 a_57739_6616.t8 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X688 a_30154_8749.t3 opcode[0].t35 VSS.t608 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X689 VDD.t59 a_37856_8106.t5 a_37916_8132.t0 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X690 VDD.t1575 a_34985_4186.t7 a_35575_3749.t3 VDD.t1574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X691 VDD.t672 a_15680_20866.t8 a_13401_n2178.t2 VDD.t671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X692 a_23081_8962.t1 a_24652_5324.t4 a_24240_5350.t4 VDD.t2576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X693 Y[5].t1 a_7464_n2148.t9 VDD.t1009 VDD.t1008 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X694 VSS.t258 A[3].t11 a_61452_20637.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X695 VDD.t686 opcode[1].t33 a_11155_10847.t2 VDD.t685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X696 VDD.t4224 a_48248_1040.t8 a_65651_n1230.t6 VDD.t4223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X697 a_22598_13724.t6 a_23777_13581.t4 a_23131_14454.t7 VDD.t2868 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X698 a_14310_5328.t2 A[5].t9 VDD.t2077 VDD.t2076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X699 a_13461_n2152.t1 a_13401_n2178.t5 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X700 VSS.t618 opcode[3].t9 a_280_n2152.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X701 a_19705_1744.t8 a_19396_11720.t5 VDD.t1269 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X702 VDD.t3582 a_57684_8194.t5 a_57739_6616.t5 VDD.t3581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X703 VDD.t2848 a_64122_11365.t5 a_70513_20044.t10 VDD.t2847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X704 VDD.t540 a_30645_3831.t14 a_62361_17053.t1 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X705 a_58326_1915.t2 a_57736_2352.t8 VDD.t3069 VDD.t3068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X706 a_53343_23888.t1 a_52753_24325.t7 VDD.t3650 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X707 a_10608_n2148.t5 a_9700_n2148.t6 a_10259_n2148.t4 VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X708 a_13711_14458.t7 a_14357_13585.t5 a_13178_13728.t3 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X709 a_4243_8992.t5 a_4183_8966.t9 a_3710_8262.t1 VDD.t4515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X710 a_39681_1042.t10 a_35575_3749.t6 VDD.t2706 VDD.t2705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X711 VDD.t2547 a_59937_9742.t5 a_60201_9159.t0 VDD.t2546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X712 a_57968_111.t1 a_54903_1041.t10 a_57731_748.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X713 a_62366_15449.t5 a_58326_16165.t7 VDD.t980 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X714 a_37916_8132.t1 a_37856_8106.t6 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X715 a_39952_20442.t1 A[0].t8 a_39715_21079.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X716 a_59223_16436.t4 a_30645_3831.t15 a_61120_15037.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X717 a_67135_3808.t0 a_64185_771.t4 VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X718 VDD.t79 a_6202_20866.t8 a_3923_n2178.t0 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 a_29952_5843.t11 B[3].t6 VDD.t2660 VDD.t2659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X720 a_19357_21596.t5 opcode[0].t36 VDD.t3866 VDD.t3865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X721 a_46818_20639.t2 a_46228_21076.t7 VDD.t3172 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X722 VDD.t2586 a_30645_10037.t14 a_46233_22680.t4 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X723 a_11133_n2633.t0 a_10576_1744.t8 VSS.t411 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X724 VDD.t2156 a_18824_20866.t9 a_16545_n2178.t1 VDD.t2155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X725 VDD.t2320 A[0].t9 a_24157_16385.t5 VDD.t2319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X726 VDD.t634 a_6832_13724.t9 a_6774_14454.t2 VDD.t633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X727 a_13778_1740.t5 a_14303_1255.t4 a_13429_1740.t9 VDD.t2686 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X728 a_45821_15761.t7 a_46176_16428.t12 VDD.t4507 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X729 VDD.t688 opcode[1].t34 a_70509_n1998.t8 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X730 a_59090_7603.t2 a_54713_3294.t6 VDD.t2401 VDD.t2400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X731 a_19987_14454.t2 opcode[0].t37 VDD.t3824 VDD.t3823 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X732 a_14367_8119.t3 opcode[0].t38 VSS.t535 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X733 VSS.t619 opcode[3].t10 a_3424_n2152.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X734 a_54567_3877.t5 a_51704_1914.t4 a_54449_3877.t2 VDD.t3596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X735 a_45050_6179.t2 a_44460_6616.t7 VDD.t1254 VDD.t1253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X736 a_10509_11720.t7 opcode[1].t35 VDD.t690 VDD.t689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X737 a_22598_10990.t3 a_23777_10847.t5 a_23131_11720.t7 VDD.t1766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 VDD.t281 A[4].t16 a_16213_21596.t8 VDD.t280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X739 a_61197_9746.t0 a_58334_7783.t4 a_61079_9746.t3 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X740 a_48418_21344.t0 A[1].t9 VDD.t1925 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X741 VDD.t3496 a_55469_11532.t6 a_57730_9870.t2 VDD.t3495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X742 a_10227_1744.t1 a_9918_11720.t5 VDD.t321 VDD.t320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X743 a_44445_4000.t2 a_42301_n1318.t9 VDD.t4089 VDD.t4088 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X744 VSS.t48 A[4].t17 a_7995_15753.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X745 VDD.t3619 a_41705_6822.t9 a_65649_10704.t9 VDD.t3618 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X746 VDD.t3014 A[6].t5 a_35001_1426.t2 VDD.t3013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X747 a_29950_1706.t2 B[5].t4 VDD.t4113 VDD.t4112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X748 VDD.t3890 opcode[3].t11 a_16046_n2152.t2 VDD.t3889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X749 a_40101_3874.t0 a_38493_311.t4 a_40219_3874.t2 VDD.t751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X750 a_6735_21596.t5 opcode[0].t39 VDD.t3338 VDD.t3337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X751 VDD.t4115 B[5].t5 a_13358_6047.t2 VDD.t4114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X752 a_50316_21344.t2 a_43319_23626.t8 VDD.t2570 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X753 a_43319_23626.t3 a_43055_24209.t7 VSS.t60 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 a_41493_21373.t4 a_41905_21347.t5 a_41611_21373.t5 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X755 VDD.t3365 a_30645_n306.t9 a_47719_15761.t11 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X756 a_70509_10624.t11 opcode[1].t36 VDD.t692 VDD.t691 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 VDD.t2928 opcode[2].t8 a_6524_1744.t2 VDD.t2927 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X758 a_807_1740.t8 opcode[2].t9 VDD.t2930 VDD.t2929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X759 VSS.t27 a_41507_3295.t7 a_45811_7603.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X760 a_49832_23623.t0 a_49568_24206.t5 VSS.t407 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X761 VDD.t1627 a_53312_9674.t6 a_53576_9091.t2 VDD.t1626 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X762 a_57981_7583.t0 a_57684_8194.t6 a_57744_8220.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X763 VDD.t3745 A[7].t7 a_9761_5354.t11 VDD.t3744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X764 VDD.t4561 a_59223_16436.t10 a_59280_15743.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X765 a_30647_7968.t4 a_30154_7310.t6 a_29954_7911.t5 VDD.t1422 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X766 a_70513_7304.t5 a_70459_8189.t5 a_71846_8013.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X767 a_7365_11720.t5 a_6774_14454.t4 a_6832_10990.t2 VDD.t1571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X768 VDD.t3822 opcode[0].t40 a_39720_22683.t2 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X769 a_3710_8262.t4 a_4889_8119.t4 a_4243_8992.t8 VDD.t3647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X770 a_16922_1740.t7 a_16014_1740.t4 a_16573_1740.t9 VDD.t3519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X771 VDD.t760 a_30645_5900.t15 a_59325_22679.t2 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X772 a_3710_8262.t5 a_4889_8119.t5 a_4834_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X773 a_40373_9071.t3 a_40109_9654.t5 VSS.t570 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X774 a_66005_5881.t0 a_64188_3841.t4 a_65769_6613.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X775 a_11155_10847.t1 opcode[1].t37 VDD.t694 VDD.t693 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X776 VDD.t479 a_13178_10994.t8 a_13120_11724.t0 VDD.t478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X777 a_62361_17053.t3 a_58326_16165.t8 a_63010_16442.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X778 a_51114_6548.t2 a_51059_8126.t8 VDD.t4291 VDD.t4290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X779 VSS.t302 a_46809_23893.t4 a_48426_24202.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X780 VDD.t3606 a_24157_16385.t7 a_23071_14428.t0 VDD.t3605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X781 a_14538_10391.t1 opcode[1].t38 a_13178_10994.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X782 VDD.t2858 a_53571_3290.t4 a_54567_3877.t2 VDD.t2857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X783 a_22172_5352.t7 a_22584_5326.t5 a_19937_8962.t3 VDD.t3150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X784 VDD.t3957 A[2].t8 a_54540_21365.t8 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X785 a_62361_17053.t0 a_30645_3831.t16 VDD.t2508 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X786 VSS.t652 a_44399_2324.t6 a_48484_308.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X787 a_20054_1744.t6 a_20579_1259.t4 a_19705_1744.t11 VDD.t4597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X788 a_16922_1740.t2 a_17447_1255.t5 a_16573_1740.t5 VDD.t3575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X789 a_59635_6910.t6 a_59090_7603.t4 a_59517_6910.t11 VDD.t4151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X790 VDD.t327 a_60201_9159.t5 a_61197_9746.t4 VDD.t326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X791 a_12478_20862.t2 A[3].t12 a_13011_21592.t4 VDD.t3283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X792 a_38493_311.t1 a_37903_748.t8 VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X793 a_41573_15739.t2 a_30643_n2374.t8 VDD.t3813 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X794 a_42301_n1318.t0 a_41711_n1755.t7 VDD.t2352 VDD.t2351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X795 VDD.t4441 a_48265_n1750.t7 a_48855_n1313.t3 VDD.t4440 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X796 a_41243_3878.t4 a_38498_1915.t4 VSS.t119 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X797 a_47417_18593.t2 a_47357_18567.t4 VDD.t1757 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X798 a_52674_17946.t3 a_53103_18576.t4 a_52809_18602.t2 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X799 a_48815_11511.t0 a_48225_11948.t7 VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X800 a_9761_5354.t5 B[7].t3 VDD.t1549 VDD.t1548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X801 a_47282_17937.t0 a_47357_18567.t5 VSS.t284 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X802 VDD.t213 a_35591_989.t9 a_39681_1042.t1 VDD.t212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X803 a_8011_13581.t2 opcode[0].t41 VDD.t1005 VDD.t1004 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X804 VDD.t4378 A[3].t13 a_63527_9231.t6 VDD.t4377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X805 VDD.t283 A[4].t18 a_15966_5352.t6 VDD.t282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X806 VSS.t368 A[0].t10 a_12672_15792.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X807 a_20578_10387.t1 a_19396_14454.t4 VSS.t384 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X808 VDD.t4450 a_6071_6357.t4 a_13721_8992.t9 VDD.t4449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X809 a_53312_9674.t1 a_51704_6111.t4 VSS.t522 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X810 VDD.t696 opcode[1].t39 a_19987_11720.t11 VDD.t695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X811 VDD.t1559 a_55469_11532.t7 a_59517_6910.t5 VDD.t1558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X812 a_60884_15037.t0 a_61178_15743.t4 a_59223_16436.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X813 VSS.t102 a_20611_n2633.t4 a_20558_n3481.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X814 VSS.t473 opcode[2].t10 a_248_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X815 VSS.t192 a_64117_5761.t6 a_66005_5881.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X816 a_18824_20866.t0 a_20003_20723.t4 a_19357_21596.t0 VDD.t353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X817 a_40310_22246.t2 a_39720_22683.t7 VDD.t3595 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X818 VDD.t3173 a_46228_21076.t8 a_46818_20639.t1 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_46823_22243.t2 a_46233_22680.t7 VDD.t876 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X820 VDD.t1927 A[1].t10 a_25633_21592.t5 VDD.t1926 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X821 a_59915_22242.t2 a_59325_22679.t7 VDD.t4200 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X822 a_39957_22046.t0 opcode[0].t42 a_39720_22683.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X823 a_16545_n2178.t0 a_18824_20866.t10 VDD.t2158 VDD.t2157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X824 a_6774_14454.t1 a_6832_13724.t10 VDD.t636 VDD.t635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X825 a_10459_8962.t5 a_15426_6045.t5 a_15966_5352.t3 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X826 a_71842_n1407.t0 a_39381_15765.t9 VSS.t100 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X827 VDD.t4547 a_51114_6548.t7 a_51704_6111.t2 VDD.t4546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X828 VDD.t903 a_48254_6910.t11 a_52465_7535.t1 VDD.t902 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X829 a_30154_8749.t2 opcode[0].t43 VDD.t4059 VDD.t4058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X830 a_71842_1973.t1 opcode[1].t40 a_70509_1028.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X831 a_59915_22242.t3 a_59325_22679.t8 VSS.t659 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X832 a_16213_21596.t7 A[4].t19 VDD.t285 VDD.t284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X833 a_16805_8966.t0 a_20515_5324.t4 a_20103_5350.t1 VDD.t1041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X834 a_46238_6910.t7 a_46650_6884.t6 a_46356_6910.t5 VDD.t331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X835 a_35004_7464.t3 B[3].t7 VDD.t2662 VDD.t2661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X836 a_7464_n2148.t3 opcode[3].t12 a_7700_n3481.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X837 a_16046_n2152.t1 opcode[3].t13 VDD.t3892 VDD.t3891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X838 VSS.t309 a_37848_2326.t7 a_38140_111.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X839 a_23198_1744.t3 a_23723_1259.t4 a_22849_1744.t5 VDD.t3101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X840 VDD.t4044 opcode[0].t44 a_6735_21596.t4 VDD.t4043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X841 a_59562_22042.t1 a_56366_23618.t6 a_59325_22679.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X842 a_56511_18089.t0 a_30643_1763.t8 VSS.t379 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X843 a_64185_771.t1 a_63595_1208.t8 VDD.t1793 VDD.t1792 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X844 a_16322_13728.t6 a_17501_13585.t4 a_16855_14458.t11 VDD.t1989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X845 a_53425_3873.t4 a_51699_310.t5 a_53307_3873.t3 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X846 a_70509_10506.t3 a_70455_11391.t4 a_71842_11215.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X847 a_56556_21365.t4 a_56011_22058.t4 a_56556_20633.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X848 a_60055_9742.t5 a_58329_6179.t4 a_59937_9742.t4 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X849 a_4857_n2637.t1 a_4300_1740.t9 VDD.t2131 VDD.t2130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X850 VDD.t2309 a_16322_13728.t8 a_16264_14458.t2 VDD.t2308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X851 a_30645_n306.t7 a_30152_475.t4 a_29952_n363.t11 VDD.t3370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X852 a_59280_15743.t0 a_59223_16436.t11 VDD.t4565 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X853 VDD.t531 a_22598_10990.t8 a_22540_11720.t2 VDD.t530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X854 VDD.t3119 a_40101_3874.t6 a_40365_3291.t1 VDD.t3118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X855 a_14538_13125.t1 opcode[0].t45 a_13178_13728.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X856 a_6832_10990.t1 a_6774_14454.t5 a_7365_11720.t4 VDD.t3567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X857 VSS.t464 a_53571_3290.t5 a_54449_3877.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X858 a_39720_22683.t1 opcode[0].t46 VDD.t1787 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X859 VDD.t4386 A[3].t14 a_61098_21369.t10 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X860 VDD.t1695 a_6813_6359.t5 a_16865_8992.t5 VDD.t1694 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X861 VSS.t55 a_60201_9159.t6 a_61079_9746.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X862 VDD.t3894 opcode[3].t14 a_19737_n2148.t11 VDD.t3893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X863 VDD.t1055 a_64188_3841.t5 a_67135_7303.t1 VDD.t1054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X864 a_59325_22679.t1 a_30645_5900.t16 VDD.t761 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X865 a_46922_9159.t3 a_46658_9742.t6 VSS.t179 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X866 VDD.t2419 B[3].t8 a_17495_6045.t1 VDD.t2418 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X867 a_44465_8220.t2 a_41507_3295.t8 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X868 a_59517_6910.t1 a_54713_3294.t7 VDD.t2403 VDD.t2402 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X869 VDD.t698 opcode[1].t41 a_8011_10847.t2 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X870 a_13120_11724.t1 a_13178_10994.t9 VDD.t481 VDD.t480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X871 a_54903_1041.t0 a_55197_1015.t5 a_54785_1041.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X872 VDD.t1098 a_5331_6357.t6 a_10519_8988.t8 VDD.t1097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X873 VDD.t4464 a_55504_n1325.t7 a_57722_4002.t2 VDD.t4463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X874 a_11101_1259.t1 a_70513_7304.t9 VDD.t2892 VDD.t2891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X875 VDD.t1961 a_56366_23618.t7 a_59320_21075.t6 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X876 a_48690_23619.t3 a_48426_24202.t5 VSS.t688 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X877 a_23071_14428.t1 a_24157_16385.t8 VDD.t3608 VDD.t3607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X878 VSS.t313 a_13130_8992.t6 a_14538_10391.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X879 VDD.t4239 a_63602_n1637.t7 a_64192_n2074.t3 VDD.t4238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X880 a_10576_1744.t2 a_9668_1744.t4 a_10227_1744.t5 VDD.t610 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X881 a_54540_21365.t7 A[2].t9 VDD.t3958 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X882 a_20633_13581.t2 opcode[0].t47 VDD.t1780 VDD.t1779 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X883 VDD.t2421 B[3].t9 a_35004_7464.t2 VDD.t2420 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X884 a_58868_15769.t9 a_58328_16462.t4 a_58986_15769.t5 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X885 a_70509_13768.t0 a_56556_21365.t8 a_70509_13650.t0 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X886 a_17479_n2637.t3 a_16922_1740.t8 VSS.t17 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X887 a_66063_6587.t3 a_64117_5761.t7 VSS.t193 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X888 a_54790_6842.t2 a_55202_6816.t4 a_54908_6842.t4 VDD.t786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X889 a_13011_21592.t3 A[3].t15 a_12478_20862.t1 VDD.t4385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X890 a_41587_6822.t7 a_39807_6822.t8 VDD.t3225 VDD.t3224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X891 VDD.t2354 a_41711_n1755.t8 a_42301_n1318.t1 VDD.t2353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X892 VDD.t2079 A[5].t10 a_4593_6357.t2 VDD.t2078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X893 a_39807_6822.t7 a_40101_6796.t5 a_39689_6822.t11 VDD.t4281 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X894 VDD.t1758 a_47357_18567.t6 a_47417_18593.t1 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X895 a_7365_14454.t2 a_6887_15819.t4 VDD.t3373 VDD.t3372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X896 a_30152_10818.t1 opcode[0].t48 VDD.t3919 VDD.t3918 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X897 VSS.t310 a_37848_2326.t8 a_41933_310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X898 a_46650_6884.t1 a_42266_11512.t7 VSS.t604 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X899 a_18389_4620.t1 B[3].t10 VSS.t383 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X900 a_52809_18602.t1 a_53103_18576.t5 a_52674_17946.t0 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X901 a_7315_8962.t5 a_13358_6047.t4 a_13898_5354.t10 VDD.t3635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X902 a_65769_2386.t0 a_66063_3092.t4 VSS.t90 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X903 a_51109_747.t6 a_48064_9163.t6 VDD.t976 VDD.t975 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X904 VSS.t158 a_42770_18699.t8 a_40799_18571.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X905 VDD.t223 a_49319_15441.t7 a_47711_18567.t2 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X906 VDD.t2108 a_37911_6528.t7 a_38501_6091.t0 VDD.t2107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X907 a_19454_10990.t0 a_20633_10847.t4 a_20578_10387.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X908 a_65649_10704.t11 a_66061_10678.t4 a_65767_10704.t7 VDD.t2864 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X909 VDD.t771 a_48064_9163.t7 a_51100_4001.t2 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X910 a_19987_11720.t10 opcode[1].t42 VDD.t700 VDD.t699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X911 a_52887_1041.t9 a_53299_1015.t4 a_53005_1041.t5 VDD.t4471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X912 a_10227_1744.t11 a_11101_1259.t5 a_10576_1744.t7 VDD.t788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X913 a_39943_23696.t1 A[0].t11 a_39706_24333.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X914 a_61216_21369.t2 a_60671_22062.t4 a_61098_21369.t2 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X915 a_63024_18092.t0 a_30645_3831.t17 VSS.t399 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X916 VDD.t2932 opcode[2].t11 a_7083_1744.t5 VDD.t2931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X917 a_37856_8106.t2 a_67135_7303.t7 VDD.t600 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X918 VDD.t4466 a_55504_n1325.t8 a_59082_1735.t2 VDD.t4465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X919 a_19357_21596.t1 a_20003_20723.t5 a_18824_20866.t1 VDD.t354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X920 a_40305_20642.t2 a_39715_21079.t7 VDD.t3349 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X921 a_23131_11720.t9 a_22540_14454.t4 a_22598_10990.t5 VDD.t4584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X922 a_51105_9802.t5 a_48815_11511.t7 VDD.t2267 VDD.t2266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X923 VDD.t1641 a_57676_2326.t5 a_61407_1042.t0 VDD.t1640 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X924 a_70513_4278.t1 a_52473_15766.t9 a_70513_4160.t1 VDD.t663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X925 VDD.t3697 a_39720_22683.t8 a_40310_22246.t1 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X926 a_63769_11165.t1 B[3].t11 a_63532_11802.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X927 a_59901_23892.t3 a_59311_24329.t7 VSS.t169 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X928 a_25633_21592.t4 A[1].t11 VDD.t1929 VDD.t1928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X929 VDD.t1606 a_61525_1042.t8 a_70513_4278.t3 VDD.t1605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X930 a_53010_6842.t5 a_52465_7535.t5 a_52892_6842.t11 VDD.t3695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X931 a_29952_9980.t7 a_30152_9379.t5 a_30645_10037.t1 VDD.t2151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X932 a_14303_1255.t0 a_70509_10506.t8 VDD.t2338 VDD.t2337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X933 a_7365_11720.t11 opcode[1].t43 VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X934 VDD.t3415 a_46922_9159.t5 a_47918_9746.t4 VDD.t3414 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X935 VDD.t287 A[4].t20 a_16213_21596.t6 VDD.t286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X936 a_59910_20638.t0 a_59320_21075.t7 VDD.t2525 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X937 a_13898_5354.t11 a_13358_6047.t5 a_7315_8962.t6 VDD.t3636 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X938 a_23958_13121.t0 opcode[0].t49 a_22598_13724.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X939 a_65767_10704.t0 a_65222_11397.t4 a_65767_9972.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X940 VSS.t490 a_70509_n2116.t9 a_1681_1255.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X941 a_7936_n3481.t0 a_6556_n2148.t4 a_7464_n2148.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X942 Cout.t2 a_39582_17945.t5 VDD.t614 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X943 a_71846_17727.t0 opcode[1].t44 a_70513_16782.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X944 VDD.t3896 opcode[3].t15 a_16046_n2152.t0 VDD.t3895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X945 VSS.t474 opcode[2].t12 a_16014_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X946 VSS.t40 a_44405_8194.t8 a_44697_5979.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X947 a_52753_24325.t3 A[2].t10 VDD.t3959 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X948 a_6735_21596.t3 opcode[0].t50 VDD.t1736 VDD.t1735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X949 VSS.t130 a_30645_5900.t17 a_59562_22042.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X950 VDD.t4475 a_12732_15818.t4 a_23131_14454.t9 VDD.t4474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X951 a_56792_20633.t0 a_54658_21365.t10 a_56556_21365.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X952 a_13461_n2152.t11 a_12902_n2152.t4 a_13810_n2152.t3 VDD.t4489 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X953 a_59509_1042.t11 a_54903_1041.t11 VDD.t1021 VDD.t1020 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X954 a_16264_14458.t1 a_16322_13728.t9 VDD.t2311 VDD.t2310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X955 a_49314_17045.t6 a_30645_n306.t10 VDD.t3366 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X956 VDD.t1067 a_51059_8126.t9 a_51119_8152.t2 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X957 a_16954_n2152.t2 a_17479_n2637.t4 a_16605_n2152.t2 VDD.t4240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X958 VDD.t2934 opcode[2].t13 a_12870_1740.t2 VDD.t2933 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X959 a_19357_21596.t4 opcode[0].t51 VDD.t1768 VDD.t1767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X960 VSS.t550 a_9228_15824.t4 a_14538_13125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X961 a_7365_11720.t3 a_6774_14454.t6 a_6832_10990.t0 VDD.t2870 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X962 VDD.t4091 a_42301_n1318.t10 a_46232_1040.t5 VDD.t4090 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X963 VDD.t762 a_30645_5900.t18 a_59325_22679.t0 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X964 VSS.t115 a_55469_11532.t8 a_59871_6178.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X965 a_13711_14458.t2 a_9228_15824.t5 VDD.t3420 VDD.t3419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X966 VDD.t4573 a_54908_6842.t11 a_66063_3092.t2 VDD.t4572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X967 a_16954_n2152.t3 opcode[3].t16 a_17190_n3485.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X968 a_8011_10847.t1 opcode[1].t45 VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X969 VDD.t2112 a_63532_11802.t7 a_64122_11365.t2 VDD.t2111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X970 VDD.t4226 a_48248_1040.t9 a_67135_n540.t2 VDD.t4225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X971 a_23230_n2148.t2 a_23755_n2633.t4 a_22881_n2148.t2 VDD.t4480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X972 a_70509_1028.t5 a_70455_1913.t5 a_70509_1146.t8 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X973 a_70513_7422.t1 a_58986_15769.t8 a_70513_7304.t1 VDD.t1113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X974 a_59320_21075.t5 a_56366_23618.t8 VDD.t1962 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X975 a_18824_20866.t2 a_20003_20723.t6 a_19948_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X976 VDD.t3960 A[2].t11 a_54540_21365.t6 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X977 VDD.t3610 a_24157_16385.t9 a_23071_14428.t2 VDD.t3609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X978 a_64192_n2074.t0 a_63602_n1637.t8 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X979 VDD.t3803 opcode[0].t52 a_29954_7911.t3 VDD.t3802 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X980 a_29952_5843.t9 a_30152_5242.t5 a_30645_5900.t2 VDD.t2515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X981 a_58986_15769.t6 a_58328_16462.t5 a_58868_15769.t10 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X982 a_46275_18597.t4 a_46215_18571.t4 VDD.t607 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X983 a_42301_n1318.t2 a_41711_n1755.t9 VDD.t2356 VDD.t2355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X984 a_41579_1042.t2 a_39799_1042.t9 VDD.t1754 VDD.t1753 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X985 VDD.t2423 B[3].t12 a_63527_6198.t4 VDD.t2422 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X986 VSS.t362 a_48815_11511.t8 a_53246_6110.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X987 a_47417_18593.t0 a_47357_18567.t7 VDD.t1759 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X988 VDD.t3375 a_6887_15819.t5 a_7365_14454.t1 VDD.t3374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X989 a_61178_15743.t2 a_30645_3831.t18 VDD.t2509 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X990 a_17447_1255.t2 a_70509_13650.t8 VDD.t1036 VDD.t1035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X991 a_4183_8966.t0 a_11289_6045.t5 a_11829_5352.t8 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X992 a_43405_16438.t0 a_30643_n2374.t9 VSS.t605 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X993 VDD.t4588 a_61071_3878.t5 a_57684_8194.t1 VDD.t4587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X994 a_47711_18567.t1 a_49319_15441.t8 VDD.t224 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X995 a_20814_10387.t1 opcode[1].t46 a_19454_10990.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X996 a_52767_15740.t2 a_52710_16433.t10 VDD.t1374 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X997 a_19454_10990.t1 a_20633_10847.t5 a_19987_11720.t3 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X998 VDD.t1721 a_16332_8262.t9 a_16274_8992.t0 VDD.t1720 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X999 a_24240_5350.t3 B[0].t8 VDD.t2205 VDD.t2204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1000 a_29952_9980.t1 B[1].t4 VDD.t4143 VDD.t4142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1001 a_45049_1913.t2 a_44459_2350.t7 VDD.t3529 VDD.t3528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1002 a_54540_21365.t10 a_54952_21339.t5 a_54658_21365.t6 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1003 a_52892_6842.t5 a_48815_11511.t9 VDD.t2269 VDD.t2268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1004 a_61098_21369.t1 a_60671_22062.t5 a_61216_21369.t1 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1005 VDD.t3856 opcode[0].t53 a_29952_3774.t7 VDD.t3855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1006 a_30645_5900.t7 a_30152_6681.t5 a_29952_5843.t5 VDD.t3287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1007 a_18824_20866.t3 a_20003_20723.t7 a_19357_21596.t2 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1008 a_23141_8988.t10 a_23081_8962.t9 a_22608_8258.t6 VDD.t293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1009 a_42761_15445.t3 A[7].t8 a_43410_14834.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1010 VSS.t257 A[3].t16 a_63769_11165.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1011 VDD.t2936 opcode[2].t14 a_16014_1740.t1 VDD.t2935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1012 a_30645_3831.t2 a_30152_3173.t5 a_29952_3774.t4 VDD.t1133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1013 a_61525_1042.t4 a_60980_1735.t5 a_61407_1042.t7 VDD.t2841 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1014 a_48690_23619.t0 a_48426_24202.t6 VDD.t416 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1015 a_16855_14458.t0 a_10397_15824.t4 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1016 VSS.t216 B[6].t7 a_11289_6045.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1017 VDD.t2404 a_30643_1763.t9 a_54665_15740.t1 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1018 VDD.t399 a_16322_10994.t8 a_16264_11724.t2 VDD.t398 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1019 a_51059_8126.t2 a_67135_n540.t9 VDD.t2998 VDD.t2997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1020 a_16855_14458.t6 a_16795_14432.t4 a_16322_13728.t1 VDD.t1986 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1021 VSS.t691 a_6071_6357.t5 a_14548_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1022 a_7956_10387.t0 a_6774_14454.t7 VSS.t345 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1023 a_48248_1040.t0 a_47703_1733.t4 a_48130_1040.t0 VDD.t3405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1024 VDD.t706 opcode[1].t47 a_7365_11720.t10 VDD.t705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1025 VSS.t398 a_55862_18700.t7 a_53891_18572.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1026 a_41913_11312.t0 B[4].t4 a_41676_11949.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1027 a_1099_8992.t7 a_1745_8119.t5 a_566_8262.t5 VDD.t649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1028 VDD.t215 a_35591_989.t10 a_39254_1735.t1 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1029 a_61827_6884.t3 a_57684_8194.t7 VSS.t568 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1030 a_3591_21596.t6 A[6].t6 a_3058_20866.t3 VDD.t3015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1031 VDD.t4301 a_18243_16385.t7 a_10449_14428.t2 VDD.t4300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1032 a_38492_9345.t2 a_37902_9782.t7 VDD.t3340 VDD.t3339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1033 VSS.t508 a_7989_n2633.t4 a_7936_n3481.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1034 a_38723_16458.t2 a_38721_16161.t8 VDD.t3540 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1035 a_19406_8988.t2 a_19464_8258.t8 VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1036 VSS.t548 a_4825_1255.t4 a_4772_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1037 a_41243_3878.t1 a_38498_1915.t5 a_41361_3878.t5 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1038 a_30645_n306.t1 a_30152_n964.t6 a_29952_n363.t4 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1039 VDD.t1734 opcode[0].t54 a_16865_8992.t7 VDD.t1733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1040 a_23131_14454.t10 a_12732_15818.t5 VDD.t4477 VDD.t4476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1041 VDD.t4228 a_48248_1040.t10 a_65651_n1230.t5 VDD.t4227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1042 VDD.t3898 opcode[3].t17 a_13461_n2152.t7 VDD.t3897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1043 a_44460_6616.t1 a_42266_11512.t8 VDD.t3793 VDD.t3792 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1044 VSS.t164 a_49832_23623.t6 a_56792_20633.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1045 a_4237_20723.t2 opcode[0].t55 VDD.t1011 VDD.t1010 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1046 a_11155_10847.t3 opcode[1].t48 VSS.t124 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1047 a_53312_9674.t2 a_51704_6111.t5 a_53430_9674.t1 VDD.t3240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1048 VDD.t3016 A[6].t7 a_49319_15441.t2 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1049 VDD.t4468 a_55504_n1325.t9 a_59509_1042.t8 VDD.t4467 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1050 a_65651_6613.t5 a_64188_3841.t6 VDD.t1057 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1051 VDD.t3584 a_57684_8194.t8 a_57739_6616.t6 VDD.t3583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1052 a_38492_9345.t3 a_37902_9782.t8 VSS.t537 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1053 a_63598_4278.t3 B[4].t5 VDD.t927 VDD.t926 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1054 a_59915_22242.t1 a_59325_22679.t9 VDD.t4201 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1055 a_16855_11724.t8 opcode[1].t49 VDD.t708 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1056 VDD.t3422 a_9228_15824.t6 a_13711_14458.t1 VDD.t3421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1057 VSS.t49 A[4].t21 a_41948_n1318.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1058 a_17426_n3485.t1 a_16046_n2152.t4 a_16954_n2152.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1059 VSS.t38 a_49319_15441.t9 a_47711_18567.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1060 a_31379_7968.t0 a_30154_8749.t4 a_30647_7968.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1061 VSS.t122 a_15680_20866.t9 a_13401_n2178.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1062 a_1690_7659.t0 a_1039_8966.t8 VSS.t86 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1063 a_18035_5352.t5 A[3].t17 VDD.t4384 VDD.t4383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1064 a_41493_21373.t5 a_41905_21347.t6 a_41611_21373.t6 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1065 a_50316_21344.t1 a_43319_23626.t9 VDD.t2571 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1066 VSS.t151 B[4].t6 a_30152_3173.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1067 a_29952_9980.t5 opcode[0].t56 VDD.t2881 VDD.t2880 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1068 a_22881_n2148.t1 a_23755_n2633.t5 a_23230_n2148.t1 VDD.t4481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1069 VDD.t1963 a_56366_23618.t9 a_59320_21075.t4 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1070 a_45050_6179.t3 a_44460_6616.t8 VSS.t200 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1071 a_20184_20263.t0 opcode[0].t57 a_18824_20866.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1072 VSS.t147 a_48254_6910.t12 a_51342_9165.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1073 a_39263_15765.t5 a_39675_15739.t4 a_39381_15765.t1 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1074 a_58868_15769.t5 a_59280_15743.t5 a_58986_15769.t3 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1075 VDD.t1373 a_19763_16387.t7 a_13651_14432.t2 VDD.t1372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1076 VDD.t2587 a_30645_10037.t15 a_46219_24330.t6 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1077 VDD.t608 a_46215_18571.t5 a_46275_18597.t3 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1078 a_9228_15824.t2 a_9168_15798.t6 VDD.t221 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1079 a_16855_11724.t1 a_16264_14458.t4 a_16322_10994.t7 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1080 VDD.t1390 B[6].t8 a_15297_16387.t2 VDD.t1389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1081 VDD.t2510 a_30645_3831.t19 a_61178_15743.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1082 a_41361_3878.t2 a_40365_3291.t4 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1083 a_61636_24201.t1 a_59901_23892.t5 VDD.t497 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1084 a_22709_16385.t2 B[1].t5 VDD.t4145 VDD.t4144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1085 a_18035_5352.t0 a_17495_6045.t4 a_13661_8966.t0 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1086 a_42756_17049.t6 a_38721_16161.t9 a_43405_16438.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1087 a_51054_2325.t0 a_54454_9678.t5 VDD.t4195 VDD.t4194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1088 a_59517_6910.t8 a_59929_6884.t5 a_59635_6910.t0 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1089 VDD.t225 a_49319_15441.t10 a_47711_18567.t0 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1090 VSS.t116 a_62375_18703.t7 a_60404_18575.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1091 VSS.t7 a_19406_8988.t4 a_20814_10387.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1092 a_13778_1740.t6 a_14303_1255.t5 a_13429_1740.t10 VDD.t2687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1093 a_19987_11720.t4 a_20633_10847.t6 a_19454_10990.t2 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1094 a_54454_9678.t4 a_51709_7715.t4 VSS.t267 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1095 a_70509_n2116.t6 a_70455_n1231.t4 a_70509_n1998.t11 VDD.t4131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1096 a_58326_1915.t1 a_57736_2352.t9 VDD.t3071 VDD.t3070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1097 a_31379_12105.t0 a_30154_12886.t5 a_30647_12105.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1098 a_70513_4278.t6 a_70459_5045.t5 a_70513_4160.t5 VDD.t1958 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1099 a_70513_19926.t0 a_70459_20811.t4 a_70513_20044.t0 VDD.t655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1100 a_41999_6796.t2 a_37856_8106.t7 VDD.t2250 VDD.t2249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1101 VDD.t3018 A[6].t8 a_3855_6357.t2 VDD.t3017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1102 VDD.t4382 A[3].t18 a_63598_4278.t5 VDD.t4381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1103 VDD.t2588 a_30645_10037.t16 a_47579_22063.t2 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1104 a_61216_21369.t0 a_60671_22062.t6 a_61098_21369.t0 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1105 VSS.t274 a_40296_23896.t4 a_41913_24205.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1106 a_7326_20263.t1 A[5].t11 VSS.t329 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1107 VDD.t2081 A[5].t12 a_16795_16385.t6 VDD.t2080 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1108 VDD.t2100 a_59929_3874.t6 a_60193_3291.t2 VDD.t2099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1109 VDD.t3900 opcode[3].t18 a_22881_n2148.t7 VDD.t3899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1110 VDD.t2938 opcode[2].t15 a_13429_1740.t4 VDD.t2937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1111 a_19146_1744.t2 opcode[2].t16 VDD.t2940 VDD.t2939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1112 a_30150_2544.t3 opcode[0].t58 VSS.t555 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1113 VDD.t445 a_10397_15824.t5 a_16855_14458.t1 VDD.t444 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1114 a_31375_1999.t0 B[5].t6 VSS.t288 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1115 a_46650_6884.t2 a_42266_11512.t9 VDD.t3795 VDD.t3794 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1116 a_37908_2352.t5 a_37848_2326.t9 VDD.t1940 VDD.t1939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1117 VSS.t84 a_13178_10994.t10 a_13120_11724.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1118 a_65767_10704.t1 a_65222_11397.t5 a_65649_10704.t5 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1119 a_60201_9159.t1 a_59937_9742.t6 VSS.t410 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1120 a_41160_7515.t2 a_39807_6822.t9 VDD.t3227 VDD.t3226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1121 a_51114_2351.t6 a_48855_n1313.t7 VDD.t1231 VDD.t1230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1122 a_58328_16462.t2 a_58326_16165.t9 VDD.t981 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1123 a_56497_16439.t0 a_30643_1763.t10 VSS.t380 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1124 a_11048_411.t0 a_9668_1744.t5 a_10576_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1125 a_19705_1744.t2 opcode[2].t17 VDD.t2942 VDD.t2941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1126 VSS.t487 A[6].t9 a_41913_11312.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1127 a_3710_8262.t6 a_4889_8119.t6 a_4243_8992.t9 VDD.t3648 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1128 a_10449_14428.t1 a_18243_16385.t8 VDD.t4303 VDD.t4302 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1129 a_19763_16387.t1 A[3].t19 VDD.t4380 VDD.t4379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1130 a_1089_11724.t0 a_498_14458.t4 a_556_10994.t0 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1131 a_9867_21592.t1 A[6].t10 VDD.t3020 VDD.t3019 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1132 VSS.t527 a_45279_16157.t10 a_45281_16454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1133 a_13461_n2152.t6 opcode[3].t19 VDD.t3902 VDD.t3901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1134 a_3855_6357.t1 A[6].t11 VDD.t3022 VDD.t3021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1135 Y[0].t2 a_23230_n2148.t8 VDD.t4212 VDD.t4211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1136 a_17394_407.t1 a_16014_1740.t5 a_16922_1740.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1137 a_14016_4622.t1 a_14310_5328.t4 a_7315_8962.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1138 VDD.t2879 opcode[0].t59 a_4237_20723.t1 VDD.t2878 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1139 a_49319_15441.t1 A[6].t12 VDD.t3023 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1140 a_1039_8966.t0 a_10173_5328.t4 a_9761_5354.t0 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1141 VDD.t3025 A[6].t13 a_35001_1426.t1 VDD.t3024 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1142 VDD.t4018 a_38484_3565.t4 a_40219_3874.t5 VDD.t4017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1143 VDD.t295 a_3923_n2178.t5 a_3983_n2152.t0 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1144 VDD.t710 opcode[1].t50 a_16855_11724.t7 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1145 a_63595_1208.t5 A[4].t22 VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1146 VSS.t666 a_17479_n2637.t5 a_17426_n3485.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1147 a_65651_3118.t0 a_64185_771.t5 VDD.t361 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1148 a_41507_3295.t1 a_41243_3878.t5 VSS.t655 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1149 a_20103_5350.t11 B[2].t2 VDD.t3727 VDD.t3726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1150 VDD.t2572 a_43319_23626.t10 a_50316_21344.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1151 a_13178_10994.t2 a_14357_10851.t4 a_13711_11724.t6 VDD.t2674 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1152 a_7375_8988.t11 a_8021_8115.t4 a_6842_8258.t7 VDD.t4293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1153 a_9761_5354.t4 B[7].t4 VDD.t1551 VDD.t1550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1154 a_23230_n2148.t0 a_23755_n2633.t6 a_22881_n2148.t0 VDD.t4482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1155 VDD.t3578 a_51114_2351.t7 a_51704_1914.t2 VDD.t3577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1156 VDD.t2944 opcode[2].t18 a_16573_1740.t8 VDD.t2943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1157 VSS.t388 B[1].t6 a_21632_6045.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1158 VSS.t591 a_35594_7027.t5 a_39262_7515.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1159 VSS.t256 A[3].t20 a_20184_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1160 a_10472_16406.t2 B[2].t3 VDD.t3729 VDD.t3728 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1161 a_70509_1146.t10 opcode[1].t51 VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1162 a_41705_6822.t4 a_41160_7515.t4 a_41587_6822.t9 VDD.t3611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1163 a_41579_1042.t10 a_41991_1016.t6 a_41697_1042.t0 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1164 a_48426_24202.t2 a_46818_20639.t4 a_48544_24202.t2 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1165 a_30154_7310.t3 B[2].t4 VDD.t3731 VDD.t3730 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1166 a_46809_23893.t2 a_46219_24330.t8 VDD.t2637 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1167 a_46275_18597.t2 a_46215_18571.t6 VDD.t609 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1168 a_15297_16387.t1 B[6].t9 VDD.t1392 VDD.t1391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1169 a_29952_9980.t11 a_30152_10818.t5 a_30645_10037.t3 VDD.t3833 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1170 a_61178_15743.t0 a_30645_3831.t20 VDD.t2511 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1171 VDD.t2715 a_59901_23892.t6 a_61636_24201.t2 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1172 VDD.t2455 B[1].t7 a_22709_16385.t1 VDD.t2454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1173 VSS.t330 A[5].t13 a_35241_6827.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1174 a_22849_1744.t2 opcode[2].t19 VDD.t2946 VDD.t2945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1175 VDD.t961 a_42770_18699.t9 a_40799_18571.t1 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1176 a_57730_9870.t5 a_54713_3294.t8 VDD.t4519 VDD.t4518 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1177 VDD.t4093 a_42301_n1318.t11 a_45805_1733.t2 VDD.t4092 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1178 VDD.t2852 a_44445_4000.t7 a_45035_3563.t2 VDD.t2851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1179 a_22172_5352.t8 a_22584_5326.t6 a_19937_8962.t4 VDD.t3175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1180 a_49319_15441.t6 a_45279_16157.t11 VDD.t3295 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1181 a_70509_n1998.t10 a_70455_n1231.t5 a_70509_n2116.t5 VDD.t4132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1182 a_13849_16387.t1 B[7].t5 VDD.t2598 VDD.t2597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1183 a_19454_10990.t3 a_20633_10847.t7 a_19987_11720.t5 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1184 a_48502_n1313.t0 B[5].t7 a_48265_n1750.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1185 a_7115_n2148.t9 a_6556_n2148.t5 a_7464_n2148.t5 VDD.t4178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1186 a_59635_6910.t3 a_59090_7603.t5 a_59517_6910.t9 VDD.t3653 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1187 VSS.t81 a_13178_13728.t8 a_13120_14458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1188 a_10459_8962.t1 a_16378_5326.t4 a_15966_5352.t8 VDD.t1953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1189 VDD.t2643 a_46356_6910.t8 a_48136_6910.t6 VDD.t2642 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1190 a_29950_n2431.t2 B[7].t6 VDD.t2600 VDD.t2599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1191 a_1713_n2637.t2 a_1156_1740.t8 VDD.t2126 VDD.t2125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1192 VDD.t1599 opcode[0].t60 a_7381_20723.t1 VDD.t1598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1193 a_6202_20866.t3 a_7381_20723.t4 a_7326_20263.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1194 a_47579_22063.t1 a_30645_10037.t17 VDD.t2589 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1195 VDD.t3904 opcode[3].t20 a_12902_n2152.t2 VDD.t3903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1196 a_29952_5843.t3 opcode[0].t61 VDD.t1800 VDD.t1799 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1197 VDD.t1812 B[5].t8 a_63527_9231.t2 VDD.t1811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1198 a_48855_n1313.t0 a_48265_n1750.t8 VDD.t420 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1199 a_9867_21592.t4 opcode[0].t62 VDD.t1802 VDD.t1801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1200 VDD.t4354 a_35012_10049.t8 a_35602_9612.t1 VDD.t4353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1201 a_8130_16410.t2 B[4].t7 VDD.t929 VDD.t928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1202 a_54879_11969.t6 A[6].t14 VDD.t3027 VDD.t3026 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1203 a_13810_n2152.t7 a_14335_n2637.t4 a_13461_n2152.t10 VDD.t4247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1204 a_53425_3873.t2 a_51690_3564.t5 VDD.t2664 VDD.t2663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1205 a_65649_10704.t6 a_65222_11397.t6 a_65767_10704.t2 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1206 a_71846_8249.t0 opcode[1].t52 a_70513_7304.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1207 a_60055_9742.t2 a_58320_9433.t4 VDD.t2990 VDD.t2989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1208 VDD.t982 a_58326_16165.t10 a_58328_16462.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1209 VDD.t1902 a_70513_4160.t10 a_7957_1259.t1 VDD.t1901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1210 a_55848_17050.t3 a_51813_16162.t5 a_56497_16439.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1211 VDD.t3586 a_57684_8194.t9 a_57744_8220.t6 VDD.t3585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1212 VDD.t2481 a_12478_20862.t8 a_10199_n2174.t2 VDD.t2480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1213 a_23755_n2633.t2 a_23198_1744.t8 VDD.t2545 VDD.t2544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1214 VDD.t3324 a_70513_16782.t9 a_20579_1259.t1 VDD.t3323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1215 a_29950_1706.t10 a_30150_2544.t6 a_30643_1763.t6 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1216 a_556_10994.t1 a_498_14458.t5 a_1089_11724.t1 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1217 a_4300_1740.t5 a_4825_1255.t5 a_3951_1740.t9 VDD.t3402 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1218 VDD.t3029 A[6].t15 a_9867_21592.t0 VDD.t3028 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1219 VDD.t3954 a_16795_16385.t8 a_7305_14428.t1 VDD.t3953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1220 VDD.t3906 opcode[3].t21 a_3424_n2152.t1 VDD.t3905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1221 VSS.t34 a_35591_989.t11 a_38131_3365.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1222 VDD.t3738 a_61782_23618.t4 a_62778_24205.t5 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1223 VSS.t479 a_53343_23888.t5 a_54960_24197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1224 VDD.t3030 A[6].t16 a_49319_15441.t0 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1225 VDD.t1426 a_57722_4002.t8 a_58312_3565.t2 VDD.t1425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1226 a_55197_1015.t2 a_51054_2325.t10 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1227 a_39799_1042.t6 a_40093_1016.t4 a_39681_1042.t5 VDD.t4503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1228 VDD.t2948 opcode[2].t20 a_10227_1744.t7 VDD.t2947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1229 a_56438_21365.t2 a_54658_21365.t11 VDD.t880 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1230 a_49328_18695.t3 A[6].t17 a_49977_18084.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1231 VDD.t2083 A[5].t14 a_35004_7464.t6 VDD.t2082 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1232 VSS.t713 a_41611_21373.t9 a_42964_22066.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1233 a_3642_14458.t1 a_3700_13728.t9 VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1234 a_54790_6842.t1 a_55202_6816.t5 a_54908_6842.t5 VDD.t787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1235 a_61827_6884.t2 a_57684_8194.t10 VDD.t2810 VDD.t2809 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1236 a_41587_6822.t8 a_39807_6822.t10 VDD.t3229 VDD.t3228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1237 VDD.t2085 A[5].t15 a_4593_6357.t1 VDD.t2084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1238 a_13011_21592.t2 opcode[0].t63 VDD.t1340 VDD.t1339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1239 VDD.t34 a_19406_8988.t5 a_19987_11720.t0 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1240 VDD.t3746 A[7].t9 a_40621_16458.t2 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1241 VDD.t3733 B[2].t5 a_10472_16406.t1 VDD.t3732 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1242 a_4243_8992.t0 a_3855_6357.t4 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1243 a_16954_n2152.t1 a_17479_n2637.t6 a_16605_n2152.t1 VDD.t4241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1244 a_46238_6910.t11 a_41507_3295.t9 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1245 a_42031_24205.t2 a_40305_20642.t4 a_41913_24205.t3 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1246 a_48544_24202.t1 a_46818_20639.t5 a_48426_24202.t1 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1247 VSS.t395 a_22598_13724.t8 a_22540_14454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1248 a_44459_2350.t2 a_44399_2324.t7 VDD.t4153 VDD.t4152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1249 VDD.t2638 a_46219_24330.t9 a_46809_23893.t1 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1250 a_56556_21365.t2 a_56011_22058.t5 a_56438_21365.t5 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1251 a_4889_8119.t3 opcode[0].t64 VSS.t640 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1252 Y[7].t3 a_1188_n2152.t8 VSS.t242 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1253 a_55078_24197.t3 a_53352_20634.t4 a_54960_24197.t1 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1254 VSS.t347 a_21956_20862.t8 a_19677_n2174.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1255 VDD.t4470 a_55504_n1325.t10 a_59082_1735.t3 VDD.t4469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1256 VDD.t4155 a_44399_2324.t8 a_44454_746.t1 VDD.t4154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1257 a_6735_21596.t8 A[5].t16 a_6202_20866.t7 VDD.t2086 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1258 a_42770_18699.t5 a_30643_n2374.t10 VDD.t3869 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1259 VSS.t530 a_61343_9163.t5 a_71842_n1171.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1260 VDD.t3296 a_45279_16157.t12 a_49319_15441.t5 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1261 a_7464_n2148.t6 a_6556_n2148.t6 a_7115_n2148.t10 VDD.t4179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1262 a_48130_1040.t3 a_44399_2324.t9 VDD.t4157 VDD.t4156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1263 a_61071_3878.t3 a_58326_1915.t4 a_61189_3878.t0 VDD.t3074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1264 VDD.t3748 A[7].t10 a_13849_16387.t5 VDD.t3747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1265 VSS.t488 A[6].t18 a_48502_n1313.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1266 VDD.t2602 B[7].t7 a_30150_n3032.t2 VDD.t2601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1267 a_11640_16408.t3 A[1].t12 a_11505_15751.t1 VDD.t1930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1268 VDD.t4042 opcode[0].t65 a_19997_8988.t2 VDD.t4041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1269 VDD.t4307 opcode[3].t22 a_16605_n2152.t5 VDD.t4306 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1270 VSS.t148 a_48254_6910.t13 a_51356_7515.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1271 VSS.t475 opcode[2].t21 a_12870_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1272 a_7381_20723.t0 opcode[0].t66 VDD.t3938 VDD.t3937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1273 VDD.t2590 a_30645_10037.t18 a_47579_22063.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1274 a_58986_15769.t7 a_58328_16462.t6 a_58868_15769.t11 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1275 a_13130_8992.t0 a_13188_8262.t8 VDD.t2677 VDD.t2676 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1276 VDD.t2252 a_37856_8106.t8 a_41587_6822.t2 VDD.t2251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1277 a_70513_20044.t7 opcode[1].t53 VDD.t714 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1278 VDD.t3417 a_46922_9159.t6 a_47918_9746.t5 VDD.t3416 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1279 a_35602_9612.t0 a_35012_10049.t9 VDD.t4356 VDD.t4355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1280 VDD.t2444 a_22709_16385.t8 a_19927_14428.t0 VDD.t2443 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1281 a_59223_16436.t5 a_60226_16462.t4 a_60766_15769.t9 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1282 a_20633_13581.t3 opcode[0].t67 VSS.t622 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1283 a_15297_16387.t6 A[6].t19 a_15946_15776.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1284 VDD.t94 a_51054_2325.t11 a_51109_747.t3 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1285 a_22584_5326.t3 A[1].t13 VSS.t307 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1286 VDD.t1394 B[6].t10 a_54879_11969.t2 VDD.t1393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1287 a_39681_1042.t6 a_39254_1735.t4 a_39799_1042.t2 VDD.t1968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1288 a_58868_15769.t6 a_58326_16165.t11 VDD.t983 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1289 a_65767_10704.t3 a_65222_11397.t7 a_65649_10704.t7 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1290 a_52887_1041.t10 a_53299_1015.t5 a_53005_1041.t6 VDD.t4472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1291 VDD.t2831 a_44465_8220.t7 a_45055_7783.t0 VDD.t2830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1292 VDD.t4262 a_53005_1041.t10 a_54358_1734.t2 VDD.t4261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1293 a_52473_15766.t2 a_51815_16459.t6 a_52355_15766.t3 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1294 a_35222_3549.t1 A[5].t17 a_34985_4186.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1295 a_65224_7306.t2 a_64188_3841.t7 VDD.t1059 VDD.t1058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1296 VDD.t886 a_59635_6910.t10 a_60988_7603.t2 VDD.t885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1297 a_11829_5352.t2 B[6].t11 VDD.t1396 VDD.t1395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1298 a_14046_n3485.t0 a_13401_n2178.t6 VSS.t23 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1299 a_21211_16387.t2 B[2].t6 VDD.t3735 VDD.t3734 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1300 VDD.t1744 opcode[0].t68 a_4879_13585.t2 VDD.t1743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1301 Y[2].t2 a_16954_n2152.t8 VDD.t1971 VDD.t1970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1302 a_53010_6842.t1 a_53304_6816.t4 a_52892_6842.t8 VDD.t2518 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1303 a_10509_14454.t0 a_10449_14428.t4 a_9976_13724.t0 VDD.t404 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1304 a_1089_11724.t2 a_498_14458.t6 a_556_10994.t3 VDD.t504 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1305 VSS.t662 a_19454_10990.t11 a_19396_11720.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1306 a_9304_16408.t2 A[3].t21 a_9168_15798.t2 VDD.t4387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1307 a_13721_8992.t3 opcode[0].t69 VDD.t3815 VDD.t3814 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1308 a_19997_8988.t4 a_20643_8115.t6 a_19464_8258.t6 VDD.t145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1309 a_13898_5354.t9 a_14310_5328.t5 a_7315_8962.t1 VDD.t3058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1310 VDD.t4309 opcode[3].t23 a_280_n2152.t2 VDD.t4308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1311 a_55224_23614.t3 a_54960_24197.t5 VSS.t170 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1312 a_13711_11724.t9 a_13120_14458.t4 a_13178_10994.t5 VDD.t3928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1313 a_30154_11447.t2 B[0].t9 VDD.t2207 VDD.t2206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1314 VDD.t1023 a_54903_1041.t12 a_57731_748.t5 VDD.t1022 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1315 a_47794_3876.t4 a_45049_1913.t6 a_47912_3876.t4 VDD.t4246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1316 VDD.t881 a_54658_21365.t12 a_56438_21365.t1 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1317 VDD.t291 A[4].t23 a_35012_10049.t5 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1318 VDD.t363 a_64185_771.t6 a_65224_3811.t0 VDD.t362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1319 a_65767_9972.t1 a_66061_10678.t5 VSS.t454 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1320 a_10458_20259.t0 A[4].t24 VSS.t320 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1321 VDD.t375 a_3700_13728.t10 a_3642_14458.t0 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1322 VDD.t313 a_9976_13724.t8 a_9918_14454.t2 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1323 a_14357_10851.t2 opcode[1].t54 VDD.t716 VDD.t715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1324 a_4183_8966.t4 a_12241_5326.t4 a_11829_5352.t9 VDD.t2257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1325 VDD.t3872 opcode[0].t70 a_13011_21592.t1 VDD.t3871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1326 VSS.t359 a_37856_8106.t9 a_38148_5891.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1327 a_23777_13581.t3 opcode[0].t71 VSS.t609 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1328 VDD.t905 a_48254_6910.t14 a_51119_8152.t6 VDD.t904 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1329 VDD.t2604 B[7].t8 a_9221_6047.t2 VDD.t2603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1330 VDD.t1670 a_41697_1042.t10 a_46232_1040.t11 VDD.t1669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1331 a_46356_6910.t0 a_45811_7603.t4 a_46356_6178.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1332 a_40621_16458.t1 A[7].t11 VDD.t3749 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1333 VDD.t383 a_1964_13805.t7 a_1089_14458.t9 VDD.t382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1334 a_566_8262.t0 a_1039_8966.t9 a_1099_8992.t0 VDD.t498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1335 a_16605_n2152.t0 a_17479_n2637.t7 a_16954_n2152.t0 VDD.t4242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1336 a_57736_2352.t3 a_57676_2326.t6 VDD.t1643 VDD.t1642 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1337 a_22849_1744.t6 a_22540_11720.t4 VDD.t3167 VDD.t3166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1338 a_24240_5350.t2 B[0].t10 VDD.t2209 VDD.t2208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1339 VDD.t1965 a_40296_23896.t5 a_42031_24205.t5 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1340 a_39689_6822.t8 a_35594_7027.t6 VDD.t3703 VDD.t3702 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1341 a_61510_21343.t3 A[3].t22 VSS.t255 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1342 VDD.t3424 a_9228_15824.t7 a_13711_14458.t0 VDD.t3423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1343 VDD.t2211 B[0].t11 a_29954_12048.t4 VDD.t2210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1344 a_61415_6910.t3 a_60988_7603.t4 a_61533_6910.t1 VDD.t1857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1345 a_54960_24197.t2 a_53352_20634.t5 a_55078_24197.t4 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1346 a_41573_15739.t3 a_30643_n2374.t11 VSS.t617 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1347 a_39807_6822.t3 a_39262_7515.t5 a_39807_6090.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1348 VDD.t3870 a_30643_n2374.t12 a_42770_18699.t6 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1349 a_4300_1740.t0 opcode[2].t22 a_4536_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1350 a_4233_11724.t2 a_3642_14458.t4 a_3700_10994.t6 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1351 a_61525_1042.t2 a_61819_1016.t4 a_61407_1042.t3 VDD.t1771 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1352 a_7989_n2633.t3 a_7432_1744.t10 VSS.t431 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1353 a_34985_4186.t5 A[5].t18 VDD.t2088 VDD.t2087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1354 a_13849_16387.t4 A[7].t12 VDD.t3751 VDD.t3750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1355 a_4233_14458.t8 opcode[0].t72 VDD.t3847 VDD.t3846 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1356 a_70513_20044.t4 a_43509_21373.t9 a_70513_19926.t5 VDD.t2695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1357 a_11505_15751.t2 A[1].t14 a_11640_16408.t4 VDD.t1931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1358 a_41579_1042.t1 a_39799_1042.t10 VDD.t3661 VDD.t3660 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1359 a_54572_9678.t1 a_53576_9091.t5 VDD.t2626 VDD.t2625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1360 a_55504_n1325.t3 a_54914_n1762.t7 VSS.t486 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1361 VDD.t3621 a_41705_6822.t10 a_65222_11397.t2 VDD.t3620 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1362 a_44682_3363.t0 a_41697_1042.t11 a_44445_4000.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1363 a_64117_5761.t1 a_63527_6198.t8 VDD.t1275 VDD.t1274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1364 a_5331_6357.t1 A[4].t25 VDD.t1993 VDD.t1992 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1365 VDD.t3474 a_58312_3565.t4 a_60047_3874.t5 VDD.t3473 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1366 a_38492_9345.t1 a_37902_9782.t9 VDD.t3342 VDD.t3341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1367 a_56366_23618.t3 a_56102_24201.t6 VSS.t211 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1368 a_19927_14428.t1 a_22709_16385.t9 VDD.t2446 VDD.t2445 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1369 a_54879_11969.t1 B[6].t12 VDD.t1398 VDD.t1397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1370 a_46770_3872.t0 a_45044_309.t4 a_46652_3872.t0 VDD.t1484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1371 VDD.t4564 a_59223_16436.t12 a_58868_15769.t2 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1372 a_57684_8194.t2 a_61071_3878.t6 VSS.t712 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1373 a_44460_6616.t2 a_42266_11512.t10 VDD.t3797 VDD.t3796 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1374 a_59901_23892.t2 a_59311_24329.t8 VDD.t1013 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1375 a_55862_18700.t0 a_30643_1763.t11 VDD.t2405 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1376 a_52355_15766.t9 a_52767_15740.t4 a_52473_15766.t5 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1377 a_29952_n363.t2 B[6].t13 VDD.t1400 VDD.t1399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1378 VDD.t1025 a_54903_1041.t13 a_59509_1042.t10 VDD.t1024 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1379 a_38140_111.t1 a_35575_3749.t7 a_37903_748.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1380 a_3392_1740.t1 opcode[2].t23 VDD.t2950 VDD.t2949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1381 VDD.t4204 a_4491_15753.t5 a_1964_13805.t0 VDD.t4203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1382 a_4879_13585.t1 opcode[0].t73 VDD.t3828 VDD.t3827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1383 VSS.t337 a_4593_6357.t5 a_8202_7655.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1384 a_61407_1042.t4 a_61819_1016.t5 a_61525_1042.t1 VDD.t1772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1385 VDD.t1973 a_16954_n2152.t9 Y[2].t1 VDD.t1972 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1386 a_38493_311.t3 a_37903_748.t9 VSS.t68 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1387 a_22489_21592.t0 opcode[0].t74 VDD.t3826 VDD.t3825 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1388 a_23358_15774.t0 B[1].t8 VSS.t389 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1389 a_9976_13724.t1 a_10449_14428.t5 a_10509_14454.t1 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1390 a_20086_n2148.t2 a_20611_n2633.t5 a_19737_n2148.t2 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1391 VSS.t415 a_53010_6842.t11 a_54363_7535.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1392 VDD.t417 a_48426_24202.t7 a_48690_23619.t1 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1393 a_63602_n1637.t2 B[6].t14 VDD.t1402 VDD.t1401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1394 a_48248_1040.t1 a_47703_1733.t5 a_48130_1040.t1 VDD.t3406 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1395 a_9168_15798.t1 A[3].t23 a_9304_16408.t1 VDD.t4395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1396 a_1926_7659.t1 opcode[0].t75 a_566_8262.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1397 VDD.t1740 opcode[0].t76 a_29950_n2431.t1 VDD.t1739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1398 a_17501_13585.t2 opcode[0].t77 VDD.t1789 VDD.t1788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1399 VDD.t2425 B[3].t13 a_29952_5843.t7 VDD.t2424 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1400 a_70513_7422.t4 a_65769_3118.t8 VDD.t2698 VDD.t2697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1401 a_280_n2152.t1 opcode[3].t24 VDD.t4311 VDD.t4310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1402 VSS.t476 opcode[2].t24 a_6524_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1403 a_41711_n1755.t3 B[5].t9 VDD.t1814 VDD.t1813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1404 a_22608_8258.t3 a_23787_8115.t4 a_23141_8988.t5 VDD.t598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1405 VSS.t678 opcode[3].t25 a_6556_n2148.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1406 a_48225_11948.t6 A[5].t19 VDD.t2090 VDD.t2089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1407 a_839_n2152.t10 opcode[3].t26 VDD.t4313 VDD.t4312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1408 VDD.t4257 a_53005_1041.t11 a_54785_1041.t10 VDD.t4256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1409 VDD.t1283 a_556_13728.t9 a_498_14458.t2 VDD.t1282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1410 a_16332_8262.t4 a_17511_8119.t5 a_16865_8992.t9 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1411 VSS.t62 a_64185_771.t7 a_67372_3171.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1412 a_60226_16462.t2 A[4].t26 VDD.t1994 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1413 VDD.t1589 a_10199_n2174.t4 a_10259_n2148.t0 VDD.t1588 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1414 a_57959_3365.t0 a_54903_1041.t14 a_57722_4002.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1415 a_70459_5045.t3 opcode[1].t55 VSS.t125 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1416 a_13011_21592.t0 opcode[0].t78 VDD.t3821 VDD.t3820 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1417 VSS.t348 a_30152_9379.t6 a_31377_10037.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1418 a_70509_10506.t6 a_63114_21369.t8 a_70509_10624.t8 VDD.t3532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1419 VDD.t582 a_51695_9365.t5 a_53430_9674.t4 VDD.t581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1420 a_30152_475.t1 opcode[0].t79 VDD.t3819 VDD.t3818 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1421 a_807_1740.t10 a_498_11724.t5 VDD.t587 VDD.t586 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1422 VDD.t68 a_57739_6616.t9 a_58329_6179.t1 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1423 VDD.t2812 a_57684_8194.t11 a_61415_6910.t6 VDD.t2811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1424 a_18035_5352.t2 a_18447_5326.t5 a_13661_8966.t3 VDD.t1624 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1425 a_7375_8988.t10 a_7315_8962.t9 a_6842_8258.t5 VDD.t3289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1426 VDD.t239 a_44405_8194.t9 a_44460_6616.t5 VDD.t238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1427 VDD.t159 a_41507_3295.t10 a_45811_7603.t1 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1428 a_51054_2325.t1 a_54454_9678.t6 VSS.t670 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1429 VSS.t19 a_11133_n2633.t5 a_11080_n3481.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1430 a_60047_3874.t1 a_58321_311.t4 a_59929_3874.t3 VDD.t3512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1431 VDD.t2645 a_46356_6910.t9 a_47709_7603.t0 VDD.t2644 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1432 a_42031_24205.t4 a_40296_23896.t6 VDD.t1966 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1433 a_30643_1763.t3 a_30150_1105.t5 a_29950_1706.t8 VDD.t3668 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1434 a_53357_22238.t2 a_52767_22675.t7 VDD.t4134 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1435 a_55078_24197.t5 a_53352_20634.t6 a_54960_24197.t3 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1436 a_46176_16428.t2 a_47179_16454.t6 a_47719_15761.t6 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1437 VSS.t553 a_58312_3565.t5 a_59929_3874.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1438 a_42770_18699.t0 a_30643_n2374.t13 VDD.t3104 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1439 VDD.t1107 a_46140_17941.t6 a_38721_16161.t1 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1440 VDD.t3843 opcode[0].t80 a_4233_14458.t7 VDD.t3842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1441 a_38506_7695.t1 a_37916_8132.t8 VDD.t2904 VDD.t2903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1442 VDD.t3753 A[7].t13 a_13849_16387.t3 VDD.t3752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1443 VDD.t3845 opcode[0].t81 a_10509_14454.t5 VDD.t3844 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1444 a_17158_407.t1 a_16264_11724.t4 VSS.t82 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1445 VDD.t424 a_40109_9654.t6 a_40373_9071.t2 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1446 a_38501_6091.t1 a_37911_6528.t8 VSS.t336 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1447 a_16322_10994.t6 a_16264_14458.t5 a_16855_11724.t2 VDD.t506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1448 VDD.t346 a_43055_24209.t8 a_43319_23626.t0 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1449 a_54785_1041.t2 a_51054_2325.t12 VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1450 a_53713_16459.t1 A[5].t20 VDD.t2091 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1451 a_14250_407.t0 a_12870_1740.t4 a_13778_1740.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1452 VSS.t35 a_35591_989.t12 a_38145_1715.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1453 VDD.t1141 a_64117_5761.t8 a_65651_6613.t8 VDD.t1140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1454 VDD.t2448 a_22709_16385.t10 a_19927_14428.t2 VDD.t2447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1455 VDD.t3569 a_9986_8258.t9 a_9928_8988.t2 VDD.t3568 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1456 a_70459_20811.t3 opcode[1].t56 VSS.t126 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1457 VDD.t984 a_58326_16165.t12 a_62361_17053.t6 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1458 a_58868_15769.t1 a_59223_16436.t13 VDD.t4563 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1459 VDD.t718 opcode[1].t57 a_17501_10851.t1 VDD.t717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1460 a_54665_15740.t2 a_30643_1763.t12 VSS.t381 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1461 a_30152_6681.t2 opcode[0].t82 VDD.t1797 VDD.t1796 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1462 a_50258_20638.t0 a_48124_21370.t12 a_50022_21370.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1463 a_61197_9746.t3 a_60201_9159.t7 VDD.t329 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1464 VDD.t2406 a_30643_1763.t13 a_55862_18700.t1 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1465 a_70513_16900.t7 a_70459_17667.t4 a_70513_16782.t5 VDD.t3418 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1466 a_52473_15766.t6 a_52767_15740.t5 a_52355_15766.t10 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1467 VDD.t4206 a_22550_8988.t5 a_23131_11720.t5 VDD.t4205 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1468 VSS.t331 A[5].t21 a_4593_6357.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1469 VSS.t414 a_30645_10037.t19 a_47579_22063.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1470 VDD.t1983 a_35001_1426.t9 a_35591_989.t1 VDD.t1982 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1471 a_64188_3841.t3 a_63598_4278.t8 VSS.t455 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1472 VSS.t703 a_54713_3294.t9 a_59090_7603.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1473 VDD.t4020 a_38484_3565.t5 a_40219_3874.t4 VDD.t4019 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1474 a_48136_6910.t1 a_47709_7603.t5 a_48254_6910.t1 VDD.t2160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1475 a_1964_13805.t1 a_4491_15753.t6 VDD.t4297 VDD.t4296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1476 a_52887_1041.t7 a_48855_n1313.t8 VDD.t1233 VDD.t1232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1477 VDD.t2952 opcode[2].t25 a_6524_1744.t1 VDD.t2951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1478 a_21956_20862.t2 a_23135_20719.t5 a_22489_21592.t6 VDD.t2806 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1479 a_10509_14454.t2 a_10449_14428.t6 a_9976_13724.t2 VDD.t406 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1480 a_44702_7583.t1 a_44405_8194.t10 a_44465_8220.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1481 a_63532_11802.t4 B[3].t14 VDD.t2427 VDD.t2426 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1482 VSS.t575 a_41705_6822.t11 a_65222_11397.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1483 a_65651_3118.t7 a_54908_6842.t12 VDD.t4575 VDD.t4574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1484 VDD.t1404 B[6].t15 a_63602_n1637.t1 VDD.t1403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1485 a_54879_11969.t5 A[6].t20 VDD.t3032 VDD.t3031 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1486 VSS.t489 A[6].t21 a_3855_6357.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1487 VSS.t10 a_3855_6357.t5 a_5070_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1488 VDD.t4315 opcode[3].t27 a_280_n2152.t0 VDD.t4314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1489 VDD.t2685 a_57731_748.t7 a_58321_311.t2 VDD.t2684 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1490 a_54253_15766.t2 a_54665_15740.t5 a_52710_16433.t1 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1491 a_30150_2544.t2 opcode[0].t83 VDD.t1746 VDD.t1745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1492 a_3700_10994.t0 a_4879_10851.t4 a_4233_11724.t6 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1493 a_40724_17941.t1 a_41153_18571.t6 a_40859_18597.t5 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1494 VDD.t4317 opcode[3].t28 a_839_n2152.t11 VDD.t4316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1495 a_51114_6548.t5 a_48815_11511.t10 VDD.t2271 VDD.t2270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1496 a_62375_18703.t4 A[4].t27 VDD.t1995 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1497 a_498_14458.t1 a_556_13728.t10 VDD.t2730 VDD.t2729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1498 a_48484_308.t0 a_46350_1040.t9 a_48248_1040.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1499 VDD.t638 a_6832_13724.t11 a_6774_14454.t0 VDD.t637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1500 VDD.t1996 A[4].t28 a_60226_16462.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1501 a_10259_n2148.t1 a_10199_n2174.t5 VDD.t1591 VDD.t1590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1502 VDD.t2322 A[0].t12 a_24652_5324.t2 VDD.t2321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1503 a_20588_7655.t0 a_19937_8962.t9 VSS.t343 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1504 VDD.t1942 a_37848_2326.t10 a_37903_748.t2 VDD.t1941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1505 a_61533_6178.t1 a_61827_6884.t5 VSS.t505 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1506 VDD.t1944 a_37848_2326.t11 a_41991_1016.t1 VDD.t1943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1507 a_20457_4618.t0 B[2].t7 VSS.t595 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1508 a_59311_24329.t6 A[3].t24 VDD.t4394 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1509 a_9976_10990.t7 a_11155_10847.t4 a_11100_10387.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1510 a_70513_20044.t1 a_70459_20811.t5 a_70513_19926.t1 VDD.t656 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1511 a_41161_15765.t8 A[7].t14 VDD.t3754 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1512 a_10509_11720.t6 opcode[1].t58 VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1513 a_58320_9433.t1 a_57730_9870.t8 VDD.t544 VDD.t543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1514 a_46356_6910.t3 a_45811_7603.t5 a_46238_6910.t2 VDD.t1860 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1515 VDD.t2340 a_70509_10506.t9 a_14303_1255.t1 VDD.t2339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1516 a_10513_20719.t2 opcode[0].t84 VDD.t1806 VDD.t1805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1517 VDD.t2787 a_65769_6613.t9 a_70513_16900.t4 VDD.t2786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1518 VDD.t3932 a_19454_13724.t8 a_19396_14454.t2 VDD.t3931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1519 VSS.t409 a_3710_8262.t9 a_3652_8992.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1520 a_59509_1042.t3 a_59082_1735.t5 a_59627_1042.t4 VDD.t2497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1521 VDD.t1967 a_40296_23896.t7 a_42031_24205.t3 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1522 VDD.t2324 A[0].t13 a_8289_6359.t1 VDD.t2323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1523 VDD.t4135 a_52767_22675.t8 a_53357_22238.t3 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1524 a_3983_n2152.t1 a_3923_n2178.t6 VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1525 VDD.t217 a_35591_989.t13 a_37908_2352.t1 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1526 a_21211_16387.t6 A[2].t12 a_21860_15776.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1527 VDD.t1717 a_1974_8339.t6 a_1099_8992.t4 VDD.t1716 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1528 VDD.t2974 a_53343_23888.t6 a_55078_24197.t1 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1529 a_47719_15761.t0 a_48131_15735.t4 a_46176_16428.t3 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1530 VSS.t98 a_1681_1255.t6 a_1628_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1531 VDD.t2213 B[0].t12 a_23700_6043.t1 VDD.t2212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1532 VDD.t4341 a_35602_9612.t7 a_37911_6528.t2 VDD.t4340 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1533 a_38721_16161.t2 a_46140_17941.t7 VDD.t1108 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1534 Y[7].t2 a_1188_n2152.t9 VDD.t1537 VDD.t1536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1535 a_4233_14458.t6 opcode[0].t85 VDD.t4061 VDD.t4060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1536 VDD.t106 a_16922_1740.t9 a_17479_n2637.t2 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1537 VDD.t2954 opcode[2].t26 a_9668_1744.t1 VDD.t2953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1538 a_3951_1740.t6 a_3392_1740.t5 a_4300_1740.t2 VDD.t2289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1539 a_53352_20634.t2 a_52762_21071.t7 VDD.t4532 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1540 a_23141_8988.t8 a_8289_6359.t4 VDD.t4065 VDD.t4064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1541 VDD.t3962 A[2].t13 a_20103_5350.t6 VDD.t3961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1542 a_54952_21339.t1 A[2].t14 VDD.t3963 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1543 a_48360_20638.t1 a_30645_10037.t20 a_48124_21370.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1544 a_1745_8119.t2 opcode[0].t86 VDD.t3998 VDD.t3997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1545 a_18447_5326.t3 A[3].t25 VSS.t254 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1546 a_13838_20259.t0 opcode[0].t87 a_12478_20862.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1547 VSS.t113 a_7551_6363.t4 a_20824_7655.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1548 a_54785_1041.t8 a_54358_1734.t5 a_54903_1041.t5 VDD.t1553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1549 a_55151_n1325.t0 B[6].t16 a_54914_n1762.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1550 VDD.t241 a_44405_8194.t11 a_48136_6910.t10 VDD.t240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1551 a_62361_17053.t5 a_58326_16165.t13 VDD.t985 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1552 a_17501_10851.t0 opcode[1].t59 VDD.t722 VDD.t721 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1553 a_11640_16408.t1 B[1].t9 VDD.t2457 VDD.t2456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1554 a_55862_18700.t2 a_30643_1763.t14 VDD.t2407 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1555 a_23198_1744.t2 a_23723_1259.t5 a_22849_1744.t4 VDD.t4420 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1556 a_70513_19926.t2 a_70459_20811.t6 a_71846_20635.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1557 a_44696_1713.t0 a_44399_2324.t10 a_44459_2350.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1558 a_64117_8794.t1 a_63527_9231.t8 VDD.t2070 VDD.t2069 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1559 a_37911_6528.t1 a_35602_9612.t8 VDD.t4343 VDD.t4342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1560 a_22489_21592.t7 a_23135_20719.t6 a_21956_20862.t3 VDD.t2807 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1561 VDD.t3691 a_42177_23622.t5 a_43173_24209.t4 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1562 VDD.t2429 B[3].t15 a_63532_11802.t5 VDD.t2428 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1563 VSS.t627 A[2].t15 a_10337_15751.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1564 a_59223_16436.t6 a_60226_16462.t5 a_60766_15769.t10 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1565 a_39263_15765.t1 a_38721_16161.t10 VDD.t1655 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1566 VDD.t3034 A[6].t22 a_54879_11969.t4 VDD.t3033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1567 a_40093_1016.t1 a_35575_3749.t8 VDD.t2708 VDD.t2707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1568 VDD.t1143 a_64117_5761.t9 a_67135_7303.t5 VDD.t1142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1569 a_70459_8189.t2 opcode[1].t60 VDD.t724 VDD.t723 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1570 a_10173_5328.t3 A[7].t15 VSS.t597 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1571 VSS.t582 a_6202_20866.t9 a_3923_n2178.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1572 a_57744_8220.t1 a_54713_3294.t10 VDD.t4521 VDD.t4520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1573 a_56850_21339.t1 a_49832_23623.t7 VDD.t994 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1574 a_46238_6910.t10 a_41507_3295.t11 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1575 VDD.t1088 a_41913_24205.t5 a_42177_23622.t0 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1576 a_60766_15769.t6 A[4].t29 VDD.t1997 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1577 a_54908_6842.t1 a_54363_7535.t5 a_54908_6110.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1578 VDD.t4244 a_556_13728.t11 a_498_14458.t0 VDD.t4243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1579 a_8011_10847.t3 opcode[1].t61 VSS.t127 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1580 a_30645_10037.t2 a_30152_9379.t7 a_29952_9980.t8 VDD.t2152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1581 VDD.t3915 opcode[0].t88 a_8021_8115.t1 VDD.t3914 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1582 a_4300_1740.t6 a_4825_1255.t6 a_3951_1740.t10 VDD.t3403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1583 a_11336_10387.t1 opcode[1].t62 a_9976_10990.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1584 a_41933_310.t0 a_39799_1042.t11 a_41697_1042.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1585 a_9976_10990.t4 a_11155_10847.t5 a_10509_11720.t9 VDD.t4074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1586 VDD.t773 a_48064_9163.t8 a_51109_747.t1 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1587 a_7305_14428.t0 a_16795_16385.t9 VDD.t3956 VDD.t3955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1588 a_54960_24197.t4 a_53352_20634.t7 VSS.t643 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1589 VDD.t3921 opcode[0].t89 a_10513_20719.t1 VDD.t3920 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1590 a_19396_14454.t1 a_19454_13724.t9 VDD.t3934 VDD.t3933 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1591 VDD.t2093 A[5].t22 a_35004_7464.t5 VDD.t2092 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1592 a_61827_6884.t1 a_57684_8194.t12 VDD.t2814 VDD.t2813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1593 a_29950_1706.t1 B[5].t10 VDD.t1816 VDD.t1815 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1594 a_53357_22238.t0 a_52767_22675.t9 VDD.t3557 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1595 VDD.t931 B[4].t8 a_30152_3173.t2 VDD.t930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1596 a_57976_5979.t1 a_55469_11532.t9 a_57739_6616.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1597 a_42761_15445.t2 a_38721_16161.t11 VDD.t1654 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1598 a_4824_10391.t0 a_3642_14458.t5 VSS.t25 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1599 a_46916_3289.t1 a_46652_3872.t6 VDD.t3147 VDD.t3146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1600 a_55078_24197.t0 a_53343_23888.t7 VDD.t2975 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1601 VSS.t576 a_41705_6822.t12 a_67370_10757.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1602 a_70509_10624.t10 opcode[1].t63 VDD.t726 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1603 a_25633_21592.t7 a_26279_20719.t5 a_25100_20862.t2 VDD.t2183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1604 VDD.t1539 a_1188_n2152.t10 Y[7].t1 VDD.t1538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1605 a_46652_3872.t1 a_45044_309.t5 VSS.t234 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1606 a_19464_8258.t2 a_19937_8962.t10 a_19997_8988.t7 VDD.t2128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1607 a_37856_8106.t1 a_67135_7303.t8 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1608 a_17444_15774.t0 B[5].t11 VSS.t289 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1609 a_16378_5326.t3 A[4].t30 VSS.t321 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1610 a_44459_2350.t1 a_44399_2324.t11 VDD.t4159 VDD.t4158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1611 VDD.t2459 B[1].t10 a_30152_9379.t2 VDD.t2458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1612 a_55144_6110.t1 a_53010_6842.t12 a_54908_6842.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1613 VSS.t304 a_40724_17941.t5 a_39657_18575.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1614 a_1735_13585.t2 opcode[0].t90 VDD.t3835 VDD.t3834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1615 a_70455_11391.t2 opcode[1].t64 VDD.t728 VDD.t727 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1616 a_51105_9802.t1 a_48254_6910.t15 VDD.t907 VDD.t906 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1617 VDD.t3817 opcode[0].t91 a_29950_1706.t5 VDD.t3816 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1618 VDD.t3633 a_47282_17937.t6 a_46215_18571.t1 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1619 a_15680_20866.t7 a_16859_20723.t5 a_16213_21596.t10 VDD.t1964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1620 VDD.t775 a_48064_9163.t9 a_53299_1015.t2 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1621 a_4626_16408.t2 B[7].t9 VDD.t2606 VDD.t2605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1622 VSS.t332 A[5].t23 a_13838_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1623 a_48006_21370.t2 a_48418_21344.t4 a_48124_21370.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1624 a_22584_5326.t2 A[1].t15 VDD.t1933 VDD.t1932 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1625 VDD.t651 a_55469_11532.t10 a_59929_6884.t2 VDD.t650 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1626 VDD.t652 a_62375_18703.t8 a_60404_18575.t2 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1627 VSS.t33 a_47179_16454.t7 a_47837_15029.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1628 VDD.t3705 a_35594_7027.t7 a_39262_7515.t2 VDD.t3704 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1629 a_10576_1744.t4 opcode[2].t27 a_10812_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1630 a_11505_15751.t3 A[1].t16 a_11640_16408.t5 VDD.t1934 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1631 a_1089_11724.t10 opcode[1].t65 VDD.t730 VDD.t729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1632 a_20643_8115.t3 opcode[0].t92 VSS.t606 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1633 VSS.t457 a_57684_8194.t13 a_57976_5979.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1634 a_57973_1715.t0 a_57676_2326.t7 a_57736_2352.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1635 VDD.t2094 A[5].t24 a_55862_18700.t4 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1636 a_13898_5354.t8 a_14310_5328.t6 a_7315_8962.t2 VDD.t3059 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1637 VDD.t1235 a_48855_n1313.t9 a_52460_1734.t1 VDD.t1234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1638 VSS.t189 a_21632_6045.t4 a_22290_4620.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1639 VDD.t3180 opcode[0].t93 a_13657_20719.t1 VDD.t3179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1640 a_37902_9782.t2 a_35602_9612.t9 VDD.t4345 VDD.t4344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1641 a_7551_6363.t1 A[1].t17 VDD.t3389 VDD.t3388 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1642 a_1660_n3485.t1 a_280_n2152.t4 a_1188_n2152.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1643 a_21956_20862.t4 a_23135_20719.t7 a_22489_21592.t8 VDD.t2808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1644 a_60766_15769.t11 a_60226_16462.t6 a_59223_16436.t7 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1645 a_51690_3564.t1 a_51100_4001.t8 VDD.t2190 VDD.t2189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1646 a_12732_15818.t2 a_12672_15792.t5 VDD.t3237 VDD.t3236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1647 VDD.t933 B[4].t9 a_15426_6045.t2 VDD.t932 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1648 VDD.t909 a_48254_6910.t16 a_51119_8152.t5 VDD.t908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1649 a_70509_13768.t11 opcode[1].t66 VDD.t732 VDD.t731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1650 a_38153_7495.t0 a_37856_8106.t10 a_37916_8132.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1651 VDD.t1298 a_4332_n2152.t8 Y[6].t2 VDD.t1297 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1652 VDD.t1672 a_41697_1042.t12 a_46232_1040.t10 VDD.t1671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1653 a_59635_6910.t4 a_59090_7603.t6 a_59635_6178.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1654 VDD.t3036 A[6].t23 a_11829_5352.t5 VDD.t3035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1655 a_53299_1015.t1 a_48064_9163.t10 VDD.t777 VDD.t776 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1656 VDD.t1343 a_51105_9802.t7 a_51695_9365.t0 VDD.t1342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1657 VDD.t2512 a_30645_3831.t21 a_60766_15769.t2 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1658 a_11133_n2633.t1 a_10576_1744.t9 VDD.t2553 VDD.t2552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1659 a_4879_13585.t0 opcode[0].t94 VDD.t1482 VDD.t1481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1660 a_39689_6822.t1 a_35602_9612.t10 VDD.t4347 VDD.t4346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1661 a_56850_21339.t3 a_49832_23623.t8 VSS.t165 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1662 a_42756_17049.t2 a_30643_n2374.t14 VDD.t3105 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1663 a_4824_13125.t1 a_4173_14432.t4 VSS.t168 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1664 a_11100_13121.t1 a_10449_14428.t7 VSS.t73 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1665 a_1735_10851.t0 opcode[1].t67 VDD.t734 VDD.t733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1666 a_65769_6613.t6 a_65224_7306.t5 a_65651_6613.t10 VDD.t1332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1667 VSS.t232 a_23700_6043.t5 a_24358_4618.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1668 VDD.t3482 a_64192_n2074.t8 a_67135_n540.t5 VDD.t3481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1669 VSS.t481 a_51813_16162.t6 a_51815_16459.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1670 a_10509_11720.t10 a_11155_10847.t6 a_9976_10990.t5 VDD.t4075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1671 VSS.t315 a_9928_8988.t4 a_11336_10387.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1672 VSS.t85 a_55504_n1325.t11 a_57973_1715.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1673 a_12672_15792.t3 A[0].t14 a_12808_16408.t4 VDD.t2325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1674 a_46644_1014.t3 a_41697_1042.t13 VSS.t271 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1675 a_34985_4186.t2 B[4].t10 VDD.t935 VDD.t934 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1676 VDD.t3936 a_19454_13724.t10 a_19396_14454.t0 VDD.t3935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1677 a_19737_n2148.t6 a_19677_n2174.t4 VDD.t2825 VDD.t2824 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1678 VDD.t462 a_16264_11724.t5 a_16573_1740.t0 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1679 a_30643_n2374.t1 a_30150_n3032.t4 a_29950_n2431.t6 VDD.t4116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1680 VDD.t1653 a_38721_16161.t12 a_42761_15445.t1 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1681 a_35012_10049.t4 A[4].t31 VDD.t1999 VDD.t1998 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1682 a_57731_748.t4 a_54903_1041.t15 VDD.t616 VDD.t615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1683 a_3700_10994.t1 a_4879_10851.t5 a_4824_10391.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1684 a_23787_8115.t3 opcode[0].t95 VSS.t621 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1685 VDD.t2608 B[7].t10 a_9221_6047.t1 VDD.t2607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1686 VDD.t3476 a_58312_3565.t6 a_60047_3874.t4 VDD.t3475 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1687 a_25100_20862.t3 a_26279_20719.t6 a_25633_21592.t8 VDD.t2184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1688 VSS.t677 a_49328_18695.t7 a_47357_18567.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1689 Y[7].t0 a_1188_n2152.t11 VDD.t1541 VDD.t1540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1690 a_57736_2352.t2 a_57676_2326.t8 VDD.t1699 VDD.t1698 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1691 a_65769_3118.t4 a_65224_3811.t5 a_65651_3118.t2 VDD.t377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1692 a_24240_5350.t7 A[0].t15 VDD.t2327 VDD.t2326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1693 a_46770_3872.t1 a_45044_309.t6 a_46652_3872.t2 VDD.t2495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1694 VDD.t593 a_25100_20862.t8 a_22821_n2174.t2 VDD.t592 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1695 VDD.t2956 opcode[2].t28 a_16014_1740.t0 VDD.t2955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1696 a_40724_17941.t0 a_40799_18571.t6 VSS.t658 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1697 VDD.t4063 opcode[0].t96 a_1735_13585.t3 VDD.t4062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1698 VDD.t2142 a_41251_9658.t6 a_37848_2326.t1 VDD.t2141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1699 a_40109_9654.t4 a_38501_6091.t5 a_40227_9654.t5 VDD.t1103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1700 VDD.t2753 a_70509_1028.t8 a_4825_1255.t2 VDD.t2752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1701 a_65651_6613.t3 a_66063_6587.t5 a_65769_6613.t1 VDD.t2054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1702 a_30154_12886.t3 opcode[0].t97 VSS.t638 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1703 VDD.t1742 opcode[0].t98 a_29952_9980.t4 VDD.t1741 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1704 a_37856_8106.t3 a_67135_7303.t9 VSS.t105 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1705 VDD.t2610 B[7].t11 a_4626_16408.t1 VDD.t2609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1706 a_70513_4278.t9 opcode[1].t68 VDD.t736 VDD.t735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1707 a_48124_21370.t1 a_48418_21344.t5 a_48006_21370.t3 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1708 a_13188_8262.t6 a_14367_8119.t6 a_14312_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1709 a_24358_4618.t0 a_24652_5324.t5 a_23081_8962.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1710 a_9867_21592.t5 A[4].t32 a_9334_20862.t3 VDD.t2000 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1711 a_60404_18575.t1 a_62375_18703.t9 VDD.t653 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1712 a_4772_407.t0 a_3392_1740.t6 a_4300_1740.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1713 a_22290_1744.t1 opcode[2].t29 VDD.t2958 VDD.t2957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1714 a_55853_15446.t2 a_51813_16162.t7 VDD.t2976 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1715 a_10519_8988.t4 a_10459_8962.t9 a_9986_8258.t6 VDD.t1977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1716 a_23131_14454.t8 a_23777_13581.t5 a_22598_13724.t7 VDD.t2869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1717 VDD.t1946 a_37848_2326.t12 a_41579_1042.t7 VDD.t1945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1718 a_64117_5761.t0 a_63527_6198.t9 VDD.t1277 VDD.t1276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1719 a_70509_13768.t1 a_56556_21365.t9 a_70509_13650.t1 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1720 VDD.t738 opcode[1].t69 a_1089_11724.t9 VDD.t737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1721 VDD.t1701 a_57676_2326.t9 a_61819_1016.t1 VDD.t1700 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1722 a_13657_20719.t0 opcode[0].t99 VDD.t4053 VDD.t4052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1723 a_41611_21373.t0 a_41066_22066.t4 a_41611_20641.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1724 a_30152_10818.t3 opcode[0].t100 VDD.t4055 VDD.t4054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1725 a_16332_8262.t6 a_17511_8119.t6 a_16865_8992.t8 VDD.t4292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1726 VDD.t485 a_55504_n1325.t12 a_57736_2352.t6 VDD.t484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1727 VDD.t2886 a_47794_3876.t7 a_44405_8194.t2 VDD.t2885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1728 VSS.t441 a_53816_17942.t6 a_52749_18576.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1729 VDD.t2634 a_45035_3563.t5 a_46770_3872.t4 VDD.t2633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1730 VDD.t570 a_59627_1042.t11 a_60980_1735.t1 VDD.t569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1731 VSS.t369 A[0].t16 a_8289_6359.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1732 a_51351_1714.t0 a_51054_2325.t13 a_51114_2351.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1733 Y[6].t1 a_4332_n2152.t9 VDD.t1300 VDD.t1299 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1734 a_67133_11394.t1 a_64117_8794.t5 VDD.t2557 VDD.t2556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1735 a_18035_5352.t9 B[3].t16 VDD.t2434 VDD.t2433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1736 a_13429_1740.t3 opcode[2].t30 VDD.t2960 VDD.t2959 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1737 VDD.t4038 opcode[0].t101 a_11155_13581.t1 VDD.t4037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1738 a_3700_13728.t0 a_4879_13585.t4 a_4824_13125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1739 VDD.t3707 a_35594_7027.t8 a_39689_6822.t7 VDD.t3706 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1740 VDD.t3799 a_42266_11512.t11 a_46650_6884.t3 VDD.t3798 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1741 a_43419_18088.t0 a_30643_n2374.t15 VSS.t499 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1742 a_12808_16408.t3 A[0].t17 a_12672_15792.t2 VDD.t2328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1743 a_66063_n1256.t3 a_48248_1040.t11 VSS.t663 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1744 VSS.t676 a_18243_16385.t9 a_10449_14428.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1745 VSS.t104 a_38723_16458.t4 a_39381_15033.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1746 a_16332_8262.t3 a_17511_8119.t7 a_17456_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1747 VDD.t2827 a_19677_n2174.t5 a_19737_n2148.t7 VDD.t2826 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1748 VDD.t528 a_61216_21369.t9 a_62996_21369.t1 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1749 a_41999_6796.t3 a_37856_8106.t11 VSS.t360 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1750 a_42761_15445.t0 a_38721_16161.t13 VDD.t1652 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1751 a_4243_8992.t11 opcode[0].t102 VDD.t4040 VDD.t4039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1752 a_44454_746.t5 a_41697_1042.t14 VDD.t1674 VDD.t1673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1753 VSS.t625 a_16795_16385.t10 a_7305_14428.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1754 VDD.t3390 A[1].t18 a_48006_21370.t11 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1755 a_65649_10704.t8 a_41705_6822.t13 VDD.t3623 VDD.t3622 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1756 a_65769_3118.t0 a_66063_3092.t5 a_65651_3118.t3 VDD.t514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1757 VDD.t1676 a_41697_1042.t15 a_44445_4000.t4 VDD.t1675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1758 a_16213_21596.t5 A[2].t16 a_15680_20866.t3 VDD.t3964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1759 a_63114_21369.t6 a_62569_22062.t4 a_63114_20637.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1760 VDD.t4539 a_49328_18695.t8 a_47357_18567.t2 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1761 a_45939_15761.t0 a_45281_16454.t4 a_45821_15761.t0 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1762 a_14367_8119.t2 opcode[0].t103 VDD.t4002 VDD.t4001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1763 VDD.t1145 a_64117_5761.t10 a_65651_6613.t7 VDD.t1144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1764 VDD.t4393 A[3].t26 a_63598_4278.t4 VDD.t4392 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1765 VDD.t1437 A[6].t24 a_12241_5326.t2 VDD.t1436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1766 a_508_8992.t2 a_566_8262.t9 VDD.t1564 VDD.t1563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1767 a_29954_7911.t8 a_30154_8749.t5 a_30647_7968.t2 VDD.t3643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1768 a_9761_5354.t1 a_10173_5328.t5 a_1039_8966.t1 VDD.t51 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1769 a_46232_1040.t6 a_46644_1014.t5 a_46350_1040.t5 VDD.t1689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1770 VSS.t574 a_39582_17945.t6 Cout.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1771 a_55848_17050.t4 a_30643_1763.t15 VDD.t3130 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1772 VDD.t2977 a_51813_16162.t8 a_51815_16459.t2 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1773 VDD.t3737 B[2].t8 a_19563_6043.t3 VDD.t3736 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1774 a_59921_1016.t2 a_54903_1041.t16 VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1775 VDD.t4427 a_46350_1040.t10 a_47703_1733.t2 VDD.t4426 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1776 a_14335_n2637.t1 a_13778_1740.t9 VDD.t1854 VDD.t1853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1777 a_1156_1740.t1 a_248_1740.t5 a_807_1740.t1 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1778 VDD.t4592 a_7551_6363.t5 a_19997_8988.t9 VDD.t4591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1779 VDD.t3392 A[1].t19 a_22172_5352.t5 VDD.t3391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1780 a_30150_1105.t1 B[5].t12 VDD.t1818 VDD.t1817 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1781 a_248_1740.t1 opcode[2].t31 VDD.t2962 VDD.t2961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1782 a_38506_7695.t0 a_37916_8132.t9 VDD.t2906 VDD.t2905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1783 VDD.t1406 B[6].t17 a_11289_6045.t1 VDD.t1405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1784 a_52887_1041.t6 a_48855_n1313.t10 VDD.t1237 VDD.t1236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1785 a_51114_2351.t1 a_51054_2325.t14 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1786 a_48136_6910.t4 a_48548_6884.t5 a_48254_6910.t5 VDD.t4024 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1787 a_48006_21370.t4 a_48418_21344.t6 a_48124_21370.t2 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1788 VDD.t62 a_55224_23614.t4 a_56220_24201.t0 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1789 VDD.t3049 a_54960_24197.t6 a_55224_23614.t2 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1790 a_9334_20862.t2 A[4].t33 a_9867_21592.t6 VDD.t2001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1791 a_29952_n363.t6 a_30152_475.t5 a_30645_n306.t3 VDD.t532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1792 VDD.t2978 a_51813_16162.t9 a_55853_15446.t1 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1793 VDD.t426 a_40109_9654.t7 a_40373_9071.t1 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1794 VDD.t430 B[2].t9 a_30154_7310.t0 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1795 a_61819_1016.t3 a_57676_2326.t10 VSS.t276 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1796 VDD.t1948 a_37848_2326.t13 a_37903_748.t1 VDD.t1947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1797 a_1713_n2637.t3 a_1156_1740.t9 VSS.t341 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1798 a_16573_1740.t11 a_16014_1740.t6 a_16922_1740.t6 VDD.t3520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1799 a_39717_18601.t2 a_40011_18575.t5 a_39582_17945.t2 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1800 a_10509_14454.t4 opcode[0].t104 VDD.t4004 VDD.t4003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1801 a_22598_13724.t0 a_23777_13581.t6 a_23131_14454.t0 VDD.t260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1802 a_29952_3774.t10 a_30152_4612.t5 a_30645_3831.t5 VDD.t1432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1803 a_70509_1146.t1 a_45939_15761.t9 a_70509_1028.t1 VDD.t630 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1804 a_41697_1042.t2 a_41152_1735.t5 a_41579_1042.t4 VDD.t1580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1805 a_16922_1740.t3 opcode[2].t32 a_17158_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1806 a_807_1740.t5 a_1681_1255.t7 a_1156_1740.t4 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1807 VDD.t4391 A[3].t27 a_6071_6357.t1 VDD.t4390 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1808 a_13401_n2178.t1 a_15680_20866.t10 VDD.t674 VDD.t673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1809 a_41847_20641.t0 a_30647_12105.t12 a_41611_21373.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1810 a_19937_8962.t0 a_21632_6045.t5 a_22172_5352.t3 VDD.t1126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1811 a_61216_20637.t1 a_61510_21343.t4 VSS.t571 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1812 a_1039_8966.t6 a_9221_6047.t5 a_9761_5354.t7 VDD.t3363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1813 VDD.t4319 opcode[3].t29 a_10259_n2148.t11 VDD.t4318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1814 a_14252_4622.t0 B[5].t13 VSS.t290 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1815 a_53816_17942.t0 a_53891_18572.t6 VSS.t44 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1816 VDD.t163 a_41507_3295.t12 a_44451_9870.t5 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1817 VDD.t4175 a_41243_3878.t6 a_41507_3295.t2 VDD.t4174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1818 VSS.t160 a_58326_16165.t14 a_58328_16462.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1819 VDD.t1102 a_3652_8992.t4 a_4233_11724.t3 VDD.t1101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1820 a_64188_3841.t1 a_63598_4278.t9 VDD.t4014 VDD.t4013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1821 a_7365_14454.t11 a_7305_14428.t4 a_6832_13724.t0 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1822 a_12902_n2152.t1 opcode[3].t30 VDD.t4321 VDD.t4320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1823 a_57731_748.t3 a_54903_1041.t17 VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1824 a_20103_5350.t10 a_19563_6043.t6 a_16805_8966.t7 VDD.t3387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1825 VDD.t3651 a_52753_24325.t8 a_53343_23888.t2 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1826 a_15966_5352.t0 B[4].t11 VDD.t937 VDD.t936 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1827 VSS.t637 opcode[0].t105 a_43745_20641.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1828 a_70509_10624.t5 a_70455_11391.t5 a_70509_10506.t2 VDD.t2837 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1829 VDD.t3625 a_41705_6822.t14 a_67133_11394.t2 VDD.t3624 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1830 a_53304_6816.t0 a_48815_11511.t11 VDD.t2273 VDD.t2272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1831 VSS.t434 a_65769_3118.t9 a_71846_8249.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1832 VDD.t219 a_35591_989.t14 a_37908_2352.t0 VDD.t218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1833 VSS.t393 a_12478_20862.t9 a_10199_n2174.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1834 a_11155_13581.t0 opcode[0].t106 VDD.t4046 VDD.t4045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1835 VDD.t455 a_13178_13728.t9 a_13120_14458.t2 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1836 VDD.t1719 a_1974_8339.t7 a_1099_8992.t5 VDD.t1718 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1837 VDD.t779 a_48064_9163.t11 a_52887_1041.t0 VDD.t778 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1838 a_46818_20639.t0 a_46228_21076.t9 VDD.t3174 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1839 a_39717_18601.t0 a_39657_18575.t4 VDD.t2862 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1840 VSS.t4 a_10337_15751.t5 a_10397_15824.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1841 a_42770_18699.t4 A[7].t16 a_43419_18088.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1842 a_39617_15033.t0 a_38721_16161.t14 VSS.t248 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1843 a_25633_21592.t10 VSS.t717 a_25100_20862.t6 VDD.t4601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1844 VDD.t1916 a_30647_7968.t9 a_54113_22058.t2 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1845 a_58321_311.t1 a_57731_748.t8 VDD.t1063 VDD.t1062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1846 a_35575_3749.t0 a_34985_4186.t8 VSS.t260 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1847 a_62996_21369.t0 a_61216_21369.t10 VDD.t529 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1848 a_22849_1744.t10 a_22290_1744.t5 a_23198_1744.t5 VDD.t3115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1849 a_20221_4618.t0 a_20515_5324.t5 a_16805_8966.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1850 a_58320_9433.t0 a_57730_9870.t9 VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1851 a_46356_6910.t2 a_45811_7603.t6 a_46238_6910.t1 VDD.t1861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1852 a_15680_20866.t2 A[2].t17 a_16213_21596.t4 VDD.t3965 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1853 a_63350_20637.t1 a_61216_21369.t11 a_63114_21369.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1854 a_47357_18567.t1 a_49328_18695.t9 VDD.t4540 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1855 a_45821_15761.t1 a_45281_16454.t5 a_45939_15761.t1 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1856 a_17511_8119.t3 opcode[0].t107 VSS.t639 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1857 VDD.t4057 opcode[0].t108 a_19987_14454.t1 VDD.t4056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1858 VDD.t4048 opcode[0].t109 a_30152_6681.t1 VDD.t4047 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1859 a_4183_8966.t3 A[6].t25 a_12183_4620.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1860 a_52355_15766.t8 a_51813_16162.t10 VDD.t2979 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1861 a_59509_1042.t6 a_59921_1016.t5 a_59627_1042.t1 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1862 a_53304_6816.t3 a_48815_11511.t12 VSS.t363 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1863 a_18447_5326.t1 A[3].t28 VDD.t4389 VDD.t4388 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1864 VDD.t1408 B[6].t18 a_63595_1208.t1 VDD.t1407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1865 a_41941_6090.t1 a_39807_6822.t11 a_41705_6822.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1866 VDD.t3131 a_30643_1763.t16 a_55848_17050.t5 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1867 a_51815_16459.t1 a_51813_16162.t11 VDD.t2980 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1868 VDD.t4230 a_48248_1040.t12 a_66063_n1256.t2 VDD.t4229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1869 VDD.t740 opcode[1].t70 a_70513_16900.t10 VDD.t739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1870 VSS.t303 a_30647_7968.t10 a_54113_22058.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1871 VSS.t385 B[3].t17 a_30152_5242.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1872 VDD.t1083 a_46658_9742.t7 a_46922_9159.t1 VDD.t1082 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1873 a_31379_8204.t0 B[2].t10 VSS.t76 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1874 VSS.t190 a_30152_3173.t6 a_31377_3831.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1875 a_45041_9433.t3 a_44451_9870.t7 VSS.t459 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1876 a_3951_1740.t8 opcode[2].t33 VDD.t2964 VDD.t2963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1877 a_38498_1915.t1 a_37908_2352.t9 VDD.t1635 VDD.t1634 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1878 a_61343_9163.t0 a_61079_9746.t5 VDD.t2537 VDD.t2536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1879 VSS.t114 a_11505_15751.t8 a_11565_15824.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1880 a_70509_13768.t7 a_70455_14535.t5 a_70509_13650.t5 VDD.t3129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1881 a_29952_9980.t0 B[1].t11 VDD.t2461 VDD.t2460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1882 a_56220_24201.t1 a_55224_23614.t5 VDD.t63 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1883 a_55224_23614.t1 a_54960_24197.t7 VDD.t3050 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1884 VDD.t742 opcode[1].t71 a_70459_17667.t1 VDD.t741 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1885 a_41587_6822.t4 a_41999_6796.t5 a_41705_6822.t1 VDD.t4147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1886 a_5108_13805.t2 a_5659_15753.t5 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1887 a_55853_15446.t0 a_51813_16162.t12 VDD.t2981 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1888 a_29950_n2431.t10 a_30150_n1593.t5 a_30643_n2374.t7 VDD.t1749 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1889 VDD.t3523 a_61343_9163.t6 a_70509_n1998.t5 VDD.t3522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1890 a_46228_21076.t2 A[1].t20 VDD.t3393 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1891 a_39582_17945.t1 a_40011_18575.t6 a_39717_18601.t4 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1892 VDD.t243 a_44405_8194.t12 a_44465_8220.t5 VDD.t242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1893 a_40093_1016.t0 a_35575_3749.t9 VDD.t2710 VDD.t2709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1894 VSS.t573 a_24157_16385.t10 a_23071_14428.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1895 a_61407_1042.t1 a_57676_2326.t11 VDD.t1703 VDD.t1702 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1896 a_31377_3831.t1 a_30152_4612.t6 a_30645_3831.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1897 VSS.t107 a_54245_18572.t7 a_53816_17942.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1898 VDD.t2492 a_22598_13724.t9 a_22540_14454.t2 VDD.t2491 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1899 a_4233_11724.t7 a_3652_8992.t5 VDD.t2254 VDD.t2253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1900 a_13429_1740.t7 a_13120_11724.t5 VDD.t2281 VDD.t2280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1901 a_18824_20866.t6 A[1].t21 a_19357_21596.t10 VDD.t3394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1902 VDD.t1438 A[6].t26 a_49328_18695.t2 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1903 a_6832_13724.t1 a_7305_14428.t5 a_7365_14454.t10 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1904 VDD.t4050 opcode[0].t110 a_11165_8115.t0 VDD.t4049 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1905 a_10173_5328.t2 A[7].t17 VDD.t3756 VDD.t3755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1906 VSS.t468 a_7957_1259.t5 a_7904_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1907 a_64117_8794.t0 a_63527_9231.t9 VDD.t2072 VDD.t2071 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1908 VDD.t4323 opcode[3].t31 a_12902_n2152.t0 VDD.t4322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1909 a_53343_23888.t3 a_52753_24325.t9 VDD.t3652 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1910 a_49904_21370.t0 a_50316_21344.t4 a_50022_21370.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1911 VDD.t2002 A[4].t34 a_62366_15449.t1 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1912 VSS.t615 a_65769_n1230.t9 a_71842_11451.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1913 VSS.t679 opcode[3].t32 a_12902_n2152.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1914 VDD.t3638 a_54449_3877.t5 a_54713_3294.t0 VDD.t3637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1915 a_37911_6528.t5 a_37856_8106.t12 VDD.t2171 VDD.t2170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1916 a_43509_20641.t1 a_43803_21347.t5 VSS.t171 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1917 VDD.t3177 a_30643_n2374.t16 a_41573_15739.t1 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1918 VSS.t61 a_19464_8258.t9 a_19406_8988.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1919 a_48855_n1313.t1 a_48265_n1750.t9 VDD.t422 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1920 a_70513_20044.t5 a_43509_21373.t10 a_70513_19926.t6 VDD.t2696 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1921 a_67133_11394.t3 a_41705_6822.t15 VDD.t3627 VDD.t3626 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1922 a_7375_8988.t3 a_4593_6357.t6 VDD.t1613 VDD.t1612 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1923 a_64185_771.t3 a_63595_1208.t9 VSS.t287 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1924 a_13120_14458.t1 a_13178_13728.t10 VDD.t457 VDD.t456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1925 VDD.t744 opcode[1].t72 a_70459_20811.t1 VDD.t743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1926 VDD.t3837 opcode[0].t111 a_8011_13581.t1 VDD.t3836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1927 VDD.t449 a_65767_10704.t8 a_70509_13768.t3 VDD.t448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1928 VDD.t2863 a_39657_18575.t5 a_39717_18601.t1 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1929 VDD.t1820 B[5].t14 a_13898_5354.t1 VDD.t1819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1930 VDD.t3396 A[1].t22 a_25633_21592.t3 VDD.t3395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1931 a_10337_15751.t0 B[2].t11 VSS.t77 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1932 a_48131_15735.t3 a_30645_n306.t11 VSS.t541 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1933 a_39381_15765.t4 a_39618_16432.t8 a_39617_15033.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1934 a_42266_11512.t1 a_41676_11949.t7 VSS.t18 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1935 a_46916_3289.t3 a_46652_3872.t7 VSS.t507 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1936 a_46238_6910.t4 a_42266_11512.t12 VDD.t3801 VDD.t3800 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1937 a_25100_20862.t5 VSS.t718 a_25633_21592.t9 VDD.t4602 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1938 VDD.t1303 a_56366_23618.t10 a_62996_21369.t5 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1939 a_56366_23618.t1 a_56102_24201.t7 VDD.t1349 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1940 a_13188_8262.t2 a_13661_8966.t10 a_13721_8992.t4 VDD.t4237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1941 VSS.t533 a_49314_17045.t7 a_46569_18571.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1942 VDD.t877 a_46233_22680.t8 a_46823_22243.t1 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1943 a_48130_1040.t7 a_46350_1040.t11 VDD.t4429 VDD.t4428 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1944 a_53307_3873.t2 a_51699_310.t6 VSS.t20 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1945 VDD.t4541 a_49328_18695.t10 a_47357_18567.t0 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1946 VSS.t696 a_12732_15818.t6 a_23958_13121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1947 a_7432_1744.t2 a_7957_1259.t6 a_7083_1744.t7 VDD.t2899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1948 VDD.t1896 a_60193_3291.t5 a_61189_3878.t4 VDD.t1895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1949 a_19987_14454.t0 opcode[0].t112 VDD.t3839 VDD.t3838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1950 a_16378_5326.t0 A[4].t35 VDD.t2004 VDD.t2003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1951 a_22584_5326.t1 A[1].t23 VDD.t3398 VDD.t3397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1952 VDD.t2982 a_51813_16162.t13 a_52355_15766.t7 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1953 a_70509_n1998.t1 a_39381_15765.t10 a_70509_n2116.t0 VDD.t577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1954 VDD.t3709 a_35594_7027.t9 a_39262_7515.t1 VDD.t3708 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1955 a_63839_n2274.t0 B[6].t19 a_63602_n1637.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1956 a_63527_6198.t1 A[4].t36 VDD.t2006 VDD.t2005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1957 a_23131_14454.t5 a_23071_14428.t5 a_22598_13724.t4 VDD.t1136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1958 VDD.t2770 a_22608_8258.t9 a_22550_8988.t1 VDD.t2769 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1959 VSS.t28 a_41507_3295.t13 a_44688_9233.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1960 a_10115_4622.t0 B[7].t12 VSS.t416 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1961 a_70513_7422.t10 opcode[1].t73 VDD.t1161 VDD.t1160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1962 a_55862_18700.t6 A[5].t25 a_56511_18089.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1963 VDD.t3514 a_62366_15449.t7 a_60758_18575.t0 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1964 a_41251_9658.t4 a_38506_7695.t6 a_41369_9658.t4 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1965 VSS.t680 opcode[3].t33 a_16046_n2152.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1966 VSS.t80 a_65767_10704.t9 a_71842_14595.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1967 a_10608_n2148.t1 a_11133_n2633.t6 a_10259_n2148.t7 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1968 a_11505_15751.t0 B[1].t12 VSS.t390 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1969 a_13898_5354.t5 A[5].t26 VDD.t2096 VDD.t2095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1970 VDD.t64 a_55224_23614.t6 a_56220_24201.t2 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1971 VDD.t3051 a_54960_24197.t8 a_55224_23614.t0 w_54924_24135# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1972 a_54908_6110.t0 a_55202_6816.t6 VSS.t326 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1973 VDD.t303 a_5659_15753.t6 a_5108_13805.t1 VDD.t302 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1974 VDD.t3442 A[5].t27 a_55853_15446.t5 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1975 a_46658_9742.t1 a_45050_6179.t5 a_46776_9742.t4 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1976 VDD.t3399 A[1].t24 a_46228_21076.t1 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1977 a_7365_14454.t5 opcode[0].t113 VDD.t3852 VDD.t3851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1978 a_46233_22680.t1 a_43319_23626.t11 VDD.t2573 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1979 VSS.t430 a_14303_1255.t6 a_14250_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1980 a_47800_9746.t2 a_45055_7783.t5 VSS.t706 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1981 a_61533_6910.t2 a_60988_7603.t5 a_61415_6910.t4 VDD.t1858 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1982 a_59187_17949.t3 a_59616_18579.t5 a_59322_18605.t2 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1983 VDD.t1069 a_51059_8126.t10 a_54790_6842.t7 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1984 a_52674_17946.t4 a_52749_18576.t4 VSS.t657 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1985 a_19987_11720.t8 a_19396_14454.t5 a_19454_10990.t4 VDD.t2430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1986 Y[3].t3 a_13810_n2152.t8 VSS.t656 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1987 VDD.t2778 a_46916_3289.t5 a_47912_3876.t1 VDD.t2777 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1988 a_13721_8992.t8 a_14367_8119.t7 a_13188_8262.t7 VDD.t3472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1989 a_19357_21596.t11 A[1].t25 a_18824_20866.t5 VDD.t3400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1990 a_49328_18695.t1 A[6].t27 VDD.t1439 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1991 a_7365_14454.t9 a_7305_14428.t6 a_6832_13724.t2 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1992 a_29954_12048.t10 a_30154_11447.t5 a_30647_12105.t5 VDD.t3908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1993 a_29950_n2431.t5 opcode[0].t114 VDD.t3854 VDD.t3853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1994 VDD.t365 a_64185_771.t8 a_65224_3811.t1 VDD.t364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1995 a_37894_4002.t6 a_35591_989.t15 VDD.t3559 VDD.t3558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1996 a_29952_5843.t8 B[3].t18 VDD.t2436 VDD.t2435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1997 a_50022_21370.t1 a_50316_21344.t5 a_49904_21370.t1 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1998 a_30152_3173.t1 B[4].t12 VDD.t939 VDD.t938 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1999 a_41573_15739.t0 a_30643_n2374.t17 VDD.t3178 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2000 VDD.t3711 a_35594_7027.t10 a_37902_9782.t6 VDD.t3710 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2001 VDD.t3629 a_41705_6822.t16 a_67133_11394.t4 VDD.t3628 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2002 a_39689_6822.t4 a_39262_7515.t6 a_39807_6822.t1 VDD.t3222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2003 a_52674_17946.t2 a_53103_18576.t6 a_52809_18602.t0 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2004 a_41369_9658.t1 a_40373_9071.t4 VDD.t1123 VDD.t1122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2005 VDD.t911 a_48254_6910.t17 a_52892_6842.t1 VDD.t910 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2006 a_9168_15798.t4 B[3].t19 VSS.t386 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2007 a_48064_9163.t0 a_47800_9746.t7 VDD.t971 VDD.t970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2008 a_8011_13581.t0 opcode[0].t115 VDD.t1776 VDD.t1775 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2009 VDD.t941 B[4].t13 a_15426_6045.t1 VDD.t940 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2010 a_43391_21373.t3 a_41611_21373.t10 VDD.t520 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2011 a_39717_18601.t5 a_39657_18575.t6 VDD.t3234 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2012 a_65767_10704.t6 a_66061_10678.t6 a_65649_10704.t3 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2013 VDD.t1410 B[6].t20 a_29952_n363.t1 VDD.t1409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2014 VDD.t1441 A[6].t28 a_11829_5352.t4 VDD.t1440 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2015 a_39381_15033.t1 a_39675_15739.t5 a_39381_15765.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2016 a_4536_407.t0 a_3642_11724.t5 VSS.t244 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2017 a_62996_21369.t4 a_56366_23618.t11 VDD.t1304 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2018 a_5794_16410.t2 B[6].t21 VDD.t1412 VDD.t1411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2019 VDD.t3862 a_65769_n1230.t10 a_70509_10624.t1 VDD.t3861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2020 a_19997_8988.t6 a_19937_8962.t11 a_19464_8258.t3 VDD.t2129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2021 a_29950_1706.t4 opcode[0].t116 VDD.t1778 VDD.t1777 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2022 VDD.t1350 a_56102_24201.t8 a_56366_23618.t0 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2023 a_21211_16387.t5 A[2].t18 VDD.t3967 VDD.t3966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2024 a_22598_10990.t6 a_22540_14454.t5 a_23131_11720.t10 VDD.t4585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2025 a_6832_10990.t4 a_8011_10847.t4 a_7956_10387.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2026 a_7365_11720.t9 opcode[1].t74 VDD.t1163 VDD.t1162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2027 a_26224_20259.t1 VSS.t403 VSS.t404 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2028 a_19737_n2148.t1 a_20611_n2633.t6 a_20086_n2148.t1 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2029 VDD.t3184 opcode[0].t117 a_1099_8992.t9 VDD.t3183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2030 VDD.t3000 a_67135_n540.t10 a_51059_8126.t3 VDD.t2999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2031 a_65651_6613.t2 a_66063_6587.t6 a_65769_6613.t0 VDD.t2055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2032 VDD.t2758 a_62361_17053.t8 a_59616_18579.t2 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2033 VDD.t3186 opcode[0].t118 a_29952_n363.t10 VDD.t3185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2034 a_49328_18695.t5 a_30645_n306.t12 VDD.t3367 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2035 a_37916_8132.t2 a_37856_8106.t13 VDD.t2173 VDD.t2172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2036 a_35575_3749.t1 a_34985_4186.t9 VDD.t1568 VDD.t1567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2037 a_43509_21373.t3 a_42964_22066.t5 a_43391_21373.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2038 VDD.t3541 a_38721_16161.t15 a_38723_16458.t1 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2039 a_19454_13724.t1 a_20633_13581.t4 a_19987_14454.t3 VDD.t1955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2040 a_50022_21370.t6 a_49477_22063.t6 a_49904_21370.t10 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2041 a_52355_15766.t6 a_51813_16162.t14 VDD.t2983 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2042 VSS.t253 A[3].t29 a_6071_6357.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2043 VSS.t131 a_30645_5900.t19 a_59548_23692.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2044 a_65651_n1230.t7 a_66063_n1256.t4 a_65769_n1230.t6 VDD.t4172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2045 a_3951_1740.t4 a_3642_11724.t6 VDD.t1051 VDD.t1050 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2046 a_24240_5350.t5 a_24652_5324.t6 a_23081_8962.t3 VDD.t2577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2047 a_23141_8988.t1 opcode[0].t119 VDD.t3948 VDD.t3947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2048 VDD.t1443 A[6].t29 a_41676_11949.t5 VDD.t1442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2049 a_65651_n1230.t10 a_64192_n2074.t9 VDD.t3484 VDD.t3483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2050 VSS.t252 A[3].t30 a_63839_n2274.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2051 VDD.t4553 a_37894_4002.t8 a_38484_3565.t2 VDD.t4552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2052 a_70509_10624.t3 a_63114_21369.t9 a_70509_10506.t4 VDD.t2682 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2053 a_31377_10273.t0 B[1].t13 VSS.t391 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2054 VSS.t187 a_40621_16458.t4 a_41279_15033.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2055 a_60758_18575.t1 a_62366_15449.t8 VDD.t3515 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2056 a_51709_7715.t1 a_51119_8152.t9 VDD.t1288 VDD.t1287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2057 VSS.t545 A[1].t26 a_11505_15751.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2058 VDD.t2313 a_16322_13728.t10 a_16264_14458.t0 VDD.t2312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2059 VDD.t487 a_55504_n1325.t13 a_57736_2352.t5 VDD.t486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2060 a_5108_13805.t0 a_5659_15753.t7 VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2061 VDD.t1165 opcode[1].t75 a_70509_13768.t10 VDD.t1164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2062 VDD.t1913 a_46809_23893.t5 a_48544_24202.t5 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2063 VDD.t3950 opcode[0].t120 a_19357_21596.t3 VDD.t3949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2064 VDD.t3917 opcode[0].t121 a_7365_14454.t4 VDD.t3916 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2065 VDD.t2574 a_43319_23626.t12 a_46233_22680.t0 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2066 VDD.t408 a_38492_9345.t4 a_40227_9654.t2 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2067 Y[0].t3 a_23230_n2148.t9 VSS.t660 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2068 a_59322_18605.t1 a_59616_18579.t6 a_59187_17949.t4 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2069 a_37848_2326.t2 a_41251_9658.t7 VSS.t346 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2070 a_30645_5900.t1 opcode[0].t122 a_31377_6136.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2071 a_44454_746.t4 a_41697_1042.t16 VDD.t1678 VDD.t1677 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2072 VDD.t2612 B[7].t13 a_30150_n3032.t1 VDD.t2611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2073 VDD.t367 a_64185_771.t9 a_67135_3808.t1 VDD.t366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2074 VDD.t1763 a_70513_19926.t9 a_23723_1259.t1 VDD.t1762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2075 VDD.t2803 a_6842_8258.t10 a_6784_8988.t1 VDD.t2802 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2076 a_7375_8988.t2 opcode[0].t123 VDD.t1725 VDD.t1724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2077 VDD.t1444 A[6].t30 a_49328_18695.t0 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2078 VSS.t435 a_35575_3749.t10 a_40035_310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2079 a_49904_21370.t2 a_50316_21344.t6 a_50022_21370.t2 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2080 a_16855_14458.t5 opcode[0].t124 VDD.t1727 VDD.t1726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2081 a_44399_2324.t1 a_67133_11394.t9 VDD.t4543 VDD.t4542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2082 VDD.t4251 a_54454_9678.t7 a_51054_2325.t2 VDD.t4250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2083 a_51699_310.t2 a_51109_747.t7 VDD.t3357 VDD.t3356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2084 VDD.t2636 a_45035_3563.t6 a_46770_3872.t3 VDD.t2635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2085 a_20578_13121.t1 a_19927_14428.t6 VSS.t66 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2086 a_14310_5328.t1 A[5].t28 VDD.t3444 VDD.t3443 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2087 a_19705_1744.t7 a_19396_11720.t6 VDD.t3346 VDD.t3345 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2088 VDD.t4523 a_54713_3294.t11 a_59090_7603.t1 VDD.t4522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2089 a_42177_23622.t1 a_41913_24205.t6 VSS.t224 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2090 VSS.t251 A[3].t31 a_9168_15798.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2091 VDD.t1256 a_44460_6616.t9 a_45050_6179.t1 VDD.t1255 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2092 a_3591_21596.t2 opcode[0].t125 VDD.t1738 VDD.t1737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2093 VSS.t291 B[5].t15 a_63764_8594.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2094 a_45044_309.t2 a_44454_746.t7 VDD.t1585 VDD.t1584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2095 a_66063_3092.t3 a_54908_6842.t13 VSS.t708 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2096 a_7381_20723.t3 opcode[0].t126 VSS.t282 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2097 VDD.t521 a_41611_21373.t11 a_43391_21373.t4 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2098 a_61098_21369.t5 a_30645_5900.t20 VDD.t763 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2099 a_70513_16782.t4 a_70459_17667.t5 a_70513_16900.t8 VDD.t3505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2100 a_65649_10704.t4 a_66061_10678.t7 a_65767_10704.t5 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2101 a_6887_15819.t2 a_6827_15753.t6 VDD.t3379 VDD.t3378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2102 a_51690_3564.t3 a_51100_4001.t9 VSS.t351 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2103 VDD.t4095 a_42301_n1318.t12 a_44445_4000.t1 VDD.t4094 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2104 a_35001_1426.t4 B[3].t20 VDD.t2438 VDD.t2437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2105 a_20054_1744.t7 a_20579_1259.t5 a_19705_1744.t10 VDD.t4598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2106 a_40219_3874.t1 a_38493_311.t5 a_40101_3874.t1 VDD.t752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2107 VDD.t1305 a_56366_23618.t12 a_63408_21343.t2 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2108 a_54658_20633.t1 a_54952_21339.t6 VSS.t478 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2109 VDD.t1414 B[6].t22 a_5794_16410.t1 VDD.t1413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2110 a_16855_14458.t7 a_16795_14432.t5 a_16322_13728.t2 VDD.t1987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2111 a_13358_6047.t1 B[5].t16 VDD.t1822 VDD.t1821 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2112 VDD.t3969 A[2].t19 a_21211_16387.t4 VDD.t3968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2113 a_8192_10387.t1 opcode[1].t76 a_6832_10990.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2114 VDD.t2549 a_59937_9742.t7 a_60201_9159.t2 VDD.t2548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2115 a_59921_1016.t1 a_54903_1041.t18 VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2116 VDD.t4431 a_46350_1040.t12 a_47703_1733.t1 VDD.t4430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2117 VDD.t2966 opcode[2].t34 a_807_1740.t7 VDD.t2965 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2118 a_6832_10990.t5 a_8011_10847.t5 a_7365_11720.t7 VDD.t2523 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2119 VDD.t4594 a_7551_6363.t6 a_19997_8988.t10 VDD.t4593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2120 VDD.t432 B[2].t12 a_19563_6043.t0 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2121 a_25100_20862.t4 a_26279_20719.t7 a_26224_20259.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2122 a_9761_5354.t10 A[7].t18 VDD.t3758 VDD.t3757 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2123 VDD.t418 a_48426_24202.t8 a_48690_23619.t2 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2124 a_20054_1744.t1 a_19146_1744.t4 a_19705_1744.t3 VDD.t2533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2125 VDD.t4452 a_6071_6357.t6 a_13721_8992.t10 VDD.t4451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2126 VDD.t4456 a_64185_771.t10 a_65651_3118.t10 VDD.t4455 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2127 a_54665_15740.t3 a_30643_1763.t17 VDD.t3132 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2128 a_57676_2326.t2 a_67135_3808.t8 VDD.t4069 VDD.t4068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2129 a_43391_21373.t1 a_42964_22066.t6 a_43509_21373.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2130 VDD.t1748 a_59187_17949.t7 a_51813_16162.t2 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2131 a_19987_14454.t4 a_20633_13581.t5 a_19454_13724.t2 VDD.t1956 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2132 VDD.t4161 a_44399_2324.t12 a_48542_1014.t1 VDD.t4160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2133 a_13778_1740.t4 opcode[2].t35 a_14014_407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2134 a_4834_7659.t0 a_4183_8966.t10 VSS.t702 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2135 a_62996_21369.t10 a_63408_21343.t5 a_63114_21369.t5 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2136 a_29954_12048.t1 opcode[0].t127 VDD.t1808 VDD.t1807 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2137 a_65769_n1230.t7 a_66063_n1256.t5 a_65651_n1230.t8 VDD.t4173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2138 a_65769_6613.t4 a_65224_7306.t6 a_65769_5881.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2139 a_42266_11512.t2 a_41676_11949.t8 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2140 VSS.t387 B[3].t21 a_63764_5561.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2141 a_3058_20866.t2 A[6].t31 a_3591_21596.t0 VDD.t1445 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2142 VDD.t1071 a_51059_8126.t11 a_51114_6548.t1 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2143 a_14367_8119.t1 opcode[0].t128 VDD.t1810 VDD.t1809 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2144 a_41515_15033.t1 A[7].t19 VSS.t598 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2145 a_19937_8962.t6 a_21632_6045.t6 a_22172_5352.t10 VDD.t4447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2146 a_56556_20633.t1 a_56850_21339.t4 VSS.t11 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2147 a_19705_1744.t9 a_20579_1259.t6 a_20054_1744.t5 VDD.t3696 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2148 a_54567_3877.t4 a_51704_1914.t5 a_54449_3877.t1 VDD.t3597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2149 a_61197_9746.t1 a_58334_7783.t5 a_61079_9746.t2 VDD.t502 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2150 VSS.t175 a_64188_3841.t8 a_65224_7306.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2151 a_71842_14359.t1 a_56556_21365.t10 VSS.t21 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2152 VSS.t592 a_35594_7027.t11 a_38139_9145.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2153 a_4879_10851.t3 opcode[1].t77 VSS.t195 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2154 VSS.t133 a_48064_9163.t12 a_53241_309.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2155 VDD.t4177 a_41243_3878.t7 a_41507_3295.t3 VDD.t4176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2156 VDD.t4325 opcode[3].t34 a_22322_n2148.t1 VDD.t4324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2157 a_31375_n2138.t0 B[7].t14 VSS.t417 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2158 a_63527_9231.t5 A[3].t32 VDD.t4401 VDD.t4400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2159 a_58321_311.t0 a_57731_748.t9 VDD.t1065 VDD.t1064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2160 a_46644_1014.t2 a_41697_1042.t17 VDD.t1680 VDD.t1679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2161 a_13721_8992.t11 a_6071_6357.t7 VDD.t4454 VDD.t4453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2162 a_15966_5352.t5 A[4].t37 VDD.t2008 VDD.t2007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2163 a_59187_17949.t0 a_59616_18579.t7 a_59322_18605.t0 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2164 a_1089_14458.t3 a_1029_14432.t4 a_556_13728.t0 VDD.t1582 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2165 a_54903_1041.t6 a_54358_1734.t6 a_54903_309.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2166 a_59517_6910.t4 a_55469_11532.t11 VDD.t3413 VDD.t3412 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2167 VDD.t3971 A[2].t20 a_22489_21592.t5 VDD.t3970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2168 VDD.t1447 A[6].t32 a_15297_16387.t5 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2169 a_29954_7911.t0 B[2].t13 VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2170 a_48248_1040.t2 a_47703_1733.t6 a_48248_308.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2171 a_59910_20638.t1 a_59320_21075.t8 VDD.t3524 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2172 a_37903_748.t0 a_37848_2326.t14 VDD.t1950 VDD.t1949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2173 a_58986_15769.t2 a_59280_15743.t6 a_58868_15769.t4 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2174 VSS.t616 a_53713_16459.t4 a_54371_15034.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2175 a_30154_12886.t1 opcode[0].t129 VDD.t3911 VDD.t3910 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2176 VDD.t3913 opcode[0].t130 a_16855_14458.t4 VDD.t3912 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2177 a_15966_5352.t4 a_15426_6045.t6 a_10459_8962.t4 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2178 VDD.t4327 opcode[3].t35 a_9700_n2148.t2 VDD.t4326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2179 a_45805_1733.t1 a_42301_n1318.t13 VDD.t4097 VDD.t4096 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2180 VSS.t477 opcode[2].t36 a_19146_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2181 a_51704_6111.t1 a_51114_6548.t8 VDD.t4549 VDD.t4548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2182 a_19454_13724.t3 a_20633_13581.t6 a_20578_13121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2183 VDD.t3330 a_49314_17045.t8 a_46569_18571.t2 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2184 VDD.t4008 opcode[0].t131 a_3591_21596.t8 VDD.t4007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2185 a_45041_9433.t2 a_44451_9870.t8 VDD.t2821 VDD.t2820 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2186 a_10259_n2148.t3 a_9700_n2148.t7 a_10608_n2148.t4 VDD.t4494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2187 a_43391_21373.t5 a_41611_21373.t12 VDD.t522 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2188 VDD.t764 a_30645_5900.t21 a_61098_21369.t4 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2189 a_13178_13728.t2 a_14357_13585.t6 a_13711_14458.t6 VDD.t2744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2190 a_29952_3774.t1 B[4].t14 VDD.t1864 VDD.t1863 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2191 a_20103_5350.t2 a_20515_5324.t6 a_16805_8966.t2 VDD.t1042 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2192 a_46356_6910.t4 a_46650_6884.t7 a_46238_6910.t6 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2193 a_59325_22679.t6 a_56366_23618.t13 VDD.t1306 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2194 a_71846_20871.t0 opcode[1].t78 a_70513_19926.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2195 a_1628_407.t0 a_248_1740.t6 a_1156_1740.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2196 a_63408_21343.t1 a_56366_23618.t14 VDD.t1307 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2197 a_5794_16410.t0 B[6].t23 VDD.t1416 VDD.t1415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2198 VSS.t355 B[0].t13 a_23700_6043.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2199 VSS.t698 a_6784_8988.t4 a_8192_10387.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2200 VDD.t1824 B[5].t17 a_30150_1105.t0 VDD.t1823 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2201 a_7365_11720.t8 a_8011_10847.t6 a_6832_10990.t6 VDD.t2524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2202 a_59937_9742.t3 a_58329_6179.t5 a_60055_9742.t4 VDD.t175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2203 a_66005_2386.t0 a_64185_771.t11 a_65769_3118.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2204 VDD.t3040 a_70509_n2116.t10 a_1681_1255.t1 VDD.t3039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2205 a_40365_3291.t0 a_40101_3874.t7 VDD.t3121 VDD.t3120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2206 VSS.t675 a_4491_15753.t7 a_1964_13805.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2207 VDD.t1167 opcode[1].t79 a_70459_8189.t1 VDD.t1166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2208 a_54449_3877.t4 a_51704_1914.t6 VSS.t580 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2209 a_43509_21373.t1 a_42964_22066.t7 a_43391_21373.t0 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2210 a_51813_16162.t3 a_59187_17949.t8 VDD.t3158 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2211 a_19454_13724.t4 a_20633_13581.t7 a_19987_14454.t5 VDD.t1957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2212 a_16865_8992.t6 a_6813_6359.t6 VDD.t1697 VDD.t1696 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2213 a_61079_9746.t0 a_58334_7783.t6 VSS.t87 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2214 a_30150_n1593.t3 opcode[0].t132 VDD.t4010 VDD.t4009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2215 a_4879_13585.t3 opcode[0].t133 VSS.t632 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2216 VSS.t117 a_45041_9433.t5 a_46658_9742.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2217 VDD.t3486 a_64192_n2074.t10 a_65224_n537.t1 VDD.t3485 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2218 a_63114_21369.t4 a_63408_21343.t6 a_62996_21369.t9 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2219 a_38506_7695.t3 a_37916_8132.t10 VSS.t470 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2220 VSS.t634 a_38484_3565.t6 a_40101_3874.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2221 VDD.t4508 a_46176_16428.t13 a_45821_15761.t6 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2222 VDD.t165 a_41507_3295.t14 a_44465_8220.t1 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2223 VDD.t114 a_41676_11949.t9 a_42266_11512.t3 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2224 a_3591_21596.t1 A[6].t33 a_3058_20866.t1 VDD.t1448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2225 a_9867_21592.t7 A[4].t38 a_9334_20862.t1 VDD.t2009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2226 VDD.t4305 a_18243_16385.t10 a_10449_14428.t0 VDD.t4304 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2227 a_57722_4002.t0 a_55504_n1325.t14 VDD.t489 VDD.t488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2228 a_39618_16432.t0 a_30643_n2374.t18 a_41515_15033.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2229 a_29954_12048.t7 a_30154_12886.t6 a_30647_12105.t2 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2230 VDD.t4329 opcode[3].t36 a_13461_n2152.t5 VDD.t4328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2231 a_20322_n3481.t0 a_19677_n2174.t6 VSS.t460 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2232 a_10227_1744.t4 a_9668_1744.t6 a_10576_1744.t1 VDD.t562 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2233 a_48418_21344.t3 A[1].t27 VSS.t546 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2234 a_3983_n2152.t2 a_3923_n2178.t7 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2235 a_65769_n1230.t4 a_65224_n537.t4 a_65651_n1230.t3 VDD.t3061 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2236 a_10173_5328.t1 A[7].t20 VDD.t3760 VDD.t3759 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2237 VSS.t709 a_54908_6842.t14 a_66005_2386.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2238 VSS.t250 A[3].t33 a_63835_3641.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2239 a_38501_6091.t2 a_37911_6528.t9 VDD.t2163 VDD.t2162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2240 a_16859_20723.t2 opcode[0].t134 VDD.t4000 VDD.t3999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2241 VDD.t1826 B[5].t18 a_6962_16408.t2 VDD.t1825 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2242 a_556_13728.t1 a_1029_14432.t5 a_1089_14458.t4 VDD.t1583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2243 a_4857_n2637.t2 a_4300_1740.t10 VDD.t2133 VDD.t2132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2244 a_46809_23893.t0 a_46219_24330.t10 VDD.t2639 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2245 a_16605_n2152.t11 a_16545_n2178.t4 VDD.t3527 VDD.t3526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2246 a_22489_21592.t4 A[2].t21 VDD.t3973 VDD.t3972 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2247 a_15297_16387.t4 A[6].t34 VDD.t1450 VDD.t1449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2248 a_39675_15739.t0 a_39618_16432.t9 VDD.t1265 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2249 VDD.t1061 a_64188_3841.t9 a_67135_7303.t2 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2250 VDD.t1169 opcode[1].t80 a_70455_11391.t1 VDD.t1168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2251 VDD.t2968 opcode[2].t37 a_12870_1740.t1 VDD.t2967 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2252 a_7083_1744.t9 a_6524_1744.t4 a_7432_1744.t4 VDD.t3603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2253 VDD.t3925 opcode[0].t135 a_30152_4612.t1 VDD.t3924 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2254 VSS.t217 B[6].t24 a_63832_571.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2255 a_54607_15034.t1 A[5].t29 VSS.t552 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2256 a_58334_7783.t1 a_57744_8220.t8 VDD.t3155 VDD.t3154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2257 Y[3].t2 a_13810_n2152.t9 VDD.t4182 VDD.t4181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2258 a_41697_1042.t3 a_41152_1735.t6 a_41697_310.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2259 a_46140_17941.t0 a_46569_18571.t4 a_46275_18597.t0 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2260 a_51109_747.t2 a_48064_9163.t13 VDD.t781 VDD.t780 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2261 a_14335_n2637.t3 a_13778_1740.t10 VSS.t294 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2262 a_52892_6842.t10 a_52465_7535.t6 a_53010_6842.t6 VDD.t4422 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2263 a_9700_n2148.t1 opcode[3].t37 VDD.t4331 VDD.t4330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2264 a_22709_16385.t0 B[1].t14 VDD.t2463 VDD.t2462 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2265 a_20814_13121.t0 opcode[0].t136 a_19454_13724.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2266 a_53951_18598.t3 a_53891_18572.t7 VDD.t259 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2267 a_46569_18571.t1 a_49314_17045.t9 VDD.t4187 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2268 a_13429_1740.t8 a_13120_11724.t6 VDD.t2283 VDD.t2282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2269 a_3591_21596.t7 opcode[0].t137 VDD.t3927 VDD.t3926 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2270 a_60464_18601.t5 a_60404_18575.t5 VDD.t3187 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2271 VDD.t1728 opcode[0].t138 a_43391_21373.t8 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2272 a_22608_8258.t4 a_23787_8115.t5 a_23732_7655.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2273 VDD.t1308 a_56366_23618.t15 a_59325_22679.t5 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2274 VDD.t2747 a_11565_15824.t4 a_19987_14454.t8 VDD.t2746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2275 VSS.t557 a_62366_15449.t9 a_60758_18575.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2276 VDD.t1292 a_9928_8988.t5 a_10509_11720.t3 VDD.t1291 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2277 a_23466_n3481.t0 a_22821_n2174.t4 VSS.t531 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2278 a_70513_16900.t9 opcode[1].t81 VDD.t1171 VDD.t1170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2279 VSS.t173 a_70509_13650.t9 a_17447_1255.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2280 a_44697_5979.t0 a_42266_11512.t13 a_44460_6616.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2281 a_18153_4620.t0 a_18447_5326.t6 a_13661_8966.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2282 VDD.t1730 opcode[0].t139 a_9867_21592.t3 VDD.t1729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2283 VDD.t1239 a_48855_n1313.t11 a_51100_4001.t6 VDD.t1238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2284 a_59320_21075.t2 A[3].t34 VDD.t4399 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2285 a_29952_n363.t9 opcode[0].t140 VDD.t1732 VDD.t1731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2286 a_51119_8152.t1 a_51059_8126.t12 VDD.t1073 VDD.t1072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2287 a_13810_n2152.t4 opcode[3].t38 a_14046_n3485.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2288 a_12870_1740.t0 opcode[2].t38 VDD.t2970 VDD.t2969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2289 a_19948_20263.t0 A[1].t28 VSS.t547 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2290 VDD.t1866 B[4].t15 a_8130_16410.t1 VDD.t1865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2291 a_39381_15765.t5 a_38723_16458.t5 a_39263_15765.t7 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2292 a_35249_9412.t1 A[4].t39 a_35012_10049.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2293 a_46232_1040.t4 a_42301_n1318.t14 VDD.t4099 VDD.t4098 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2294 a_7956_13121.t1 a_7305_14428.t7 VSS.t32 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2295 a_30152_n964.t1 B[6].t25 VDD.t1418 VDD.t1417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2296 a_46219_24330.t2 A[1].t29 VDD.t3401 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2297 a_51105_9802.t4 a_48815_11511.t13 VDD.t2275 VDD.t2274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2298 a_51704_1914.t3 a_51114_2351.t8 VSS.t174 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2299 a_66063_3092.t1 a_54908_6842.t15 VDD.t4577 VDD.t4576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2300 a_62996_21369.t8 a_63408_21343.t7 a_63114_21369.t3 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2301 a_54658_21365.t1 a_54113_22058.t6 a_54658_20633.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2302 a_42266_11512.t0 a_41676_11949.t10 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2303 a_18243_16385.t2 B[4].t16 VDD.t1868 VDD.t1867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2304 VSS.t521 a_12672_15792.t6 a_12732_15818.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2305 VDD.t1173 opcode[1].t82 a_70455_14535.t1 VDD.t1172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2306 a_10812_411.t0 a_9918_11720.t6 VSS.t54 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2307 a_53571_3290.t3 a_53307_3873.t7 VSS.t510 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2308 a_48490_6178.t0 a_46356_6910.t10 a_48254_6910.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2309 a_41279_15033.t1 a_41573_15739.t4 a_39618_16432.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2310 a_67135_n540.t1 a_48248_1040.t13 VDD.t4232 VDD.t4231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2311 a_11155_13581.t3 opcode[0].t141 VSS.t611 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2312 a_20086_n2148.t7 opcode[3].t39 a_20322_n3481.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2313 VDD.t3297 a_45279_16157.t13 a_49314_17045.t2 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2314 a_16795_16385.t2 B[5].t19 VDD.t1828 VDD.t1827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2315 a_29950_n2431.t7 a_30150_n3032.t5 a_30643_n2374.t2 VDD.t4117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2316 a_63527_6198.t2 A[4].t40 VDD.t2011 VDD.t2010 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2317 a_10513_20719.t3 opcode[0].t142 VSS.t612 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2318 a_22881_n2148.t11 a_22322_n2148.t4 a_23230_n2148.t6 VDD.t1917 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2319 a_48265_n1750.t2 B[5].t20 VDD.t1830 VDD.t1829 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2320 a_24652_5324.t3 A[0].t18 VSS.t370 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2321 a_11829_5352.t7 a_11289_6045.t6 a_4183_8966.t1 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2322 a_65651_n1230.t0 a_65224_n537.t5 a_65769_n1230.t0 VDD.t1326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2323 a_22540_11720.t1 a_22598_10990.t9 VDD.t1157 VDD.t1156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2324 a_46350_308.t1 a_46644_1014.t6 VSS.t273 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2325 a_1089_14458.t5 a_1029_14432.t6 a_556_13728.t2 VDD.t2486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2326 VSS.t218 B[6].t26 a_30152_n964.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2327 a_19737_n2148.t10 opcode[3].t40 VDD.t4333 VDD.t4332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2328 a_64117_8794.t3 a_63527_9231.t10 VSS.t397 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2329 a_1974_8339.t2 A[7].t21 VDD.t3762 VDD.t3761 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2330 VDD.t2530 a_16545_n2178.t5 a_16605_n2152.t10 VDD.t2529 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2331 VDD.t1452 A[6].t35 a_15297_16387.t3 VDD.t1451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2332 VDD.t3531 a_44459_2350.t8 a_45049_1913.t3 VDD.t3530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2333 VDD.t1266 a_39618_16432.t10 a_39675_15739.t1 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2334 a_19987_11720.t1 a_19406_8988.t6 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2335 VSS.t445 a_9976_10990.t9 a_9918_11720.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2336 a_46776_9742.t1 a_45041_9433.t6 VDD.t660 VDD.t659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2337 a_17446_10391.t1 a_16264_14458.t6 VSS.t89 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2338 a_10472_16406.t0 B[2].t14 VDD.t436 VDD.t435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2339 VDD.t483 a_13178_10994.t11 a_13120_11724.t3 VDD.t482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2340 a_71846_5105.t1 opcode[1].t83 a_70513_4160.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2341 a_13711_14458.t9 a_13651_14432.t4 a_13178_13728.t5 VDD.t3785 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2342 a_52710_16433.t4 a_30643_1763.t18 a_54607_15034.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2343 VDD.t1914 a_46809_23893.t6 a_48544_24202.t4 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2344 VDD.t4184 a_13810_n2152.t10 Y[3].t1 VDD.t4183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2345 a_46275_18597.t1 a_46569_18571.t5 a_46140_17941.t1 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2346 VSS.t51 a_5659_15753.t8 a_5108_13805.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2347 VDD.t3078 opcode[3].t41 a_9700_n2148.t0 VDD.t3077 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2348 a_46233_15735.t3 a_46176_16428.t14 VSS.t701 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2349 VSS.t442 a_11565_15824.t5 a_20814_13121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2350 a_54454_9678.t3 a_51709_7715.t5 a_54572_9678.t3 VDD.t2790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2351 VDD.t4188 a_49314_17045.t10 a_46569_18571.t0 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2352 a_14357_13585.t2 opcode[0].t143 VDD.t3841 VDD.t3840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2353 a_43803_21347.t2 opcode[0].t144 VDD.t3804 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2354 VDD.t3188 a_60404_18575.t6 a_60464_18601.t4 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2355 a_7115_n2148.t11 a_6556_n2148.t7 a_7464_n2148.t7 VDD.t4180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2356 a_566_8262.t4 a_1745_8119.t6 a_1099_8992.t6 VDD.t1562 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2357 a_70509_n2116.t2 a_39381_15765.t11 a_70509_n1998.t0 VDD.t578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2358 a_55116_11332.t1 A[6].t36 a_54879_11969.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2359 a_10509_11720.t4 a_9928_8988.t6 VDD.t1294 VDD.t1293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2360 VDD.t3713 a_35594_7027.t12 a_37902_9782.t5 VDD.t3712 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2361 a_23230_n2148.t3 opcode[3].t42 a_23466_n3481.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2362 a_35575_3749.t2 a_34985_4186.t10 VDD.t1570 VDD.t1569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2363 VDD.t350 a_19464_8258.t10 a_19406_8988.t1 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2364 a_16865_8992.t11 opcode[0].t145 VDD.t3806 VDD.t3805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2365 a_70509_n1998.t7 opcode[1].t84 VDD.t1175 VDD.t1174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2366 a_64117_5761.t3 a_63527_6198.t10 VSS.t204 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2367 a_24240_5350.t0 a_24652_5324.t7 a_23081_8962.t0 VDD.t1421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2368 a_48548_6884.t1 a_44405_8194.t13 VDD.t245 VDD.t244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2369 a_70513_7304.t6 a_70459_8189.t6 a_70513_7422.t7 VDD.t3243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2370 a_13711_11724.t0 opcode[1].t85 VDD.t1177 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2371 VDD.t4590 a_61071_3878.t7 a_57684_8194.t3 VDD.t4589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2372 a_65651_n1230.t4 a_48248_1040.t14 VDD.t4234 VDD.t4233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2373 a_6735_21596.t11 A[7].t22 VDD.t3764 VDD.t3763 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2374 a_41161_15765.t5 a_41573_15739.t5 a_39618_16432.t7 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2375 a_60766_15769.t5 a_61178_15743.t5 a_59223_16436.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2376 a_14282_n3485.t0 a_12902_n2152.t5 a_13810_n2152.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2377 a_59509_1042.t0 a_55504_n1325.t15 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2378 a_4233_14458.t3 a_4173_14432.t5 a_3700_13728.t4 VDD.t1012 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2379 VSS.t686 a_23723_1259.t6 a_23670_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2380 a_40310_22246.t0 a_39720_22683.t9 VDD.t3698 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2381 VSS.t198 a_48855_n1313.t12 a_51351_1714.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2382 VDD.t187 A[1].t30 a_46219_24330.t1 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2383 a_6887_15819.t1 a_6827_15753.t7 VDD.t3381 VDD.t3380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2384 VDD.t2451 a_15297_16387.t7 a_4173_14432.t2 VDD.t2450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2385 a_49686_24206.t4 a_48690_23619.t6 VDD.t3601 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2386 a_54894_20633.t1 a_30647_7968.t11 a_54658_21365.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2387 a_70509_10506.t1 a_70455_11391.t6 a_70509_10624.t6 VDD.t2838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2388 VDD.t410 a_38492_9345.t5 a_40227_9654.t1 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2389 a_47709_7603.t1 a_46356_6910.t11 VDD.t2647 VDD.t2646 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2390 a_59262_18579.t2 a_60329_17945.t6 VDD.t1032 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2391 VDD.t3975 A[2].t22 a_21211_16387.t3 VDD.t3974 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2392 a_70455_1913.t0 opcode[1].t86 VDD.t1179 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2393 a_13778_1740.t1 a_12870_1740.t5 a_13429_1740.t0 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2394 a_66061_10678.t2 a_64117_8794.t6 VDD.t2559 VDD.t2558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2395 VDD.t3614 a_39582_17945.t7 Cout.t1 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2396 VDD.t3976 A[2].t23 a_52753_24325.t2 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2397 a_6202_20866.t2 a_7381_20723.t5 a_6735_21596.t2 VDD.t4148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2398 a_49314_17045.t1 a_45279_16157.t14 VDD.t3298 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2399 VDD.t1832 B[5].t21 a_16795_16385.t1 VDD.t1831 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2400 a_17446_13125.t0 a_16795_14432.t6 VSS.t318 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2401 VSS.t664 a_48248_1040.t15 a_66005_n1962.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2402 a_13178_10994.t6 a_13120_14458.t5 a_13711_11724.t10 VDD.t3929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2403 VDD.t1834 B[5].t22 a_48265_n1750.t1 VDD.t1833 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2404 VDD.t2440 B[3].t22 a_30152_5242.t1 VDD.t2439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2405 a_65769_n1230.t1 a_65224_n537.t6 a_65651_n1230.t1 VDD.t1327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2406 a_54785_1041.t9 a_53005_1041.t12 VDD.t4255 VDD.t4254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2407 a_40035_310.t0 a_35591_989.t16 a_39799_1042.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2408 VDD.t4202 a_59325_22679.t10 a_59915_22242.t0 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2409 a_56438_21365.t0 a_54658_21365.t13 VDD.t882 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2410 a_35012_10049.t3 A[4].t41 VDD.t2013 VDD.t2012 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2411 VDD.t6 a_40365_3291.t5 a_41361_3878.t1 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2412 a_61415_6910.t1 a_59635_6910.t11 VDD.t888 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2413 a_4182_20263.t0 A[6].t37 VSS.t225 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2414 VDD.t1159 a_22598_10990.t10 a_22540_11720.t0 VDD.t1158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2415 VDD.t2888 a_47794_3876.t8 a_44405_8194.t3 VDD.t2887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2416 a_59635_6910.t1 a_59929_6884.t6 a_59517_6910.t7 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2417 a_10519_8988.t1 opcode[0].t146 VDD.t3808 VDD.t3807 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2418 VSS.t428 a_13188_8262.t9 a_13130_8992.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2419 VDD.t3571 a_9986_8258.t10 a_9928_8988.t1 VDD.t3570 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2420 VDD.t3080 opcode[3].t43 a_19737_n2148.t9 VDD.t3079 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2421 VDD.t3073 a_57736_2352.t10 a_58326_1915.t0 VDD.t3072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2422 a_16605_n2152.t9 a_16545_n2178.t6 VDD.t2532 VDD.t2531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2423 VDD.t2175 a_37856_8106.t14 a_41999_6796.t1 VDD.t2174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2424 VDD.t38 a_19406_8988.t7 a_19987_11720.t2 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2425 a_63598_4278.t2 B[4].t17 VDD.t1870 VDD.t1869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2426 a_3710_8262.t0 a_4183_8966.t11 a_4243_8992.t4 VDD.t4516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2427 a_60193_3291.t1 a_59929_3874.t7 VDD.t4511 VDD.t4510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2428 a_10337_15751.t4 A[2].t24 a_10472_16406.t4 VDD.t3977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2429 VDD.t2465 B[1].t15 a_30152_9379.t1 VDD.t2464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2430 a_54371_15034.t0 a_54665_15740.t6 a_52710_16433.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2431 a_48544_24202.t3 a_46809_23893.t7 VDD.t2640 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2432 VDD.t3715 a_35594_7027.t13 a_37916_8132.t5 VDD.t3714 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2433 VDD.t2972 opcode[2].t39 a_19146_1744.t1 VDD.t2971 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2434 a_13429_1740.t1 a_12870_1740.t6 a_13778_1740.t2 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2435 a_5659_15753.t0 B[6].t27 VSS.t219 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2436 a_64122_11365.t1 a_63532_11802.t8 VDD.t2114 VDD.t2113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2437 a_24157_16385.t2 B[0].t14 VDD.t2215 VDD.t2214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2438 a_42301_n1318.t3 a_41711_n1755.t10 VSS.t373 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2439 VSS.t484 a_58320_9433.t5 a_59937_9742.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2440 VDD.t3123 a_39807_6822.t12 a_41160_7515.t1 VDD.t3122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2441 a_22881_n2148.t8 a_22821_n2174.t5 VDD.t3320 VDD.t3319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2442 VDD.t2764 a_9976_10990.t10 a_9918_11720.t1 VDD.t2763 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2443 VDD.t1241 a_48855_n1313.t13 a_51114_2351.t5 VDD.t1240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2444 a_61510_21343.t2 A[3].t35 VDD.t4398 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2445 VDD.t3848 opcode[0].t147 a_43803_21347.t1 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2446 a_60464_18601.t3 a_60404_18575.t7 VDD.t3189 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2447 a_23131_11720.t2 opcode[1].t87 VDD.t1181 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2448 VDD.t3082 opcode[3].t44 a_7115_n2148.t5 VDD.t3081 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2449 VDD.t1682 a_41697_1042.t18 a_44454_746.t3 VDD.t1681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2450 VDD.t3445 A[5].t30 a_53713_16459.t0 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2451 VDD.t838 opcode[2].t40 a_19705_1744.t1 VDD.t837 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2452 a_47282_17937.t2 a_47711_18567.t5 a_47417_18593.t5 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2453 VSS.t220 B[6].t28 a_55116_11332.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2454 a_4243_8992.t10 a_4889_8119.t7 a_3710_8262.t7 VDD.t3649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2455 Y[1].t2 a_20086_n2148.t8 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2456 a_23702_n3481.t1 a_22322_n2148.t5 a_23230_n2148.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2457 a_43803_21347.t3 opcode[0].t148 VSS.t613 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2458 VDD.t4484 a_6784_8988.t5 a_7365_11720.t2 VDD.t4483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2459 a_65222_11397.t1 a_41705_6822.t17 VDD.t3631 VDD.t3630 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2460 VDD.t3850 opcode[0].t149 a_10519_8988.t0 VDD.t3849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2461 VDD.t1375 a_52710_16433.t11 a_52767_15740.t1 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2462 a_39799_310.t0 a_40093_1016.t5 VSS.t700 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2463 a_41611_21373.t3 a_41066_22066.t5 a_41493_21373.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2464 a_47719_15761.t4 A[6].t38 VDD.t1453 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2465 VDD.t1183 opcode[1].t88 a_13711_11724.t1 VDD.t1182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2466 a_52355_15766.t11 a_52767_15740.t6 a_52473_15766.t7 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2467 a_40310_22246.t3 a_39720_22683.t10 VSS.t590 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2468 a_59223_16436.t2 a_61178_15743.t6 a_60766_15769.t4 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2469 a_57730_9870.t1 a_55469_11532.t12 VDD.t1561 VDD.t1560 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2470 a_9761_5354.t2 a_10173_5328.t6 a_1039_8966.t2 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2471 VSS.t669 a_14335_n2637.t5 a_14282_n3485.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2472 a_35001_1426.t0 A[6].t39 VDD.t1455 VDD.t1454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2473 a_20515_5324.t3 A[2].t25 VSS.t628 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2474 a_54567_3877.t1 a_53571_3290.t6 VDD.t2860 VDD.t2859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2475 a_46219_24330.t0 A[1].t31 VDD.t188 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2476 VDD.t3383 a_6827_15753.t8 a_6887_15819.t0 VDD.t3382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2477 VSS.t620 a_30154_11447.t6 a_31379_12105.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2478 VDD.t2467 B[1].t16 a_22172_5352.t2 VDD.t2466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2479 VDD.t840 opcode[2].t41 a_807_1740.t6 VDD.t839 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2480 a_63408_21343.t0 a_56366_23618.t16 VDD.t1309 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2481 a_71842_11451.t1 opcode[1].t89 a_70509_10506.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2482 a_53576_9091.t1 a_53312_9674.t7 VDD.t1629 VDD.t1628 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2483 a_37903_748.t5 a_35575_3749.t11 VDD.t2712 VDD.t2711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2484 VSS.t1 a_40365_3291.t6 a_41243_3878.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2485 VSS.t629 A[2].t26 a_54894_20633.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2486 a_16322_13728.t3 a_16795_14432.t7 a_16855_14458.t8 VDD.t1988 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2487 a_23777_10847.t2 opcode[1].t90 VDD.t1185 VDD.t1184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2488 VDD.t1033 a_60329_17945.t7 a_59262_18579.t1 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2489 a_6842_8258.t2 a_8021_8115.t5 a_7375_8988.t6 VDD.t2745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2490 Y[2].t0 a_16954_n2152.t10 VDD.t1975 VDD.t1974 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2491 a_29952_n363.t7 a_30152_475.t6 a_30645_n306.t4 VDD.t533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2492 a_51704_1914.t1 a_51114_2351.t9 VDD.t1045 VDD.t1044 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2493 a_16573_1740.t10 a_16014_1740.t7 a_16922_1740.t5 VDD.t3521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2494 VSS.t439 a_51695_9365.t6 a_53312_9674.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2495 a_16605_n2152.t8 a_16046_n2152.t5 a_16954_n2152.t7 VDD.t3645 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2496 a_23723_1259.t0 a_70513_19926.t10 VDD.t1765 VDD.t1764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2497 a_40101_6796.t1 a_35602_9612.t11 VDD.t4349 VDD.t4348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2498 VDD.t4034 opcode[0].t150 a_17501_13585.t1 VDD.t4033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2499 a_41697_1042.t1 a_41991_1016.t7 a_41579_1042.t9 VDD.t769 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2500 a_6735_21596.t1 a_7381_20723.t6 a_6202_20866.t1 VDD.t4149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2501 a_16795_16385.t0 B[5].t23 VDD.t1836 VDD.t1835 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2502 a_65769_n1962.t1 a_66063_n1256.t6 VSS.t264 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2503 a_13711_11724.t11 a_13120_14458.t6 a_13178_10994.t7 VDD.t3930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2504 VDD.t1838 B[5].t24 a_41711_n1755.t2 VDD.t1837 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2505 a_48265_n1750.t0 B[5].t25 VDD.t1840 VDD.t1839 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2506 VDD.t3447 A[5].t31 a_54914_n1762.t4 VDD.t3446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2507 a_61518_24201.t1 a_59910_20638.t5 VSS.t70 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2508 VDD.t4479 a_12732_15818.t7 a_23131_14454.t11 VDD.t4478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2509 a_70513_16900.t1 a_50022_21370.t9 a_70513_16782.t1 VDD.t1270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2510 VDD.t1842 B[5].t26 a_48225_11948.t2 VDD.t1841 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2511 VDD.t4036 opcode[0].t151 a_1745_8119.t3 VDD.t4035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2512 VDD.t4525 a_54713_3294.t12 a_57730_9870.t6 VDD.t4524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2513 VSS.t687 a_46350_1040.t13 a_47703_1733.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2514 VDD.t2894 a_70513_7304.t10 a_11101_1259.t0 VDD.t2893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2515 a_3058_20866.t4 a_4237_20723.t4 a_4182_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2516 a_19937_8962.t5 a_22584_5326.t7 a_22172_5352.t9 VDD.t3176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2517 a_15966_5352.t9 a_16378_5326.t5 a_10459_8962.t2 VDD.t1954 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2518 VDD.t1128 a_53571_3290.t7 a_54567_3877.t0 VDD.t1127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2519 a_51704_6111.t0 a_51114_6548.t9 VDD.t3502 VDD.t3501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2520 a_12478_20862.t5 a_13657_20719.t5 a_13011_21592.t6 VDD.t2033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2521 VDD.t2850 a_64122_11365.t6 a_70513_20044.t9 VDD.t2849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2522 VDD.t1577 a_1156_1740.t10 a_1713_n2637.t0 VDD.t1576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2523 VDD.t1631 a_53312_9674.t8 a_53576_9091.t0 VDD.t1630 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2524 a_63595_1208.t4 A[4].t42 VDD.t2015 VDD.t2014 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2525 a_70459_5045.t0 opcode[1].t91 VDD.t1187 VDD.t1186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2526 a_10472_16406.t3 A[2].t27 a_10337_15751.t3 VDD.t3978 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2527 VDD.t3599 a_21211_16387.t7 a_16795_14432.t3 VDD.t3598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2528 a_63527_9231.t4 A[3].t36 VDD.t4397 VDD.t4396 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2529 a_53005_309.t1 a_53299_1015.t6 VSS.t695 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2530 a_30152_4612.t3 opcode[0].t152 VSS.t636 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2531 a_46644_1014.t1 a_41697_1042.t19 VDD.t1684 VDD.t1683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2532 a_3700_13728.t1 a_4879_13585.t5 a_4233_14458.t0 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2533 a_20103_5350.t0 B[2].t15 VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2534 a_70459_17667.t0 opcode[1].t92 VDD.t1189 VDD.t1188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2535 a_23198_1744.t0 opcode[2].t42 a_23434_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2536 VDD.t2666 a_51690_3564.t6 a_53425_3873.t1 VDD.t2665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2537 VDD.t2992 a_58320_9433.t6 a_60055_9742.t1 VDD.t2991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2538 VSS.t671 a_53005_1041.t13 a_54358_1734.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2539 VDD.t842 opcode[2].t43 a_16573_1740.t7 VDD.t841 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2540 VDD.t3765 A[7].t23 a_42770_18699.t2 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2541 a_23722_10387.t0 a_22540_14454.t6 VSS.t711 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2542 VDD.t1191 opcode[1].t93 a_23131_11720.t1 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2543 a_7115_n2148.t4 opcode[3].t45 VDD.t3084 VDD.t3083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2544 a_41705_6822.t5 a_41160_7515.t5 a_41587_6822.t10 VDD.t3612 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2545 a_10509_14454.t3 opcode[0].t153 VDD.t3942 VDD.t3941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2546 a_70513_4160.t2 a_52473_15766.t10 a_70513_4278.t2 VDD.t664 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2547 VDD.t3944 opcode[0].t154 a_29954_12048.t0 VDD.t3943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2548 VDD.t4218 a_20086_n2148.t9 Y[1].t1 VDD.t4217 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2549 VSS.t697 a_23755_n2633.t7 a_23702_n3481.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2550 a_70513_4278.t4 a_61525_1042.t9 VDD.t1608 VDD.t1607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2551 a_52767_15740.t0 a_52710_16433.t12 VDD.t1376 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2552 VDD.t2520 a_49568_24206.t6 a_49832_23623.t1 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2553 a_13711_11724.t2 opcode[1].t94 VDD.t1193 VDD.t1192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2554 a_45041_9433.t1 a_44451_9870.t9 VDD.t2823 VDD.t2822 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2555 VDD.t2342 a_70509_10506.t10 a_14303_1255.t2 VDD.t2341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2556 a_20003_20723.t2 opcode[0].t155 VDD.t3946 VDD.t3945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2557 a_61098_21369.t11 a_61510_21343.t5 a_61216_21369.t7 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2558 a_1188_n2152.t4 a_1713_n2637.t5 a_839_n2152.t7 VDD.t2358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2559 a_41705_6090.t1 a_41999_6796.t6 VSS.t159 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2560 VDD.t4562 a_59223_16436.t14 a_58868_15769.t0 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2561 a_62366_15449.t0 A[4].t43 a_63015_14838.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2562 VDD.t3663 a_39799_1042.t12 a_41152_1735.t1 VDD.t3662 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2563 VSS.t451 a_65769_6613.t10 a_71846_17727.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2564 a_48815_11511.t1 a_48225_11948.t8 VSS.t689 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2565 a_58321_311.t3 a_57731_748.t10 VSS.t176 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2566 a_58320_9433.t3 a_57730_9870.t10 VSS.t96 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2567 VDD.t3686 a_16274_8992.t5 a_16855_11724.t10 VDD.t3685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2568 a_4593_6357.t0 A[5].t32 VDD.t3449 VDD.t3448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2569 a_59262_18579.t0 a_60329_17945.t8 VDD.t1034 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2570 VSS.t456 a_19454_13724.t11 a_19396_14454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2571 VDD.t3672 a_13849_16387.t7 a_1029_14432.t2 VDD.t3671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2572 a_48462_11311.t1 A[5].t33 a_48225_11948.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2573 VDD.t440 B[2].t16 a_29954_7911.t1 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2574 VDD.t3980 A[2].t28 a_6813_6359.t1 VDD.t3979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2575 a_16954_n2152.t6 a_16046_n2152.t6 a_16605_n2152.t7 VDD.t3646 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2576 a_63602_n1637.t0 B[6].t29 VDD.t1420 VDD.t1419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2577 VDD.t47 a_3855_6357.t6 a_4243_8992.t1 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2578 VDD.t4403 A[3].t37 a_19763_16387.t0 VDD.t4402 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2579 a_17501_13585.t0 opcode[0].t156 VDD.t1782 VDD.t1781 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2580 a_23755_n2633.t1 a_23198_1744.t9 VDD.t3789 VDD.t3788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2581 a_70513_7422.t9 opcode[1].t95 VDD.t1195 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2582 a_41711_n1755.t1 B[5].t27 VDD.t1844 VDD.t1843 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2583 a_54914_n1762.t5 A[5].t34 VDD.t3451 VDD.t3450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2584 a_4233_11724.t5 a_4879_10851.t6 a_3700_10994.t2 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2585 a_59082_1735.t0 a_55504_n1325.t16 VDD.t493 VDD.t492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2586 a_53352_20634.t3 a_52762_21071.t8 VSS.t498 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2587 VDD.t4214 a_23230_n2148.t10 Y[0].t1 VDD.t4213 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2588 a_4237_20723.t0 opcode[0].t157 VDD.t1784 VDD.t1783 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2589 a_48225_11948.t1 B[5].t28 VDD.t1846 VDD.t1845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2590 a_7904_411.t0 a_6524_1744.t5 a_7432_1744.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2591 a_70513_7304.t2 a_58986_15769.t9 a_70513_7422.t2 VDD.t1114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2592 VDD.t2016 A[4].t44 a_62375_18703.t3 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2593 a_61189_3878.t1 a_58326_1915.t5 a_61071_3878.t2 VDD.t3075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2594 a_4889_8119.t2 opcode[0].t158 VDD.t1786 VDD.t1785 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2595 VSS.t566 a_51815_16459.t7 a_52473_15034.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2596 a_29954_7911.t2 opcode[0].t159 VDD.t2037 VDD.t2036 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2597 a_13011_21592.t7 a_13657_20719.t6 a_12478_20862.t6 VDD.t2034 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2598 a_16855_11724.t6 opcode[1].t96 VDD.t1197 VDD.t1196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2599 VDD.t4413 A[3].t38 a_59311_24329.t5 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2600 VSS.t462 a_64122_11365.t7 a_71846_20871.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2601 a_29954_7911.t6 a_30154_7310.t7 a_30647_7968.t3 VDD.t1423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2602 VDD.t1038 a_70509_13650.t10 a_17447_1255.t1 VDD.t1037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2603 a_55197_1015.t1 a_51054_2325.t15 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2604 VDD.t1147 a_64117_5761.t11 a_66063_6587.t1 VDD.t1146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2605 a_57967_9233.t1 a_55469_11532.t13 a_57730_9870.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2606 a_48131_15735.t2 a_30645_n306.t13 VDD.t3106 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2607 a_9304_16408.t5 B[3].t23 VDD.t2442 VDD.t2441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2608 a_39799_1042.t3 a_39254_1735.t5 a_39681_1042.t7 VDD.t1969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2609 a_46176_16428.t4 a_48131_15735.t5 a_47719_15761.t1 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2610 a_53005_1041.t7 a_53299_1015.t7 a_52887_1041.t11 VDD.t4473 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2611 a_6962_16408.t1 B[5].t29 VDD.t1848 VDD.t1847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2612 VDD.t1587 a_44454_746.t8 a_45044_309.t1 VDD.t1586 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2613 VDD.t604 a_67135_7303.t10 a_37856_8106.t0 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2614 a_42770_18699.t1 A[7].t24 VDD.t3766 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2615 a_22598_10990.t2 a_23777_10847.t6 a_23722_10387.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2616 a_45055_7783.t1 a_44465_8220.t8 VDD.t2833 VDD.t2832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2617 a_61525_310.t0 a_61819_1016.t6 VSS.t286 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2618 a_54358_1734.t1 a_53005_1041.t14 VDD.t4266 VDD.t4265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2619 VSS.t153 a_35602_9612.t12 a_40043_6090.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2620 a_29952_5843.t4 a_30152_6681.t6 a_30645_5900.t4 VDD.t2641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2621 a_23131_11720.t0 opcode[1].t97 VDD.t1199 VDD.t1198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2622 a_60988_7603.t1 a_59635_6910.t12 VDD.t890 VDD.t889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2623 VDD.t3102 a_52762_21071.t9 a_53352_20634.t1 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2624 a_9976_13724.t6 a_11155_13581.t5 a_10509_14454.t7 VDD.t3565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2625 a_556_10994.t5 a_1735_10851.t4 a_1089_11724.t7 VDD.t3165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2626 a_45044_309.t3 a_44454_746.t9 VSS.t262 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2627 Y[1].t0 a_20086_n2148.t10 VDD.t4220 VDD.t4219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2628 a_29952_3774.t11 a_30152_4612.t7 a_30645_3831.t7 VDD.t1433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2629 VSS.t31 A[1].t32 a_48360_20638.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2630 a_52892_6842.t7 a_53304_6816.t5 a_53010_6842.t2 VDD.t2519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2631 a_66063_3092.t0 a_54908_6842.t16 VDD.t4579 VDD.t4578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2632 a_48073_15029.t0 A[6].t40 VSS.t226 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2633 VSS.t583 a_39799_1042.t13 a_41152_1735.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2634 a_49832_23623.t2 a_49568_24206.t7 VDD.t2521 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2635 a_19357_21596.t7 A[3].t39 VDD.t4412 VDD.t4411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2636 a_51351_5911.t1 a_48815_11511.t14 a_51114_6548.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2637 VDD.t1898 a_60193_3291.t6 a_61189_3878.t3 VDD.t1897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2638 a_48254_6178.t1 a_48548_6884.t6 VSS.t644 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2639 VDD.t2039 opcode[0].t160 a_20003_20723.t1 VDD.t2038 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2640 a_30154_8749.t1 opcode[0].t161 VDD.t2041 VDD.t2040 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2641 a_7562_20263.t0 opcode[0].t162 a_6202_20866.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2642 VDD.t3864 a_65769_n1230.t11 a_70509_10624.t0 VDD.t3863 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2643 a_19464_8258.t5 a_20643_8115.t7 a_19997_8988.t3 VDD.t4533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2644 a_71842_1737.t0 a_45939_15761.t10 VSS.t112 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2645 a_34985_4186.t4 A[5].t35 VDD.t3453 VDD.t3452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2646 a_31377_n306.t1 a_30152_475.t7 a_30645_n306.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2647 a_47912_3876.t3 a_45049_1913.t7 a_47794_3876.t0 VDD.t2728 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2648 VDD.t2177 a_37856_8106.t15 a_41587_6822.t1 VDD.t2176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2649 VSS.t704 a_54713_3294.t13 a_57967_9233.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2650 a_20515_5324.t1 A[2].t29 VDD.t3982 VDD.t3981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2651 a_29952_n363.t3 a_30152_n964.t7 a_30645_n306.t0 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2652 VDD.t2714 a_35575_3749.t12 a_37894_4002.t5 VDD.t2713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2653 a_63527_6198.t5 B[3].t24 VDD.t4120 VDD.t4119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2654 a_13461_n2152.t9 a_14335_n2637.t6 a_13810_n2152.t6 VDD.t4248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2655 VDD.t624 a_54903_1041.t19 a_59509_1042.t9 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2656 VDD.t1243 a_48855_n1313.t14 a_51100_4001.t5 VDD.t1242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2657 VSS.t292 B[5].t30 a_48462_11311.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2658 a_1099_8992.t1 a_1039_8966.t10 a_566_8262.t1 VDD.t499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2659 VDD.t4410 A[3].t40 a_63602_n1637.t6 VDD.t4409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2660 a_54540_21365.t0 a_30647_7968.t12 VDD.t333 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2661 VDD.t1267 a_39618_16432.t11 a_39263_15765.t0 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2662 a_53241_309.t0 a_48855_n1313.t15 a_53005_1041.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2663 VSS.t97 a_61533_6910.t9 a_71842_1973.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2664 a_30152_4612.t0 opcode[0].t163 VDD.t2043 VDD.t2042 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2665 VDD.t2217 B[0].t15 a_24240_5350.t1 VDD.t2216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2666 VSS.t236 a_30647_12105.t13 a_41066_22066.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2667 a_1089_14458.t2 opcode[0].t164 VDD.t2045 VDD.t2044 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2668 a_23755_n2633.t3 a_23198_1744.t10 VSS.t603 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2669 VSS.t293 B[5].t31 a_13358_6047.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2670 VDD.t3455 A[5].t36 a_54914_n1762.t6 VDD.t3454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2671 a_61533_6910.t3 a_60988_7603.t6 a_61415_6910.t5 VDD.t1859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2672 a_3700_10994.t3 a_4879_10851.t7 a_4233_11724.t4 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2673 a_22608_8258.t5 a_23081_8962.t10 a_23141_8988.t9 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2674 VDD.t1850 B[5].t32 a_48225_11948.t0 VDD.t1849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2675 a_67135_n540.t0 a_48248_1040.t16 VDD.t2872 VDD.t2871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2676 Y[0].t0 a_23230_n2148.t11 VDD.t4216 VDD.t4215 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2677 VDD.t1705 a_57676_2326.t12 a_57731_748.t2 VDD.t1704 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2678 a_42177_23622.t2 a_41913_24205.t7 VDD.t1434 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2679 a_61407_1042.t5 a_61819_1016.t7 a_61525_1042.t0 VDD.t1773 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2680 VDD.t3457 A[5].t37 a_34985_4186.t3 VDD.t3456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2681 a_13721_8992.t2 opcode[0].t165 VDD.t2047 VDD.t2046 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2682 VSS.t599 A[7].t25 a_1974_8339.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2683 VDD.t3665 a_39799_1042.t14 a_41579_1042.t0 VDD.t3664 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2684 a_16322_10994.t3 a_17501_10851.t4 a_16855_11724.t4 VDD.t1026 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2685 VDD.t2628 a_53576_9091.t6 a_54572_9678.t0 VDD.t2627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2686 VDD.t3984 A[2].t30 a_20515_5324.t0 VDD.t3983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2687 a_59311_24329.t4 A[3].t41 VDD.t4408 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2688 VDD.t523 a_41611_21373.t13 a_42964_22066.t0 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2689 a_5060_10391.t0 opcode[1].t98 a_3700_10994.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2690 a_54658_21365.t2 a_54113_22058.t7 a_54540_21365.t3 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2691 a_37894_4002.t0 a_35575_3749.t13 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2692 VDD.t4122 B[3].t25 a_63527_6198.t6 VDD.t4121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2693 a_53357_22238.t1 a_52767_22675.t10 VSS.t564 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2694 a_11110_7655.t1 a_10459_8962.t10 VSS.t316 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2695 VSS.t520 a_9221_6047.t6 a_9879_4622.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2696 a_65769_n1230.t2 a_65224_n537.t7 a_65769_n1962.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2697 a_10513_20719.t0 opcode[0].t166 VDD.t2049 VDD.t2048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2698 a_22608_8258.t2 a_23787_8115.t6 a_23141_8988.t4 VDD.t2123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2699 a_60047_3874.t2 a_58321_311.t5 a_59929_3874.t4 VDD.t3513 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2700 VSS.t400 a_30152_5242.t6 a_31377_5900.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2701 VDD.t3344 a_37902_9782.t10 a_38492_9345.t0 VDD.t3343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2702 VDD.t3107 a_30645_n306.t14 a_48131_15735.t1 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2703 a_66061_10678.t3 a_64117_8794.t7 VSS.t412 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2704 VDD.t4124 B[3].t26 a_9304_16408.t4 VDD.t4123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2705 VSS.t589 a_20579_1259.t7 a_20526_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2706 a_47719_15761.t5 a_48131_15735.t6 a_46176_16428.t5 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2707 a_1735_13585.t0 opcode[0].t167 VDD.t2051 VDD.t2050 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2708 VSS.t299 a_60193_3291.t7 a_61071_3878.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2709 a_70513_4160.t6 a_70459_5045.t6 a_70513_4278.t7 VDD.t1959 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2710 VSS.t569 a_42266_11512.t14 a_46592_6178.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2711 VDD.t3588 a_42266_11512.t15 a_44460_6616.t0 VDD.t3587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2712 a_70509_13768.t9 opcode[1].t99 VDD.t1201 VDD.t1200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2713 VDD.t3086 opcode[3].t46 a_3424_n2152.t0 VDD.t3085 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2714 VDD.t3739 a_61782_23618.t5 a_62778_24205.t4 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2715 a_52710_16433.t5 a_53713_16459.t5 a_54253_15766.t9 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2716 a_56438_21365.t4 a_56011_22058.t6 a_56556_21365.t1 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2717 a_53352_20634.t0 a_52762_21071.t10 VDD.t3103 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2718 a_10509_14454.t6 a_11155_13581.t6 a_9976_13724.t5 VDD.t3566 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2719 VDD.t561 a_61343_9163.t7 a_70509_n1998.t4 VDD.t560 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2720 a_1156_1740.t7 opcode[2].t44 a_1392_407.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2721 a_48124_20638.t0 a_48418_21344.t7 VSS.t207 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2722 a_839_n2152.t0 a_280_n2152.t5 a_1188_n2152.t0 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2723 a_20633_10847.t2 opcode[1].t100 VDD.t1203 VDD.t1202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2724 a_8202_7655.t0 opcode[0].t168 a_6842_8258.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2725 a_53299_1015.t3 a_48064_9163.t14 VSS.t134 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2726 a_46215_18571.t0 a_47282_17937.t7 VDD.t3634 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2727 a_46176_16428.t7 a_30645_n306.t15 a_48073_15029.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2728 a_70455_14535.t0 opcode[1].t101 VDD.t1205 VDD.t1204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2729 a_31377_5900.t1 a_30152_6681.t7 a_30645_5900.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2730 VDD.t2522 a_49568_24206.t8 a_49832_23623.t3 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2731 VDD.t4407 A[3].t42 a_19357_21596.t6 VDD.t4406 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2732 a_566_8262.t3 a_1745_8119.t7 a_1690_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2733 a_48130_1040.t2 a_47703_1733.t7 a_48248_1040.t3 VDD.t3407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2734 a_31377_4067.t0 B[4].t18 VSS.t295 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2735 a_67372_n1177.t0 a_48248_1040.t17 a_67135_n540.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2736 VSS.t600 A[7].t26 a_7562_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2737 a_3951_1740.t3 a_3642_11724.t7 VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2738 VDD.t352 a_19464_8258.t11 a_19406_8988.t0 VDD.t351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2739 a_23141_8988.t3 a_23787_8115.t7 a_22608_8258.t1 VDD.t2124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2740 VDD.t1014 a_59311_24329.t9 a_59901_23892.t1 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2741 VDD.t1279 a_3710_8262.t10 a_3652_8992.t1 VDD.t1278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2742 a_16865_8992.t3 opcode[0].t169 VDD.t1506 VDD.t1505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2743 a_67372_3171.t1 a_54908_6842.t17 a_67135_3808.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2744 a_48548_6884.t0 a_44405_8194.t14 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2745 a_55862_18700.t3 A[5].t38 VDD.t3458 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2746 a_13810_n2152.t5 a_14335_n2637.t7 a_13461_n2152.t8 VDD.t4249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2747 VSS.t375 a_1713_n2637.t6 a_1660_n3485.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2748 a_24806_15774.t0 B[0].t16 VSS.t356 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2749 a_53430_9674.t2 a_51704_6111.t6 a_53312_9674.t3 VDD.t3241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2750 a_13661_8966.t6 a_17495_6045.t5 a_18035_5352.t7 VDD.t2121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2751 a_61415_6910.t0 a_59635_6910.t13 VDD.t892 VDD.t891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2752 VDD.t3768 A[7].t27 a_6735_21596.t10 VDD.t3767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2753 a_31377_n70.t0 B[6].t30 VSS.t221 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2754 a_44460_6616.t4 a_44405_8194.t15 VDD.t249 VDD.t248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2755 VDD.t3460 A[5].t39 a_13011_21592.t11 VDD.t3459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2756 a_19677_n2174.t2 a_21956_20862.t9 VDD.t2144 VDD.t2143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2757 VDD.t334 a_30647_7968.t13 a_54540_21365.t1 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2758 a_39263_15765.t10 a_39618_16432.t12 VDD.t3517 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2759 VSS.t447 a_46916_3289.t6 a_47794_3876.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2760 a_5060_13125.t0 opcode[0].t170 a_3700_13728.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2761 VDD.t1508 opcode[0].t171 a_1089_14458.t1 VDD.t1507 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2762 a_55504_n1325.t2 a_54914_n1762.t8 VDD.t3002 VDD.t3001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2763 a_48815_11511.t2 a_48225_11948.t9 VDD.t4444 VDD.t4443 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2764 VDD.t1435 a_41913_24205.t8 a_42177_23622.t3 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2765 a_60766_15769.t1 a_30645_3831.t22 VDD.t2513 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2766 a_23777_10847.t1 opcode[1].t102 VDD.t1207 VDD.t1206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2767 a_53343_23888.t0 a_52753_24325.t10 VSS.t581 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2768 VDD.t3717 a_35594_7027.t14 a_37916_8132.t4 VDD.t3716 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2769 a_48248_1040.t5 a_48542_1014.t7 a_48130_1040.t9 VDD.t1542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2770 VDD.t4581 a_54908_6842.t18 a_67135_3808.t2 VDD.t4580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2771 VDD.t1600 a_30643_n2374.t19 a_42756_17049.t1 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2772 a_9976_13724.t4 a_11155_13581.t7 a_11100_13121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2773 VSS.t349 a_18824_20866.t11 a_16545_n2178.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2774 VDD.t1209 opcode[1].t103 a_70509_1146.t9 VDD.t1208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2775 a_12241_5326.t3 A[6].t41 VSS.t227 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2776 a_42964_22066.t1 a_41611_21373.t14 VDD.t524 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2777 a_16855_11724.t5 a_17501_10851.t5 a_16322_10994.t2 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2778 VDD.t3359 a_51109_747.t8 a_51699_310.t1 VDD.t3358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2779 VSS.t650 B[3].t27 a_17495_6045.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2780 a_9334_20862.t6 a_10513_20719.t4 a_10458_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2781 a_39675_15739.t3 a_39618_16432.t13 VSS.t558 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2782 a_66005_n1962.t1 a_64192_n2074.t11 a_65769_n1230.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2783 VDD.t1211 opcode[1].t104 a_14357_10851.t1 VDD.t1210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2784 VDD.t102 a_51054_2325.t16 a_54785_1041.t3 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2785 VDD.t1510 opcode[0].t172 a_20643_8115.t1 VDD.t1509 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2786 a_839_n2152.t3 a_779_n2178.t5 VDD.t2723 VDD.t2722 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2787 a_65651_6613.t0 a_64188_3841.t10 VDD.t469 VDD.t468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2788 a_43173_24209.t0 a_40310_22246.t4 a_43055_24209.t0 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2789 a_70509_n2116.t4 a_70455_n1231.t6 a_70509_n1998.t9 VDD.t4133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2790 a_48131_15735.t0 a_30645_n306.t16 VDD.t3108 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2791 VDD.t2734 a_51695_9365.t7 a_53430_9674.t3 VDD.t2733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2792 a_807_1740.t9 a_498_11724.t6 VDD.t589 VDD.t588 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2793 VSS.t58 a_30647_7968.t14 a_53004_22038.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2794 a_9304_16408.t3 B[3].t28 VDD.t4126 VDD.t4125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2795 VDD.t3769 A[7].t28 a_40621_16458.t0 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2796 a_9986_8258.t1 a_11165_8115.t6 a_10519_8988.t11 VDD.t2717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2797 a_18035_5352.t1 a_18447_5326.t7 a_13661_8966.t2 VDD.t1625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2798 a_70509_13650.t3 a_70455_14535.t6 a_71842_14359.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2799 a_7375_8988.t9 a_7315_8962.t10 a_6842_8258.t4 VDD.t3290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2800 a_30154_12886.t0 opcode[0].t173 VDD.t1512 VDD.t1511 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2801 a_62778_24205.t3 a_61782_23618.t6 VDD.t2363 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2802 VDD.t1457 A[6].t42 a_3855_6357.t0 VDD.t1456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2803 VDD.t2614 B[7].t15 a_29950_n2431.t3 VDD.t2613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2804 a_70509_1146.t7 a_70455_1913.t6 a_70509_1028.t4 VDD.t873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2805 VDD.t1514 opcode[0].t174 a_29952_5843.t2 VDD.t1513 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2806 a_56556_21365.t3 a_56011_22058.t7 a_56438_21365.t3 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2807 a_64192_n2074.t1 a_63602_n1637.t9 VSS.t22 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2808 VSS.t649 a_30150_n3032.t6 a_31375_n2374.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2809 a_16859_20723.t3 opcode[0].t175 VSS.t240 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2810 a_45279_16157.t2 a_52674_17946.t7 VDD.t396 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2811 a_35591_989.t0 a_35001_1426.t10 VDD.t1985 VDD.t1984 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2812 a_22821_n2174.t1 a_25100_20862.t9 VDD.t595 VDD.t594 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2813 a_1188_n2152.t1 a_280_n2152.t6 a_839_n2152.t1 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2814 VDD.t1516 opcode[0].t176 a_29952_3774.t6 VDD.t1515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2815 a_30645_5900.t3 a_30152_5242.t7 a_29952_5843.t10 VDD.t2516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2816 VSS.t78 B[2].t17 a_19563_6043.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2817 VSS.t503 a_41153_18571.t7 a_40724_17941.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2818 VDD.t1213 opcode[1].t105 a_20633_10847.t1 VDD.t1212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2819 VDD.t3137 a_61216_21369.t12 a_62569_22062.t2 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2820 a_57676_2326.t1 a_67135_3808.t9 VDD.t4071 VDD.t4070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2821 VSS.t554 a_64192_n2074.t12 a_67372_n1177.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2822 VDD.t844 opcode[2].t45 a_19705_1744.t0 VDD.t843 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2823 a_7957_1259.t0 a_70513_4160.t11 VDD.t1904 VDD.t1903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2824 a_6842_8258.t3 a_8021_8115.t6 a_7375_8988.t7 VDD.t3056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2825 VSS.t72 a_16322_10994.t9 a_16264_11724.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2826 a_51704_1914.t0 a_51114_2351.t10 VDD.t1047 VDD.t1046 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2827 VDD.t2062 a_6774_11720.t6 a_7083_1744.t0 VDD.t2061 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2828 a_30152_5242.t0 B[3].t29 VDD.t4128 VDD.t4127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2829 VDD.t1075 a_51059_8126.t13 a_55202_6816.t0 VDD.t1074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2830 VDD.t335 a_30647_7968.t15 a_52767_22675.t6 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2831 a_40093_1016.t3 a_35575_3749.t14 VSS.t30 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2832 a_1089_11724.t8 opcode[1].t106 VDD.t1215 VDD.t1214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2833 a_40101_6796.t0 a_35602_9612.t13 VDD.t949 VDD.t948 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2834 a_59901_23892.t0 a_59311_24329.t10 VDD.t1015 w_59157_24267# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2835 a_30643_1763.t4 a_30150_2544.t7 a_29950_1706.t9 VDD.t526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2836 VDD.t2277 a_48815_11511.t15 a_51114_6548.t4 VDD.t2276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2837 a_24652_5324.t1 A[0].t19 VDD.t2330 VDD.t2329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2838 VSS.t458 a_57684_8194.t14 a_61769_6178.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2839 a_24157_16385.t6 A[0].t20 a_24806_15774.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2840 VSS.t544 a_19563_6043.t7 a_20221_4618.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2841 a_4233_11724.t1 a_3642_14458.t6 a_3700_10994.t5 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2842 VDD.t1518 opcode[0].t177 a_23787_8115.t1 VDD.t1517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2843 a_45035_3563.t1 a_44445_4000.t8 VDD.t2854 VDD.t2853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2844 VDD.t1531 a_53010_6842.t13 a_54363_7535.t1 VDD.t1530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2845 a_13011_21592.t10 A[5].t40 VDD.t3462 VDD.t3461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2846 a_54540_21365.t2 a_30647_7968.t16 VDD.t336 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2847 a_59627_1042.t5 a_59082_1735.t6 a_59509_1042.t2 VDD.t2498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2848 a_59517_6910.t6 a_59929_6884.t7 a_59635_6910.t2 VDD.t229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2849 VDD.t2146 a_21956_20862.t10 a_19677_n2174.t1 VDD.t2145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2850 VDD.t3518 a_39618_16432.t14 a_39263_15765.t11 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2851 a_8289_6359.t0 A[0].t21 VDD.t2332 VDD.t2331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2852 VSS.t83 a_64188_3841.t11 a_67372_6666.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2853 a_22709_16385.t6 A[1].t33 a_23358_15774.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2854 a_5659_15753.t1 A[6].t43 a_5794_16410.t3 VDD.t1458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2855 VDD.t3004 a_54914_n1762.t9 a_55504_n1325.t1 VDD.t3003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2856 a_8011_13581.t3 opcode[0].t178 VSS.t241 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2857 a_4332_n2152.t6 a_3424_n2152.t6 a_3983_n2152.t10 VDD.t4558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2858 a_23700_6043.t0 B[0].t17 VDD.t2219 VDD.t2218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2859 a_61636_24201.t4 a_59910_20638.t6 a_61518_24201.t2 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2860 a_56102_24201.t4 a_53357_22238.t6 VSS.t184 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2861 VDD.t4446 a_48225_11948.t10 a_48815_11511.t3 VDD.t4445 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2862 a_63527_9231.t1 B[5].t33 VDD.t1852 VDD.t1851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2863 VDD.t3048 a_20054_1744.t10 a_20611_n2633.t0 VDD.t3047 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2864 VDD.t2514 a_30645_3831.t23 a_60766_15769.t0 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2865 VDD.t1217 opcode[1].t107 a_23777_10847.t0 VDD.t1216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2866 VDD.t1219 opcode[1].t108 a_70455_n1231.t0 VDD.t1218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2867 a_4300_1740.t1 a_3392_1740.t7 a_3951_1740.t2 VDD.t1284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2868 a_42756_17049.t0 a_30643_n2374.t20 VDD.t1601 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2869 VDD.t3674 a_13849_16387.t8 a_1029_14432.t1 VDD.t3673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2870 a_11336_13121.t0 opcode[0].t179 a_9976_13724.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2871 VDD.t4067 a_8289_6359.t5 a_23141_8988.t7 VDD.t4066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2872 a_20103_5350.t5 A[2].t31 VDD.t3986 VDD.t3985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2873 VSS.t296 B[4].t19 a_15426_6045.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2874 VSS.t495 opcode[3].t47 a_19178_n2148.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2875 a_10694_20259.t0 opcode[0].t180 a_9334_20862.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2876 VDD.t2104 a_5108_13805.t5 a_4233_14458.t10 VDD.t2103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2877 a_59937_9742.t2 a_58329_6179.t6 VSS.t29 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2878 a_59929_3874.t0 a_58321_311.t6 VSS.t233 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2879 a_12672_15792.t1 A[0].t22 a_12808_16408.t5 VDD.t2333 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2880 a_45939_15761.t2 a_45281_16454.t6 a_45821_15761.t2 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2881 a_9918_11720.t0 a_9976_10990.t11 VDD.t2766 VDD.t2765 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2882 a_14357_10851.t0 opcode[1].t109 VDD.t1221 VDD.t1220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2883 VDD.t2725 a_779_n2178.t6 a_839_n2152.t4 VDD.t2724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2884 a_43055_24209.t1 a_40310_22246.t5 a_43173_24209.t1 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2885 VDD.t3770 A[7].t29 a_42761_15445.t5 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2886 VSS.t427 a_6832_10990.t9 a_6774_11720.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2887 a_23787_8115.t0 opcode[0].t181 VDD.t1520 VDD.t1519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2888 a_15966_5352.t11 a_16378_5326.t6 a_10459_8962.t6 VDD.t2861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2889 a_71842_n1171.t1 opcode[1].t110 a_70509_n2116.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2890 a_54903_1041.t3 a_54358_1734.t7 a_54785_1041.t6 VDD.t1341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2891 a_20824_7655.t1 opcode[0].t182 a_19464_8258.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2892 VSS.t532 a_70513_16782.t10 a_20579_1259.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2893 VDD.t626 a_54903_1041.t20 a_57722_4002.t4 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2894 VDD.t2561 a_64117_8794.t8 a_65649_10704.t2 VDD.t2560 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2895 a_17511_8119.t0 opcode[0].t183 VDD.t1522 VDD.t1521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2896 a_8056_15820.t1 a_7995_15753.t6 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2897 a_56438_21365.t8 a_56850_21339.t5 a_56556_21365.t7 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2898 VDD.t1223 opcode[1].t111 a_70513_20044.t6 VDD.t1222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2899 VSS.t367 a_16322_13728.t11 a_16264_14458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2900 VDD.t397 a_52674_17946.t8 a_45279_16157.t3 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2901 VDD.t597 a_25100_20862.t10 a_22821_n2174.t0 VDD.t596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2902 a_39582_17945.t4 a_39657_18575.t7 VSS.t519 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2903 VDD.t2409 B[5].t34 a_63527_9231.t0 VDD.t2408 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2904 a_839_n2152.t2 a_280_n2152.t7 a_1188_n2152.t2 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2905 a_39681_1042.t4 a_40093_1016.t6 a_39799_1042.t7 VDD.t4517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2906 VDD.t3667 a_39799_1042.t15 a_41152_1735.t0 VDD.t3666 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2907 a_62569_22062.t1 a_61216_21369.t13 VDD.t3138 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2908 a_52767_15740.t3 a_52710_16433.t13 VSS.t214 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2909 a_67135_7303.t4 a_64117_5761.t12 VDD.t1149 VDD.t1148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2910 VDD.t846 opcode[2].t46 a_9668_1744.t0 VDD.t845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2911 a_41611_20641.t1 a_41905_21347.t7 VSS.t342 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2912 a_23670_411.t1 a_22290_1744.t6 a_23198_1744.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2913 a_62778_24205.t2 a_59915_22242.t4 a_62660_24205.t1 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2914 VDD.t4527 a_54713_3294.t14 a_57744_8220.t0 VDD.t4526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2915 VDD.t3488 a_64192_n2074.t13 a_65224_n537.t0 VDD.t3487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2916 VSS.t496 opcode[3].t48 a_22322_n2148.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2917 a_13898_5354.t0 B[5].t35 VDD.t2411 VDD.t2410 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2918 a_70513_16782.t0 a_50022_21370.t10 a_70513_16900.t2 VDD.t1271 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2919 a_556_10994.t7 a_1735_10851.t5 a_1089_11724.t11 VDD.t4442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2920 VDD.t572 a_59627_1042.t12 a_61407_1042.t9 VDD.t571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2921 a_3951_1740.t11 a_4825_1255.t7 a_4300_1740.t7 VDD.t3404 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2922 VDD.t749 a_54658_21365.t14 a_56011_22058.t1 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2923 VDD.t1493 a_30647_12105.t14 a_39706_24333.t5 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2924 a_25633_21592.t2 opcode[0].t184 VDD.t1524 VDD.t1523 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2925 VSS.t448 a_43319_23626.t13 a_50258_20638.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2926 a_3700_10994.t4 a_3642_14458.t7 a_4233_11724.t0 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2927 a_58312_3565.t1 a_57722_4002.t9 VDD.t1428 VDD.t1427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2928 VSS.t466 a_70513_7304.t11 a_11101_1259.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2929 VDD.t251 a_44405_8194.t16 a_48136_6910.t9 VDD.t250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2930 a_10259_n2148.t10 opcode[3].t49 VDD.t3088 VDD.t3087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2931 a_30643_1763.t0 opcode[0].t185 a_31375_1999.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2932 VDD.t3464 A[5].t41 a_13011_21592.t9 VDD.t3463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2933 a_1680_10391.t1 a_498_14458.t7 VSS.t88 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2934 VDD.t2221 B[0].t18 a_30154_11447.t1 VDD.t2220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2935 a_23968_7655.t0 opcode[0].t186 a_22608_8258.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2936 a_35004_7464.t4 A[5].t42 VDD.t3466 VDD.t3465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2937 a_63015_14838.t1 a_58326_16165.t15 VSS.t161 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2938 VDD.t3149 a_46652_3872.t8 a_46916_3289.t0 VDD.t3148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2939 a_3983_n2152.t11 a_3424_n2152.t7 a_4332_n2152.t7 VDD.t4559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2940 a_45035_3563.t3 a_44445_4000.t9 VSS.t463 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2941 a_61518_24201.t3 a_59910_20638.t7 a_61636_24201.t3 w_61482_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2942 a_63832_571.t1 A[4].t45 a_63595_1208.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2943 VDD.t1459 A[6].t44 a_47179_16454.t2 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2944 VDD.t49 a_3855_6357.t7 a_4243_8992.t2 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2945 VDD.t3304 B[6].t31 a_30152_n964.t0 VDD.t3303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2946 VDD.t1656 a_38721_16161.t16 a_42756_17049.t4 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2947 a_1029_14432.t0 a_13849_16387.t9 VDD.t3676 VDD.t3675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2948 VSS.t534 a_8056_15820.t5 a_11336_13121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2949 a_7083_1744.t10 a_6524_1744.t6 a_7432_1744.t6 VDD.t3604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2950 VDD.t4163 a_44399_2324.t13 a_44459_2350.t0 VDD.t4162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2951 a_46823_22243.t0 a_46233_22680.t9 VDD.t878 w_46079_22618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2952 VSS.t228 A[6].t45 a_10694_20259.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2953 a_4233_14458.t9 a_5108_13805.t6 VDD.t2106 VDD.t2105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2954 a_45055_7783.t2 a_44465_8220.t9 VDD.t2835 VDD.t2834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2955 a_58334_7783.t0 a_57744_8220.t9 VDD.t3157 VDD.t3156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2956 a_29954_12048.t3 B[0].t19 VDD.t2223 VDD.t2222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2957 a_45821_15761.t10 a_46233_15735.t6 a_45939_15761.t5 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2958 VDD.t3164 a_53307_3873.t8 a_53571_3290.t0 VDD.t3163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2959 VDD.t1610 a_61525_1042.t10 a_70513_4278.t5 VDD.t1609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2960 VDD.t471 a_64188_3841.t12 a_65224_7306.t0 VDD.t470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2961 a_1964_13805.t3 a_4491_15753.t8 VDD.t4299 VDD.t4298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2962 VDD.t3306 B[6].t32 a_11829_5352.t1 VDD.t3305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2963 a_53299_1015.t0 a_48064_9163.t15 VDD.t783 VDD.t782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2964 VDD.t1602 a_30643_n2374.t21 a_41161_15765.t4 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2965 a_42761_15445.t4 A[7].t30 VDD.t3771 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2966 a_11133_n2633.t2 a_10576_1744.t10 VDD.t2555 VDD.t2554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2967 a_59929_6884.t1 a_55469_11532.t14 VDD.t2543 VDD.t2542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2968 VDD.t848 opcode[2].t47 a_10227_1744.t6 VDD.t847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2969 VSS.t438 a_8289_6359.t6 a_23968_7655.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2970 a_65649_10704.t1 a_64117_8794.t9 VDD.t2563 VDD.t2562 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2971 a_71846_4869.t0 a_52473_15766.t11 VSS.t118 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2972 a_16213_21596.t3 A[2].t32 a_15680_20866.t1 VDD.t3987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2973 a_18892_15774.t0 B[4].t20 VSS.t297 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2974 VDD.t2798 a_35004_7464.t10 a_35594_7027.t3 VDD.t2797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2975 a_7315_8962.t3 a_14310_5328.t7 a_13898_5354.t7 VDD.t3060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2976 VSS.t641 a_40011_18575.t7 a_39582_17945.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2977 VDD.t190 A[1].t34 a_7551_6363.t0 VDD.t189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2978 a_71846_17491.t0 a_50022_21370.t11 VSS.t203 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2979 a_55848_17050.t6 a_30643_1763.t19 VDD.t3133 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2980 VDD.t3139 a_61216_21369.t14 a_62569_22062.t0 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2981 VDD.t2192 a_51100_4001.t10 a_51690_3564.t0 VDD.t2191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2982 VSS.t446 a_22608_8258.t10 a_22550_8988.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2983 a_1680_13125.t0 a_1029_14432.t7 VSS.t394 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2984 a_46232_1040.t9 a_41697_1042.t20 VDD.t1686 VDD.t1685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2985 a_20611_n2633.t3 a_20054_1744.t11 VSS.t491 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2986 a_44459_2350.t4 a_42301_n1318.t15 VDD.t4101 VDD.t4100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2987 a_62660_24205.t2 a_59915_22242.t5 a_62778_24205.t1 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2988 a_11829_5352.t0 B[6].t33 VDD.t3308 VDD.t3307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2989 a_51695_9365.t1 a_51105_9802.t8 VDD.t1345 VDD.t1344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2990 a_54790_6842.t9 a_53010_6842.t14 VDD.t1533 VDD.t1532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2991 a_1089_11724.t6 a_1735_10851.t6 a_556_10994.t4 VDD.t2897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2992 VDD.t3534 a_10576_1744.t11 a_11133_n2633.t3 VDD.t3533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2993 VSS.t372 a_70509_10506.t11 a_14303_1255.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2994 VDD.t951 a_35602_9612.t14 a_39689_6822.t0 VDD.t950 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2995 a_48006_21370.t8 a_30645_10037.t21 VDD.t2291 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2996 a_56011_22058.t0 a_54658_21365.t15 VDD.t750 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2997 a_65651_6613.t9 a_65224_7306.t7 a_65769_6613.t5 VDD.t1333 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2998 a_70513_7422.t3 a_58986_15769.t10 a_70513_7304.t3 VDD.t1115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2999 VDD.t986 a_58326_16165.t16 a_62361_17053.t4 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3000 VDD.t3326 a_70513_16782.t11 a_20579_1259.t0 VDD.t3325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3001 VDD.t1526 opcode[0].t187 a_25633_21592.t1 VDD.t1525 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3002 a_50022_20638.t0 a_50316_21344.t7 VSS.t109 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3003 VDD.t2700 a_65769_3118.t10 a_70513_7422.t5 VDD.t2699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3004 a_67135_n540.t4 a_64192_n2074.t14 VDD.t3490 VDD.t3489 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3005 VDD.t3090 opcode[3].t50 a_10259_n2148.t9 VDD.t3089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3006 VDD.t1527 opcode[0].t188 a_43391_21373.t7 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3007 a_54952_21339.t0 A[2].t33 VDD.t3988 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3008 a_29952_3774.t0 B[4].t21 VDD.t1872 VDD.t1871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3009 VDD.t1874 B[4].t22 a_34985_4186.t1 VDD.t1873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3010 VSS.t272 a_41697_1042.t21 a_46586_308.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3011 a_16573_1740.t1 a_16264_11724.t6 VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3012 a_70513_7422.t8 a_70459_8189.t7 a_70513_7304.t7 VDD.t3244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3013 a_52767_22675.t2 a_49832_23623.t9 VDD.t995 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3014 VDD.t1245 a_48855_n1313.t16 a_52460_1734.t0 VDD.t1244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3015 a_19937_8962.t1 A[1].t35 a_22526_4620.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3016 VSS.t502 a_39807_6822.t13 a_41160_7515.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3017 a_23081_8962.t6 a_23700_6043.t6 a_24240_5350.t10 VDD.t1479 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3018 a_71846_8013.t0 a_58986_15769.t11 VSS.t186 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3019 a_11346_7655.t0 opcode[0].t189 a_9986_8258.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3020 VDD.t3092 opcode[3].t51 a_3983_n2152.t7 VDD.t3091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3021 VDD.t1529 opcode[0].t190 a_30152_475.t0 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3022 a_48124_21370.t4 a_47579_22063.t6 a_48006_21370.t6 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3023 a_60047_3874.t3 a_58312_3565.t7 VDD.t3478 VDD.t3477 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3024 a_47179_16454.t1 A[6].t46 VDD.t1460 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3025 VDD.t3492 a_64192_n2074.t15 a_65651_n1230.t9 VDD.t3491 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3026 VDD.t3169 a_22540_11720.t5 a_22849_1744.t7 VDD.t3168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3027 a_19987_14454.t9 a_19927_14428.t7 a_19454_13724.t5 VDD.t386 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3028 a_42756_17049.t3 a_38721_16161.t17 VDD.t1658 w_42662_17013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3029 a_46652_3872.t3 a_45044_309.t7 a_46770_3872.t2 VDD.t2496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3030 a_11640_16408.t0 B[1].t17 VDD.t2469 VDD.t2468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3031 VDD.t1290 a_51119_8152.t10 a_51709_7715.t0 VDD.t1289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3032 VDD.t1557 a_55469_11532.t15 a_57739_6616.t0 VDD.t1556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3033 a_30150_n1593.t1 opcode[0].t191 VDD.t3191 VDD.t3190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3034 a_29950_1706.t7 a_30150_1105.t6 a_30643_1763.t2 VDD.t3669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3035 a_46233_15735.t0 a_46176_16428.t15 VDD.t4509 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3036 a_26279_20719.t3 opcode[0].t192 VSS.t513 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3037 a_40227_9654.t4 a_38501_6091.t6 a_40109_9654.t3 VDD.t1104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3038 a_45939_15761.t4 a_46233_15735.t7 a_45821_15761.t9 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3039 a_16332_8262.t2 a_16805_8966.t10 a_16865_8992.t1 VDD.t1335 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3040 a_41161_15765.t3 a_30643_n2374.t22 VDD.t1803 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3041 a_14312_7659.t0 a_13661_8966.t11 VSS.t665 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3042 a_23081_8962.t4 A[0].t23 a_24594_4618.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3043 VDD.t850 opcode[2].t48 a_22290_1744.t0 VDD.t849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3044 a_45055_7783.t3 a_44465_8220.t10 VSS.t461 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3045 VDD.t2565 a_64117_8794.t10 a_65649_10704.t0 VDD.t2564 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3046 a_41579_1042.t6 a_37848_2326.t15 VDD.t1952 VDD.t1951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3047 a_16320_4620.t0 B[4].t23 VSS.t298 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3048 a_18243_16385.t6 A[4].t46 a_18892_15774.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3049 a_61819_1016.t0 a_57676_2326.t13 VDD.t1707 VDD.t1706 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3050 VDD.t2984 a_51813_16162.t15 a_55848_17050.t2 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3051 a_22849_1744.t8 a_22540_11720.t6 VDD.t3171 VDD.t3170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3052 a_22598_13724.t3 a_23071_14428.t6 a_23131_14454.t4 VDD.t1137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3053 VDD.t1281 a_3710_8262.t11 a_3652_8992.t0 VDD.t1280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3054 a_16795_16385.t3 A[5].t43 a_17444_15774.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3055 a_7365_14454.t3 opcode[0].t193 VDD.t3193 VDD.t3192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3056 VSS.t37 a_45281_16454.t7 a_45939_15029.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3057 a_4237_20723.t3 opcode[0].t194 VSS.t514 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3058 a_65769_3118.t3 a_65224_3811.t6 a_65651_3118.t9 VDD.t4051 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3059 a_62778_24205.t0 a_59915_22242.t6 a_62660_24205.t3 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3060 VDD.t3134 a_30643_1763.t20 a_54253_15766.t7 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3061 a_55853_15446.t4 A[5].t44 VDD.t3467 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3062 a_49968_14830.t1 a_45279_16157.t15 VSS.t528 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3063 a_16865_8992.t0 a_16805_8966.t11 a_16332_8262.t0 VDD.t1336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3064 VDD.t2630 a_41251_9658.t8 a_37848_2326.t3 VDD.t2629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3065 VDD.t4130 B[3].t30 a_18035_5352.t11 VDD.t4129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3066 VDD.t2781 a_43319_23626.t14 a_49904_21370.t6 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3067 a_39689_6822.t6 a_35594_7027.t15 VDD.t3719 VDD.t3718 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3068 VSS.t180 a_3700_10994.t10 a_3642_11724.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3069 a_25633_21592.t0 opcode[0].t195 VDD.t3195 VDD.t3194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3070 a_39799_1042.t4 a_39254_1735.t6 a_39799_310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3071 VSS.t69 a_53103_18576.t7 a_52674_17946.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3072 a_20412_15776.t1 B[3].t31 VSS.t301 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3073 VSS.t277 a_57676_2326.t14 a_57968_111.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3074 a_10519_8988.t5 a_10459_8962.t11 a_9986_8258.t7 VDD.t1978 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3075 a_6784_8988.t0 a_6842_8258.t11 VDD.t2805 VDD.t2804 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3076 VSS.t424 a_46356_6910.t12 a_47709_7603.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3077 VDD.t996 a_49832_23623.t10 a_52767_22675.t1 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3078 VDD.t3197 opcode[0].t196 a_4243_8992.t7 VDD.t3196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3079 a_54952_21339.t3 A[2].t34 VSS.t630 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3080 VSS.t392 B[1].t18 a_30152_9379.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3081 a_3983_n2152.t8 opcode[3].t52 VDD.t3094 VDD.t3093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3082 a_65651_3118.t4 a_66063_3092.t6 a_65769_3118.t1 VDD.t515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3083 a_48006_21370.t7 a_47579_22063.t7 a_48124_21370.t5 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3084 a_59509_1042.t5 a_59921_1016.t6 a_59627_1042.t2 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3085 VDD.t962 a_42770_18699.t10 a_40799_18571.t0 w_42676_18663# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3086 VDD.t1461 A[6].t47 a_47179_16454.t0 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3087 a_65651_6613.t6 a_64117_5761.t13 VDD.t1151 VDD.t1150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3088 a_12241_5326.t1 A[6].t48 VDD.t1463 VDD.t1462 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3089 VDD.t574 a_59627_1042.t13 a_60980_1735.t0 VDD.t573 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3090 VSS.t149 a_48254_6910.t18 a_52465_7535.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3091 a_52762_21071.t4 A[2].t35 VDD.t3989 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3092 a_70513_16900.t5 a_65769_6613.t11 VDD.t2789 VDD.t2788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3093 a_1735_10851.t3 opcode[1].t112 VSS.t196 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3094 VDD.t1566 a_566_8262.t10 a_508_8992.t1 VDD.t1565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3095 a_46350_1040.t1 a_45805_1733.t6 a_46232_1040.t1 VDD.t1980 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3096 VDD.t180 a_35575_3749.t15 a_39681_1042.t9 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3097 VDD.t323 a_9918_11720.t7 a_10227_1744.t2 VDD.t322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3098 a_807_1740.t2 a_248_1740.t7 a_1156_1740.t3 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3099 VDD.t2148 a_21956_20862.t11 a_19677_n2174.t0 VDD.t2147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3100 VDD.t748 a_10608_n2148.t9 Y[4].t1 VDD.t747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3101 a_22172_5352.t1 B[1].t19 VDD.t2471 VDD.t2470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3102 VDD.t852 opcode[2].t49 a_248_1740.t0 VDD.t851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3103 a_45049_1913.t0 a_44459_2350.t9 VSS.t506 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3104 VDD.t1486 a_51054_2325.t17 a_51114_2351.t0 VDD.t1485 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3105 VDD.t1804 a_30643_n2374.t23 a_41161_15765.t2 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3106 VSS.t322 A[4].t47 a_60226_16462.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3107 a_9976_10990.t6 a_11155_10847.t7 a_10509_11720.t11 VDD.t4076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3108 a_12732_15818.t1 a_12672_15792.t7 VDD.t3239 VDD.t3238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3109 Y[5].t3 a_7464_n2148.t10 VSS.t167 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3110 VDD.t1087 a_3700_10994.t11 a_3642_11724.t1 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3111 a_59616_18579.t1 a_62361_17053.t9 VDD.t2759 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3112 a_40373_9071.t0 a_40109_9654.t8 VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3113 VDD.t337 a_30647_7968.t17 a_52753_24325.t6 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3114 VSS.t275 a_6813_6359.t7 a_17692_7659.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3115 a_41579_1042.t3 a_41152_1735.t7 a_41697_1042.t4 VDD.t1581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3116 VDD.t2502 a_508_8992.t6 a_1089_11724.t4 VDD.t2501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3117 a_6071_6357.t0 A[3].t43 VDD.t4405 VDD.t4404 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3118 VDD.t2816 a_57684_8194.t15 a_61415_6910.t7 VDD.t2815 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3119 VDD.t167 a_41507_3295.t15 a_45811_7603.t0 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3120 a_55848_17050.t1 a_51813_16162.t16 VDD.t2985 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3121 a_49963_16434.t1 a_30645_n306.t17 VSS.t500 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3122 VSS.t8 a_38492_9345.t6 a_40109_9654.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3123 a_9986_8258.t0 a_11165_8115.t7 a_10519_8988.t6 VDD.t2052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3124 VSS.t578 a_13358_6047.t6 a_14016_4622.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3125 a_6832_13724.t5 a_8011_13581.t5 a_7365_14454.t7 VDD.t1329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3126 VSS.t64 a_3700_13728.t11 a_3642_14458.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3127 a_57730_9870.t0 a_55469_11532.t16 VDD.t3411 VDD.t3410 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3128 VSS.t653 a_44399_2324.t14 a_44691_109.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3129 a_44451_9870.t1 a_42266_11512.t16 VDD.t3590 VDD.t3589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3130 a_53004_22038.t0 a_49832_23623.t11 a_52767_22675.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3131 VDD.t4016 a_63598_4278.t10 a_64188_3841.t0 VDD.t4015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3132 VSS.t201 a_9334_20862.t11 a_7055_n2174.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3133 a_46232_1040.t7 a_46644_1014.t7 a_46350_1040.t6 VDD.t1690 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3134 a_54253_15766.t8 a_30643_1763.t21 VDD.t3135 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3135 VDD.t3468 A[5].t45 a_55853_15446.t3 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3136 a_14335_n2637.t0 a_13778_1740.t11 VDD.t1856 VDD.t1855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3137 a_6524_1744.t0 opcode[2].t50 VDD.t854 VDD.t853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3138 VDD.t1535 a_53010_6842.t15 a_54363_7535.t0 VDD.t1534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3139 a_4626_16408.t0 B[7].t16 VDD.t2616 VDD.t2615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3140 a_40859_18597.t0 a_40799_18571.t7 VDD.t4197 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3141 VDD.t192 A[1].t36 a_22172_5352.t4 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3142 VDD.t654 a_62375_18703.t10 a_60404_18575.t0 w_62281_18667# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3143 VSS.t504 a_61216_21369.t15 a_62569_22062.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3144 VDD.t3310 B[6].t34 a_11289_6045.t0 VDD.t3309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3145 a_39681_1042.t0 a_35591_989.t17 VDD.t3561 VDD.t3560 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3146 a_48136_6910.t3 a_48548_6884.t7 a_48254_6910.t4 VDD.t4083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3147 a_22881_n2148.t3 a_22821_n2174.t6 VDD.t2910 VDD.t2909 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3148 a_52887_1041.t1 a_48064_9163.t16 VDD.t785 VDD.t784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3149 a_19763_16387.t3 A[3].t44 a_20412_15776.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3150 a_1735_13585.t1 opcode[0].t197 VSS.t515 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3151 a_23135_20719.t1 opcode[0].t198 VDD.t3199 VDD.t3198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3152 a_42031_24205.t1 a_40305_20642.t5 a_41913_24205.t2 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3153 a_24652_5324.t0 A[0].t24 VDD.t2335 VDD.t2334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3154 a_52767_22675.t0 a_49832_23623.t12 VDD.t997 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3155 a_29952_9980.t10 a_30152_10818.t6 a_30645_10037.t6 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3156 a_23198_1744.t4 a_22290_1744.t7 a_22849_1744.t9 VDD.t2193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3157 a_46818_20639.t3 a_46228_21076.t10 VSS.t512 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3158 a_16805_8966.t4 A[2].t36 a_20457_4618.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3159 a_70509_n1998.t6 opcode[1].t113 VDD.t1225 VDD.t1224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3160 VDD.t3096 opcode[3].t53 a_3983_n2152.t9 VDD.t3095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3161 a_46238_6910.t0 a_45811_7603.t7 a_46356_6910.t1 VDD.t1862 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3162 VDD.t4545 a_67133_11394.t10 a_44399_2324.t0 VDD.t4544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3163 a_56220_24201.t3 a_53357_22238.t7 a_56102_24201.t1 w_56066_24139# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3164 VDD.t169 a_41507_3295.t16 a_44451_9870.t4 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3165 a_12183_4620.t0 B[6].t35 VSS.t529 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3166 a_59627_1042.t3 a_59082_1735.t7 a_59509_1042.t1 VDD.t2073 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3167 VDD.t3990 A[2].t37 a_52762_21071.t3 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3168 a_46465_20439.t0 A[1].t37 a_46228_21076.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3169 a_63595_1208.t0 B[6].t36 VDD.t3312 VDD.t3311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3170 a_70509_1028.t3 a_70455_1913.t7 a_70509_1146.t6 VDD.t1622 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3171 a_41705_6822.t6 a_41160_7515.t6 a_41705_6090.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3172 a_66063_n1256.t1 a_48248_1040.t18 VDD.t2874 VDD.t2873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3173 VSS.t199 a_48855_n1313.t17 a_51337_3364.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3174 a_17511_8119.t1 opcode[0].t199 VDD.t3201 VDD.t3200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3175 a_23434_411.t0 a_22540_11720.t7 VSS.t511 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3176 VDD.t2413 B[5].t36 a_29950_1706.t0 VDD.t2412 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3177 a_54790_6842.t4 a_54363_7535.t6 a_54908_6842.t2 VDD.t459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3178 a_46456_23693.t0 A[1].t38 a_46219_24330.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3179 a_61216_21369.t3 a_60671_22062.t7 a_61216_20637.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3180 VDD.t1227 opcode[1].t114 a_70509_10624.t9 VDD.t1226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3181 VDD.t1637 a_37908_2352.t10 a_38498_1915.t0 VDD.t1636 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3182 VDD.t3640 a_54449_3877.t6 a_54713_3294.t1 VDD.t3639 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3183 a_53307_3873.t1 a_51699_310.t7 a_53425_3873.t3 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3184 VDD.t2539 a_61079_9746.t6 a_61343_9163.t1 VDD.t2538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3185 a_17479_n2637.t1 a_16922_1740.t10 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3186 VDD.t856 opcode[2].t51 a_3951_1740.t0 VDD.t855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3187 VDD.t2732 a_8289_6359.t7 a_23141_8988.t6 VDD.t2731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3188 VDD.t2896 a_12672_15792.t8 a_12732_15818.t0 VDD.t2895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3189 a_41705_6822.t0 a_41999_6796.t7 a_41587_6822.t3 VDD.t4146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3190 a_19737_n2148.t8 a_19677_n2174.t7 VDD.t2829 VDD.t2828 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3191 a_48548_6884.t3 a_44405_8194.t17 VSS.t41 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3192 VDD.t2760 a_62361_17053.t10 a_59616_18579.t0 w_62267_17017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3193 a_44465_8220.t4 a_44405_8194.t18 VDD.t253 VDD.t252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3194 Y[6].t0 a_4332_n2152.t10 VDD.t1302 VDD.t1301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3195 a_52753_24325.t5 a_30647_7968.t18 VDD.t338 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3196 a_52465_7535.t0 a_48254_6910.t19 VDD.t913 VDD.t912 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3197 VDD.t2505 a_55862_18700.t8 a_53891_18572.t2 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3198 a_52990_23688.t0 A[2].t38 a_52753_24325.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3199 a_1089_11724.t3 a_508_8992.t7 VDD.t2504 VDD.t2503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3200 a_67133_11394.t5 a_64117_8794.t11 VDD.t4496 VDD.t4495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3201 a_65651_n1230.t2 a_66063_n1256.t7 a_65769_n1230.t3 VDD.t1611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3202 a_26279_20719.t2 opcode[0].t200 VDD.t3203 VDD.t3202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3203 VDD.t2986 a_51813_16162.t17 a_55848_17050.t0 w_55754_17014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3204 VDD.t1709 a_57676_2326.t15 a_61407_1042.t2 VDD.t1708 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3205 a_54785_1041.t4 a_55197_1015.t6 a_54903_1041.t1 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3206 a_7365_14454.t6 a_8011_13581.t6 a_6832_13724.t6 VDD.t1330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3207 a_22849_1744.t3 a_23723_1259.t7 a_23198_1744.t1 VDD.t4421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3208 VSS.t539 a_21211_16387.t8 a_16795_14432.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3209 VDD.t1795 a_63595_1208.t10 a_64185_771.t0 VDD.t1794 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3210 VDD.t3205 opcode[0].t201 a_16859_20723.t1 VDD.t3204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3211 a_59557_20438.t0 A[3].t45 a_59320_21075.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3212 a_54908_6842.t3 a_54363_7535.t7 a_54790_6842.t5 VDD.t460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3213 VDD.t76 a_30643_1763.t22 a_54253_15766.t0 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3214 VDD.t2179 a_37856_8106.t16 a_37911_6528.t4 VDD.t2178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3215 a_47800_9746.t3 a_45055_7783.t6 a_47918_9746.t1 VDD.t4537 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3216 a_54713_3294.t2 a_54449_3877.t7 VDD.t3642 VDD.t3641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3217 a_4491_15753.t3 A[7].t31 a_4626_16408.t5 VDD.t3772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3218 VDD.t1615 a_4593_6357.t7 a_7375_8988.t4 VDD.t1614 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3219 VSS.t246 a_19763_16387.t8 a_13651_14432.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3220 VDD.t1085 a_46658_9742.t8 a_46922_9159.t0 VDD.t1084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3221 VDD.t3992 A[2].t39 a_6813_6359.t0 VDD.t3991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3222 a_30152_475.t3 opcode[0].t202 VSS.t516 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3223 a_67135_7303.t3 a_64117_5761.t14 VDD.t1153 VDD.t1152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3224 a_17495_6045.t0 B[3].t32 VDD.t1906 VDD.t1905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3225 VSS.t422 a_45035_3563.t7 a_46652_3872.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3226 VDD.t4529 a_54713_3294.t15 a_59517_6910.t0 VDD.t4528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3227 VDD.t676 a_15680_20866.t11 a_13401_n2178.t0 VDD.t675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3228 VSS.t371 A[0].t25 a_41847_20641.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3229 a_7432_1744.t0 opcode[2].t52 a_7668_411.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3230 VDD.t3592 a_42266_11512.t17 a_46238_6910.t3 VDD.t3591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3231 VDD.t3207 opcode[0].t203 a_23135_20719.t0 VDD.t3206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3232 a_10844_n3481.t0 a_10199_n2174.t6 VSS.t263 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3233 a_30150_2544.t1 opcode[0].t204 VDD.t3209 VDD.t3208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3234 a_10519_8988.t7 a_5331_6357.t7 VDD.t1100 VDD.t1099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3235 a_70509_n2116.t7 a_70455_n1231.t7 a_71842_n1407.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3236 a_53010_6842.t7 a_52465_7535.t7 a_52892_6842.t9 VDD.t4423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3237 VDD.t4433 a_46350_1040.t14 a_48130_1040.t8 VDD.t4432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3238 VDD.t3109 a_30645_n306.t18 a_47719_15761.t10 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3239 VDD.t3211 opcode[0].t205 a_30154_8749.t0 VDD.t3210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3240 VSS.t177 a_51059_8126.t14 a_51351_5911.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3241 a_39689_6822.t10 a_40101_6796.t6 a_39807_6822.t6 VDD.t4282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3242 VDD.t194 A[1].t39 a_22584_5326.t0 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3243 VSS.t449 a_43319_23626.t15 a_46465_20439.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3244 VSS.t340 a_17495_6045.t6 a_18153_4620.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3245 a_47918_9746.t0 a_45055_7783.t7 a_47800_9746.t4 VDD.t4538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3246 a_61098_21369.t3 a_30645_5900.t22 VDD.t765 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3247 VSS.t212 B[2].t18 a_30154_7310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3248 a_39262_7515.t0 a_35594_7027.t16 VDD.t3721 VDD.t3720 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3249 a_51100_4001.t0 a_48064_9163.t17 VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3250 a_44688_9233.t0 a_42266_11512.t18 a_44451_9870.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3251 VSS.t278 a_57676_2326.t16 a_61761_310.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3252 a_45044_309.t0 a_44454_746.t10 VDD.t3332 VDD.t3331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3253 a_6832_13724.t7 a_8011_13581.t7 a_7956_13121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3254 a_71842_11215.t1 a_63114_21369.t10 VSS.t429 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3255 a_41369_9658.t3 a_38506_7695.t7 a_41251_9658.t1 VDD.t1572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3256 a_16213_21596.t2 opcode[0].t206 VDD.t3213 VDD.t3212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3257 a_61452_20637.t0 a_30645_5900.t23 a_61216_21369.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3258 a_11155_10847.t0 opcode[1].t115 VDD.t4358 VDD.t4357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3259 a_10576_1744.t6 a_11101_1259.t6 a_10227_1744.t10 VDD.t789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3260 a_4183_8966.t2 a_11289_6045.t7 a_11829_5352.t6 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3261 a_53005_1041.t3 a_52460_1734.t6 a_52887_1041.t5 VDD.t2138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3262 a_6832_10990.t3 a_8011_10847.t7 a_7365_11720.t6 VDD.t2449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3263 VSS.t710 a_58328_16462.t7 a_58986_15037.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3264 VDD.t3470 A[5].t46 a_13898_5354.t4 VDD.t3469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3265 VSS.t178 a_51059_8126.t15 a_55144_6110.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3266 a_46776_9742.t3 a_45050_6179.t6 a_46658_9742.t2 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3267 VDD.t2473 B[1].t20 a_21632_6045.t1 VDD.t2472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3268 a_4491_15753.t0 B[7].t17 VSS.t418 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3269 VDD.t339 a_30647_7968.t19 a_52753_24325.t4 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3270 a_70513_19926.t3 a_70459_20811.t7 a_70513_20044.t2 VDD.t956 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3271 a_4825_1255.t1 a_70509_1028.t9 VDD.t2755 VDD.t2754 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3272 a_53891_18572.t1 a_55862_18700.t9 VDD.t2506 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3273 VDD.t3336 a_8056_15820.t6 a_10509_14454.t10 VDD.t3335 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3274 VDD.t4498 a_64117_8794.t12 a_67133_11394.t6 VDD.t4497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3275 a_59929_6884.t0 a_55469_11532.t17 VDD.t958 VDD.t957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3276 VDD.t3215 opcode[0].t207 a_26279_20719.t1 VDD.t3214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3277 a_51695_9365.t2 a_51105_9802.t9 VDD.t1347 VDD.t1346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3278 a_54790_6842.t6 a_51059_8126.t16 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3279 VSS.t146 a_59635_6910.t14 a_60988_7603.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3280 a_7432_1744.t1 a_7957_1259.t7 a_7083_1744.t6 VDD.t2900 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3281 a_70509_13650.t2 a_56556_21365.t11 a_70509_13768.t2 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3282 a_30152_6681.t3 opcode[0].t208 VSS.t517 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3283 a_16859_20723.t0 opcode[0].t209 VDD.t3217 VDD.t3216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3284 VDD.t340 a_30647_7968.t20 a_54113_22058.t0 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3285 VDD.t3219 opcode[0].t210 a_30152_10818.t0 VDD.t3218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3286 a_37902_9782.t1 a_35602_9612.t15 VDD.t953 VDD.t952 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3287 a_9879_4622.t0 a_10173_5328.t7 a_1039_8966.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3288 a_16573_1740.t2 a_16264_11724.t7 VDD.t466 VDD.t465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3289 a_53246_6110.t0 a_48254_6910.t20 a_53010_6842.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3290 a_39807_6822.t0 a_39262_7515.t7 a_39689_6822.t5 VDD.t3223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3291 VDD.t1125 a_40373_9071.t5 a_41369_9658.t2 VDD.t1124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3292 VDD.t2844 a_22608_8258.t11 a_22550_8988.t0 VDD.t2843 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3293 a_41493_21373.t10 A[0].t26 VDD.t2336 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3294 a_53005_1041.t4 a_52460_1734.t7 a_53005_309.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3295 a_52892_6842.t0 a_48254_6910.t21 VDD.t915 VDD.t914 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3296 a_15426_6045.t0 B[4].t24 VDD.t1876 VDD.t1875 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3297 a_17501_10851.t3 opcode[1].t116 VSS.t682 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3298 VSS.t692 a_64185_771.t12 a_65224_3811.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3299 a_59871_6178.t0 a_54713_3294.t16 a_59635_6910.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3300 a_6962_16408.t0 B[5].t37 VDD.t2415 VDD.t2414 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3301 a_19454_10990.t5 a_19396_14454.t6 a_19987_11720.t7 VDD.t2431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3302 VSS.t593 a_35594_7027.t17 a_38153_7495.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3303 a_23080_20259.t1 A[0].t27 VSS.t365 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3304 VDD.t3994 A[2].t40 a_22489_21592.t3 VDD.t3993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3305 a_11829_5352.t3 A[6].t49 VDD.t1465 VDD.t1464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3306 a_57731_748.t1 a_57676_2326.t17 VDD.t1711 VDD.t1710 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3307 a_30150_n1593.t2 opcode[0].t211 VSS.t518 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3308 a_61533_6910.t7 a_61827_6884.t6 a_61415_6910.t10 VDD.t3141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3309 a_61407_1042.t8 a_60980_1735.t6 a_61525_1042.t3 VDD.t2842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3310 a_1099_8992.t10 opcode[0].t212 VDD.t3221 VDD.t3220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3311 a_47719_15761.t9 a_30645_n306.t19 VDD.t3110 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3312 a_22540_14454.t1 a_22598_13724.t10 VDD.t2494 VDD.t2493 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3313 VDD.t2256 a_3652_8992.t6 a_4233_11724.t8 VDD.t2255 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3314 VDD.t1878 B[4].t25 a_34985_4186.t0 VDD.t1877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3315 VDD.t2780 a_46916_3289.t7 a_47912_3876.t0 VDD.t2779 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3316 a_14548_7659.t0 opcode[0].t213 a_13188_8262.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3317 a_3058_20866.t5 a_4237_20723.t5 a_3591_21596.t9 VDD.t4191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3318 a_23081_8962.t5 a_23700_6043.t7 a_24240_5350.t9 VDD.t1480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3319 a_43391_21373.t6 opcode[0].t214 VDD.t2365 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3320 a_40305_20642.t3 a_39715_21079.t8 VSS.t538 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3321 VDD.t3542 A[3].t46 a_61098_21369.t9 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3322 VDD.t2367 opcode[0].t215 a_23141_8988.t0 VDD.t2366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3323 a_20526_411.t0 a_19146_1744.t5 a_20054_1744.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3324 a_19987_14454.t7 a_11565_15824.t6 VDD.t2749 VDD.t2748 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3325 a_38484_3565.t1 a_37894_4002.t9 VDD.t4555 VDD.t4554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3326 a_70513_16782.t6 a_70459_17667.t6 a_71846_17491.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3327 VDD.t519 a_13178_13728.t11 a_13120_14458.t0 VDD.t518 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3328 a_16084_4620.t1 a_16378_5326.t7 a_10459_8962.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3329 a_59322_18605.t4 a_59262_18579.t6 VDD.t990 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3330 a_8192_13121.t1 opcode[0].t216 a_6832_13724.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3331 a_16274_8992.t1 a_16332_8262.t10 VDD.t1723 VDD.t1722 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3332 VDD.t2369 opcode[0].t217 a_16213_21596.t1 VDD.t2368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3333 a_1392_407.t1 a_498_11724.t7 VSS.t101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3334 VDD.t1617 a_48815_11511.t16 a_52892_6842.t4 VDD.t1616 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3335 Y[1].t3 a_20086_n2148.t11 VSS.t661 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3336 VDD.t4419 A[3].t47 a_59320_21075.t1 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3337 a_59222_15037.t1 a_58326_16165.t17 VSS.t162 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3338 a_30647_7968.t6 a_30154_8749.t6 a_29954_7911.t10 VDD.t4294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3339 a_57736_2352.t4 a_55504_n1325.t17 VDD.t495 VDD.t494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3340 a_48426_24202.t3 a_46818_20639.t6 VSS.t14 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3341 VSS.t601 A[7].t32 a_4491_15753.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3342 a_39263_15765.t8 a_38723_16458.t6 a_39381_15765.t6 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3343 a_40227_9654.t3 a_38501_6091.t7 a_40109_9654.t2 VDD.t1105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3344 a_61415_6910.t8 a_61827_6884.t7 a_61533_6910.t5 VDD.t2877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3345 a_51704_6111.t3 a_51114_6548.t10 VSS.t556 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3346 a_49904_21370.t9 a_49477_22063.t7 a_50022_21370.t5 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3347 a_10509_14454.t11 a_8056_15820.t7 VDD.t4190 VDD.t4189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3348 a_26279_20719.t0 opcode[0].t218 VDD.t2371 VDD.t2370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3349 VSS.t188 a_40373_9071.t6 a_41251_9658.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3350 a_39254_1735.t0 a_35591_989.t18 VDD.t3563 VDD.t3562 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3351 a_13711_14458.t5 opcode[0].t219 VDD.t2373 VDD.t2372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3352 a_17501_13585.t3 opcode[0].t220 VSS.t377 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3353 a_51342_9165.t1 a_48815_11511.t17 a_51105_9802.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3354 a_41361_3878.t4 a_38498_1915.t6 a_41243_3878.t3 VDD.t666 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3355 a_20558_n3481.t1 a_19178_n2148.t4 a_20086_n2148.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3356 VDD.t1040 a_70509_13650.t11 a_17447_1255.t0 VDD.t1039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3357 a_53430_9674.t0 a_51704_6111.t7 a_53312_9674.t0 VDD.t2517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3358 a_10259_n2148.t6 a_11133_n2633.t7 a_10608_n2148.t2 VDD.t661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3359 a_20643_8115.t0 opcode[0].t221 VDD.t2375 VDD.t2374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3360 VDD.t3426 A[5].t47 a_14310_5328.t0 VDD.t3425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3361 VDD.t3348 a_19396_11720.t7 a_19705_1744.t6 VDD.t3347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3362 a_13661_8966.t7 a_17495_6045.t7 a_18035_5352.t8 VDD.t2122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3363 a_57739_6616.t4 a_57684_8194.t16 VDD.t2818 VDD.t2817 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3364 a_45050_6179.t0 a_44460_6616.t10 VDD.t1258 VDD.t1257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3365 a_63764_8594.t1 A[3].t48 a_63527_9231.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3366 a_46228_21076.t0 A[1].t40 VDD.t2578 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3367 a_19987_11720.t6 a_19396_14454.t7 a_19454_10990.t6 VDD.t2432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3368 a_6827_15753.t2 A[5].t48 a_6962_16408.t5 VDD.t3427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3369 a_65651_3118.t5 a_66063_3092.t7 a_65769_3118.t2 VDD.t516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3370 VDD.t1908 B[3].t33 a_35001_1426.t3 VDD.t1907 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3371 a_30643_1763.t1 a_30150_1105.t7 a_29950_1706.t6 VDD.t3670 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3372 a_39675_15739.t2 a_39618_16432.t15 VDD.t2650 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3373 a_70509_10506.t0 a_70455_11391.t7 a_70509_10624.t7 VDD.t2839 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3374 a_61525_1042.t6 a_60980_1735.t7 a_61525_310.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3375 VDD.t2417 B[5].t38 a_13358_6047.t0 VDD.t2416 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3376 VDD.t182 a_35575_3749.t16 a_39681_1042.t8 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3377 a_60201_9159.t3 a_59937_9742.t8 VDD.t2551 VDD.t2550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3378 VDD.t628 a_54903_1041.t21 a_59921_1016.t0 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3379 VDD.t3136 a_42761_15445.t10 a_41153_18571.t0 w_42667_15409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3380 a_13178_13728.t6 a_13651_14432.t5 a_13711_14458.t10 VDD.t3786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3381 a_19997_8988.t11 a_7551_6363.t7 VDD.t4596 VDD.t4595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3382 a_19563_6043.t2 B[2].t19 VDD.t1355 VDD.t1354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3383 a_47703_1733.t0 a_46350_1040.t15 VDD.t4435 VDD.t4434 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3384 a_51699_310.t0 a_51109_747.t9 VDD.t3361 VDD.t3360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3385 a_41493_21373.t8 a_30647_12105.t15 VDD.t1494 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3386 VDD.t3774 A[7].t33 a_9761_5354.t9 VDD.t3773 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3387 a_19705_1744.t4 a_19146_1744.t6 a_20054_1744.t3 VDD.t2534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3388 VDD.t2490 a_22598_13724.t11 a_22540_14454.t0 VDD.t2489 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3389 a_65651_3118.t11 a_64185_771.t13 VDD.t4458 VDD.t4457 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3390 VDD.t4460 a_64185_771.t14 a_67135_3808.t6 VDD.t4459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3391 VSS.t565 a_35591_989.t19 a_39254_1735.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3392 a_49314_17045.t5 a_30645_n306.t20 VDD.t3111 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3393 a_70455_14535.t3 opcode[1].t117 VSS.t683 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3394 a_3591_21596.t10 a_4237_20723.t6 a_3058_20866.t6 VDD.t4192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3395 a_61098_21369.t8 A[3].t49 VDD.t4418 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3396 VDD.t2751 a_11565_15824.t7 a_19987_14454.t6 VDD.t2750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3397 a_63764_5561.t0 A[4].t48 a_63527_6198.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3398 VDD.t1296 a_9928_8988.t7 a_10509_11720.t5 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3399 a_13429_1740.t11 a_14303_1255.t7 a_13778_1740.t7 VDD.t3659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3400 VSS.t213 a_15297_16387.t8 a_4173_14432.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3401 VDD.t2377 opcode[0].t222 a_14367_8119.t0 VDD.t2376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3402 VDD.t991 a_59262_18579.t7 a_59322_18605.t3 w_59093_17960# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3403 VSS.t542 a_6887_15819.t6 a_8192_13121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3404 VDD.t4531 a_54713_3294.t17 a_59090_7603.t0 VDD.t4530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3405 a_16213_21596.t0 opcode[0].t223 VDD.t2379 VDD.t2378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3406 VSS.t378 opcode[0].t224 a_39952_20442.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3407 a_22172_5352.t11 a_21632_6045.t7 a_19937_8962.t7 VDD.t4448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3408 a_12241_5326.t0 A[6].t50 VDD.t1467 VDD.t1466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3409 a_54449_3877.t3 a_51704_1914.t7 a_54567_3877.t3 VDD.t3644 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3410 VDD.t2344 a_566_8262.t11 a_508_8992.t0 VDD.t2343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3411 a_61079_9746.t1 a_58334_7783.t7 a_61197_9746.t2 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3412 a_30152_6681.t0 opcode[0].t225 VDD.t2381 VDD.t2380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3413 a_59320_21075.t0 A[3].t50 VDD.t4417 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3414 a_58986_15769.t0 a_59223_16436.t15 a_59222_15037.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3415 a_46823_22243.t3 a_46233_22680.t10 VSS.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3416 VSS.t585 a_13849_16387.t10 a_1029_14432.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3417 VDD.t315 a_9976_13724.t9 a_9918_14454.t1 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3418 a_38139_9145.t0 a_35602_9612.t16 a_37902_9782.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3419 VDD.t4103 a_42301_n1318.t16 a_44445_4000.t0 VDD.t4102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3420 VDD.t1310 a_56366_23618.t17 a_62996_21369.t3 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3421 a_39381_15765.t7 a_38723_16458.t7 a_39263_15765.t9 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3422 a_23131_14454.t3 opcode[0].t226 VDD.t2383 VDD.t2382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3423 a_23131_11720.t11 a_22540_14454.t7 a_22598_10990.t7 VDD.t4586 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3424 a_41507_3295.t0 a_41243_3878.t8 VDD.t3369 VDD.t3368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3425 a_40219_3874.t0 a_38493_311.t6 a_40101_3874.t3 VDD.t753 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3426 a_64122_11365.t3 a_63532_11802.t9 VSS.t338 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3427 a_20086_n2148.t0 a_20611_n2633.t7 a_19737_n2148.t0 VDD.t632 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3428 a_46470_22043.t0 a_43319_23626.t16 a_46233_22680.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3429 VDD.t3377 a_6887_15819.t7 a_7365_14454.t0 VDD.t3376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3430 a_30647_7968.t0 opcode[0].t227 a_31379_8204.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3431 Y[4].t0 a_10608_n2148.t10 VDD.t875 VDD.t874 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3432 VDD.t3112 a_30645_n306.t21 a_49328_18695.t4 w_49234_18659# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3433 a_40101_6796.t3 a_35602_9612.t17 VSS.t154 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3434 a_70509_13650.t4 a_70455_14535.t7 a_70509_13768.t6 VDD.t1659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3435 VDD.t2385 opcode[0].t228 a_29952_9980.t3 VDD.t2384 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3436 VDD.t1129 a_52710_16433.t14 a_52355_15766.t0 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3437 VDD.t2387 opcode[0].t229 a_13711_14458.t4 VDD.t2386 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3438 VDD.t3098 opcode[3].t54 a_6556_n2148.t2 VDD.t3097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3439 a_30643_n2374.t5 a_30150_n1593.t6 a_29950_n2431.t9 VDD.t4350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3440 a_56438_21365.t11 a_49832_23623.t13 VDD.t998 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3441 VDD.t4500 a_64117_8794.t13 a_66061_10678.t1 VDD.t4499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3442 Cout.t0 a_39582_17945.t8 VDD.t3615 w_39488_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3443 a_52753_24325.t1 A[2].t41 VDD.t3995 w_52599_24263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3444 VDD.t3299 a_45279_16157.t16 a_49314_17045.t0 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3445 VDD.t3516 a_62366_15449.t10 a_60758_18575.t3 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3446 a_10459_8962.t3 a_15426_6045.t7 a_15966_5352.t10 VDD.t2743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3447 VSS.t142 opcode[2].t53 a_3392_1740.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3448 VDD.t4105 a_42301_n1318.t17 a_45805_1733.t0 VDD.t4104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3449 a_61533_6910.t4 a_60988_7603.t7 a_61533_6178.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3450 VDD.t1079 a_51059_8126.t17 a_51114_6548.t0 VDD.t1078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3451 a_7315_8962.t4 A[5].t49 a_14252_4622.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3452 a_7464_n2148.t0 a_7989_n2633.t5 a_7115_n2148.t2 VDD.t3151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3453 Y[6].t3 a_4332_n2152.t11 VSS.t206 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3454 VDD.t2388 opcode[0].t230 a_39715_21079.t2 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3455 a_10337_15751.t2 A[2].t42 a_10472_16406.t5 VDD.t3996 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3456 a_23777_13581.t2 opcode[0].t231 VDD.t2390 VDD.t2389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3457 VSS.t280 a_16332_8262.t11 a_16274_8992.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3458 a_45035_3563.t0 a_44445_4000.t10 VDD.t2856 VDD.t2855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3459 VDD.t2782 a_43319_23626.t17 a_46228_21076.t5 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3460 a_6962_16408.t4 A[5].t50 a_6827_15753.t3 VDD.t3428 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3461 a_48542_1014.t2 a_44399_2324.t15 VSS.t654 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3462 a_16573_1740.t4 a_17447_1255.t6 a_16922_1740.t1 VDD.t3576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3463 a_70513_4160.t7 a_70459_5045.t7 a_70513_4278.t8 VDD.t1960 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3464 a_59517_6910.t10 a_59090_7603.t7 a_59635_6910.t5 VDD.t3654 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3465 a_11947_4620.t1 a_12241_5326.t5 a_4183_8966.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3466 a_63114_21369.t7 a_62569_22062.t5 a_62996_21369.t11 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3467 VDD.t3525 a_59320_21075.t9 a_59910_20638.t2 w_59166_21013# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3468 VDD.t2618 B[7].t18 a_9761_5354.t3 VDD.t2617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3469 VSS.t270 a_37856_8106.t17 a_41941_6090.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3470 a_13711_14458.t11 a_13651_14432.t6 a_13178_13728.t7 VDD.t3787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3471 a_66063_n1256.t0 a_48248_1040.t19 VDD.t2876 VDD.t2875 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3472 VDD.t3100 opcode[3].t55 a_7115_n2148.t3 VDD.t3099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3473 a_65769_3118.t6 a_65224_3811.t7 a_65769_2386.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3474 a_70459_20811.t0 opcode[1].t118 VDD.t4360 VDD.t4359 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3475 a_70509_13768.t4 a_65767_10704.t10 VDD.t451 VDD.t450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3476 VDD.t1495 a_30647_12105.t16 a_41493_21373.t7 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3477 VDD.t2225 B[0].t20 a_24157_16385.t1 VDD.t2224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3478 VDD.t2912 a_22821_n2174.t7 a_22881_n2148.t4 VDD.t2911 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3479 VDD.t858 opcode[2].t54 a_3951_1740.t1 VDD.t857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3480 VDD.t4416 A[3].t51 a_61510_21343.t1 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3481 VDD.t3113 a_30645_n306.t22 a_49314_17045.t4 w_49220_17009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3482 a_46658_9742.t3 a_45050_6179.t7 VSS.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3483 a_65769_5881.t0 a_66063_6587.t7 VSS.t325 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3484 a_3058_20866.t7 a_4237_20723.t7 a_3591_21596.t11 VDD.t4193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3485 a_43803_21347.t0 opcode[0].t232 VDD.t2391 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3486 a_60329_17945.t3 a_60758_18575.t5 a_60464_18601.t2 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3487 VDD.t860 opcode[2].t55 a_22849_1744.t1 VDD.t859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3488 a_47417_18593.t4 a_47711_18567.t6 a_47282_17937.t3 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3489 a_57744_8220.t3 a_57684_8194.t17 VDD.t2346 VDD.t2345 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3490 a_35241_6827.t1 B[3].t34 a_35004_7464.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3491 a_40101_3874.t2 a_38493_311.t7 VSS.t128 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3492 a_40296_23896.t3 a_39706_24333.t10 VSS.t586 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3493 a_16922_1740.t0 a_17447_1255.t7 a_16573_1740.t3 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3494 VDD.t1313 a_55504_n1325.t18 a_57722_4002.t1 VDD.t1312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3495 a_48136_6910.t7 a_46356_6910.t13 VDD.t2649 VDD.t2648 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3496 a_15680_20866.t6 a_16859_20723.t6 a_16213_21596.t9 VDD.t3057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3497 a_839_n2152.t5 a_779_n2178.t7 VDD.t2727 VDD.t2726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3498 a_41493_21373.t1 a_41066_22066.t6 a_41611_21373.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3499 VDD.t1468 A[6].t51 a_47719_15761.t3 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3500 a_20103_5350.t3 a_20515_5324.t7 a_16805_8966.t3 VDD.t1043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3501 VDD.t3503 a_55853_15446.t9 a_54245_18572.t1 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3502 a_39263_15765.t6 a_39675_15739.t6 a_39381_15765.t3 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3503 VDD.t2393 opcode[0].t233 a_23131_14454.t2 VDD.t2392 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3504 a_30645_n306.t6 opcode[0].t234 a_31377_n70.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3505 a_13461_n2152.t0 a_13401_n2178.t7 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3506 a_39681_1042.t3 a_40093_1016.t7 a_39799_1042.t1 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3507 a_63835_3641.t0 B[4].t26 a_63598_4278.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3508 a_26460_20259.t0 opcode[0].t235 a_25100_20862.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3509 a_9228_15824.t1 a_9168_15798.t7 VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3510 VDD.t3776 A[7].t34 a_10173_5328.t0 VDD.t3775 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3511 VSS.t237 a_30647_12105.t17 a_39957_22046.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3512 VSS.t183 a_46140_17941.t8 a_38721_16161.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3513 VDD.t3536 a_61079_9746.t7 a_61343_9163.t2 VDD.t3535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3514 VSS.t419 B[7].t19 a_9221_6047.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3515 VDD.t2135 a_4300_1740.t11 a_4857_n2637.t3 VDD.t2134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3516 VDD.t2018 A[4].t49 a_41711_n1755.t6 VDD.t2017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3517 a_54713_3294.t3 a_54449_3877.t8 VSS.t579 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3518 a_13711_14458.t3 opcode[0].t236 VDD.t2395 VDD.t2394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3519 a_67135_7303.t0 a_64188_3841.t13 VDD.t473 VDD.t472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3520 VDD.t999 a_49832_23623.t14 a_56438_21365.t10 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3521 a_66061_10678.t0 a_64117_8794.t14 VDD.t4502 VDD.t4501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3522 a_61343_9163.t3 a_61079_9746.t8 VSS.t560 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3523 a_6556_n2148.t1 opcode[3].t56 VDD.t4268 VDD.t4267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3524 a_7432_1744.t7 a_6524_1744.t7 a_7083_1744.t11 VDD.t4258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3525 a_59910_20638.t3 a_59320_21075.t10 VSS.t559 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3526 VDD.t1357 B[2].t20 a_30154_7310.t2 VDD.t1356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3527 VDD.t3409 a_55469_11532.t18 a_59517_6910.t3 VDD.t3408 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3528 a_6202_20866.t0 a_7381_20723.t7 a_6735_21596.t0 VDD.t4150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3529 a_62366_15449.t4 a_58326_16165.t18 VDD.t987 w_62272_15413# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3530 a_30645_10037.t5 a_30152_10818.t7 a_29952_9980.t9 VDD.t2364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3531 VDD.t171 a_41507_3295.t17 a_44465_8220.t0 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3532 a_12478_20862.t7 a_13657_20719.t7 a_13011_21592.t8 VDD.t2035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3533 a_70509_1146.t0 a_45939_15761.t11 a_70509_1028.t0 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3534 VDD.t1470 A[6].t52 a_48265_n1750.t6 VDD.t1469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3535 a_54785_1041.t5 a_55197_1015.t7 a_54903_1041.t2 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3536 a_38131_3365.t1 a_35575_3749.t17 a_37894_4002.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3537 VDD.t3656 a_6202_20866.t10 a_3923_n2178.t2 VDD.t3655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3538 a_39618_16432.t3 a_40621_16458.t5 a_41161_15765.t7 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3539 a_18447_5326.t0 A[3].t52 VDD.t4415 VDD.t4414 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3540 a_7115_n2148.t1 a_7989_n2633.t6 a_7464_n2148.t1 VDD.t3152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3541 a_58312_3565.t0 a_57722_4002.t10 VDD.t1430 VDD.t1429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3542 VDD.t447 a_10397_15824.t6 a_16855_14458.t2 VDD.t446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3543 VDD.t554 a_61533_6910.t10 a_70509_1146.t4 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3544 a_4418_20263.t0 opcode[0].t237 a_3058_20866.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3545 a_39715_21079.t1 opcode[0].t238 VDD.t3245 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3546 a_10227_1744.t3 a_9668_1744.t7 a_10576_1744.t0 VDD.t1691 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3547 VDD.t1496 a_30647_12105.t18 a_39720_22683.t6 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3548 a_46228_21076.t4 a_43319_23626.t18 VDD.t2783 w_46074_21014# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3549 a_6827_15753.t4 A[5].t51 a_6962_16408.t3 VDD.t3429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3550 a_54665_15740.t0 a_30643_1763.t23 VDD.t77 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3551 a_35004_7464.t1 B[3].t35 VDD.t1910 VDD.t1909 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3552 VDD.t4165 a_44399_2324.t16 a_48130_1040.t4 VDD.t4164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3553 VSS.t53 a_9976_13724.t10 a_9918_14454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3554 a_23732_7655.t1 a_23081_8962.t11 VSS.t108 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3555 VSS.t420 B[7].t20 a_30150_n3032.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3556 a_54908_6842.t7 a_55202_6816.t7 a_54790_6842.t0 VDD.t2056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3557 a_56438_21365.t7 a_56850_21339.t6 a_56556_21365.t6 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3558 a_30647_12105.t6 a_30154_11447.t7 a_29954_12048.t9 VDD.t3909 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3559 VDD.t3125 a_39807_6822.t14 a_41587_6822.t6 VDD.t3124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3560 VDD.t3247 opcode[0].t239 a_29950_n2431.t4 VDD.t3246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3561 a_51356_7515.t0 a_51059_8126.t18 a_51119_8152.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3562 VDD.t3249 opcode[0].t240 a_29952_5843.t1 VDD.t3248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3563 a_39689_6822.t9 a_40101_6796.t7 a_39807_6822.t5 VDD.t4283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3564 a_62996_21369.t6 a_62569_22062.t6 a_63114_21369.t1 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3565 VDD.t2679 a_13188_8262.t10 a_13130_8992.t2 VDD.t2678 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3566 VDD.t1880 B[4].t27 a_30152_3173.t0 VDD.t1879 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3567 a_13661_8966.t5 A[3].t53 a_18389_4620.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3568 a_16804_20263.t0 A[2].t43 VSS.t631 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3569 a_16795_14432.t1 a_21211_16387.t9 VDD.t3353 VDD.t3352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3570 a_4233_14458.t1 a_4879_13585.t6 a_3700_13728.t2 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3571 a_51100_4001.t1 a_48064_9163.t18 VDD.t648 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3572 a_38501_6091.t3 a_37911_6528.t10 VDD.t2165 VDD.t2164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3573 a_41493_21373.t6 a_30647_12105.t19 VDD.t1497 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3574 a_24157_16385.t0 B[0].t21 VDD.t2227 VDD.t2226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3575 a_29952_n363.t0 B[6].t37 VDD.t3314 VDD.t3313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3576 a_10576_1744.t5 a_11101_1259.t7 a_10227_1744.t9 VDD.t790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3577 a_58868_15769.t3 a_59280_15743.t7 a_58986_15769.t1 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3578 a_7083_1744.t4 opcode[2].t56 VDD.t862 VDD.t861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3579 a_61510_21343.t0 A[3].t54 VDD.t3552 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3580 a_60464_18601.t1 a_60758_18575.t6 a_60329_17945.t2 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3581 a_16855_14458.t3 opcode[0].t241 VDD.t3251 VDD.t3250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3582 VDD.t1619 a_48815_11511.t18 a_51105_9802.t3 VDD.t1618 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3583 VDD.t3431 A[5].t52 a_13898_5354.t3 VDD.t3430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3584 a_43055_24209.t2 a_40310_22246.t6 VSS.t668 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3585 a_60055_9742.t3 a_58329_6179.t7 a_59937_9742.t1 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3586 VDD.t3253 opcode[0].t242 a_29950_1706.t3 VDD.t3252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3587 VDD.t475 a_64188_3841.t14 a_65224_7306.t1 VDD.t474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3588 a_47282_17937.t4 a_47711_18567.t7 a_47417_18593.t3 w_47188_17948# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3589 VDD.t4270 opcode[3].t57 a_22322_n2148.t0 VDD.t4269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3590 a_48254_6910.t3 a_47709_7603.t6 a_48254_6178.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3591 a_39715_21079.t5 A[0].t28 VDD.t2294 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3592 a_19997_8988.t1 opcode[0].t243 VDD.t3255 VDD.t3254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3593 a_19737_n2148.t5 a_19178_n2148.t5 a_20086_n2148.t5 VDD.t2284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3594 a_41611_21373.t1 a_41066_22066.t7 a_41493_21373.t0 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3595 a_47719_15761.t2 A[6].t53 VDD.t1471 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3596 a_13178_10994.t1 a_14357_10851.t5 a_13711_11724.t7 VDD.t2675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3597 VSS.t238 a_30647_12105.t20 a_39943_23696.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3598 a_47918_9746.t3 a_46922_9159.t7 VDD.t2120 VDD.t2119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3599 a_61216_21369.t5 a_61510_21343.t6 a_61098_21369.t6 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3600 a_10397_15824.t1 a_10337_15751.t6 VDD.t3507 VDD.t3506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3601 a_54245_18572.t0 a_55853_15446.t10 VDD.t3504 w_55759_15410# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3602 a_7315_8962.t0 a_13358_6047.t7 a_13898_5354.t6 VDD.t2908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3603 a_39381_15765.t0 a_39675_15739.t7 a_39263_15765.t4 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3604 a_23131_14454.t1 opcode[0].t244 VDD.t3257 VDD.t3256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3605 a_66003_9972.t1 a_41705_6822.t18 a_65767_10704.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3606 a_48855_n1313.t2 a_48265_n1750.t10 VSS.t75 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3607 VDD.t414 a_9168_15798.t8 a_9228_15824.t0 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3608 a_556_13728.t6 a_1735_13585.t5 a_1089_14458.t8 VDD.t2526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3609 a_30645_10037.t7 opcode[0].t245 a_31377_10273.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3610 a_14302_10391.t1 a_13120_14458.t7 VSS.t623 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3611 a_63602_n1637.t5 A[3].t55 VDD.t3551 VDD.t3550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3612 a_38493_311.t0 a_37903_748.t10 VDD.t1119 VDD.t1118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3613 a_46140_17941.t2 a_46215_18571.t7 VSS.t106 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3614 a_43391_21373.t10 a_43803_21347.t6 a_43509_21373.t6 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3615 VDD.t3778 A[7].t35 a_1974_8339.t1 VDD.t3777 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3616 a_44691_109.t1 a_41697_1042.t22 a_44454_746.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3617 a_7989_n2633.t0 a_7432_1744.t11 VDD.t2689 VDD.t2688 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3618 VDD.t864 opcode[2].t57 a_7083_1744.t3 VDD.t863 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3619 a_38148_5891.t0 a_35602_9612.t18 a_37911_6528.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3620 VDD.t307 a_40373_9071.t7 a_41369_9658.t0 VDD.t306 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3621 a_51119_8152.t0 a_51059_8126.t19 VDD.t1081 VDD.t1080 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3622 a_41711_n1755.t5 A[4].t50 VDD.t2020 VDD.t2019 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3623 a_45049_1913.t1 a_44459_2350.t10 VDD.t3143 VDD.t3142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3624 a_46232_1040.t3 a_42301_n1318.t18 VDD.t4107 VDD.t4106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3625 VDD.t4272 opcode[3].t58 a_6556_n2148.t0 VDD.t4271 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3626 a_16605_n2152.t6 a_16046_n2152.t7 a_16954_n2152.t5 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3627 a_61120_15037.t1 A[4].t51 VSS.t323 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3628 a_48265_n1750.t5 A[6].t54 VDD.t1473 VDD.t1472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3629 a_7464_n2148.t2 a_7989_n2633.t7 a_7115_n2148.t0 VDD.t3153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3630 a_46586_308.t0 a_42301_n1318.t19 a_46350_1040.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3631 a_3923_n2178.t3 a_6202_20866.t11 VDD.t3658 VDD.t3657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3632 a_52809_18602.t5 a_52749_18576.t5 VDD.t1250 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3633 a_41161_15765.t0 a_40621_16458.t6 a_39618_16432.t2 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3634 a_54572_9678.t5 a_51709_7715.t6 a_54454_9678.t2 VDD.t2791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3635 VSS.t402 VSS.t401 a_4418_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3636 VDD.t3258 opcode[0].t246 a_39715_21079.t0 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3637 a_30150_n3032.t0 B[7].t21 VDD.t2620 VDD.t2619 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3638 VSS.t382 B[5].t39 a_30150_1105.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3639 a_65224_3811.t3 a_64185_771.t15 VDD.t4462 VDD.t4461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3640 a_39720_22683.t5 a_30647_12105.t21 VDD.t1498 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3641 a_1099_8992.t11 opcode[0].t247 VDD.t3260 VDD.t3259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3642 VSS.t699 a_64117_8794.t15 a_66003_9972.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3643 a_52709_15034.t1 a_51813_16162.t18 VSS.t482 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3644 VDD.t988 a_58326_16165.t19 a_58328_16462.t0 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3645 a_37902_9782.t4 a_35594_7027.t18 VDD.t3723 VDD.t3722 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3646 VDD.t4080 a_48124_21370.t13 a_49477_22063.t2 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3647 VSS.t166 a_49832_23623.t15 a_52999_20434.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3648 a_63114_21369.t2 a_62569_22062.t7 a_62996_21369.t7 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3649 Y[2].t3 a_16954_n2152.t11 VSS.t314 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3650 a_53010_6110.t0 a_53304_6816.t6 VSS.t406 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3651 a_11829_5352.t10 a_12241_5326.t6 a_4183_8966.t6 VDD.t2258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3652 VDD.t2483 a_12478_20862.t10 a_10199_n2174.t1 VDD.t2482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3653 a_15680_20866.t5 a_16859_20723.t7 a_16804_20263.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3654 VDD.t3355 a_21211_16387.t10 a_16795_14432.t2 VDD.t3354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3655 VDD.t2022 A[4].t52 a_5331_6357.t0 VDD.t2021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3656 a_57684_8194.t0 a_61071_3878.t8 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3657 a_38484_3565.t0 a_37894_4002.t10 VDD.t4557 VDD.t4556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3658 a_3700_13728.t3 a_4879_13585.t7 a_4233_14458.t2 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3659 VDD.t2295 A[0].t29 a_41493_21373.t9 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3660 a_52749_18576.t1 a_53816_17942.t7 VDD.t2741 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3661 VDD.t2297 A[0].t30 a_24157_16385.t4 VDD.t2296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3662 VDD.t1621 a_48815_11511.t19 a_52892_6842.t3 VDD.t1620 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3663 a_48064_9163.t3 a_47800_9746.t8 VSS.t563 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3664 a_60329_17945.t1 a_60758_18575.t7 a_60464_18601.t0 w_60235_17956# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3665 a_16322_13728.t5 a_17501_13585.t5 a_16855_14458.t10 VDD.t1990 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3666 a_23958_10387.t0 opcode[1].t119 a_22598_10990.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3667 VSS.t588 a_42177_23622.t6 a_43055_24209.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3668 a_22598_10990.t1 a_23777_10847.t7 a_23131_11720.t6 VDD.t3699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3669 VDD.t2757 a_70509_1028.t10 a_4825_1255.t0 VDD.t2756 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3670 a_55469_11532.t3 a_54879_11969.t8 VSS.t333 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3671 VDD.t2580 A[1].t41 a_22709_16385.t5 VDD.t2579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3672 a_41676_11949.t3 B[4].t28 VDD.t1882 VDD.t1881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3673 a_40227_9654.t0 a_38492_9345.t7 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3674 VDD.t4437 a_46356_6910.t14 a_47709_7603.t3 VDD.t4436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3675 VDD.t2298 A[0].t31 a_39715_21079.t4 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3676 a_49319_15441.t4 a_45279_16157.t17 VDD.t3300 w_49225_15405# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3677 a_14302_13125.t0 a_13651_14432.t7 VSS.t602 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3678 a_13429_1740.t2 a_12870_1740.t7 a_13778_1740.t3 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3679 a_58334_7783.t3 a_57744_8220.t10 VSS.t509 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3680 a_39720_22683.t0 opcode[0].t248 VDD.t3261 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3681 a_20086_n2148.t4 a_19178_n2148.t6 a_19737_n2148.t4 VDD.t2285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3682 VSS.t229 A[6].t55 a_47179_16454.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3683 a_59325_22679.t4 a_56366_23618.t18 VDD.t1311 w_59171_22617# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3684 a_13711_11724.t8 a_14357_10851.t6 a_13178_10994.t0 VDD.t3128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3685 a_20003_20723.t0 opcode[0].t249 VDD.t3263 VDD.t3262 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3686 a_61098_21369.t7 a_61510_21343.t7 a_61216_21369.t6 w_60634_22000# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3687 VDD.t3509 a_10337_15751.t7 a_10397_15824.t2 VDD.t3508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3688 VDD.t2229 B[0].t22 a_30154_11447.t0 VDD.t2228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3689 VSS.t443 a_70509_1028.t11 a_4825_1255.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3690 a_48544_24202.t0 a_46818_20639.t7 a_48426_24202.t0 w_48390_24140# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3691 a_9867_21592.t11 opcode[0].t250 VDD.t3265 VDD.t3264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3692 a_41361_3878.t3 a_38498_1915.t7 a_41243_3878.t2 VDD.t667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3693 a_13178_10994.t3 a_14357_10851.t7 a_14302_10391.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3694 VDD.t3549 A[3].t56 a_63602_n1637.t4 VDD.t3548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3695 VSS.t690 a_46569_18571.t6 a_46140_17941.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3696 a_8130_16410.t0 B[4].t29 VDD.t1884 VDD.t1883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3697 a_20633_13581.t1 opcode[0].t251 VDD.t3267 VDD.t3266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3698 a_6735_21596.t7 A[5].t53 a_6202_20866.t6 VDD.t3432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3699 a_9928_8988.t0 a_9986_8258.t11 VDD.t3573 VDD.t3572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3700 a_62660_24205.t4 a_59915_22242.t7 VSS.t405 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3701 a_43509_21373.t0 a_43803_21347.t7 a_43391_21373.t9 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3702 a_59509_1042.t4 a_55504_n1325.t19 VDD.t1315 VDD.t1314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3703 a_41999_6796.t0 a_37856_8106.t18 VDD.t1662 VDD.t1661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3704 VDD.t2024 A[4].t53 a_41711_n1755.t4 VDD.t2023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3705 VDD.t3269 opcode[0].t252 a_29952_n363.t8 VDD.t3268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3706 VDD.t477 a_64188_3841.t15 a_65651_6613.t1 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3707 a_58329_6179.t0 a_57739_6616.t10 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3708 VDD.t866 opcode[2].t58 a_3392_1740.t0 VDD.t865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3709 VDD.t1886 B[4].t30 a_63598_4278.t1 VDD.t1885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3710 VSS.t577 a_47282_17937.t8 a_46215_18571.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3711 VDD.t4274 opcode[3].t59 a_16605_n2152.t4 VDD.t4273 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3712 VDD.t4513 a_59929_3874.t8 a_60193_3291.t0 VDD.t4512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3713 VDD.t1888 B[4].t31 a_18243_16385.t1 VDD.t1887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3714 VDD.t2671 a_6832_10990.t10 a_6774_11720.t1 VDD.t2670 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3715 a_12672_15792.t0 B[0].t23 VSS.t357 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3716 a_19987_11720.t9 opcode[1].t120 VDD.t4362 VDD.t4361 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3717 VDD.t3547 A[3].t57 a_18035_5352.t4 VDD.t3546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3718 VDD.t1475 A[6].t56 a_48265_n1750.t4 VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3719 VDD.t1251 a_52749_18576.t6 a_52809_18602.t4 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3720 a_39618_16432.t1 a_40621_16458.t7 a_41161_15765.t1 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3721 a_40305_20642.t1 a_39715_21079.t9 VDD.t3350 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3722 VDD.t3271 opcode[0].t253 a_7375_8988.t1 VDD.t3270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3723 VDD.t1499 a_30647_12105.t22 a_39720_22683.t4 w_39566_22621# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3724 a_23230_n2148.t5 a_22322_n2148.t6 a_22881_n2148.t10 VDD.t1918 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3725 a_19705_1744.t5 a_19146_1744.t7 a_20054_1744.t4 VDD.t2535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3726 a_52473_15766.t1 a_52710_16433.t15 a_52709_15034.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3727 VDD.t4600 VSS.t719 a_3591_21596.t3 VDD.t4599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3728 a_49477_22063.t1 a_48124_21370.t14 VDD.t4081 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3729 VSS.t361 a_3652_8992.t7 a_5060_10391.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3730 a_48542_1014.t3 a_44399_2324.t17 VDD.t4167 VDD.t4166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3731 VDD.t4199 a_40365_3291.t7 a_41361_3878.t0 VDD.t4198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3732 a_10199_n2174.t0 a_12478_20862.t11 VDD.t2485 VDD.t2484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3733 a_17040_20263.t0 opcode[0].t254 a_15680_20866.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3734 VDD.t4253 a_54454_9678.t8 a_51054_2325.t3 VDD.t4252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3735 a_21211_16387.t1 B[2].t21 VDD.t1359 VDD.t1358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3736 a_41905_21347.t2 A[0].t32 VDD.t2299 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3737 a_38145_1715.t1 a_37848_2326.t16 a_37908_2352.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3738 a_49686_24206.t2 a_46823_22243.t5 a_49568_24206.t2 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3739 a_16322_10994.t0 a_17501_10851.t6 a_17446_10391.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3740 VSS.t421 a_53576_9091.t7 a_54454_9678.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3741 VSS.t143 opcode[2].t59 a_9668_1744.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3742 a_24157_16385.t3 A[0].t33 VDD.t2301 VDD.t2300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3743 a_23777_13581.t1 opcode[0].t255 VDD.t3273 VDD.t3272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3744 a_29954_7911.t11 a_30154_8749.t7 a_30647_7968.t7 VDD.t4295 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3745 a_1039_8966.t5 a_9221_6047.t7 a_9761_5354.t6 VDD.t3235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3746 a_59627_310.t0 a_59921_1016.t7 VSS.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3747 a_7700_n3481.t1 a_7055_n2174.t7 VSS.t339 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3748 a_46350_1040.t0 a_45805_1733.t7 a_46232_1040.t0 VDD.t1981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3749 a_23722_13121.t0 a_23071_14428.t7 VSS.t191 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3750 a_59929_6884.t3 a_55469_11532.t19 VSS.t245 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3751 a_19763_16387.t4 B[3].t36 VDD.t1912 VDD.t1911 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3752 Y[3].t0 a_13810_n2152.t11 VDD.t4186 VDD.t4185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3753 a_30645_3831.t3 a_30152_3173.t7 a_29952_3774.t3 VDD.t1134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3754 a_46140_17941.t4 a_46569_18571.t7 a_46275_18597.t5 w_46046_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3755 a_16855_14458.t9 a_17501_13585.t6 a_16322_13728.t4 VDD.t1991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3756 a_54253_15766.t10 a_53713_16459.t6 a_52710_16433.t6 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3757 a_22172_5352.t0 B[1].t21 VDD.t2475 VDD.t2474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3758 VSS.t99 a_59627_1042.t14 a_60980_1735.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3759 VDD.t868 opcode[2].t60 a_19146_1744.t0 VDD.t867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3760 a_22709_16385.t4 A[1].t42 VDD.t2582 VDD.t2581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3761 VDD.t1890 B[4].t32 a_41676_11949.t2 VDD.t1889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3762 a_61761_310.t1 a_59627_1042.t15 a_61525_1042.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3763 VDD.t3275 opcode[0].t256 a_14357_13585.t1 VDD.t3274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3764 a_48254_6910.t0 a_47709_7603.t7 a_48136_6910.t0 VDD.t2161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3765 VSS.t705 a_54713_3294.t18 a_57981_7583.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3766 a_39715_21079.t3 A[0].t34 VDD.t2302 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3767 a_13178_13728.t1 a_14357_13585.t7 a_14302_13125.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3768 a_7375_8988.t0 opcode[0].t257 VDD.t3277 VDD.t3276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3769 VDD.t3127 a_39807_6822.t15 a_41160_7515.t0 VDD.t3126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3770 VDD.t548 a_37848_2326.t17 a_37908_2352.t4 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3771 a_47837_15029.t1 a_48131_15735.t7 a_46176_16428.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3772 a_70459_8189.t0 opcode[1].t121 VDD.t4364 VDD.t4363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3773 a_19737_n2148.t3 a_19178_n2148.t7 a_20086_n2148.t3 VDD.t2286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3774 a_14014_407.t0 a_13120_11724.t7 VSS.t364 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3775 VDD.t1247 a_48855_n1313.t18 a_51114_2351.t4 VDD.t1246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3776 VDD.t4073 a_67135_3808.t10 a_57676_2326.t0 VDD.t4072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3777 VDD.t606 a_65769_3118.t11 a_70513_7422.t0 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3778 a_10397_15824.t3 a_10337_15751.t8 VDD.t3511 VDD.t3510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3779 a_8011_10847.t0 opcode[1].t122 VDD.t4366 VDD.t4365 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3780 a_41913_24205.t1 a_40305_20642.t6 a_42031_24205.t0 w_41877_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3781 a_9334_20862.t7 a_10513_20719.t5 a_9867_21592.t10 VDD.t2867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3782 VDD.t3780 A[7].t36 a_6735_21596.t9 VDD.t3779 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3783 VDD.t3545 A[3].t58 a_63532_11802.t0 VDD.t3544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3784 a_1745_8119.t0 opcode[0].t258 VDD.t3279 VDD.t3278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3785 a_64192_n2074.t2 a_63602_n1637.t10 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3786 a_7995_15753.t4 A[4].t54 a_8130_16410.t5 VDD.t2025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3787 VDD.t3281 opcode[0].t259 a_20633_13581.t0 VDD.t3280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3788 VDD.t3316 B[6].t38 a_54879_11969.t0 VDD.t3315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3789 a_70509_10624.t4 a_63114_21369.t11 a_70509_10506.t5 VDD.t2683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3790 a_44451_9870.t0 a_42266_11512.t19 VDD.t3594 VDD.t3593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3791 a_6202_20866.t5 A[5].t54 a_6735_21596.t6 VDD.t3433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3792 VSS.t376 a_61782_23618.t7 a_62660_24205.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3793 a_4173_14432.t1 a_15297_16387.t9 VDD.t1365 VDD.t1364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3794 a_1713_n2637.t1 a_1156_1740.t11 VDD.t1579 VDD.t1578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3795 a_40219_3874.t3 a_38484_3565.t7 VDD.t4022 VDD.t4021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3796 VDD.t3600 a_48690_23619.t7 a_49686_24206.t3 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3797 VDD.t2027 A[4].t55 a_63595_1208.t3 VDD.t2026 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3798 a_16605_n2152.t3 opcode[3].t60 VDD.t4276 VDD.t4275 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3799 a_18243_16385.t0 B[4].t33 VDD.t1892 VDD.t1891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3800 a_6774_11720.t2 a_6832_10990.t11 VDD.t2673 VDD.t2672 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3801 VDD.t1688 a_41697_1042.t23 a_46644_1014.t0 VDD.t1687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3802 VDD.t4583 a_54908_6842.t19 a_65651_3118.t6 VDD.t4582 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3803 VSS.t335 a_5108_13805.t7 a_5060_13125.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3804 a_37908_2352.t3 a_37848_2326.t18 VDD.t550 VDD.t549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3805 a_1089_14458.t0 opcode[0].t260 VDD.t2231 VDD.t2230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3806 VDD.t1361 B[2].t22 a_20103_5350.t4 VDD.t1360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3807 a_5070_7659.t0 opcode[0].t261 a_3710_8262.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3808 a_52809_18602.t3 a_52749_18576.t7 VDD.t1252 w_52580_17957# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3809 a_41161_15765.t6 a_41573_15739.t6 a_39618_16432.t6 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3810 a_16322_13728.t7 a_17501_13585.t7 a_17446_13125.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3811 a_16573_1740.t6 opcode[2].t61 VDD.t870 VDD.t869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3812 VDD.t3351 a_39715_21079.t10 a_40305_20642.t0 w_39561_21017# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3813 a_4233_14458.t4 a_4173_14432.t6 a_3700_13728.t5 VDD.t1120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3814 a_70455_11391.t0 opcode[1].t123 VDD.t4368 VDD.t4367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3815 a_22881_n2148.t9 a_22322_n2148.t7 a_23230_n2148.t4 VDD.t1919 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3816 a_41587_6822.t11 a_41160_7515.t7 a_41705_6822.t7 VDD.t3613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3817 a_52473_15034.t1 a_52767_15740.t7 a_52473_15766.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3818 VDD.t1645 B[4].t34 a_35012_10049.t0 VDD.t1644 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3819 VDD.t525 a_41611_21373.t15 a_42964_22066.t2 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3820 VDD.t1000 a_49832_23623.t16 a_56438_21365.t9 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3821 a_16322_10994.t1 a_17501_10851.t7 a_16855_11724.t0 VDD.t394 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3822 VDD.t4082 a_48124_21370.t15 a_49477_22063.t0 w_47542_22001# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3823 VSS.t59 a_30647_7968.t21 a_52990_23688.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3824 VDD.t401 a_16322_10994.t10 a_16264_11724.t1 VDD.t400 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3825 a_39657_18575.t2 a_40724_17941.t6 VDD.t1920 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3826 a_41991_1016.t0 a_37848_2326.t19 VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3827 VDD.t872 opcode[2].t62 a_22849_1744.t0 VDD.t871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3828 VDD.t12 a_7995_15753.t7 a_8056_15820.t2 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3829 VDD.t1363 B[2].t23 a_21211_16387.t0 VDD.t1362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3830 VDD.t4260 a_54713_3294.t19 a_57730_9870.t4 VDD.t4259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3831 VSS.t285 a_70513_19926.t11 a_23723_1259.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3832 VDD.t2866 a_44451_9870.t10 a_45041_9433.t0 VDD.t2865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3833 VDD.t2303 A[0].t35 a_41905_21347.t1 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3834 a_49568_24206.t1 a_46823_22243.t6 a_49686_24206.t0 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3835 VDD.t2987 a_51813_16162.t19 a_51815_16459.t0 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3836 a_17682_10391.t0 opcode[1].t124 a_16322_10994.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3837 a_9168_15798.t3 A[3].t59 a_9304_16408.t0 VDD.t3543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3838 VDD.t2233 opcode[0].t262 a_23777_13581.t0 VDD.t2232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3839 a_4889_8119.t1 opcode[0].t263 VDD.t2235 VDD.t2234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3840 a_48136_6910.t8 a_46356_6910.t15 VDD.t4439 VDD.t4438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3841 VDD.t3063 B[3].t37 a_19763_16387.t5 VDD.t3062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3842 a_22598_13724.t1 a_23777_13581.t7 a_23722_13121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3843 a_41905_21347.t3 A[0].t36 VSS.t366 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3844 a_70513_16782.t3 a_70459_17667.t7 a_70513_16900.t6 VDD.t3371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3845 VSS.t230 A[6].t57 a_5659_15753.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3846 a_52710_16433.t7 a_53713_16459.t7 a_54253_15766.t11 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3847 VSS.t672 opcode[3].t61 a_9700_n2148.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3848 a_4626_16408.t4 A[7].t37 a_4491_15753.t2 VDD.t3781 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3849 a_45821_15761.t4 a_45279_16157.t18 VDD.t3301 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3850 a_37911_6528.t0 a_35602_9612.t19 VDD.t955 VDD.t954 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3851 VDD.t2584 A[1].t43 a_22709_16385.t3 VDD.t2583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3852 a_41676_11949.t1 B[4].t35 VDD.t1647 VDD.t1646 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3853 a_48225_11948.t5 A[5].t55 VDD.t3435 VDD.t3434 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3854 a_17479_n2637.t0 a_16922_1740.t11 VDD.t1555 VDD.t1554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3855 a_14357_13585.t0 opcode[0].t264 VDD.t2237 VDD.t2236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3856 a_9918_14454.t0 a_9976_13724.t11 VDD.t317 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3857 a_20633_10847.t0 opcode[1].t125 VDD.t4370 VDD.t4369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3858 VDD.t2668 a_51690_3564.t7 a_53425_3873.t0 VDD.t2667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3859 a_35602_9612.t3 a_35012_10049.t10 VSS.t681 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3860 VDD.t2994 a_58320_9433.t7 a_60055_9742.t0 VDD.t2993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3861 a_49977_18084.t1 a_30645_n306.t23 VSS.t501 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3862 a_13461_n2152.t3 a_12902_n2152.t6 a_13810_n2152.t2 VDD.t1769 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3863 a_7365_11720.t1 a_6784_8988.t6 VDD.t4486 VDD.t4485 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3864 a_57744_8220.t4 a_57684_8194.t18 VDD.t2348 VDD.t2347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3865 VDD.t2239 opcode[0].t265 a_30150_2544.t0 VDD.t2238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3866 a_40365_3291.t3 a_40101_3874.t8 VSS.t497 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3867 VDD.t2488 a_41705_6822.t19 a_65222_11397.t0 VDD.t2487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3868 a_17190_n3485.t1 a_16545_n2178.t7 VSS.t408 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3869 VDD.t3791 a_23198_1744.t11 a_23755_n2633.t0 VDD.t3790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3870 a_9867_21592.t8 a_10513_20719.t6 a_9334_20862.t4 VDD.t2185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3871 a_52767_22675.t5 a_30647_7968.t22 VDD.t341 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3872 a_64122_11365.t0 a_63532_11802.t10 VDD.t2116 VDD.t2115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3873 a_60766_15769.t3 a_61178_15743.t7 a_59223_16436.t3 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3874 a_8130_16410.t4 A[4].t56 a_7995_15753.t1 VDD.t2028 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3875 a_55469_11532.t1 a_54879_11969.t9 VDD.t3160 VDD.t3159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3876 VDD.t2241 opcode[0].t266 a_4889_8119.t0 VDD.t2240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3877 a_58326_16165.t3 a_62660_24205.t6 VSS.t261 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3878 VDD.t1371 a_19763_16387.t9 a_13651_14432.t1 VDD.t1370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3879 VDD.t2292 a_30645_10037.t22 a_46219_24330.t5 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3880 VDD.t1367 a_15297_16387.t10 a_4173_14432.t0 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3881 a_30643_n2374.t3 a_30150_n3032.t7 a_29950_n2431.t8 VDD.t4118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3882 VDD.t1001 a_49832_23623.t17 a_52762_21071.t1 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3883 VDD.t1488 a_51054_2325.t18 a_55197_1015.t0 VDD.t1487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3884 a_66063_6587.t0 a_64117_5761.t15 VDD.t1155 VDD.t1154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3885 VDD.t2030 A[4].t57 a_18243_16385.t3 VDD.t2029 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3886 VDD.t4169 a_44399_2324.t18 a_44454_746.t0 VDD.t4168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3887 VDD.t2350 a_57684_8194.t19 a_61827_6884.t0 VDD.t2349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3888 a_63408_21343.t3 a_56366_23618.t19 VSS.t208 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3889 a_556_13728.t5 a_1735_13585.t6 a_1089_14458.t7 VDD.t2527 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3890 VDD.t453 a_65767_10704.t11 a_70509_13768.t5 VDD.t452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3891 a_55504_n1325.t0 a_54914_n1762.t10 VDD.t3006 VDD.t3005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3892 a_7668_411.t0 a_6774_11720.t7 VSS.t327 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3893 a_54658_21365.t7 a_54952_21339.t7 a_54540_21365.t11 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3894 VSS.t12 a_55224_23614.t7 a_56102_24201.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3895 a_39618_16432.t5 a_41573_15739.t7 a_41161_15765.t11 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3896 VDD.t3437 A[5].t56 a_16795_16385.t5 VDD.t3436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3897 a_17682_13125.t1 opcode[0].t267 a_16322_13728.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3898 VDD.t4264 a_53005_1041.t15 a_54358_1734.t0 VDD.t4263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3899 a_3700_13728.t6 a_4173_14432.t7 a_4233_14458.t5 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3900 VDD.t4278 opcode[3].t62 a_22881_n2148.t6 VDD.t4277 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3901 VDD.t173 a_41507_3295.t18 a_46238_6910.t9 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3902 VSS.t436 a_59901_23892.t7 a_61518_24201.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3903 a_43410_14834.t0 a_38721_16161.t18 VSS.t247 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3904 VDD.t894 a_59635_6910.t15 a_60988_7603.t0 VDD.t893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3905 a_35012_10049.t1 B[4].t36 VDD.t1649 VDD.t1648 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3906 a_8021_8115.t0 opcode[0].t268 VDD.t2243 VDD.t2242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3907 VSS.t92 a_61525_1042.t11 a_71846_5105.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3908 VDD.t2507 a_55862_18700.t10 a_53891_18572.t0 w_55768_18664# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3909 VDD.t4208 a_22550_8988.t6 a_23131_11720.t4 VDD.t4207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3910 VSS.t110 a_54903_1041.t22 a_59863_310.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3911 VDD.t3230 a_62660_24205.t7 a_58326_16165.t1 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3912 a_16264_11724.t0 a_16322_10994.t11 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3913 VDD.t917 a_48254_6910.t22 a_51105_9802.t0 VDD.t916 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3914 VDD.t1028 a_40724_17941.t7 a_39657_18575.t1 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3915 a_8056_15820.t3 a_7995_15753.t8 VDD.t2181 VDD.t2180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3916 VDD.t4171 a_44399_2324.t19 a_48130_1040.t5 VDD.t4170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3917 a_61189_3878.t2 a_58326_1915.t6 a_61071_3878.t1 VDD.t3076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3918 VSS.t45 a_44405_8194.t19 a_48490_6178.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3919 a_43173_24209.t2 a_40310_22246.t7 a_43055_24209.t3 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3920 a_41905_21347.t0 A[0].t37 VDD.t2304 w_41029_22004# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3921 a_49686_24206.t1 a_46823_22243.t7 a_49568_24206.t0 w_49532_24144# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3922 VSS.t103 a_25100_20862.t11 a_22821_n2174.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3923 VSS.t587 a_16274_8992.t6 a_17682_10391.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3924 a_19997_8988.t0 opcode[0].t269 VDD.t2245 VDD.t2244 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3925 a_31375_n2374.t1 a_30150_n1593.t7 a_30643_n2374.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3926 Y[4].t3 a_10608_n2148.t11 VSS.t144 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3927 a_13711_11724.t3 a_13130_8992.t7 VDD.t1094 VDD.t1093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3928 a_19763_16387.t6 B[3].t38 VDD.t3065 VDD.t3064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3929 VDD.t1657 a_38721_16161.t19 a_38723_16458.t0 w_38687_16396# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3930 VDD.t2681 a_13188_8262.t11 a_13130_8992.t3 VDD.t2680 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3931 a_51695_9365.t3 a_51105_9802.t10 VSS.t210 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3932 a_41587_6822.t0 a_37856_8106.t19 VDD.t1664 VDD.t1663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3933 a_56556_21365.t5 a_56850_21339.t7 a_56438_21365.t6 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3934 a_54253_15766.t4 a_54665_15740.t7 a_52710_16433.t0 w_51779_16397# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3935 a_71846_20635.t0 a_43509_21373.t11 VSS.t433 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3936 a_37894_4002.t2 a_35575_3749.t18 VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3937 a_4491_15753.t1 A[7].t38 a_4626_16408.t3 VDD.t3782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3938 VDD.t3302 a_45279_16157.t19 a_45821_15761.t3 w_45245_16392# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3939 VDD.t3439 A[5].t57 a_48225_11948.t4 VDD.t3438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3940 a_51100_4001.t4 a_48855_n1313.t19 VDD.t1249 VDD.t1248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3941 VDD.t1477 A[6].t58 a_41676_11949.t4 VDD.t1476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3942 VDD.t2031 A[4].t58 a_60226_16462.t0 w_58292_16400# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3943 VSS.t268 B[4].t37 a_35249_9412.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3944 a_10259_n2148.t2 a_10199_n2174.t7 VDD.t1593 VDD.t1592 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3945 a_39799_1042.t5 a_39254_1735.t7 a_39681_1042.t11 VDD.t2836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3946 VDD.t2477 B[1].t22 a_21632_6045.t0 VDD.t2476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3947 VSS.t235 a_51054_2325.t19 a_55139_309.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3948 VDD.t3042 a_70509_n2116.t11 a_1681_1255.t0 VDD.t3041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3949 a_50316_21344.t3 a_43319_23626.t19 VSS.t450 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3950 a_52749_18576.t0 a_53816_17942.t8 VDD.t2742 w_53722_17953# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3951 a_13810_n2152.t1 a_12902_n2152.t7 a_13461_n2152.t4 VDD.t1770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3952 VSS.t269 B[4].t38 a_35222_3549.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3953 VDD.t4488 a_6784_8988.t7 a_7365_11720.t0 VDD.t4487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3954 a_59921_1016.t3 a_54903_1041.t23 VSS.t111 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3955 a_23135_20719.t3 opcode[0].t270 VSS.t358 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3956 a_9334_20862.t5 a_10513_20719.t7 a_9867_21592.t9 VDD.t2186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3957 a_52892_6842.t6 a_53304_6816.t7 a_53010_6842.t3 VDD.t2669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3958 VDD.t342 a_30647_7968.t23 a_52767_22675.t4 w_52613_22613# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3959 VDD.t2288 a_54879_11969.t10 a_55469_11532.t0 VDD.t2287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3960 a_7966_7655.t1 a_7315_8962.t11 VSS.t524 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3961 VDD.t186 a_35575_3749.t19 a_37903_748.t4 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3962 a_7995_15753.t3 A[4].t59 a_8130_16410.t3 VDD.t2032 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3963 VSS.t551 A[5].t58 a_55151_n1325.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3964 a_51346_110.t1 a_48064_9163.t19 a_51109_747.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3965 a_70509_1146.t3 a_61533_6910.t11 VDD.t556 VDD.t555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3966 a_13651_14432.t0 a_19763_16387.t10 VDD.t1369 VDD.t1368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3967 a_51699_310.t3 a_51109_747.t10 VSS.t540 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3968 a_39706_24333.t4 a_30647_12105.t23 VDD.t1500 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3969 a_46219_24330.t4 a_30645_10037.t23 VDD.t2293 w_46065_24268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3970 VDD.t2247 opcode[0].t271 a_13721_8992.t1 VDD.t2246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3971 a_15297_16387.t0 B[6].t39 VDD.t3318 VDD.t3317 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3972 a_29954_12048.t6 a_30154_12886.t7 a_30647_12105.t3 VDD.t201 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3973 a_54572_9678.t4 a_51709_7715.t7 a_54454_9678.t1 VDD.t2792 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3974 a_52762_21071.t2 a_49832_23623.t18 VDD.t1002 w_52608_21009# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3975 VSS.t194 a_22598_10990.t11 a_22540_11720.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3976 a_16855_11724.t9 a_16274_8992.t7 VDD.t3688 VDD.t3687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3977 a_556_10994.t2 a_1735_10851.t7 a_1680_10391.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3978 Y[5].t0 a_7464_n2148.t11 VDD.t3182 VDD.t3181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3979 a_59929_3874.t1 a_58321_311.t7 a_60047_3874.t0 VDD.t1483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3980 a_13849_16387.t0 B[7].t22 VDD.t2622 VDD.t2621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3981 a_16855_11724.t3 a_16264_14458.t7 a_16322_10994.t5 VDD.t507 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3982 a_1089_14458.t6 a_1735_13585.t7 a_556_13728.t4 VDD.t2528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3983 a_63532_11802.t6 B[3].t39 VDD.t3067 VDD.t3066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3984 VDD.t3784 A[7].t39 a_1974_8339.t0 VDD.t3783 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3985 a_11829_5352.t11 a_12241_5326.t7 a_4183_8966.t7 VDD.t2259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3986 VDD.t1713 a_57676_2326.t18 a_57731_748.t0 VDD.t1712 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3987 a_51119_8152.t4 a_48254_6910.t23 VDD.t919 VDD.t918 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3988 a_61071_3878.t0 a_58326_1915.t7 VSS.t494 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3989 VDD.t965 a_45041_9433.t7 a_46776_9742.t2 VDD.t964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3990 a_9221_6047.t0 B[7].t23 VDD.t2624 VDD.t2623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3991 a_46592_6178.t1 a_41507_3295.t19 a_46356_6910.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3992 a_41913_24205.t0 a_40305_20642.t7 VSS.t67 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3993 a_16795_16385.t4 A[5].t59 VDD.t3441 VDD.t3440 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3994 VSS.t79 a_10397_15824.t7 a_17682_13125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3995 a_1099_8992.t2 a_1039_8966.t11 a_566_8262.t2 VDD.t500 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3996 a_1188_n2152.t3 a_1713_n2637.t7 a_839_n2152.t6 VDD.t2359 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3997 a_22881_n2148.t5 opcode[3].t63 VDD.t4280 VDD.t4279 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X3998 VDD.t3694 a_57676_2326.t19 a_57736_2352.t1 VDD.t3693 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3999 VDD.t2306 A[0].t38 a_24240_5350.t6 VDD.t2305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4000 a_61782_23618.t3 a_61518_24201.t8 VSS.t157 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4001 VDD.t1003 a_49832_23623.t19 a_56850_21339.t0 w_54076_21996# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4002 a_30152_9379.t0 B[1].t23 VDD.t2479 VDD.t2478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4003 VDD.t1651 B[4].t39 a_35012_10049.t2 VDD.t1650 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4004 a_23131_11720.t3 a_22550_8988.t7 VDD.t4210 VDD.t4209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4005 a_20633_10847.t3 opcode[1].t126 VSS.t684 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4006 a_6842_8258.t0 a_8021_8115.t7 a_7966_7655.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4007 a_58326_16165.t0 a_62660_24205.t8 VDD.t3231 w_62624_24143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4008 a_39657_18575.t0 a_40724_17941.t8 VDD.t1029 w_40630_17952# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4009 a_70459_17667.t3 opcode[1].t127 VSS.t685 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4010 a_40043_6090.t1 a_35594_7027.t19 a_39807_6822.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4011 a_39706_24333.t2 A[0].t39 VDD.t2307 w_39552_24271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4012 VSS.t624 a_60226_16462.t7 a_60884_15037.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4013 VSS.t231 A[6].t59 a_35238_789.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4014 a_20054_1744.t0 opcode[2].t63 a_20290_411.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4015 VDD.t3692 a_42177_23622.t7 a_43173_24209.t3 w_43019_24147# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
R0 a_48690_23619.t4 a_48690_23619.t5 800.071
R1 a_48690_23619.n3 a_48690_23619.n2 672.951
R2 a_48690_23619.n1 a_48690_23619.t7 285.109
R3 a_48690_23619.n2 a_48690_23619.t4 193.602
R4 a_48690_23619.n1 a_48690_23619.t6 160.666
R5 a_48690_23619.n2 a_48690_23619.n1 91.507
R6 a_48690_23619.n0 a_48690_23619.t1 28.57
R7 a_48690_23619.n4 a_48690_23619.t2 28.565
R8 a_48690_23619.t0 a_48690_23619.n4 28.565
R9 a_48690_23619.n0 a_48690_23619.t3 17.638
R10 a_48690_23619.n4 a_48690_23619.n3 0.69
R11 a_48690_23619.n3 a_48690_23619.n0 0.6
R12 a_49686_24206.n0 a_49686_24206.t5 14.282
R13 a_49686_24206.n0 a_49686_24206.t1 14.282
R14 a_49686_24206.n1 a_49686_24206.t3 14.282
R15 a_49686_24206.n1 a_49686_24206.t4 14.282
R16 a_49686_24206.t0 a_49686_24206.n3 14.282
R17 a_49686_24206.n3 a_49686_24206.t2 14.282
R18 a_49686_24206.n3 a_49686_24206.n2 2.546
R19 a_49686_24206.n2 a_49686_24206.n1 2.367
R20 a_49686_24206.n2 a_49686_24206.n0 0.001
R21 VDD.t4601 VDD.t596 95474.9
R22 VDD.t2000 VDD.t1263 95474.9
R23 VDD.t3282 VDD.t2480 95474.9
R24 VDD.t898 VDD.t2145 95474.9
R25 VDD.t1921 VDD.t2153 95474.9
R26 VDD.t3964 VDD.t675 95474.9
R27 VDD.t3432 VDD.t78 95474.9
R28 VDD.t3015 VDD.t946 95474.9
R29 VDD.t631 VDD.t2756 95474.9
R30 VDD.t663 VDD.t1899 95474.9
R31 VDD.t1113 VDD.t2893 95474.9
R32 VDD.t2683 VDD.t2341 95474.9
R33 VDD.t576 VDD.t3041 95474.9
R34 VDD.t121 VDD.t1037 95474.9
R35 VDD.t1270 VDD.t3323 95474.9
R36 VDD.t2695 VDD.t1760 95474.9
R37 VDD.t3289 VDD.t2802 95474.9
R38 VDD.t1977 VDD.t3570 95474.9
R39 VDD.t293 VDD.t2843 95474.9
R40 VDD.t2129 VDD.t351 95474.9
R41 VDD.t1334 VDD.t1720 95474.9
R42 VDD.t4235 VDD.t2680 95474.9
R43 VDD.t4515 VDD.t1280 95474.9
R44 VDD.t499 VDD.t2343 95474.9
R45 VDD.t1571 VDD.t3328 95474.9
R46 VDD.t2819 VDD.t2761 95474.9
R47 VDD.t4584 VDD.t1158 95474.9
R48 VDD.t2430 VDD.t4221 95474.9
R49 VDD.t507 VDD.t398 95474.9
R50 VDD.t3928 VDD.t482 95474.9
R51 VDD.t143 VDD.t2692 95474.9
R52 VDD.t26 VDD.t1594 95474.9
R53 VDD.t1986 VDD.t2312 95474.9
R54 VDD.t3785 VDD.t518 95474.9
R55 VDD.t1582 VDD.t4243 95474.9
R56 VDD.t1120 VDD.t374 95474.9
R57 VDD.t195 VDD.t637 95474.9
R58 VDD.t404 VDD.t312 95474.9
R59 VDD.t386 VDD.t3935 95474.9
R60 VDD.t1136 VDD.t2489 95474.9
R61 VDD.t4482 VDD.t4211 95474.9
R62 VDD.t2358 VDD.t1536 95474.9
R63 VDD.t2739 VDD.t1301 95474.9
R64 VDD.t4249 VDD.t4181 95474.9
R65 VDD.t4240 VDD.t1970 95474.9
R66 VDD.t632 VDD.t1 95474.9
R67 VDD.t115 VDD.t874 95474.9
R68 VDD.t3153 VDD.t3181 95474.9
R69 VDD.t3101 VDD.t2544 95474.9
R70 VDD.t558 VDD.t1578 95474.9
R71 VDD.t3403 VDD.t2130 95474.9
R72 VDD.t2687 VDD.t1853 95474.9
R73 VDD.t222 VDD.t1554 95474.9
R74 VDD.t4597 VDD.t3043 95474.9
R75 VDD.t790 VDD.t2554 95474.9
R76 VDD.t2900 VDD.t2688 95474.9
R77 VDD.t4348 VDD.t4338 2079.61
R78 VDD.t3794 VDD.t512 2079.61
R79 VDD.t2272 VDD.t1620 2079.61
R80 VDD.t2542 VDD.t1558 2079.61
R81 VDD.t617 VDD.t623 2079.61
R82 VDD.t782 VDD.t778 2079.61
R83 VDD.t1679 VDD.t1671 2079.61
R84 VDD.t2707 VDD.t181 2079.61
R85 VDD.n2745 VDD.n2744 1412.62
R86 VDD.n3193 VDD.n3192 1412.62
R87 VDD.n456 VDD.n455 1412.59
R88 VDD.n368 VDD.n356 1408.41
R89 VDD.n3075 VDD.n3074 1404.25
R90 VDD.n524 VDD.n523 1239.11
R91 VDD.n3005 VDD.n3004 1235.85
R92 VDD.n2808 VDD.n2807 1235.85
R93 VDD.n2779 VDD.n2778 1033.17
R94 VDD.n2985 VDD.n2979 1033.13
R95 VDD.n3137 VDD.n3131 1033.13
R96 VDD.n3161 VDD.n3160 1033.13
R97 VDD.n334 VDD.n333 1033.13
R98 VDD.n3113 VDD.n3107 1033.12
R99 VDD.n489 VDD.n488 1029.24
R100 VDD.n2970 VDD.n2966 1029.22
R101 VDD.n2719 VDD.n2718 1029.21
R102 VDD.n2832 VDD.n2831 1029.21
R103 VDD.n428 VDD.n427 1025.33
R104 VDD.n321 VDD.n317 1025.3
R105 VDD.t3122 VDD.t948 999.845
R106 VDD.t4436 VDD.t508 999.845
R107 VDD.t1530 VDD.t2264 999.845
R108 VDD.t893 VDD.t957 999.845
R109 VDD.t569 VDD.t621 999.845
R110 VDD.t4263 VDD.t776 999.845
R111 VDD.t4426 VDD.t1683 999.845
R112 VDD.t3662 VDD.t2709 999.845
R113 VDD.n2787 VDD.n2781 880.922
R114 VDD.n2712 VDD.n2711 874.899
R115 VDD.n3148 VDD.n3142 874.857
R116 VDD.n3046 VDD.n3042 874.804
R117 VDD.n542 VDD.n541 871.829
R118 VDD.n2896 VDD.n2890 871.811
R119 VDD.n436 VDD.n430 871.81
R120 VDD.n501 VDD.n496 871.809
R121 VDD.n3248 VDD.n3247 871.808
R122 VDD.n2862 VDD.n2861 871.808
R123 VDD.n3226 VDD.n3225 871.808
R124 VDD.n3055 VDD.n3054 871.808
R125 VDD.n2853 VDD.n2852 809.201
R126 VDD.n3215 VDD.n3214 805.926
R127 VDD.n3239 VDD.n3238 805.926
R128 VDD.n3102 VDD.n3101 805.925
R129 VDD.n556 VDD.n555 802.65
R130 VDD.n2822 VDD.n2821 687.118
R131 VDD.n2884 VDD.n2882 687.068
R132 VDD.n3127 VDD.n3125 684.693
R133 VDD.n600 VDD.n599 600.209
R134 VDD.n730 VDD.n729 600.209
R135 VDD.n586 VDD.n585 600.207
R136 VDD.n264 VDD.n263 600.207
R137 VDD.n1199 VDD.n1198 565.289
R138 VDD.n1169 VDD.n1168 563.326
R139 VDD.n1184 VDD.n1183 561.363
R140 VDD.n1214 VDD.n1213 559.4
R141 VDD.n1127 VDD.n1126 557.438
R142 VDD.n1142 VDD.n1141 553.512
R143 VDD.t433 VDD.t429 541.402
R144 VDD.t4142 VDD.t2458 541.402
R145 VDD.t2196 VDD.t2220 541.402
R146 VDD.t1546 VDD.t2611 541.402
R147 VDD.t3313 VDD.t1387 541.402
R148 VDD.t1815 VDD.t1823 541.402
R149 VDD.t1871 VDD.t1879 541.402
R150 VDD.t2659 VDD.t2653 541.402
R151 VDD.n2918 VDD.n2917 491.958
R152 VDD.n3120 VDD.t4194 479.007
R153 VDD.n3199 VDD.t970 479.007
R154 VDD.n2873 VDD.t3368 479.006
R155 VDD.n3232 VDD.t2139 479.006
R156 VDD.n2846 VDD.t2883 479.006
R157 VDD.n534 VDD.t3641 479.006
R158 VDD.n1250 VDD.t3062 473.001
R159 VDD.n1246 VDD.t1544 473.001
R160 VDD.n1248 VDD.t1831 473.001
R161 VDD.n1249 VDD.t1887 473.001
R162 VDD.n1252 VDD.t2454 473.001
R163 VDD.n371 VDD.t2536 424.731
R164 VDD.t2176 VDD.t1661 422.41
R165 VDD.t250 VDD.t244 422.41
R166 VDD.t1068 VDD.t4284 422.41
R167 VDD.t2815 VDD.t2809 422.41
R168 VDD.t1640 VDD.t1706 422.41
R169 VDD.t85 VDD.t91 422.41
R170 VDD.t4170 VDD.t2063 422.41
R171 VDD.t1945 VDD.t551 422.41
R172 VDD.n563 VDD.t31 422.371
R173 VDD.t1395 VDD.t3309 413.681
R174 VDD.t3726 VDD.t431 413.681
R175 VDD.t2204 VDD.t2212 413.681
R176 VDD.t2474 VDD.t2472 413.681
R177 VDD.t2651 VDD.t2418 413.681
R178 VDD.t920 VDD.t940 413.681
R179 VDD.t2410 VDD.t4114 413.681
R180 VDD.t1548 VDD.t2607 413.681
R181 VDD.t3508 VDD.t3510 406.159
R182 VDD.t641 VDD.t643 406.159
R183 VDD.n1140 VDD.t3506 402.717
R184 VDD.n1125 VDD.t639 402.717
R185 VDD.t11 VDD.t2180 397.517
R186 VDD.t4203 VDD.t4296 397.517
R187 VDD.t302 VDD.t304 396.113
R188 VDD.t3382 VDD.t3378 396.113
R189 VDD.t4231 VDD.t2875 394.32
R190 VDD.t4566 VDD.t4578 394.32
R191 VDD.t1148 VDD.t1138 394.32
R192 VDD.t4495 VDD.t4501 394.32
R193 VDD.n1167 VDD.t9 394.148
R194 VDD.n1212 VDD.t4298 394.148
R195 VDD.n1197 VDD.t300 392.756
R196 VDD.n1182 VDD.t3380 392.756
R197 VDD.t3395 VDD.t3202 382.217
R198 VDD.t3028 VDD.t1805 382.217
R199 VDD.t3463 VDD.t3677 382.217
R200 VDD.t3993 VDD.t3198 382.217
R201 VDD.t4406 VDD.t3945 382.217
R202 VDD.t286 VDD.t3999 382.217
R203 VDD.t3779 VDD.t4534 382.217
R204 VDD.t4599 VDD.t1010 382.217
R205 VDD.t3857 VDD.t795 382.217
R206 VDD.t1609 VDD.t1186 382.217
R207 VDD.t2699 VDD.t723 382.217
R208 VDD.t3861 VDD.t727 382.217
R209 VDD.t560 VDD.t821 382.217
R210 VDD.t452 VDD.t683 382.217
R211 VDD.t2784 VDD.t801 382.217
R212 VDD.t2847 VDD.t809 382.217
R213 VDD.t2109 VDD.t2242 382.217
R214 VDD.t1097 VDD.t3867 382.217
R215 VDD.t2731 VDD.t1352 382.217
R216 VDD.t4593 VDD.t3689 382.217
R217 VDD.t1694 VDD.t1521 382.217
R218 VDD.t4449 VDD.t4001 382.217
R219 VDD.t48 VDD.t2234 382.217
R220 VDD.t1718 VDD.t3278 382.217
R221 VDD.t4487 VDD.t4365 382.217
R222 VDD.t1295 VDD.t4357 382.217
R223 VDD.t4205 VDD.t1206 382.217
R224 VDD.t37 VDD.t1202 382.217
R225 VDD.t3683 VDD.t815 382.217
R226 VDD.t1089 VDD.t715 382.217
R227 VDD.t2255 VDD.t831 382.217
R228 VDD.t2499 VDD.t827 382.217
R229 VDD.t444 VDD.t1788 382.217
R230 VDD.t3421 VDD.t3840 382.217
R231 VDD.t382 VDD.t3834 382.217
R232 VDD.t2101 VDD.t1481 382.217
R233 VDD.t3374 VDD.t1004 382.217
R234 VDD.t3333 VDD.t3829 382.217
R235 VDD.t2750 VDD.t3266 382.217
R236 VDD.t4478 VDD.t3272 382.217
R237 VDD.t3319 VDD.t4324 382.217
R238 VDD.t2722 VDD.t4314 382.217
R239 VDD.t296 VDD.t3905 382.217
R240 VDD.t132 VDD.t4322 382.217
R241 VDD.t3526 VDD.t3895 382.217
R242 VDD.t2824 VDD.t3885 382.217
R243 VDD.t1592 VDD.t3077 382.217
R244 VDD.t2771 VDD.t4271 382.217
R245 VDD.t3166 VDD.t2921 382.217
R246 VDD.t586 VDD.t2925 382.217
R247 VDD.t1050 VDD.t2913 382.217
R248 VDD.t2280 VDD.t2933 382.217
R249 VDD.t463 VDD.t2935 382.217
R250 VDD.t1268 VDD.t867 382.217
R251 VDD.t318 VDD.t845 382.217
R252 VDD.t2057 VDD.t2927 382.217
R253 VDD.t4379 VDD.t4402 359.294
R254 VDD.t1324 VDD.t4379 359.294
R255 VDD.t3064 VDD.t1324 359.294
R256 VDD.t3062 VDD.t3064 359.294
R257 VDD.t3062 VDD.t1911 359.294
R258 VDD.t1911 VDD.t1372 359.294
R259 VDD.t1372 VDD.t1368 359.294
R260 VDD.t1368 VDD.t1370 359.294
R261 VDD.t3750 VDD.t3752 359.294
R262 VDD.t3747 VDD.t3750 359.294
R263 VDD.t2597 VDD.t3747 359.294
R264 VDD.t1544 VDD.t2597 359.294
R265 VDD.t1544 VDD.t2621 359.294
R266 VDD.t2621 VDD.t3671 359.294
R267 VDD.t3671 VDD.t3675 359.294
R268 VDD.t3675 VDD.t3673 359.294
R269 VDD.t3440 VDD.t2080 359.294
R270 VDD.t3436 VDD.t3440 359.294
R271 VDD.t1835 VDD.t3436 359.294
R272 VDD.t1831 VDD.t1835 359.294
R273 VDD.t1831 VDD.t1827 359.294
R274 VDD.t1827 VDD.t3953 359.294
R275 VDD.t3953 VDD.t3955 359.294
R276 VDD.t3955 VDD.t3951 359.294
R277 VDD.t269 VDD.t276 359.294
R278 VDD.t2029 VDD.t269 359.294
R279 VDD.t1891 VDD.t2029 359.294
R280 VDD.t1887 VDD.t1891 359.294
R281 VDD.t1887 VDD.t1867 359.294
R282 VDD.t1867 VDD.t4304 359.294
R283 VDD.t4304 VDD.t4302 359.294
R284 VDD.t4302 VDD.t4300 359.294
R285 VDD.t2581 VDD.t2583 359.294
R286 VDD.t2579 VDD.t2581 359.294
R287 VDD.t2462 VDD.t2579 359.294
R288 VDD.t2454 VDD.t2462 359.294
R289 VDD.t2454 VDD.t4144 359.294
R290 VDD.t4144 VDD.t2447 359.294
R291 VDD.t2447 VDD.t2445 359.294
R292 VDD.t2445 VDD.t2443 359.294
R293 VDD.t4227 VDD.t2873 352.102
R294 VDD.t4568 VDD.t4576 352.102
R295 VDD.t1144 VDD.t1154 352.102
R296 VDD.t2564 VDD.t2558 352.102
R297 VDD.t596 VDD.t594 345.987
R298 VDD.t594 VDD.t592 345.987
R299 VDD.t3214 VDD.t2370 345.987
R300 VDD.t3202 VDD.t3214 345.987
R301 VDD.t1263 VDD.t1261 345.987
R302 VDD.t1261 VDD.t1259 345.987
R303 VDD.t3920 VDD.t2048 345.987
R304 VDD.t1805 VDD.t3920 345.987
R305 VDD.t2480 VDD.t2484 345.987
R306 VDD.t2484 VDD.t2482 345.987
R307 VDD.t3179 VDD.t4052 345.987
R308 VDD.t3677 VDD.t3179 345.987
R309 VDD.t2145 VDD.t2143 345.987
R310 VDD.t2143 VDD.t2147 345.987
R311 VDD.t3206 VDD.t3831 345.987
R312 VDD.t3198 VDD.t3206 345.987
R313 VDD.t2153 VDD.t2157 345.987
R314 VDD.t2157 VDD.t2155 345.987
R315 VDD.t2038 VDD.t3262 345.987
R316 VDD.t3945 VDD.t2038 345.987
R317 VDD.t675 VDD.t673 345.987
R318 VDD.t673 VDD.t671 345.987
R319 VDD.t3204 VDD.t3216 345.987
R320 VDD.t3999 VDD.t3204 345.987
R321 VDD.t78 VDD.t3657 345.987
R322 VDD.t3657 VDD.t3655 345.987
R323 VDD.t1598 VDD.t3937 345.987
R324 VDD.t4534 VDD.t1598 345.987
R325 VDD.t946 VDD.t944 345.987
R326 VDD.t944 VDD.t942 345.987
R327 VDD.t2878 VDD.t1783 345.987
R328 VDD.t1010 VDD.t2878 345.987
R329 VDD.t3343 VDD.t3341 345.987
R330 VDD.t3339 VDD.t3343 345.987
R331 VDD.t3712 VDD.t3339 345.987
R332 VDD.t3722 VDD.t3712 345.987
R333 VDD.t3710 VDD.t952 345.987
R334 VDD.t952 VDD.t4336 345.987
R335 VDD.t4336 VDD.t4344 345.987
R336 VDD.t4552 VDD.t4556 345.987
R337 VDD.t4554 VDD.t4552 345.987
R338 VDD.t208 VDD.t4554 345.987
R339 VDD.t3558 VDD.t208 345.987
R340 VDD.t204 VDD.t177 345.987
R341 VDD.t177 VDD.t2713 345.987
R342 VDD.t2713 VDD.t183 345.987
R343 VDD.t2851 VDD.t2853 345.987
R344 VDD.t2855 VDD.t2851 345.987
R345 VDD.t4102 VDD.t2855 345.987
R346 VDD.t4088 VDD.t4102 345.987
R347 VDD.t4094 VDD.t1667 345.987
R348 VDD.t1667 VDD.t1675 345.987
R349 VDD.t1675 VDD.t1665 345.987
R350 VDD.t2191 VDD.t2189 345.987
R351 VDD.t2187 VDD.t2191 345.987
R352 VDD.t1242 VDD.t2187 345.987
R353 VDD.t1248 VDD.t1242 345.987
R354 VDD.t1238 VDD.t647 345.987
R355 VDD.t647 VDD.t770 345.987
R356 VDD.t770 VDD.t645 345.987
R357 VDD.t1425 VDD.t1427 345.987
R358 VDD.t1429 VDD.t1425 345.987
R359 VDD.t4463 VDD.t1429 345.987
R360 VDD.t488 VDD.t4463 345.987
R361 VDD.t1312 VDD.t1018 345.987
R362 VDD.t1018 VDD.t625 345.987
R363 VDD.t625 VDD.t1016 345.987
R364 VDD.t2353 VDD.t2355 345.987
R365 VDD.t2351 VDD.t2353 345.987
R366 VDD.t2023 VDD.t2351 345.987
R367 VDD.t2019 VDD.t2023 345.987
R368 VDD.t2017 VDD.t1843 345.987
R369 VDD.t1843 VDD.t1837 345.987
R370 VDD.t1837 VDD.t1813 345.987
R371 VDD.t541 VDD.t545 345.987
R372 VDD.t543 VDD.t541 345.987
R373 VDD.t4259 VDD.t543 345.987
R374 VDD.t4518 VDD.t4259 345.987
R375 VDD.t4524 VDD.t1560 345.987
R376 VDD.t1560 VDD.t3495 345.987
R377 VDD.t3495 VDD.t3410 345.987
R378 VDD.t1342 VDD.t1346 345.987
R379 VDD.t1344 VDD.t1342 345.987
R380 VDD.t2166 VDD.t1344 345.987
R381 VDD.t906 VDD.t2166 345.987
R382 VDD.t916 VDD.t2274 345.987
R383 VDD.t2274 VDD.t1618 345.987
R384 VDD.t1618 VDD.t2266 345.987
R385 VDD.t2865 VDD.t2822 345.987
R386 VDD.t2820 VDD.t2865 345.987
R387 VDD.t168 VDD.t2820 345.987
R388 VDD.t152 VDD.t168 345.987
R389 VDD.t162 VDD.t3589 345.987
R390 VDD.t3589 VDD.t510 345.987
R391 VDD.t510 VDD.t3593 345.987
R392 VDD.t3126 VDD.t3226 345.987
R393 VDD.t3226 VDD.t3122 345.987
R394 VDD.t948 VDD.t4334 345.987
R395 VDD.t4334 VDD.t4348 345.987
R396 VDD.t2174 VDD.t2249 345.987
R397 VDD.t1661 VDD.t2174 345.987
R398 VDD.t2901 VDD.t2905 345.987
R399 VDD.t2903 VDD.t2901 345.987
R400 VDD.t3716 VDD.t2903 345.987
R401 VDD.t3700 VDD.t3716 345.987
R402 VDD.t3714 VDD.t60 345.987
R403 VDD.t60 VDD.t58 345.987
R404 VDD.t58 VDD.t2172 345.987
R405 VDD.t2107 VDD.t2164 345.987
R406 VDD.t2162 VDD.t2107 345.987
R407 VDD.t56 VDD.t2162 345.987
R408 VDD.t2170 VDD.t56 345.987
R409 VDD.t2178 VDD.t4342 345.987
R410 VDD.t4342 VDD.t4340 345.987
R411 VDD.t4340 VDD.t954 345.987
R412 VDD.t2644 VDD.t2646 345.987
R413 VDD.t2646 VDD.t4436 345.987
R414 VDD.t508 VDD.t3798 345.987
R415 VDD.t3798 VDD.t3794 345.987
R416 VDD.t230 VDD.t246 345.987
R417 VDD.t244 VDD.t230 345.987
R418 VDD.t2830 VDD.t2834 345.987
R419 VDD.t2832 VDD.t2830 345.987
R420 VDD.t170 VDD.t2832 345.987
R421 VDD.t154 VDD.t170 345.987
R422 VDD.t164 VDD.t236 345.987
R423 VDD.t236 VDD.t242 345.987
R424 VDD.t242 VDD.t252 345.987
R425 VDD.t1255 VDD.t1253 345.987
R426 VDD.t1257 VDD.t1255 345.987
R427 VDD.t238 VDD.t1257 345.987
R428 VDD.t248 VDD.t238 345.987
R429 VDD.t232 VDD.t3796 345.987
R430 VDD.t3796 VDD.t3587 345.987
R431 VDD.t3587 VDD.t3792 345.987
R432 VDD.t1534 VDD.t2595 345.987
R433 VDD.t2595 VDD.t1530 345.987
R434 VDD.t2264 VDD.t2262 345.987
R435 VDD.t2262 VDD.t2272 345.987
R436 VDD.t1074 VDD.t4286 345.987
R437 VDD.t4284 VDD.t1074 345.987
R438 VDD.t1289 VDD.t1287 345.987
R439 VDD.t1285 VDD.t1289 345.987
R440 VDD.t908 VDD.t1285 345.987
R441 VDD.t918 VDD.t908 345.987
R442 VDD.t904 VDD.t1080 345.987
R443 VDD.t1080 VDD.t1066 345.987
R444 VDD.t1066 VDD.t1072 345.987
R445 VDD.t4546 VDD.t3501 345.987
R446 VDD.t4548 VDD.t4546 345.987
R447 VDD.t1078 VDD.t4548 345.987
R448 VDD.t4290 VDD.t1078 345.987
R449 VDD.t1070 VDD.t2270 345.987
R450 VDD.t2270 VDD.t2276 345.987
R451 VDD.t2276 VDD.t2260 345.987
R452 VDD.t829 VDD.t1178 345.987
R453 VDD.t795 VDD.t829 345.987
R454 VDD.t2756 VDD.t2754 345.987
R455 VDD.t2754 VDD.t2752 345.987
R456 VDD.t805 VDD.t681 345.987
R457 VDD.t1186 VDD.t805 345.987
R458 VDD.t1899 VDD.t1903 345.987
R459 VDD.t1903 VDD.t1901 345.987
R460 VDD.t1166 VDD.t4363 345.987
R461 VDD.t723 VDD.t1166 345.987
R462 VDD.t2893 VDD.t2891 345.987
R463 VDD.t2891 VDD.t2889 345.987
R464 VDD.t1168 VDD.t4367 345.987
R465 VDD.t727 VDD.t1168 345.987
R466 VDD.t2341 VDD.t2337 345.987
R467 VDD.t2337 VDD.t2339 345.987
R468 VDD.t1218 VDD.t803 345.987
R469 VDD.t821 VDD.t1218 345.987
R470 VDD.t3041 VDD.t3037 345.987
R471 VDD.t3037 VDD.t3039 345.987
R472 VDD.t1172 VDD.t1204 345.987
R473 VDD.t683 VDD.t1172 345.987
R474 VDD.t1037 VDD.t1035 345.987
R475 VDD.t1035 VDD.t1039 345.987
R476 VDD.t741 VDD.t1188 345.987
R477 VDD.t801 VDD.t741 345.987
R478 VDD.t3323 VDD.t3321 345.987
R479 VDD.t3321 VDD.t3325 345.987
R480 VDD.t743 VDD.t4359 345.987
R481 VDD.t809 VDD.t743 345.987
R482 VDD.t1760 VDD.t1764 345.987
R483 VDD.t1764 VDD.t1762 345.987
R484 VDD.t885 VDD.t889 345.987
R485 VDD.t889 VDD.t893 345.987
R486 VDD.t957 VDD.t650 345.987
R487 VDD.t650 VDD.t2542 345.987
R488 VDD.t2349 VDD.t2813 345.987
R489 VDD.t2809 VDD.t2349 345.987
R490 VDD.t2360 VDD.t3154 345.987
R491 VDD.t3156 VDD.t2360 345.987
R492 VDD.t2396 VDD.t3156 345.987
R493 VDD.t4520 VDD.t2396 345.987
R494 VDD.t4526 VDD.t2347 345.987
R495 VDD.t2347 VDD.t3585 345.987
R496 VDD.t3585 VDD.t2345 345.987
R497 VDD.t67 VDD.t65 345.987
R498 VDD.t69 VDD.t67 345.987
R499 VDD.t3583 VDD.t69 345.987
R500 VDD.t2817 VDD.t3583 345.987
R501 VDD.t3581 VDD.t3497 345.987
R502 VDD.t3497 VDD.t1556 345.987
R503 VDD.t1556 VDD.t3499 345.987
R504 VDD.t573 VDD.t565 345.987
R505 VDD.t565 VDD.t569 345.987
R506 VDD.t621 VDD.t627 345.987
R507 VDD.t627 VDD.t617 345.987
R508 VDD.t1700 VDD.t1638 345.987
R509 VDD.t1706 VDD.t1700 345.987
R510 VDD.t3072 VDD.t3070 345.987
R511 VDD.t3068 VDD.t3072 345.987
R512 VDD.t486 VDD.t3068 345.987
R513 VDD.t494 VDD.t486 345.987
R514 VDD.t484 VDD.t1698 345.987
R515 VDD.t1698 VDD.t3693 345.987
R516 VDD.t3693 VDD.t1642 345.987
R517 VDD.t2684 VDD.t1062 345.987
R518 VDD.t1064 VDD.t2684 345.987
R519 VDD.t1704 VDD.t1064 345.987
R520 VDD.t1710 VDD.t1704 345.987
R521 VDD.t1712 VDD.t615 345.987
R522 VDD.t615 VDD.t1022 345.987
R523 VDD.t1022 VDD.t619 345.987
R524 VDD.t4261 VDD.t4265 345.987
R525 VDD.t4265 VDD.t4263 345.987
R526 VDD.t776 VDD.t774 345.987
R527 VDD.t774 VDD.t782 345.987
R528 VDD.t1487 VDD.t99 345.987
R529 VDD.t91 VDD.t1487 345.987
R530 VDD.t3577 VDD.t1046 345.987
R531 VDD.t1044 VDD.t3577 345.987
R532 VDD.t1246 VDD.t1044 345.987
R533 VDD.t1230 VDD.t1246 345.987
R534 VDD.t1240 VDD.t97 345.987
R535 VDD.t97 VDD.t1485 345.987
R536 VDD.t1485 VDD.t87 345.987
R537 VDD.t3358 VDD.t3356 345.987
R538 VDD.t3360 VDD.t3358 345.987
R539 VDD.t83 VDD.t3360 345.987
R540 VDD.t89 VDD.t83 345.987
R541 VDD.t93 VDD.t975 345.987
R542 VDD.t975 VDD.t772 345.987
R543 VDD.t772 VDD.t780 345.987
R544 VDD.t4430 VDD.t4434 345.987
R545 VDD.t4434 VDD.t4426 345.987
R546 VDD.t1683 VDD.t1687 345.987
R547 VDD.t1687 VDD.t1679 345.987
R548 VDD.t4160 VDD.t4166 345.987
R549 VDD.t2063 VDD.t4160 345.987
R550 VDD.t3530 VDD.t3528 345.987
R551 VDD.t3142 VDD.t3530 345.987
R552 VDD.t4086 VDD.t3142 345.987
R553 VDD.t4100 VDD.t4086 345.987
R554 VDD.t4084 VDD.t4158 345.987
R555 VDD.t4158 VDD.t4162 345.987
R556 VDD.t4162 VDD.t4152 345.987
R557 VDD.t1586 VDD.t1584 345.987
R558 VDD.t3331 VDD.t1586 345.987
R559 VDD.t4168 VDD.t3331 345.987
R560 VDD.t2065 VDD.t4168 345.987
R561 VDD.t4154 VDD.t1673 345.987
R562 VDD.t1673 VDD.t1681 345.987
R563 VDD.t1681 VDD.t1677 345.987
R564 VDD.t3666 VDD.t1751 345.987
R565 VDD.t1751 VDD.t3662 345.987
R566 VDD.t2709 VDD.t2701 345.987
R567 VDD.t2701 VDD.t2707 345.987
R568 VDD.t1943 VDD.t1935 345.987
R569 VDD.t551 VDD.t1943 345.987
R570 VDD.t1636 VDD.t1634 345.987
R571 VDD.t1632 VDD.t1636 345.987
R572 VDD.t218 VDD.t1632 345.987
R573 VDD.t202 VDD.t218 345.987
R574 VDD.t216 VDD.t549 345.987
R575 VDD.t549 VDD.t547 345.987
R576 VDD.t547 VDD.t1939 345.987
R577 VDD.t389 VDD.t1118 345.987
R578 VDD.t391 VDD.t389 345.987
R579 VDD.t1941 VDD.t391 345.987
R580 VDD.t1949 VDD.t1941 345.987
R581 VDD.t1947 VDD.t2711 345.987
R582 VDD.t2711 VDD.t185 345.987
R583 VDD.t185 VDD.t2703 345.987
R584 VDD.t3210 VDD.t4058 345.987
R585 VDD.t2040 VDD.t3210 345.987
R586 VDD.t429 VDD.t3730 345.987
R587 VDD.t3730 VDD.t1356 345.987
R588 VDD.t3218 VDD.t3918 345.987
R589 VDD.t4054 VDD.t3218 345.987
R590 VDD.t2458 VDD.t2478 345.987
R591 VDD.t2478 VDD.t2464 345.987
R592 VDD.t1030 VDD.t3910 345.987
R593 VDD.t1511 VDD.t1030 345.987
R594 VDD.t2220 VDD.t2206 345.987
R595 VDD.t2206 VDD.t2228 345.987
R596 VDD.t3309 VDD.t1385 345.987
R597 VDD.t1385 VDD.t1405 345.987
R598 VDD.t1436 VDD.t1466 345.987
R599 VDD.t1462 VDD.t1436 345.987
R600 VDD.t431 VDD.t1354 345.987
R601 VDD.t1354 VDD.t3736 345.987
R602 VDD.t3983 VDD.t4030 345.987
R603 VDD.t3981 VDD.t3983 345.987
R604 VDD.t2212 VDD.t2218 345.987
R605 VDD.t2218 VDD.t2194 345.987
R606 VDD.t2321 VDD.t2334 345.987
R607 VDD.t2329 VDD.t2321 345.987
R608 VDD.t2472 VDD.t4140 345.987
R609 VDD.t4140 VDD.t2476 345.987
R610 VDD.t193 VDD.t3397 345.987
R611 VDD.t1932 VDD.t193 345.987
R612 VDD.t2418 VDD.t1905 345.987
R613 VDD.t1905 VDD.t2657 345.987
R614 VDD.t4371 VDD.t4414 345.987
R615 VDD.t4388 VDD.t4371 345.987
R616 VDD.t940 VDD.t1875 345.987
R617 VDD.t1875 VDD.t932 345.987
R618 VDD.t272 VDD.t278 345.987
R619 VDD.t2003 VDD.t272 345.987
R620 VDD.t4114 VDD.t1821 345.987
R621 VDD.t1821 VDD.t2416 345.987
R622 VDD.t3425 VDD.t3443 345.987
R623 VDD.t2076 VDD.t3425 345.987
R624 VDD.t2607 VDD.t2623 345.987
R625 VDD.t2623 VDD.t2603 345.987
R626 VDD.t3775 VDD.t3759 345.987
R627 VDD.t3755 VDD.t3775 345.987
R628 VDD.t2802 VDD.t2804 345.987
R629 VDD.t2804 VDD.t1503 345.987
R630 VDD.t3914 VDD.t3809 345.987
R631 VDD.t2242 VDD.t3914 345.987
R632 VDD.t3570 VDD.t3572 345.987
R633 VDD.t3572 VDD.t3568 345.987
R634 VDD.t4049 VDD.t1603 345.987
R635 VDD.t3867 VDD.t4049 345.987
R636 VDD.t2843 VDD.t2767 345.987
R637 VDD.t2767 VDD.t2769 345.987
R638 VDD.t1517 VDD.t1519 345.987
R639 VDD.t1352 VDD.t1517 345.987
R640 VDD.t351 VDD.t347 345.987
R641 VDD.t347 VDD.t349 345.987
R642 VDD.t1509 VDD.t2374 345.987
R643 VDD.t3689 VDD.t1509 345.987
R644 VDD.t1720 VDD.t1722 345.987
R645 VDD.t1722 VDD.t3873 345.987
R646 VDD.t3939 VDD.t3200 345.987
R647 VDD.t1521 VDD.t3939 345.987
R648 VDD.t2680 VDD.t2676 345.987
R649 VDD.t2676 VDD.t2678 345.987
R650 VDD.t2376 VDD.t1809 345.987
R651 VDD.t4001 VDD.t2376 345.987
R652 VDD.t1280 VDD.t2540 345.987
R653 VDD.t2540 VDD.t1278 345.987
R654 VDD.t2240 VDD.t1785 345.987
R655 VDD.t2234 VDD.t2240 345.987
R656 VDD.t2343 VDD.t1563 345.987
R657 VDD.t1563 VDD.t1565 345.987
R658 VDD.t4035 VDD.t3997 345.987
R659 VDD.t3278 VDD.t4035 345.987
R660 VDD.t3328 VDD.t2672 345.987
R661 VDD.t2672 VDD.t2670 345.987
R662 VDD.t697 VDD.t703 345.987
R663 VDD.t4365 VDD.t697 345.987
R664 VDD.t2761 VDD.t2765 345.987
R665 VDD.t2765 VDD.t2763 345.987
R666 VDD.t685 VDD.t693 345.987
R667 VDD.t4357 VDD.t685 345.987
R668 VDD.t1158 VDD.t1156 345.987
R669 VDD.t1156 VDD.t530 345.987
R670 VDD.t1216 VDD.t1184 345.987
R671 VDD.t1206 VDD.t1216 345.987
R672 VDD.t4221 VDD.t4492 345.987
R673 VDD.t4492 VDD.t4490 345.987
R674 VDD.t1212 VDD.t4369 345.987
R675 VDD.t1202 VDD.t1212 345.987
R676 VDD.t398 VDD.t402 345.987
R677 VDD.t402 VDD.t400 345.987
R678 VDD.t717 VDD.t721 345.987
R679 VDD.t815 VDD.t717 345.987
R680 VDD.t482 VDD.t480 345.987
R681 VDD.t480 VDD.t478 345.987
R682 VDD.t1210 VDD.t1220 345.987
R683 VDD.t715 VDD.t1210 345.987
R684 VDD.t2692 VDD.t2690 345.987
R685 VDD.t2690 VDD.t1086 345.987
R686 VDD.t797 VDD.t813 345.987
R687 VDD.t831 VDD.t797 345.987
R688 VDD.t1594 VDD.t3555 345.987
R689 VDD.t3555 VDD.t3553 345.987
R690 VDD.t835 VDD.t733 345.987
R691 VDD.t827 VDD.t835 345.987
R692 VDD.t2312 VDD.t2310 345.987
R693 VDD.t2310 VDD.t2308 345.987
R694 VDD.t4033 VDD.t1781 345.987
R695 VDD.t1788 VDD.t4033 345.987
R696 VDD.t518 VDD.t456 345.987
R697 VDD.t456 VDD.t454 345.987
R698 VDD.t3274 VDD.t2236 345.987
R699 VDD.t3840 VDD.t3274 345.987
R700 VDD.t4243 VDD.t2729 345.987
R701 VDD.t2729 VDD.t1282 345.987
R702 VDD.t4062 VDD.t2050 345.987
R703 VDD.t3834 VDD.t4062 345.987
R704 VDD.t374 VDD.t372 345.987
R705 VDD.t372 VDD.t370 345.987
R706 VDD.t1743 VDD.t3827 345.987
R707 VDD.t1481 VDD.t1743 345.987
R708 VDD.t637 VDD.t635 345.987
R709 VDD.t635 VDD.t633 345.987
R710 VDD.t3836 VDD.t1775 345.987
R711 VDD.t1004 VDD.t3836 345.987
R712 VDD.t312 VDD.t316 345.987
R713 VDD.t316 VDD.t314 345.987
R714 VDD.t4037 VDD.t4045 345.987
R715 VDD.t3829 VDD.t4037 345.987
R716 VDD.t3935 VDD.t3933 345.987
R717 VDD.t3933 VDD.t3931 345.987
R718 VDD.t3280 VDD.t1779 345.987
R719 VDD.t3266 VDD.t3280 345.987
R720 VDD.t2489 VDD.t2493 345.987
R721 VDD.t2493 VDD.t2491 345.987
R722 VDD.t2232 VDD.t2389 345.987
R723 VDD.t3272 VDD.t2232 345.987
R724 VDD.t1596 VDD.t3190 345.987
R725 VDD.t4009 VDD.t1596 345.987
R726 VDD.t2611 VDD.t2619 345.987
R727 VDD.t2619 VDD.t2601 345.987
R728 VDD.t1528 VDD.t3493 345.987
R729 VDD.t3818 VDD.t1528 345.987
R730 VDD.t1387 VDD.t1417 345.987
R731 VDD.t1417 VDD.t3303 345.987
R732 VDD.t2238 VDD.t1745 345.987
R733 VDD.t3208 VDD.t2238 345.987
R734 VDD.t1823 VDD.t1817 345.987
R735 VDD.t1817 VDD.t4108 345.987
R736 VDD.t3924 VDD.t2042 345.987
R737 VDD.t103 VDD.t3924 345.987
R738 VDD.t1879 VDD.t938 345.987
R739 VDD.t938 VDD.t930 345.987
R740 VDD.t4047 VDD.t2380 345.987
R741 VDD.t1796 VDD.t4047 345.987
R742 VDD.t2653 VDD.t4127 345.987
R743 VDD.t4127 VDD.t2439 345.987
R744 VDD.t4324 VDD.t3887 345.987
R745 VDD.t3887 VDD.t4269 345.987
R746 VDD.t4213 VDD.t4215 345.987
R747 VDD.t4211 VDD.t4213 345.987
R748 VDD.t4314 VDD.t4310 345.987
R749 VDD.t4310 VDD.t4308 345.987
R750 VDD.t1538 VDD.t1540 345.987
R751 VDD.t1536 VDD.t1538 345.987
R752 VDD.t3905 VDD.t4550 345.987
R753 VDD.t4550 VDD.t3085 345.987
R754 VDD.t1297 VDD.t1299 345.987
R755 VDD.t1301 VDD.t1297 345.987
R756 VDD.t4322 VDD.t4320 345.987
R757 VDD.t4320 VDD.t3903 345.987
R758 VDD.t4183 VDD.t4185 345.987
R759 VDD.t4181 VDD.t4183 345.987
R760 VDD.t3895 VDD.t3891 345.987
R761 VDD.t3891 VDD.t3889 345.987
R762 VDD.t1972 VDD.t1974 345.987
R763 VDD.t1970 VDD.t1972 345.987
R764 VDD.t3885 VDD.t3881 345.987
R765 VDD.t3881 VDD.t3879 345.987
R766 VDD.t4217 VDD.t4219 345.987
R767 VDD.t1 VDD.t4217 345.987
R768 VDD.t3077 VDD.t4330 345.987
R769 VDD.t4330 VDD.t4326 345.987
R770 VDD.t747 VDD.t745 345.987
R771 VDD.t874 VDD.t747 345.987
R772 VDD.t4271 VDD.t4267 345.987
R773 VDD.t4267 VDD.t3097 345.987
R774 VDD.t1006 VDD.t1008 345.987
R775 VDD.t3181 VDD.t1006 345.987
R776 VDD.t2921 VDD.t2957 345.987
R777 VDD.t2957 VDD.t849 345.987
R778 VDD.t3790 VDD.t3788 345.987
R779 VDD.t2544 VDD.t3790 345.987
R780 VDD.t2925 VDD.t2961 345.987
R781 VDD.t2961 VDD.t851 345.987
R782 VDD.t1576 VDD.t2125 345.987
R783 VDD.t1578 VDD.t1576 345.987
R784 VDD.t2913 VDD.t2949 345.987
R785 VDD.t2949 VDD.t865 345.987
R786 VDD.t2134 VDD.t2132 345.987
R787 VDD.t2130 VDD.t2134 345.987
R788 VDD.t2933 VDD.t2969 345.987
R789 VDD.t2969 VDD.t2967 345.987
R790 VDD.t1116 VDD.t1855 345.987
R791 VDD.t1853 VDD.t1116 345.987
R792 VDD.t2935 VDD.t2919 345.987
R793 VDD.t2919 VDD.t2955 345.987
R794 VDD.t105 VDD.t107 345.987
R795 VDD.t1554 VDD.t105 345.987
R796 VDD.t867 VDD.t2939 345.987
R797 VDD.t2939 VDD.t2971 345.987
R798 VDD.t3047 VDD.t3045 345.987
R799 VDD.t3043 VDD.t3047 345.987
R800 VDD.t845 VDD.t2915 345.987
R801 VDD.t2915 VDD.t2953 345.987
R802 VDD.t3533 VDD.t2552 345.987
R803 VDD.t2554 VDD.t3533 345.987
R804 VDD.t2927 VDD.t853 345.987
R805 VDD.t853 VDD.t2951 345.987
R806 VDD.t3052 VDD.t3054 345.987
R807 VDD.t2688 VDD.t3052 345.987
R808 VDD.n2917 VDD.t2017 343.055
R809 VDD.t3611 VDD.t3126 312.28
R810 VDD.t2161 VDD.t2644 312.28
R811 VDD.t458 VDD.t1534 312.28
R812 VDD.t1859 VDD.t885 312.28
R813 VDD.t2840 VDD.t573 312.28
R814 VDD.t1341 VDD.t4261 312.28
R815 VDD.t3405 VDD.t4430 312.28
R816 VDD.t2149 VDD.t3666 312.28
R817 VDD.t4295 VDD.t2040 312.28
R818 VDD.t3833 VDD.t4054 312.28
R819 VDD.t200 VDD.t1511 312.28
R820 VDD.t2259 VDD.t1462 312.28
R821 VDD.t1043 VDD.t3981 312.28
R822 VDD.t1421 VDD.t2329 312.28
R823 VDD.t3175 VDD.t1932 312.28
R824 VDD.t1625 VDD.t4388 312.28
R825 VDD.t2861 VDD.t2003 312.28
R826 VDD.t3059 VDD.t2076 312.28
R827 VDD.t51 VDD.t3755 312.28
R828 VDD.t1749 VDD.t4009 312.28
R829 VDD.t533 VDD.t3818 312.28
R830 VDD.t138 VDD.t3208 312.28
R831 VDD.t1432 VDD.t103 312.28
R832 VDD.t2641 VDD.t1796 312.28
R833 VDD.t1523 VDD.t4603 276.597
R834 VDD.t1801 VDD.t2009 276.597
R835 VDD.t1339 VDD.t4385 276.597
R836 VDD.t3811 VDD.t2315 276.597
R837 VDD.t1767 VDD.t3400 276.597
R838 VDD.t3212 VDD.t3987 276.597
R839 VDD.t3337 VDD.t2086 276.597
R840 VDD.t1737 VDD.t1448 276.597
R841 VDD.t711 VDD.t630 276.597
R842 VDD.t833 VDD.t662 276.597
R843 VDD.t1194 VDD.t1115 276.597
R844 VDD.t725 VDD.t2682 276.597
R845 VDD.t1174 VDD.t577 276.597
R846 VDD.t731 VDD.t120 276.597
R847 VDD.t799 VDD.t134 276.597
R848 VDD.t713 VDD.t2696 276.597
R849 VDD.t1724 VDD.t3290 276.597
R850 VDD.t3807 VDD.t1978 276.597
R851 VDD.t3875 VDD.t292 276.597
R852 VDD.t3254 VDD.t2127 276.597
R853 VDD.t3805 VDD.t1336 276.597
R854 VDD.t3814 VDD.t4236 276.597
R855 VDD.t1337 VDD.t4514 276.597
R856 VDD.t3220 VDD.t500 276.597
R857 VDD.t701 VDD.t2870 276.597
R858 VDD.t689 VDD.t369 276.597
R859 VDD.t1180 VDD.t4586 276.597
R860 VDD.t4361 VDD.t2432 276.597
R861 VDD.t707 VDD.t505 276.597
R862 VDD.t1176 VDD.t3930 276.597
R863 VDD.t807 VDD.t142 276.597
R864 VDD.t729 VDD.t504 276.597
R865 VDD.t1726 VDD.t1987 276.597
R866 VDD.t2372 VDD.t3787 276.597
R867 VDD.t2044 VDD.t2486 276.597
R868 VDD.t3846 VDD.t1012 276.597
R869 VDD.t3851 VDD.t197 276.597
R870 VDD.t4003 VDD.t406 276.597
R871 VDD.t3823 VDD.t385 276.597
R872 VDD.t2382 VDD.t1135 276.597
R873 VDD.t3899 VDD.t4480 276.597
R874 VDD.t4316 VDD.t2359 276.597
R875 VDD.t3095 VDD.t2737 276.597
R876 VDD.t4328 VDD.t4247 276.597
R877 VDD.t4306 VDD.t4241 276.597
R878 VDD.t3079 VDD.t590 276.597
R879 VDD.t3089 VDD.t116 276.597
R880 VDD.t3099 VDD.t3151 276.597
R881 VDD.t871 VDD.t4420 276.597
R882 VDD.t839 VDD.t557 276.597
R883 VDD.t857 VDD.t3402 276.597
R884 VDD.t2923 VDD.t2686 276.597
R885 VDD.t841 VDD.t3575 276.597
R886 VDD.t843 VDD.t4598 276.597
R887 VDD.t847 VDD.t789 276.597
R888 VDD.t863 VDD.t2899 276.597
R889 VDD.t2184 VDD.t1926 269.594
R890 VDD.t2186 VDD.t3007 269.594
R891 VDD.t2035 VDD.t3459 269.594
R892 VDD.t2808 VDD.t3970 269.594
R893 VDD.t355 VDD.t1316 269.594
R894 VDD.t1964 VDD.t280 269.594
R895 VDD.t4150 VDD.t3767 269.594
R896 VDD.t4193 VDD.t4606 269.594
R897 VDD.t1622 VDD.t553 269.594
R898 VDD.t1959 VDD.t1605 269.594
R899 VDD.t3242 VDD.t605 269.594
R900 VDD.t2839 VDD.t3863 269.594
R901 VDD.t4131 VDD.t3522 269.594
R902 VDD.t1659 VDD.t448 269.594
R903 VDD.t3505 VDD.t2786 269.594
R904 VDD.t956 VDD.t2849 269.594
R905 VDD.t3056 VDD.t1614 269.594
R906 VDD.t2052 VDD.t1095 269.594
R907 VDD.t598 VDD.t4066 269.594
R908 VDD.t583 VDD.t4591 269.594
R909 VDD.t4292 VDD.t1692 269.594
R910 VDD.t3471 VDD.t4451 269.594
R911 VDD.t3648 VDD.t46 269.594
R912 VDD.t1774 VDD.t1716 269.594
R913 VDD.t2449 VDD.t4483 269.594
R914 VDD.t4076 VDD.t1291 269.594
R915 VDD.t1766 VDD.t4207 269.594
R916 VDD.t129 VDD.t33 269.594
R917 VDD.t394 VDD.t3685 269.594
R918 VDD.t2674 VDD.t1091 269.594
R919 VDD.t55 VDD.t1101 269.594
R920 VDD.t3165 VDD.t2501 269.594
R921 VDD.t1989 VDD.t446 269.594
R922 VDD.t2744 VDD.t3423 269.594
R923 VDD.t2526 VDD.t378 269.594
R924 VDD.t141 VDD.t2103 269.594
R925 VDD.t1328 VDD.t3376 269.594
R926 VDD.t3564 VDD.t3335 269.594
R927 VDD.t1957 VDD.t2746 269.594
R928 VDD.t260 VDD.t4474 269.594
R929 VDD.t1917 VDD.t2909 269.594
R930 VDD.t73 VDD.t2726 269.594
R931 VDD.t575 VDD.t298 269.594
R932 VDD.t1769 VDD.t130 269.594
R933 VDD.t3645 VDD.t2531 269.594
R934 VDD.t2284 VDD.t2828 269.594
R935 VDD.t3574 VDD.t1590 269.594
R936 VDD.t4178 VDD.t2117 269.594
R937 VDD.t3114 VDD.t3170 269.594
R938 VDD.t82 VDD.t588 269.594
R939 VDD.t2290 VDD.t1048 269.594
R940 VDD.t25 VDD.t2282 269.594
R941 VDD.t3520 VDD.t465 269.594
R942 VDD.t2534 VDD.t3345 269.594
R943 VDD.t562 VDD.t320 269.594
R944 VDD.t3604 VDD.t2059 269.594
R945 VDD.n1050 VDD.n1047 258.915
R946 VDD.n925 VDD.n922 258.915
R947 VDD.n950 VDD.n947 258.915
R948 VDD.n1025 VDD.n1022 258.915
R949 VDD.n1000 VDD.n997 258.915
R950 VDD.n975 VDD.n972 258.915
R951 VDD.n900 VDD.n897 258.915
R952 VDD.n876 VDD.n873 258.915
R953 VDD.n634 VDD.n632 258.915
R954 VDD.n652 VDD.n650 258.915
R955 VDD.n670 VDD.n668 258.915
R956 VDD.n687 VDD.n685 258.915
R957 VDD.n616 VDD.n614 258.915
R958 VDD.n747 VDD.n745 258.915
R959 VDD.n765 VDD.n763 258.915
R960 VDD.n783 VDD.n781 258.915
R961 VDD.n1739 VDD.n1737 258.915
R962 VDD.n1764 VDD.n1762 258.915
R963 VDD.n1869 VDD.n1867 258.915
R964 VDD.n1844 VDD.n1842 258.915
R965 VDD.n1814 VDD.n1812 258.915
R966 VDD.n1789 VDD.n1787 258.915
R967 VDD.n1714 VDD.n1712 258.915
R968 VDD.n1690 VDD.n1688 258.915
R969 VDD.n1544 VDD.n1542 258.915
R970 VDD.n1569 VDD.n1567 258.915
R971 VDD.n1669 VDD.n1667 258.915
R972 VDD.n1644 VDD.n1642 258.915
R973 VDD.n1619 VDD.n1617 258.915
R974 VDD.n1594 VDD.n1592 258.915
R975 VDD.n1519 VDD.n1517 258.915
R976 VDD.n1495 VDD.n1493 258.915
R977 VDD.n1394 VDD.n1392 258.915
R978 VDD.n1369 VDD.n1367 258.915
R979 VDD.n1270 VDD.n1268 258.915
R980 VDD.n1294 VDD.n1292 258.915
R981 VDD.n1319 VDD.n1317 258.915
R982 VDD.n1344 VDD.n1342 258.915
R983 VDD.n1419 VDD.n1417 258.915
R984 VDD.n1444 VDD.n1442 258.915
R985 VDD.n2600 VDD.n2598 258.915
R986 VDD.n2461 VDD.n2459 258.915
R987 VDD.n2480 VDD.n2478 258.915
R988 VDD.n2540 VDD.n2538 258.915
R989 VDD.n2560 VDD.n2558 258.915
R990 VDD.n2580 VDD.n2578 258.915
R991 VDD.n2520 VDD.n2518 258.915
R992 VDD.n2500 VDD.n2498 258.915
R993 VDD.n2396 VDD.n2394 258.915
R994 VDD.n2252 VDD.n2250 258.915
R995 VDD.n2271 VDD.n2269 258.915
R996 VDD.n2336 VDD.n2334 258.915
R997 VDD.n2356 VDD.n2354 258.915
R998 VDD.n2376 VDD.n2374 258.915
R999 VDD.n2311 VDD.n2309 258.915
R1000 VDD.n2291 VDD.n2289 258.915
R1001 VDD.n1041 VDD.n1040 258.161
R1002 VDD.n916 VDD.n915 258.161
R1003 VDD.n941 VDD.n940 258.161
R1004 VDD.n1016 VDD.n1015 258.161
R1005 VDD.n991 VDD.n990 258.161
R1006 VDD.n966 VDD.n965 258.161
R1007 VDD.n891 VDD.n890 258.161
R1008 VDD.n867 VDD.n866 258.161
R1009 VDD.n637 VDD.n636 258.161
R1010 VDD.n655 VDD.n654 258.161
R1011 VDD.n673 VDD.n672 258.161
R1012 VDD.n690 VDD.n689 258.161
R1013 VDD.n619 VDD.n618 258.161
R1014 VDD.n750 VDD.n749 258.161
R1015 VDD.n768 VDD.n767 258.161
R1016 VDD.n786 VDD.n785 258.161
R1017 VDD.n1742 VDD.n1741 258.161
R1018 VDD.n1767 VDD.n1766 258.161
R1019 VDD.n1860 VDD.n1859 258.161
R1020 VDD.n1835 VDD.n1834 258.161
R1021 VDD.n1817 VDD.n1816 258.161
R1022 VDD.n1792 VDD.n1791 258.161
R1023 VDD.n1717 VDD.n1716 258.161
R1024 VDD.n1693 VDD.n1692 258.161
R1025 VDD.n1535 VDD.n1534 258.161
R1026 VDD.n1560 VDD.n1559 258.161
R1027 VDD.n1660 VDD.n1659 258.161
R1028 VDD.n1635 VDD.n1634 258.161
R1029 VDD.n1610 VDD.n1609 258.161
R1030 VDD.n1585 VDD.n1584 258.161
R1031 VDD.n1510 VDD.n1509 258.161
R1032 VDD.n1486 VDD.n1485 258.161
R1033 VDD.n1385 VDD.n1384 258.161
R1034 VDD.n1360 VDD.n1359 258.161
R1035 VDD.n1261 VDD.n1260 258.161
R1036 VDD.n1285 VDD.n1284 258.161
R1037 VDD.n1310 VDD.n1309 258.161
R1038 VDD.n1335 VDD.n1334 258.161
R1039 VDD.n1410 VDD.n1409 258.161
R1040 VDD.n1435 VDD.n1434 258.161
R1041 VDD.n2603 VDD.n2602 258.161
R1042 VDD.n2464 VDD.n2463 258.161
R1043 VDD.n2483 VDD.n2482 258.161
R1044 VDD.n2543 VDD.n2542 258.161
R1045 VDD.n2563 VDD.n2562 258.161
R1046 VDD.n2583 VDD.n2582 258.161
R1047 VDD.n2523 VDD.n2522 258.161
R1048 VDD.n2503 VDD.n2502 258.161
R1049 VDD.n2387 VDD.n2386 258.161
R1050 VDD.n2255 VDD.n2254 258.161
R1051 VDD.n2274 VDD.n2273 258.161
R1052 VDD.n2327 VDD.n2326 258.161
R1053 VDD.n2347 VDD.n2346 258.161
R1054 VDD.n2367 VDD.n2366 258.161
R1055 VDD.n2314 VDD.n2313 258.161
R1056 VDD.n2294 VDD.n2293 258.161
R1057 VDD.n3247 VDD.t3710 240.432
R1058 VDD.n2890 VDD.t204 240.432
R1059 VDD.n2861 VDD.t4094 240.432
R1060 VDD.n2831 VDD.t1238 240.432
R1061 VDD.n541 VDD.t1312 240.432
R1062 VDD.n3107 VDD.t4524 240.432
R1063 VDD.n3131 VDD.t916 240.432
R1064 VDD.n3225 VDD.t162 240.432
R1065 VDD.n2979 VDD.t3714 240.432
R1066 VDD.n2966 VDD.t2178 240.432
R1067 VDD.n3160 VDD.t164 240.432
R1068 VDD.n3142 VDD.t232 240.432
R1069 VDD.n3054 VDD.t904 240.432
R1070 VDD.n3042 VDD.t1070 240.432
R1071 VDD.n333 VDD.t4526 240.432
R1072 VDD.n317 VDD.t3581 240.432
R1073 VDD.n430 VDD.t484 240.432
R1074 VDD.n427 VDD.t1712 240.432
R1075 VDD.n496 VDD.t1240 240.432
R1076 VDD.n488 VDD.t93 240.432
R1077 VDD.n2781 VDD.t4084 240.432
R1078 VDD.n2778 VDD.t4154 240.432
R1079 VDD.n2718 VDD.t216 240.432
R1080 VDD.n2711 VDD.t1947 240.432
R1081 VDD.t3223 VDD.t3708 218.264
R1082 VDD.t1860 VDD.t166 218.264
R1083 VDD.t4423 VDD.t902 218.264
R1084 VDD.t4151 VDD.t4530 218.264
R1085 VDD.t2498 VDD.t4469 218.264
R1086 VDD.t2136 VDD.t1244 218.264
R1087 VDD.t1981 VDD.t4092 218.264
R1088 VDD.t1969 VDD.t214 218.264
R1089 VDD.t4021 VDD.t4017 213.931
R1090 VDD.t4017 VDD.t753 213.931
R1091 VDD.t753 VDD.t751 213.931
R1092 VDD.t751 VDD.t752 213.931
R1093 VDD.t3 VDD.t5 213.931
R1094 VDD.t5 VDD.t667 213.931
R1095 VDD.t667 VDD.t665 213.931
R1096 VDD.t665 VDD.t666 213.931
R1097 VDD.t2631 VDD.t2633 213.931
R1098 VDD.t2633 VDD.t2495 213.931
R1099 VDD.t2495 VDD.t2496 213.931
R1100 VDD.t2496 VDD.t1484 213.931
R1101 VDD.t2775 VDD.t2777 213.931
R1102 VDD.t2777 VDD.t4245 213.931
R1103 VDD.t4245 VDD.t4246 213.931
R1104 VDD.t4246 VDD.t2728 213.931
R1105 VDD.t2663 VDD.t2665 213.931
R1106 VDD.t2665 VDD.t118 213.931
R1107 VDD.t118 VDD.t119 213.931
R1108 VDD.t119 VDD.t117 213.931
R1109 VDD.t2859 VDD.t2857 213.931
R1110 VDD.t2857 VDD.t3597 213.931
R1111 VDD.t3597 VDD.t3644 213.931
R1112 VDD.t3644 VDD.t3596 213.931
R1113 VDD.t3477 VDD.t3473 213.931
R1114 VDD.t3473 VDD.t3513 213.931
R1115 VDD.t3513 VDD.t1483 213.931
R1116 VDD.t1483 VDD.t3512 213.931
R1117 VDD.t1893 VDD.t1897 213.931
R1118 VDD.t1897 VDD.t3076 213.931
R1119 VDD.t3076 VDD.t3074 213.931
R1120 VDD.t3074 VDD.t3075 213.931
R1121 VDD.t2989 VDD.t2991 213.931
R1122 VDD.t2991 VDD.t174 213.931
R1123 VDD.t174 VDD.t175 213.931
R1124 VDD.t175 VDD.t176 213.931
R1125 VDD.t328 VDD.t326 213.931
R1126 VDD.t326 VDD.t502 213.931
R1127 VDD.t502 VDD.t503 213.931
R1128 VDD.t503 VDD.t501 213.931
R1129 VDD.t579 VDD.t581 213.931
R1130 VDD.t581 VDD.t3241 213.931
R1131 VDD.t3241 VDD.t3240 213.931
R1132 VDD.t3240 VDD.t2517 213.931
R1133 VDD.t2625 VDD.t2627 213.931
R1134 VDD.t2627 VDD.t2792 213.931
R1135 VDD.t2792 VDD.t2790 213.931
R1136 VDD.t2790 VDD.t2791 213.931
R1137 VDD.t659 VDD.t657 213.931
R1138 VDD.t657 VDD.t20 213.931
R1139 VDD.t20 VDD.t21 213.931
R1140 VDD.t21 VDD.t22 213.931
R1141 VDD.t39 VDD.t407 213.931
R1142 VDD.t407 VDD.t1105 213.931
R1143 VDD.t1105 VDD.t1103 213.931
R1144 VDD.t1103 VDD.t1104 213.931
R1145 VDD.t1122 VDD.t1124 213.931
R1146 VDD.t1124 VDD.t767 213.931
R1147 VDD.t767 VDD.t768 213.931
R1148 VDD.t768 VDD.t1572 213.931
R1149 VDD.t3708 VDD.t3720 213.931
R1150 VDD.t3720 VDD.t3704 213.931
R1151 VDD.t2119 VDD.t3414 213.931
R1152 VDD.t3414 VDD.t4538 213.931
R1153 VDD.t4538 VDD.t4537 213.931
R1154 VDD.t4537 VDD.t4536 213.931
R1155 VDD.t166 VDD.t71 213.931
R1156 VDD.t71 VDD.t158 213.931
R1157 VDD.t902 VDD.t912 213.931
R1158 VDD.t912 VDD.t2168 213.931
R1159 VDD.t4530 VDD.t2400 213.931
R1160 VDD.t2400 VDD.t4522 213.931
R1161 VDD.t4469 VDD.t492 213.931
R1162 VDD.t492 VDD.t4465 213.931
R1163 VDD.t1244 VDD.t1228 213.931
R1164 VDD.t1228 VDD.t1234 213.931
R1165 VDD.t4092 VDD.t4096 213.931
R1166 VDD.t4096 VDD.t4104 213.931
R1167 VDD.t214 VDD.t3562 213.931
R1168 VDD.t3562 VDD.t210 213.931
R1169 VDD.t17 VDD.t2487 205.749
R1170 VDD.t3061 VDD.t3485 205.749
R1171 VDD.t377 VDD.t362 205.749
R1172 VDD.t1331 VDD.t470 205.749
R1173 VDD.t2487 VDD.t3630 197.707
R1174 VDD.t3630 VDD.t3620 197.707
R1175 VDD.t3485 VDD.t3479 197.707
R1176 VDD.t3479 VDD.t3487 197.707
R1177 VDD.t2875 VDD.t4229 197.707
R1178 VDD.t362 VDD.t4461 197.707
R1179 VDD.t4461 VDD.t364 197.707
R1180 VDD.t4578 VDD.t4572 197.707
R1181 VDD.t470 VDD.t1058 197.707
R1182 VDD.t1058 VDD.t474 197.707
R1183 VDD.t1138 VDD.t1146 197.707
R1184 VDD.t4501 VDD.t4499 197.707
R1185 VDD.t4353 VDD.t4355 196.666
R1186 VDD.t4351 VDD.t4353 196.666
R1187 VDD.t1650 VDD.t4351 196.666
R1188 VDD.t1648 VDD.t1650 196.666
R1189 VDD.t1644 VDD.t1648 196.666
R1190 VDD.t2012 VDD.t290 196.666
R1191 VDD.t290 VDD.t1998 196.666
R1192 VDD.t1982 VDD.t2735 196.666
R1193 VDD.t1984 VDD.t1982 196.666
R1194 VDD.t3024 VDD.t1984 196.666
R1195 VDD.t1454 VDD.t3024 196.666
R1196 VDD.t3013 VDD.t1454 196.666
R1197 VDD.t2437 VDD.t1907 196.666
R1198 VDD.t1907 VDD.t2655 196.666
R1199 VDD.t1574 VDD.t1569 196.666
R1200 VDD.t1567 VDD.t1574 196.666
R1201 VDD.t1877 VDD.t1567 196.666
R1202 VDD.t934 VDD.t1877 196.666
R1203 VDD.t1873 VDD.t934 196.666
R1204 VDD.t2087 VDD.t3456 196.666
R1205 VDD.t3456 VDD.t3452 196.666
R1206 VDD.t2797 VDD.t2795 196.666
R1207 VDD.t2793 VDD.t2797 196.666
R1208 VDD.t2092 VDD.t2793 196.666
R1209 VDD.t3465 VDD.t2092 196.666
R1210 VDD.t2082 VDD.t3465 196.666
R1211 VDD.t1909 VDD.t2420 196.666
R1212 VDD.t2420 VDD.t2661 196.666
R1213 VDD.t3003 VDD.t3005 196.666
R1214 VDD.t3001 VDD.t3003 196.666
R1215 VDD.t3454 VDD.t3001 196.666
R1216 VDD.t3450 VDD.t3454 196.666
R1217 VDD.t3446 VDD.t3450 196.666
R1218 VDD.t1377 VDD.t1383 196.666
R1219 VDD.t1383 VDD.t1381 196.666
R1220 VDD.t4440 VDD.t421 196.666
R1221 VDD.t419 VDD.t4440 196.666
R1222 VDD.t1474 VDD.t419 196.666
R1223 VDD.t1472 VDD.t1474 196.666
R1224 VDD.t1469 VDD.t1472 196.666
R1225 VDD.t1839 VDD.t1833 196.666
R1226 VDD.t1833 VDD.t1829 196.666
R1227 VDD.t2067 VDD.t2071 196.666
R1228 VDD.t2069 VDD.t2067 196.666
R1229 VDD.t2408 VDD.t2069 196.666
R1230 VDD.t1851 VDD.t2408 196.666
R1231 VDD.t1811 VDD.t1851 196.666
R1232 VDD.t4396 VDD.t4377 196.666
R1233 VDD.t4377 VDD.t4400 196.666
R1234 VDD.t1272 VDD.t1276 196.666
R1235 VDD.t1274 VDD.t1272 196.666
R1236 VDD.t4121 VDD.t1274 196.666
R1237 VDD.t4119 VDD.t4121 196.666
R1238 VDD.t2422 VDD.t4119 196.666
R1239 VDD.t2010 VDD.t274 196.666
R1240 VDD.t274 VDD.t2005 196.666
R1241 VDD.t1794 VDD.t1792 196.666
R1242 VDD.t1790 VDD.t1794 196.666
R1243 VDD.t1407 VDD.t1790 196.666
R1244 VDD.t3311 VDD.t1407 196.666
R1245 VDD.t1379 VDD.t3311 196.666
R1246 VDD.t2014 VDD.t2026 196.666
R1247 VDD.t2026 VDD.t288 196.666
R1248 VDD.t4238 VDD.t123 196.666
R1249 VDD.t125 VDD.t4238 196.666
R1250 VDD.t3548 VDD.t125 196.666
R1251 VDD.t3550 VDD.t3548 196.666
R1252 VDD.t4409 VDD.t3550 196.666
R1253 VDD.t1419 VDD.t1403 196.666
R1254 VDD.t1403 VDD.t1401 196.666
R1255 VDD.t4445 VDD.t343 196.666
R1256 VDD.t4443 VDD.t4445 196.666
R1257 VDD.t1849 VDD.t4443 196.666
R1258 VDD.t1845 VDD.t1849 196.666
R1259 VDD.t1841 VDD.t1845 196.666
R1260 VDD.t2089 VDD.t3438 196.666
R1261 VDD.t3438 VDD.t3434 196.666
R1262 VDD.t2287 VDD.t2097 196.666
R1263 VDD.t3159 VDD.t2287 196.666
R1264 VDD.t3315 VDD.t3159 196.666
R1265 VDD.t1397 VDD.t3315 196.666
R1266 VDD.t1393 VDD.t1397 196.666
R1267 VDD.t3026 VDD.t3033 196.666
R1268 VDD.t3033 VDD.t3031 196.666
R1269 VDD.t113 VDD.t7 196.666
R1270 VDD.t111 VDD.t113 196.666
R1271 VDD.t1442 VDD.t111 196.666
R1272 VDD.t3011 VDD.t1442 196.666
R1273 VDD.t1476 VDD.t3011 196.666
R1274 VDD.t1646 VDD.t1889 196.666
R1275 VDD.t1889 VDD.t1881 196.666
R1276 VDD.t2111 VDD.t2113 196.666
R1277 VDD.t2115 VDD.t2111 196.666
R1278 VDD.t3544 VDD.t2115 196.666
R1279 VDD.t1318 VDD.t3544 196.666
R1280 VDD.t1322 VDD.t1318 196.666
R1281 VDD.t3066 VDD.t2428 196.666
R1282 VDD.t2428 VDD.t2426 196.666
R1283 VDD.t2999 VDD.t2997 196.666
R1284 VDD.t2995 VDD.t2999 196.666
R1285 VDD.t3481 VDD.t2995 196.666
R1286 VDD.t3489 VDD.t3481 196.666
R1287 VDD.t1109 VDD.t3489 196.666
R1288 VDD.t2871 VDD.t4225 196.666
R1289 VDD.t4225 VDD.t4231 196.666
R1290 VDD.t4015 VDD.t4013 196.666
R1291 VDD.t2800 VDD.t4015 196.666
R1292 VDD.t4392 VDD.t2800 196.666
R1293 VDD.t1320 VDD.t4392 196.666
R1294 VDD.t4381 VDD.t1320 196.666
R1295 VDD.t1869 VDD.t1885 196.666
R1296 VDD.t1885 VDD.t926 196.666
R1297 VDD.t4072 VDD.t4070 196.666
R1298 VDD.t4068 VDD.t4072 196.666
R1299 VDD.t4459 VDD.t4068 196.666
R1300 VDD.t358 VDD.t4459 196.666
R1301 VDD.t366 VDD.t358 196.666
R1302 VDD.t4570 VDD.t4580 196.666
R1303 VDD.t4580 VDD.t4566 196.666
R1304 VDD.t603 VDD.t601 196.666
R1305 VDD.t599 VDD.t603 196.666
R1306 VDD.t1060 VDD.t599 196.666
R1307 VDD.t472 VDD.t1060 196.666
R1308 VDD.t1054 VDD.t472 196.666
R1309 VDD.t1152 VDD.t1142 196.666
R1310 VDD.t1142 VDD.t1148 196.666
R1311 VDD.t4544 VDD.t534 196.666
R1312 VDD.t4542 VDD.t4544 196.666
R1313 VDD.t3628 VDD.t4542 196.666
R1314 VDD.t3626 VDD.t3628 196.666
R1315 VDD.t3624 VDD.t3626 196.666
R1316 VDD.t2556 VDD.t4497 196.666
R1317 VDD.t4497 VDD.t4495 196.666
R1318 VDD.t3966 VDD.t3968 196.666
R1319 VDD.t3974 VDD.t3966 196.666
R1320 VDD.t3734 VDD.t1362 196.666
R1321 VDD.t1362 VDD.t1358 196.666
R1322 VDD.t1358 VDD.t3354 196.666
R1323 VDD.t3354 VDD.t3352 196.666
R1324 VDD.t3352 VDD.t3598 196.666
R1325 VDD.t1449 VDD.t1451 196.666
R1326 VDD.t1446 VDD.t1449 196.666
R1327 VDD.t1391 VDD.t1389 196.666
R1328 VDD.t1389 VDD.t3317 196.666
R1329 VDD.t3317 VDD.t1366 196.666
R1330 VDD.t1366 VDD.t1364 196.666
R1331 VDD.t1364 VDD.t2450 196.666
R1332 VDD.t2300 VDD.t2319 196.666
R1333 VDD.t2296 VDD.t2300 196.666
R1334 VDD.t2226 VDD.t2224 196.666
R1335 VDD.t2224 VDD.t2214 196.666
R1336 VDD.t2214 VDD.t3609 196.666
R1337 VDD.t3609 VDD.t3607 196.666
R1338 VDD.t3607 VDD.t3605 196.666
R1339 VDD.t3120 VDD.t3118 192.281
R1340 VDD.t3368 VDD.t4176 192.281
R1341 VDD.t3368 VDD.t4174 192.281
R1342 VDD.t3146 VDD.t3144 192.281
R1343 VDD.t2883 VDD.t2885 192.281
R1344 VDD.t2883 VDD.t2887 192.281
R1345 VDD.t13 VDD.t3161 192.281
R1346 VDD.t3641 VDD.t3637 192.281
R1347 VDD.t3641 VDD.t3639 192.281
R1348 VDD.t4510 VDD.t2099 192.281
R1349 VDD.t31 VDD.t4589 192.281
R1350 VDD.t31 VDD.t4587 192.281
R1351 VDD.t2550 VDD.t2548 192.281
R1352 VDD.t2536 VDD.t3535 192.281
R1353 VDD.t2536 VDD.t2538 192.281
R1354 VDD.t1628 VDD.t1630 192.281
R1355 VDD.t4194 VDD.t4252 192.281
R1356 VDD.t4194 VDD.t4250 192.281
R1357 VDD.t1755 VDD.t1084 192.281
R1358 VDD.t427 VDD.t425 192.281
R1359 VDD.t2139 VDD.t2629 192.281
R1360 VDD.t2139 VDD.t2141 192.281
R1361 VDD.t970 VDD.t968 192.281
R1362 VDD.t970 VDD.t966 192.281
R1363 VDD.t413 VDD.t220 191.952
R1364 VDD.t413 VDD.t411 191.952
R1365 VDD.t2895 VDD.t3236 190
R1366 VDD.t2895 VDD.t3238 190
R1367 VDD.n1043 VDD.n1042 184.375
R1368 VDD.n918 VDD.n917 184.375
R1369 VDD.n943 VDD.n942 184.375
R1370 VDD.n1018 VDD.n1017 184.375
R1371 VDD.n993 VDD.n992 184.375
R1372 VDD.n968 VDD.n967 184.375
R1373 VDD.n893 VDD.n892 184.375
R1374 VDD.n869 VDD.n868 184.375
R1375 VDD.n639 VDD.n638 184.375
R1376 VDD.n657 VDD.n656 184.375
R1377 VDD.n675 VDD.n674 184.375
R1378 VDD.n692 VDD.n691 184.375
R1379 VDD.n621 VDD.n620 184.375
R1380 VDD.n752 VDD.n751 184.375
R1381 VDD.n770 VDD.n769 184.375
R1382 VDD.n788 VDD.n787 184.375
R1383 VDD.n1744 VDD.n1743 184.375
R1384 VDD.n1769 VDD.n1768 184.375
R1385 VDD.n1862 VDD.n1861 184.375
R1386 VDD.n1837 VDD.n1836 184.375
R1387 VDD.n1819 VDD.n1818 184.375
R1388 VDD.n1794 VDD.n1793 184.375
R1389 VDD.n1719 VDD.n1718 184.375
R1390 VDD.n1695 VDD.n1694 184.375
R1391 VDD.n1537 VDD.n1536 184.375
R1392 VDD.n1562 VDD.n1561 184.375
R1393 VDD.n1662 VDD.n1661 184.375
R1394 VDD.n1637 VDD.n1636 184.375
R1395 VDD.n1612 VDD.n1611 184.375
R1396 VDD.n1587 VDD.n1586 184.375
R1397 VDD.n1512 VDD.n1511 184.375
R1398 VDD.n1488 VDD.n1487 184.375
R1399 VDD.n1387 VDD.n1386 184.375
R1400 VDD.n1362 VDD.n1361 184.375
R1401 VDD.n1263 VDD.n1262 184.375
R1402 VDD.n1287 VDD.n1286 184.375
R1403 VDD.n1312 VDD.n1311 184.375
R1404 VDD.n1337 VDD.n1336 184.375
R1405 VDD.n1412 VDD.n1411 184.375
R1406 VDD.n1437 VDD.n1436 184.375
R1407 VDD.n2605 VDD.n2604 184.375
R1408 VDD.n2466 VDD.n2465 184.375
R1409 VDD.n2485 VDD.n2484 184.375
R1410 VDD.n2545 VDD.n2544 184.375
R1411 VDD.n2565 VDD.n2564 184.375
R1412 VDD.n2585 VDD.n2584 184.375
R1413 VDD.n2525 VDD.n2524 184.375
R1414 VDD.n2505 VDD.n2504 184.375
R1415 VDD.n2389 VDD.n2388 184.375
R1416 VDD.n2257 VDD.n2256 184.375
R1417 VDD.n2276 VDD.n2275 184.375
R1418 VDD.n2329 VDD.n2328 184.375
R1419 VDD.n2349 VDD.n2348 184.375
R1420 VDD.n2369 VDD.n2368 184.375
R1421 VDD.n2316 VDD.n2315 184.375
R1422 VDD.n2296 VDD.n2295 184.375
R1423 VDD.n1046 VDD.n1045 182.117
R1424 VDD.n921 VDD.n920 182.117
R1425 VDD.n946 VDD.n945 182.117
R1426 VDD.n1021 VDD.n1020 182.117
R1427 VDD.n996 VDD.n995 182.117
R1428 VDD.n971 VDD.n970 182.117
R1429 VDD.n896 VDD.n895 182.117
R1430 VDD.n872 VDD.n871 182.117
R1431 VDD.n631 VDD.n629 182.117
R1432 VDD.n649 VDD.n647 182.117
R1433 VDD.n667 VDD.n665 182.117
R1434 VDD.n684 VDD.n682 182.117
R1435 VDD.n613 VDD.n611 182.117
R1436 VDD.n744 VDD.n742 182.117
R1437 VDD.n762 VDD.n760 182.117
R1438 VDD.n780 VDD.n778 182.117
R1439 VDD.n1736 VDD.n1734 182.117
R1440 VDD.n1761 VDD.n1759 182.117
R1441 VDD.n1866 VDD.n1864 182.117
R1442 VDD.n1841 VDD.n1839 182.117
R1443 VDD.n1811 VDD.n1809 182.117
R1444 VDD.n1786 VDD.n1784 182.117
R1445 VDD.n1711 VDD.n1709 182.117
R1446 VDD.n1687 VDD.n1685 182.117
R1447 VDD.n1541 VDD.n1539 182.117
R1448 VDD.n1566 VDD.n1564 182.117
R1449 VDD.n1666 VDD.n1664 182.117
R1450 VDD.n1641 VDD.n1639 182.117
R1451 VDD.n1616 VDD.n1614 182.117
R1452 VDD.n1591 VDD.n1589 182.117
R1453 VDD.n1516 VDD.n1514 182.117
R1454 VDD.n1492 VDD.n1490 182.117
R1455 VDD.n1391 VDD.n1389 182.117
R1456 VDD.n1366 VDD.n1364 182.117
R1457 VDD.n1267 VDD.n1265 182.117
R1458 VDD.n1291 VDD.n1289 182.117
R1459 VDD.n1316 VDD.n1314 182.117
R1460 VDD.n1341 VDD.n1339 182.117
R1461 VDD.n1416 VDD.n1414 182.117
R1462 VDD.n1441 VDD.n1439 182.117
R1463 VDD.n2597 VDD.n2595 182.117
R1464 VDD.n2458 VDD.n2456 182.117
R1465 VDD.n2477 VDD.n2475 182.117
R1466 VDD.n2537 VDD.n2535 182.117
R1467 VDD.n2557 VDD.n2555 182.117
R1468 VDD.n2577 VDD.n2575 182.117
R1469 VDD.n2517 VDD.n2515 182.117
R1470 VDD.n2497 VDD.n2495 182.117
R1471 VDD.n2393 VDD.n2391 182.117
R1472 VDD.n2249 VDD.n2247 182.117
R1473 VDD.n2268 VDD.n2266 182.117
R1474 VDD.n2333 VDD.n2331 182.117
R1475 VDD.n2353 VDD.n2351 182.117
R1476 VDD.n2373 VDD.n2371 182.117
R1477 VDD.n2308 VDD.n2306 182.117
R1478 VDD.n2288 VDD.n2286 182.117
R1479 VDD.n2084 VDD.t189 174.172
R1480 VDD.n2090 VDD.t3979 173.061
R1481 VDD.n2120 VDD.t3777 172.51
R1482 VDD.n2114 VDD.t3017 172.51
R1483 VDD.n2108 VDD.t2078 172.51
R1484 VDD.n2102 VDD.t2021 172.51
R1485 VDD.n2096 VDD.t4373 172.51
R1486 VDD.n2078 VDD.t896 172.51
R1487 VDD.n2085 VDD.t148 170.712
R1488 VDD.n2178 VDD.t3724 170.677
R1489 VDD.n2162 VDD.t2460 170.677
R1490 VDD.n1465 VDD.t2222 170.677
R1491 VDD.n2042 VDD.t3307 170.677
R1492 VDD.n1942 VDD.t437 170.677
R1493 VDD.n1892 VDD.t2208 170.677
R1494 VDD.n1917 VDD.t2470 170.677
R1495 VDD.n1967 VDD.t2433 170.677
R1496 VDD.n1992 VDD.t936 170.677
R1497 VDD.n2017 VDD.t4110 170.677
R1498 VDD.n2067 VDD.t1550 170.677
R1499 VDD.n2630 VDD.t2599 170.677
R1500 VDD.n2437 VDD.t1399 170.677
R1501 VDD.n2412 VDD.t4112 170.677
R1502 VDD.n2228 VDD.t1863 170.677
R1503 VDD.n2203 VDD.t2435 170.677
R1504 VDD.n2091 VDD.t3991 169.626
R1505 VDD.n2881 VDD.t3116 169.468
R1506 VDD.n2851 VDD.t3148 169.468
R1507 VDD.n2820 VDD.t3163 169.468
R1508 VDD.n554 VDD.t4512 169.468
R1509 VDD.n3100 VDD.t2546 169.468
R1510 VDD.n3124 VDD.t1626 169.468
R1511 VDD.n3213 VDD.t1082 169.468
R1512 VDD.n3237 VDD.t423 169.468
R1513 VDD.n2121 VDD.t3783 169.088
R1514 VDD.n2115 VDD.t1456 169.088
R1515 VDD.n2109 VDD.t2084 169.088
R1516 VDD.n2103 VDD.t261 169.088
R1517 VDD.n2097 VDD.t4390 169.088
R1518 VDD.n2079 VDD.t2323 169.088
R1519 VDD.n2179 VDD.n2178 151.673
R1520 VDD.n1466 VDD.n1465 151.673
R1521 VDD.n2438 VDD.n2437 151.673
R1522 VDD.n2413 VDD.n2412 151.673
R1523 VDD.n2229 VDD.n2228 151.673
R1524 VDD.n2204 VDD.n2203 151.673
R1525 VDD.n2163 VDD.n2162 151.671
R1526 VDD.n2631 VDD.n2630 151.671
R1527 VDD.n2043 VDD.n2042 151.379
R1528 VDD.n1943 VDD.n1942 151.379
R1529 VDD.n1893 VDD.n1892 151.379
R1530 VDD.n1918 VDD.n1917 151.379
R1531 VDD.n1968 VDD.n1967 151.379
R1532 VDD.n1993 VDD.n1992 151.379
R1533 VDD.n2018 VDD.n2017 151.379
R1534 VDD.n2068 VDD.n2067 151.379
R1535 VDD.t4387 VDD.t4395 144.087
R1536 VDD.t3543 VDD.t4387 144.087
R1537 VDD.t4125 VDD.t3543 144.087
R1538 VDD.t2028 VDD.t2032 144.087
R1539 VDD.t2025 VDD.t2028 144.087
R1540 VDD.t1883 VDD.t2025 144.087
R1541 VDD.t3009 VDD.t3010 144.087
R1542 VDD.t1458 VDD.t3009 144.087
R1543 VDD.t1415 VDD.t1458 144.087
R1544 VDD.t1930 VDD.t1931 144.087
R1545 VDD.t1934 VDD.t1930 144.087
R1546 VDD.t2456 VDD.t1934 144.087
R1547 VDD.t2328 VDD.t2333 144.087
R1548 VDD.t2325 VDD.t2328 144.087
R1549 VDD.t2202 VDD.t2325 144.087
R1550 VDD.t3781 VDD.t3782 143.717
R1551 VDD.t3772 VDD.t3781 143.717
R1552 VDD.t2615 VDD.t3772 143.717
R1553 VDD.t3428 VDD.t3429 143.717
R1554 VDD.t3427 VDD.t3428 143.717
R1555 VDD.t2414 VDD.t3427 143.717
R1556 VDD.t3978 VDD.t3996 143.717
R1557 VDD.t3977 VDD.t3978 143.717
R1558 VDD.t435 VDD.t3977 143.717
R1559 VDD.n3004 VDD.n3003 142.5
R1560 VDD.n3192 VDD.n3191 142.5
R1561 VDD.n3074 VDD.n3073 142.5
R1562 VDD.n356 VDD.n355 142.5
R1563 VDD.n455 VDD.n454 142.5
R1564 VDD.n523 VDD.n522 142.5
R1565 VDD.n2807 VDD.n2806 142.5
R1566 VDD.n2744 VDD.n2743 142.5
R1567 VDD.n1158 VDD.t4125 137.982
R1568 VDD.n1173 VDD.t1883 137.982
R1569 VDD.n1203 VDD.t1415 137.982
R1570 VDD.n1131 VDD.t2456 137.982
R1571 VDD.n1236 VDD.t2202 137.982
R1572 VDD.t1928 VDD.t3395 137.714
R1573 VDD.t1926 VDD.t1928 137.714
R1574 VDD.t2183 VDD.t2184 137.714
R1575 VDD.t1525 VDD.t1523 137.714
R1576 VDD.t4603 VDD.t4602 137.714
R1577 VDD.t4602 VDD.t4601 137.714
R1578 VDD.t3019 VDD.t3028 137.714
R1579 VDD.t3007 VDD.t3019 137.714
R1580 VDD.t2185 VDD.t2186 137.714
R1581 VDD.t1729 VDD.t1801 137.714
R1582 VDD.t2009 VDD.t2001 137.714
R1583 VDD.t2001 VDD.t2000 137.714
R1584 VDD.t3461 VDD.t3463 137.714
R1585 VDD.t3459 VDD.t3461 137.714
R1586 VDD.t2034 VDD.t2035 137.714
R1587 VDD.t3871 VDD.t1339 137.714
R1588 VDD.t4385 VDD.t3283 137.714
R1589 VDD.t3283 VDD.t3282 137.714
R1590 VDD.t3972 VDD.t3993 137.714
R1591 VDD.t3970 VDD.t3972 137.714
R1592 VDD.t2807 VDD.t2808 137.714
R1593 VDD.t3681 VDD.t3811 137.714
R1594 VDD.t2315 VDD.t2314 137.714
R1595 VDD.t2314 VDD.t898 137.714
R1596 VDD.t4411 VDD.t4406 137.714
R1597 VDD.t1316 VDD.t4411 137.714
R1598 VDD.t354 VDD.t355 137.714
R1599 VDD.t3949 VDD.t1767 137.714
R1600 VDD.t3400 VDD.t3394 137.714
R1601 VDD.t3394 VDD.t1921 137.714
R1602 VDD.t284 VDD.t286 137.714
R1603 VDD.t280 VDD.t284 137.714
R1604 VDD.t3384 VDD.t1964 137.714
R1605 VDD.t2368 VDD.t3212 137.714
R1606 VDD.t3987 VDD.t3965 137.714
R1607 VDD.t3965 VDD.t3964 137.714
R1608 VDD.t3763 VDD.t3779 137.714
R1609 VDD.t3767 VDD.t3763 137.714
R1610 VDD.t4149 VDD.t4150 137.714
R1611 VDD.t4043 VDD.t3337 137.714
R1612 VDD.t2086 VDD.t3433 137.714
R1613 VDD.t3433 VDD.t3432 137.714
R1614 VDD.t4604 VDD.t4599 137.714
R1615 VDD.t4606 VDD.t4604 137.714
R1616 VDD.t4192 VDD.t4193 137.714
R1617 VDD.t4007 VDD.t1737 137.714
R1618 VDD.t1448 VDD.t1445 137.714
R1619 VDD.t1445 VDD.t3015 137.714
R1620 VDD.t555 VDD.t3857 137.714
R1621 VDD.t553 VDD.t555 137.714
R1622 VDD.t873 VDD.t1622 137.714
R1623 VDD.t1208 VDD.t711 137.714
R1624 VDD.t630 VDD.t629 137.714
R1625 VDD.t629 VDD.t631 137.714
R1626 VDD.t1607 VDD.t1609 137.714
R1627 VDD.t1605 VDD.t1607 137.714
R1628 VDD.t1958 VDD.t1959 137.714
R1629 VDD.t791 VDD.t833 137.714
R1630 VDD.t662 VDD.t664 137.714
R1631 VDD.t664 VDD.t663 137.714
R1632 VDD.t2697 VDD.t2699 137.714
R1633 VDD.t605 VDD.t2697 137.714
R1634 VDD.t3244 VDD.t3242 137.714
R1635 VDD.t793 VDD.t1194 137.714
R1636 VDD.t1115 VDD.t1114 137.714
R1637 VDD.t1114 VDD.t1113 137.714
R1638 VDD.t3859 VDD.t3861 137.714
R1639 VDD.t3863 VDD.t3859 137.714
R1640 VDD.t2837 VDD.t2839 137.714
R1641 VDD.t1226 VDD.t725 137.714
R1642 VDD.t2682 VDD.t3532 137.714
R1643 VDD.t3532 VDD.t2683 137.714
R1644 VDD.t356 VDD.t560 137.714
R1645 VDD.t3522 VDD.t356 137.714
R1646 VDD.t4132 VDD.t4131 137.714
R1647 VDD.t687 VDD.t1174 137.714
R1648 VDD.t577 VDD.t578 137.714
R1649 VDD.t578 VDD.t576 137.714
R1650 VDD.t450 VDD.t452 137.714
R1651 VDD.t448 VDD.t450 137.714
R1652 VDD.t3129 VDD.t1659 137.714
R1653 VDD.t1164 VDD.t731 137.714
R1654 VDD.t120 VDD.t122 137.714
R1655 VDD.t122 VDD.t121 137.714
R1656 VDD.t2788 VDD.t2784 137.714
R1657 VDD.t2786 VDD.t2788 137.714
R1658 VDD.t3418 VDD.t3505 137.714
R1659 VDD.t739 VDD.t799 137.714
R1660 VDD.t134 VDD.t1271 137.714
R1661 VDD.t1271 VDD.t1270 137.714
R1662 VDD.t2845 VDD.t2847 137.714
R1663 VDD.t2849 VDD.t2845 137.714
R1664 VDD.t656 VDD.t956 137.714
R1665 VDD.t1222 VDD.t713 137.714
R1666 VDD.t2696 VDD.t2694 137.714
R1667 VDD.t2694 VDD.t2695 137.714
R1668 VDD.t1612 VDD.t2109 137.714
R1669 VDD.t1614 VDD.t1612 137.714
R1670 VDD.t4293 VDD.t3056 137.714
R1671 VDD.t3270 VDD.t1724 137.714
R1672 VDD.t3290 VDD.t3288 137.714
R1673 VDD.t3288 VDD.t3289 137.714
R1674 VDD.t1099 VDD.t1097 137.714
R1675 VDD.t1095 VDD.t1099 137.714
R1676 VDD.t2716 VDD.t2052 137.714
R1677 VDD.t3849 VDD.t3807 137.714
R1678 VDD.t1978 VDD.t1976 137.714
R1679 VDD.t1976 VDD.t1977 137.714
R1680 VDD.t4064 VDD.t2731 137.714
R1681 VDD.t4066 VDD.t4064 137.714
R1682 VDD.t2124 VDD.t598 137.714
R1683 VDD.t2366 VDD.t3875 137.714
R1684 VDD.t292 VDD.t613 137.714
R1685 VDD.t613 VDD.t293 137.714
R1686 VDD.t4595 VDD.t4593 137.714
R1687 VDD.t4591 VDD.t4595 137.714
R1688 VDD.t145 VDD.t583 137.714
R1689 VDD.t4041 VDD.t3254 137.714
R1690 VDD.t2127 VDD.t2128 137.714
R1691 VDD.t2128 VDD.t2129 137.714
R1692 VDD.t1696 VDD.t1694 137.714
R1693 VDD.t1692 VDD.t1696 137.714
R1694 VDD.t1798 VDD.t4292 137.714
R1695 VDD.t1733 VDD.t3805 137.714
R1696 VDD.t1336 VDD.t1335 137.714
R1697 VDD.t1335 VDD.t1334 137.714
R1698 VDD.t4453 VDD.t4449 137.714
R1699 VDD.t4451 VDD.t4453 137.714
R1700 VDD.t3472 VDD.t3471 137.714
R1701 VDD.t2246 VDD.t3814 137.714
R1702 VDD.t4236 VDD.t4237 137.714
R1703 VDD.t4237 VDD.t4235 137.714
R1704 VDD.t44 VDD.t48 137.714
R1705 VDD.t46 VDD.t44 137.714
R1706 VDD.t3649 VDD.t3648 137.714
R1707 VDD.t3196 VDD.t1337 137.714
R1708 VDD.t4514 VDD.t4516 137.714
R1709 VDD.t4516 VDD.t4515 137.714
R1710 VDD.t1714 VDD.t1718 137.714
R1711 VDD.t1716 VDD.t1714 137.714
R1712 VDD.t649 VDD.t1774 137.714
R1713 VDD.t3183 VDD.t3220 137.714
R1714 VDD.t500 VDD.t498 137.714
R1715 VDD.t498 VDD.t499 137.714
R1716 VDD.t4485 VDD.t4487 137.714
R1717 VDD.t4483 VDD.t4485 137.714
R1718 VDD.t2524 VDD.t2449 137.714
R1719 VDD.t705 VDD.t701 137.714
R1720 VDD.t2870 VDD.t3567 137.714
R1721 VDD.t3567 VDD.t1571 137.714
R1722 VDD.t1293 VDD.t1295 137.714
R1723 VDD.t1291 VDD.t1293 137.714
R1724 VDD.t4075 VDD.t4076 137.714
R1725 VDD.t819 VDD.t689 137.714
R1726 VDD.t369 VDD.t368 137.714
R1727 VDD.t368 VDD.t2819 137.714
R1728 VDD.t4209 VDD.t4205 137.714
R1729 VDD.t4207 VDD.t4209 137.714
R1730 VDD.t2362 VDD.t1766 137.714
R1731 VDD.t1190 VDD.t1180 137.714
R1732 VDD.t4586 VDD.t4585 137.714
R1733 VDD.t4585 VDD.t4584 137.714
R1734 VDD.t35 VDD.t37 137.714
R1735 VDD.t33 VDD.t35 137.714
R1736 VDD.t128 VDD.t129 137.714
R1737 VDD.t695 VDD.t4361 137.714
R1738 VDD.t2432 VDD.t2431 137.714
R1739 VDD.t2431 VDD.t2430 137.714
R1740 VDD.t3687 VDD.t3683 137.714
R1741 VDD.t3685 VDD.t3687 137.714
R1742 VDD.t1027 VDD.t394 137.714
R1743 VDD.t709 VDD.t707 137.714
R1744 VDD.t505 VDD.t506 137.714
R1745 VDD.t506 VDD.t507 137.714
R1746 VDD.t1093 VDD.t1089 137.714
R1747 VDD.t1091 VDD.t1093 137.714
R1748 VDD.t3128 VDD.t2674 137.714
R1749 VDD.t1182 VDD.t1176 137.714
R1750 VDD.t3930 VDD.t3929 137.714
R1751 VDD.t3929 VDD.t3928 137.714
R1752 VDD.t2253 VDD.t2255 137.714
R1753 VDD.t1101 VDD.t2253 137.714
R1754 VDD.t54 VDD.t55 137.714
R1755 VDD.t817 VDD.t807 137.714
R1756 VDD.t142 VDD.t144 137.714
R1757 VDD.t144 VDD.t143 137.714
R1758 VDD.t2503 VDD.t2499 137.714
R1759 VDD.t2501 VDD.t2503 137.714
R1760 VDD.t2897 VDD.t3165 137.714
R1761 VDD.t737 VDD.t729 137.714
R1762 VDD.t504 VDD.t27 137.714
R1763 VDD.t27 VDD.t26 137.714
R1764 VDD.t442 VDD.t444 137.714
R1765 VDD.t446 VDD.t442 137.714
R1766 VDD.t1991 VDD.t1989 137.714
R1767 VDD.t3912 VDD.t1726 137.714
R1768 VDD.t1987 VDD.t1988 137.714
R1769 VDD.t1988 VDD.t1986 137.714
R1770 VDD.t3419 VDD.t3421 137.714
R1771 VDD.t3423 VDD.t3419 137.714
R1772 VDD.t388 VDD.t2744 137.714
R1773 VDD.t2386 VDD.t2372 137.714
R1774 VDD.t3787 VDD.t3786 137.714
R1775 VDD.t3786 VDD.t3785 137.714
R1776 VDD.t380 VDD.t382 137.714
R1777 VDD.t378 VDD.t380 137.714
R1778 VDD.t2528 VDD.t2526 137.714
R1779 VDD.t1507 VDD.t2044 137.714
R1780 VDD.t2486 VDD.t1583 137.714
R1781 VDD.t1583 VDD.t1582 137.714
R1782 VDD.t2105 VDD.t2101 137.714
R1783 VDD.t2103 VDD.t2105 137.714
R1784 VDD.t140 VDD.t141 137.714
R1785 VDD.t3842 VDD.t3846 137.714
R1786 VDD.t1012 VDD.t1121 137.714
R1787 VDD.t1121 VDD.t1120 137.714
R1788 VDD.t3372 VDD.t3374 137.714
R1789 VDD.t3376 VDD.t3372 137.714
R1790 VDD.t1330 VDD.t1328 137.714
R1791 VDD.t3916 VDD.t3851 137.714
R1792 VDD.t197 VDD.t196 137.714
R1793 VDD.t196 VDD.t195 137.714
R1794 VDD.t4189 VDD.t3333 137.714
R1795 VDD.t3335 VDD.t4189 137.714
R1796 VDD.t3566 VDD.t3564 137.714
R1797 VDD.t3844 VDD.t4003 137.714
R1798 VDD.t406 VDD.t405 137.714
R1799 VDD.t405 VDD.t404 137.714
R1800 VDD.t2748 VDD.t2750 137.714
R1801 VDD.t2746 VDD.t2748 137.714
R1802 VDD.t1956 VDD.t1957 137.714
R1803 VDD.t4056 VDD.t3823 137.714
R1804 VDD.t385 VDD.t384 137.714
R1805 VDD.t384 VDD.t386 137.714
R1806 VDD.t4476 VDD.t4478 137.714
R1807 VDD.t4474 VDD.t4476 137.714
R1808 VDD.t2869 VDD.t260 137.714
R1809 VDD.t2392 VDD.t2382 137.714
R1810 VDD.t1135 VDD.t1137 137.714
R1811 VDD.t1137 VDD.t1136 137.714
R1812 VDD.t4481 VDD.t4482 137.714
R1813 VDD.t4480 VDD.t4481 137.714
R1814 VDD.t4279 VDD.t3899 137.714
R1815 VDD.t1918 VDD.t1917 137.714
R1816 VDD.t2909 VDD.t2911 137.714
R1817 VDD.t2911 VDD.t3319 137.714
R1818 VDD.t2357 VDD.t2358 137.714
R1819 VDD.t2359 VDD.t2357 137.714
R1820 VDD.t4312 VDD.t4316 137.714
R1821 VDD.t74 VDD.t73 137.714
R1822 VDD.t2726 VDD.t2724 137.714
R1823 VDD.t2724 VDD.t2722 137.714
R1824 VDD.t2738 VDD.t2739 137.714
R1825 VDD.t2737 VDD.t2738 137.714
R1826 VDD.t3093 VDD.t3095 137.714
R1827 VDD.t4558 VDD.t575 137.714
R1828 VDD.t298 VDD.t294 137.714
R1829 VDD.t294 VDD.t296 137.714
R1830 VDD.t4248 VDD.t4249 137.714
R1831 VDD.t4247 VDD.t4248 137.714
R1832 VDD.t3901 VDD.t4328 137.714
R1833 VDD.t1770 VDD.t1769 137.714
R1834 VDD.t130 VDD.t2452 137.714
R1835 VDD.t2452 VDD.t132 137.714
R1836 VDD.t4242 VDD.t4240 137.714
R1837 VDD.t4241 VDD.t4242 137.714
R1838 VDD.t4275 VDD.t4306 137.714
R1839 VDD.t3646 VDD.t3645 137.714
R1840 VDD.t2531 VDD.t2529 137.714
R1841 VDD.t2529 VDD.t3526 137.714
R1842 VDD.t591 VDD.t632 137.714
R1843 VDD.t590 VDD.t591 137.714
R1844 VDD.t4332 VDD.t3079 137.714
R1845 VDD.t2285 VDD.t2284 137.714
R1846 VDD.t2828 VDD.t2826 137.714
R1847 VDD.t2826 VDD.t2824 137.714
R1848 VDD.t661 VDD.t115 137.714
R1849 VDD.t116 VDD.t661 137.714
R1850 VDD.t3087 VDD.t3089 137.714
R1851 VDD.t226 VDD.t3574 137.714
R1852 VDD.t1590 VDD.t1588 137.714
R1853 VDD.t1588 VDD.t1592 137.714
R1854 VDD.t3152 VDD.t3153 137.714
R1855 VDD.t3151 VDD.t3152 137.714
R1856 VDD.t3083 VDD.t3099 137.714
R1857 VDD.t4179 VDD.t4178 137.714
R1858 VDD.t2117 VDD.t2773 137.714
R1859 VDD.t2773 VDD.t2771 137.714
R1860 VDD.t4421 VDD.t3101 137.714
R1861 VDD.t4420 VDD.t4421 137.714
R1862 VDD.t2945 VDD.t871 137.714
R1863 VDD.t2193 VDD.t3114 137.714
R1864 VDD.t3170 VDD.t3168 137.714
R1865 VDD.t3168 VDD.t3166 137.714
R1866 VDD.t559 VDD.t558 137.714
R1867 VDD.t557 VDD.t559 137.714
R1868 VDD.t2929 VDD.t839 137.714
R1869 VDD.t81 VDD.t82 137.714
R1870 VDD.t588 VDD.t584 137.714
R1871 VDD.t584 VDD.t586 137.714
R1872 VDD.t3404 VDD.t3403 137.714
R1873 VDD.t3402 VDD.t3404 137.714
R1874 VDD.t2963 VDD.t857 137.714
R1875 VDD.t1284 VDD.t2290 137.714
R1876 VDD.t1048 VDD.t1052 137.714
R1877 VDD.t1052 VDD.t1050 137.714
R1878 VDD.t3659 VDD.t2687 137.714
R1879 VDD.t2686 VDD.t3659 137.714
R1880 VDD.t2959 VDD.t2923 137.714
R1881 VDD.t23 VDD.t25 137.714
R1882 VDD.t2282 VDD.t2278 137.714
R1883 VDD.t2278 VDD.t2280 137.714
R1884 VDD.t3576 VDD.t222 137.714
R1885 VDD.t3575 VDD.t3576 137.714
R1886 VDD.t869 VDD.t841 137.714
R1887 VDD.t3519 VDD.t3520 137.714
R1888 VDD.t465 VDD.t461 137.714
R1889 VDD.t461 VDD.t463 137.714
R1890 VDD.t3696 VDD.t4597 137.714
R1891 VDD.t4598 VDD.t3696 137.714
R1892 VDD.t2941 VDD.t843 137.714
R1893 VDD.t2533 VDD.t2534 137.714
R1894 VDD.t3345 VDD.t3347 137.714
R1895 VDD.t3347 VDD.t1268 137.714
R1896 VDD.t788 VDD.t790 137.714
R1897 VDD.t789 VDD.t788 137.714
R1898 VDD.t2917 VDD.t847 137.714
R1899 VDD.t610 VDD.t562 137.714
R1900 VDD.t320 VDD.t322 137.714
R1901 VDD.t322 VDD.t318 137.714
R1902 VDD.t2898 VDD.t2900 137.714
R1903 VDD.t2899 VDD.t2898 137.714
R1904 VDD.t861 VDD.t863 137.714
R1905 VDD.t4258 VDD.t3604 137.714
R1906 VDD.t2059 VDD.t2061 137.714
R1907 VDD.t2061 VDD.t2057 137.714
R1908 VDD.n1218 VDD.t2615 137.628
R1909 VDD.n1188 VDD.t2414 137.628
R1910 VDD.n1146 VDD.t435 137.628
R1911 VDD.n642 VDD.t873 136.641
R1912 VDD.n660 VDD.t1958 136.641
R1913 VDD.n678 VDD.t3244 136.641
R1914 VDD.n695 VDD.t2837 136.641
R1915 VDD.n624 VDD.t4132 136.641
R1916 VDD.n755 VDD.t3129 136.641
R1917 VDD.n773 VDD.t3418 136.641
R1918 VDD.n791 VDD.t656 136.641
R1919 VDD.n1038 VDD.t2183 136.641
R1920 VDD.n913 VDD.t2185 136.641
R1921 VDD.n938 VDD.t2034 136.641
R1922 VDD.n1013 VDD.t2807 136.641
R1923 VDD.n988 VDD.t354 136.641
R1924 VDD.n963 VDD.t3384 136.641
R1925 VDD.n888 VDD.t4149 136.641
R1926 VDD.n864 VDD.t4192 136.641
R1927 VDD.n1732 VDD.t4293 136.641
R1928 VDD.n1757 VDD.t2716 136.641
R1929 VDD.n1857 VDD.t2124 136.641
R1930 VDD.n1832 VDD.t145 136.641
R1931 VDD.n1807 VDD.t1798 136.641
R1932 VDD.n1782 VDD.t3472 136.641
R1933 VDD.n1707 VDD.t3649 136.641
R1934 VDD.n1683 VDD.t649 136.641
R1935 VDD.n1532 VDD.t2524 136.641
R1936 VDD.n1557 VDD.t4075 136.641
R1937 VDD.n1657 VDD.t2362 136.641
R1938 VDD.n1632 VDD.t128 136.641
R1939 VDD.n1607 VDD.t1027 136.641
R1940 VDD.n1582 VDD.t3128 136.641
R1941 VDD.n1507 VDD.t54 136.641
R1942 VDD.n1483 VDD.t2897 136.641
R1943 VDD.n1382 VDD.t1991 136.641
R1944 VDD.n1357 VDD.t388 136.641
R1945 VDD.n1258 VDD.t2528 136.641
R1946 VDD.n1282 VDD.t140 136.641
R1947 VDD.n1307 VDD.t1330 136.641
R1948 VDD.n1332 VDD.t3566 136.641
R1949 VDD.n1407 VDD.t1956 136.641
R1950 VDD.n1432 VDD.t2869 136.641
R1951 VDD.n2590 VDD.t1918 136.641
R1952 VDD.n2451 VDD.t74 136.641
R1953 VDD.n2470 VDD.t4558 136.641
R1954 VDD.n2530 VDD.t1770 136.641
R1955 VDD.n2550 VDD.t3646 136.641
R1956 VDD.n2570 VDD.t2285 136.641
R1957 VDD.n2510 VDD.t226 136.641
R1958 VDD.n2490 VDD.t4179 136.641
R1959 VDD.n2381 VDD.t2193 136.641
R1960 VDD.n2242 VDD.t81 136.641
R1961 VDD.n2261 VDD.t1284 136.641
R1962 VDD.n2321 VDD.t23 136.641
R1963 VDD.n2341 VDD.t3519 136.641
R1964 VDD.n2361 VDD.t2533 136.641
R1965 VDD.n2301 VDD.t610 136.641
R1966 VDD.n2281 VDD.t4258 136.641
R1967 VDD.t3368 VDD.t3 135.973
R1968 VDD.t2883 VDD.t2775 135.973
R1969 VDD.t3641 VDD.t2859 135.973
R1970 VDD.t31 VDD.t1893 135.973
R1971 VDD.t2536 VDD.t328 135.973
R1972 VDD.t4194 VDD.t2625 135.973
R1973 VDD.t2139 VDD.t1122 135.973
R1974 VDD.t970 VDD.t2119 135.973
R1975 VDD.n643 VDD.t1208 121.615
R1976 VDD.n661 VDD.t791 121.615
R1977 VDD.n679 VDD.t793 121.615
R1978 VDD.n696 VDD.t1226 121.615
R1979 VDD.n625 VDD.t687 121.615
R1980 VDD.n756 VDD.t1164 121.615
R1981 VDD.n774 VDD.t739 121.615
R1982 VDD.n792 VDD.t1222 121.615
R1983 VDD.n1036 VDD.t1525 120.208
R1984 VDD.n911 VDD.t1729 120.208
R1985 VDD.n936 VDD.t3871 120.208
R1986 VDD.n1011 VDD.t3681 120.208
R1987 VDD.n986 VDD.t3949 120.208
R1988 VDD.n961 VDD.t2368 120.208
R1989 VDD.n886 VDD.t4043 120.208
R1990 VDD.n862 VDD.t4007 120.208
R1991 VDD.n1730 VDD.t3270 120.208
R1992 VDD.n1755 VDD.t3849 120.208
R1993 VDD.n1855 VDD.t2366 120.208
R1994 VDD.n1830 VDD.t4041 120.208
R1995 VDD.n1805 VDD.t1733 120.208
R1996 VDD.n1780 VDD.t2246 120.208
R1997 VDD.n1705 VDD.t3196 120.208
R1998 VDD.n1681 VDD.t3183 120.208
R1999 VDD.n1530 VDD.t705 120.208
R2000 VDD.n1555 VDD.t819 120.208
R2001 VDD.n1655 VDD.t1190 120.208
R2002 VDD.n1630 VDD.t695 120.208
R2003 VDD.n1605 VDD.t709 120.208
R2004 VDD.n1580 VDD.t1182 120.208
R2005 VDD.n1505 VDD.t817 120.208
R2006 VDD.n1481 VDD.t737 120.208
R2007 VDD.n1380 VDD.t3912 120.208
R2008 VDD.n1355 VDD.t2386 120.208
R2009 VDD.n1256 VDD.t1507 120.208
R2010 VDD.n1280 VDD.t3842 120.208
R2011 VDD.n1305 VDD.t3916 120.208
R2012 VDD.n1330 VDD.t3844 120.208
R2013 VDD.n1405 VDD.t4056 120.208
R2014 VDD.n1430 VDD.t2392 120.208
R2015 VDD.n2593 VDD.t4279 120.208
R2016 VDD.n2454 VDD.t4312 120.208
R2017 VDD.n2473 VDD.t3093 120.208
R2018 VDD.n2533 VDD.t3901 120.208
R2019 VDD.n2553 VDD.t4275 120.208
R2020 VDD.n2573 VDD.t4332 120.208
R2021 VDD.n2513 VDD.t3087 120.208
R2022 VDD.n2493 VDD.t3083 120.208
R2023 VDD.n2384 VDD.t2945 120.208
R2024 VDD.n2245 VDD.t2929 120.208
R2025 VDD.n2264 VDD.t2963 120.208
R2026 VDD.n2324 VDD.t2959 120.208
R2027 VDD.n2344 VDD.t869 120.208
R2028 VDD.n2364 VDD.t2941 120.208
R2029 VDD.n2304 VDD.t2917 120.208
R2030 VDD.n2284 VDD.t861 120.208
R2031 VDD.n2178 VDD.n2175 115.932
R2032 VDD.n2162 VDD.n2159 115.932
R2033 VDD.n1465 VDD.n1462 115.932
R2034 VDD.n2042 VDD.n2039 115.932
R2035 VDD.n1942 VDD.n1939 115.932
R2036 VDD.n1892 VDD.n1889 115.932
R2037 VDD.n1917 VDD.n1914 115.932
R2038 VDD.n1967 VDD.n1964 115.932
R2039 VDD.n1992 VDD.n1989 115.932
R2040 VDD.n2017 VDD.n2014 115.932
R2041 VDD.n2067 VDD.n2064 115.932
R2042 VDD.n2630 VDD.n2627 115.932
R2043 VDD.n2437 VDD.n2434 115.932
R2044 VDD.n2412 VDD.n2409 115.932
R2045 VDD.n2228 VDD.n2225 115.932
R2046 VDD.n2203 VDD.n2200 115.932
R2047 VDD.n2881 VDD.t4021 110.591
R2048 VDD.n2851 VDD.t2631 110.591
R2049 VDD.n2820 VDD.t2663 110.591
R2050 VDD.n554 VDD.t3477 110.591
R2051 VDD.n3100 VDD.t2989 110.591
R2052 VDD.n3124 VDD.t579 110.591
R2053 VDD.n3213 VDD.t659 110.591
R2054 VDD.n3237 VDD.t39 110.591
R2055 VDD.n3247 VDD.t3722 105.555
R2056 VDD.n2890 VDD.t3558 105.555
R2057 VDD.n2861 VDD.t4088 105.555
R2058 VDD.n2831 VDD.t1248 105.555
R2059 VDD.n541 VDD.t488 105.555
R2060 VDD.n3107 VDD.t4518 105.555
R2061 VDD.n3131 VDD.t906 105.555
R2062 VDD.n3225 VDD.t152 105.555
R2063 VDD.n2979 VDD.t3700 105.555
R2064 VDD.n2966 VDD.t2170 105.555
R2065 VDD.n3160 VDD.t154 105.555
R2066 VDD.n3142 VDD.t248 105.555
R2067 VDD.n3054 VDD.t918 105.555
R2068 VDD.n3042 VDD.t4290 105.555
R2069 VDD.n333 VDD.t4520 105.555
R2070 VDD.n317 VDD.t2817 105.555
R2071 VDD.n430 VDD.t494 105.555
R2072 VDD.n427 VDD.t1710 105.555
R2073 VDD.n496 VDD.t1230 105.555
R2074 VDD.n488 VDD.t89 105.555
R2075 VDD.n2781 VDD.t4100 105.555
R2076 VDD.n2778 VDD.t2065 105.555
R2077 VDD.n2718 VDD.t202 105.555
R2078 VDD.n2711 VDD.t1949 105.555
R2079 VDD.t4019 VDD.n2881 103.339
R2080 VDD.t2635 VDD.n2851 103.339
R2081 VDD.t2667 VDD.n2820 103.339
R2082 VDD.t3475 VDD.n554 103.339
R2083 VDD.t2993 VDD.n3100 103.339
R2084 VDD.t2733 VDD.n3124 103.339
R2085 VDD.t964 VDD.n3213 103.339
R2086 VDD.t409 VDD.n3237 103.339
R2087 VDD.n1049 VDD.n1048 85.695
R2088 VDD.n924 VDD.n923 85.695
R2089 VDD.n949 VDD.n948 85.695
R2090 VDD.n1024 VDD.n1023 85.695
R2091 VDD.n999 VDD.n998 85.695
R2092 VDD.n974 VDD.n973 85.695
R2093 VDD.n899 VDD.n898 85.695
R2094 VDD.n875 VDD.n874 85.695
R2095 VDD.t3368 VDD.t4198 77.958
R2096 VDD.t2883 VDD.t2779 77.958
R2097 VDD.t3641 VDD.t1127 77.958
R2098 VDD.t31 VDD.t1895 77.958
R2099 VDD.t2536 VDD.t324 77.958
R2100 VDD.t4194 VDD.t308 77.958
R2101 VDD.t2139 VDD.t306 77.958
R2102 VDD.t970 VDD.t3416 77.958
R2103 VDD.n1159 VDD.t4123 61.054
R2104 VDD.n1174 VDD.t1865 61.054
R2105 VDD.n1204 VDD.t1413 61.054
R2106 VDD.n1132 VDD.t4136 61.054
R2107 VDD.n1237 VDD.t2200 61.054
R2108 VDD.n1219 VDD.t2609 60.898
R2109 VDD.n1189 VDD.t1825 60.898
R2110 VDD.n1147 VDD.t3732 60.898
R2111 VDD.n1037 VDD.t3194 58.354
R2112 VDD.n912 VDD.t3264 58.354
R2113 VDD.n937 VDD.t3820 58.354
R2114 VDD.n1012 VDD.t3825 58.354
R2115 VDD.n987 VDD.t3865 58.354
R2116 VDD.n962 VDD.t2378 58.354
R2117 VDD.n887 VDD.t1735 58.354
R2118 VDD.n863 VDD.t3926 58.354
R2119 VDD.t972 VDD.t2251 53.244
R2120 VDD.t3224 VDD.t3611 53.244
R2121 VDD.t4024 VDD.t240 53.244
R2122 VDD.t2648 VDD.t2161 53.244
R2123 VDD.t786 VDD.t4288 53.244
R2124 VDD.t2591 VDD.t458 53.244
R2125 VDD.t3140 VDD.t2811 53.244
R2126 VDD.t887 VDD.t1859 53.244
R2127 VDD.t1773 VDD.t1708 53.244
R2128 VDD.t563 VDD.t2840 53.244
R2129 VDD.t109 VDD.t101 53.244
R2130 VDD.t4254 VDD.t1341 53.244
R2131 VDD.t2575 VDD.t4164 53.244
R2132 VDD.t4424 VDD.t3405 53.244
R2133 VDD.t2988 VDD.t1937 53.244
R2134 VDD.t1753 VDD.t2149 53.244
R2135 VDD.t3877 VDD.t4295 53.244
R2136 VDD.t1741 VDD.t3833 53.244
R2137 VDD.t3943 VDD.t200 53.244
R2138 VDD.t1440 VDD.t2259 53.244
R2139 VDD.t3961 VDD.t1043 53.244
R2140 VDD.t2316 VDD.t1421 53.244
R2141 VDD.t191 VDD.t3175 53.244
R2142 VDD.t3546 VDD.t1625 53.244
R2143 VDD.t282 VDD.t2861 53.244
R2144 VDD.t3430 VDD.t3059 53.244
R2145 VDD.t3744 VDD.t51 53.244
R2146 VDD.t1739 VDD.t1749 53.244
R2147 VDD.t3268 VDD.t533 53.244
R2148 VDD.t3252 VDD.t138 53.244
R2149 VDD.t3855 VDD.t1432 53.244
R2150 VDD.t1513 VDD.t2641 53.244
R2151 VDD.t1663 VDD.n2999 47.617
R2152 VDD.t2251 VDD.n3000 47.617
R2153 VDD.n3002 VDD.t3124 47.617
R2154 VDD.n3001 VDD.t3224 47.617
R2155 VDD.t234 VDD.n3187 47.617
R2156 VDD.t240 VDD.n3188 47.617
R2157 VDD.n3190 VDD.t2642 47.617
R2158 VDD.n3189 VDD.t2648 47.617
R2159 VDD.t1076 VDD.n3069 47.617
R2160 VDD.t4288 VDD.n3070 47.617
R2161 VDD.n3072 VDD.t2593 47.617
R2162 VDD.n3071 VDD.t2591 47.617
R2163 VDD.t3579 VDD.n351 47.617
R2164 VDD.t2811 VDD.n352 47.617
R2165 VDD.n354 VDD.t883 47.617
R2166 VDD.n353 VDD.t887 47.617
R2167 VDD.t1702 VDD.n450 47.617
R2168 VDD.t1708 VDD.n451 47.617
R2169 VDD.n453 VDD.t571 47.617
R2170 VDD.n452 VDD.t563 47.617
R2171 VDD.t95 VDD.n518 47.617
R2172 VDD.t101 VDD.n519 47.617
R2173 VDD.n521 VDD.t4256 47.617
R2174 VDD.n520 VDD.t4254 47.617
R2175 VDD.t4156 VDD.n2802 47.617
R2176 VDD.t4164 VDD.n2803 47.617
R2177 VDD.n2805 VDD.t4432 47.617
R2178 VDD.n2804 VDD.t4424 47.617
R2179 VDD.t1951 VDD.n2739 47.617
R2180 VDD.t1937 VDD.n2740 47.617
R2181 VDD.n2742 VDD.t3664 47.617
R2182 VDD.n2741 VDD.t1753 47.617
R2183 VDD.t4283 VDD.t4346 47.617
R2184 VDD.t4281 VDD.t950 47.617
R2185 VDD.t4282 VDD.t3702 47.617
R2186 VDD.t2882 VDD.t3706 47.617
R2187 VDD.t3222 VDD.t3718 47.617
R2188 VDD.t331 VDD.t3800 47.617
R2189 VDD.t332 VDD.t3591 47.617
R2190 VDD.t330 VDD.t160 47.617
R2191 VDD.t1861 VDD.t172 47.617
R2192 VDD.t1862 VDD.t156 47.617
R2193 VDD.t2669 VDD.t2268 47.617
R2194 VDD.t2518 VDD.t1616 47.617
R2195 VDD.t2519 VDD.t900 47.617
R2196 VDD.t3695 VDD.t910 47.617
R2197 VDD.t4422 VDD.t914 47.617
R2198 VDD.t227 VDD.t3412 47.617
R2199 VDD.t228 VDD.t3408 47.617
R2200 VDD.t229 VDD.t2402 47.617
R2201 VDD.t3653 VDD.t4528 47.617
R2202 VDD.t3654 VDD.t2398 47.617
R2203 VDD.t30 VDD.t1020 47.617
R2204 VDD.t28 VDD.t1024 47.617
R2205 VDD.t29 VDD.t1314 47.617
R2206 VDD.t2073 VDD.t4467 47.617
R2207 VDD.t2497 VDD.t490 47.617
R2208 VDD.t4472 VDD.t784 47.617
R2209 VDD.t4473 VDD.t973 47.617
R2210 VDD.t4471 VDD.t1236 47.617
R2211 VDD.t2138 VDD.t679 47.617
R2212 VDD.t2137 VDD.t1232 47.617
R2213 VDD.t1690 VDD.t1685 47.617
R2214 VDD.t3327 VDD.t1669 47.617
R2215 VDD.t1689 VDD.t4106 47.617
R2216 VDD.t1980 VDD.t4090 47.617
R2217 VDD.t1979 VDD.t4098 47.617
R2218 VDD.t4517 VDD.t2705 47.617
R2219 VDD.t4503 VDD.t179 47.617
R2220 VDD.t146 VDD.t206 47.617
R2221 VDD.t2836 VDD.t212 47.617
R2222 VDD.t1968 VDD.t3560 47.617
R2223 VDD.n2882 VDD.t4019 47.137
R2224 VDD.n2852 VDD.t2635 47.137
R2225 VDD.n2821 VDD.t2667 47.137
R2226 VDD.n555 VDD.t3475 47.137
R2227 VDD.n3101 VDD.t2993 47.137
R2228 VDD.n3125 VDD.t2733 47.137
R2229 VDD.n3214 VDD.t964 47.137
R2230 VDD.n3238 VDD.t409 47.137
R2231 VDD.n1141 VDD.n1140 47.107
R2232 VDD.n1126 VDD.n1125 47.107
R2233 VDD.t4233 VDD.t1611 45.992
R2234 VDD.t4223 VDD.t4173 45.992
R2235 VDD.t1327 VDD.t3491 45.992
R2236 VDD.t1326 VDD.t1111 45.992
R2237 VDD.t4574 VDD.t516 45.992
R2238 VDD.t4582 VDD.t514 45.992
R2239 VDD.t4051 VDD.t4455 45.992
R2240 VDD.t376 VDD.t4457 45.992
R2241 VDD.t1150 VDD.t2055 45.992
R2242 VDD.t1140 VDD.t2053 45.992
R2243 VDD.t1332 VDD.t476 45.992
R2244 VDD.t1333 VDD.t1056 45.992
R2245 VDD.t2562 VDD.t16 45.992
R2246 VDD.t2560 VDD.t15 45.992
R2247 VDD.t19 VDD.t3618 45.992
R2248 VDD.t18 VDD.t3616 45.992
R2249 VDD.n3000 VDD.t1663 44.495
R2250 VDD.t3228 VDD.n3002 44.495
R2251 VDD.t3124 VDD.n3001 44.495
R2252 VDD.n2999 VDD.t2176 44.495
R2253 VDD.n3188 VDD.t234 44.495
R2254 VDD.t4438 VDD.n3190 44.495
R2255 VDD.t2642 VDD.n3189 44.495
R2256 VDD.n3187 VDD.t250 44.495
R2257 VDD.n3070 VDD.t1076 44.495
R2258 VDD.t1532 VDD.n3072 44.495
R2259 VDD.t2593 VDD.n3071 44.495
R2260 VDD.n3069 VDD.t1068 44.495
R2261 VDD.n352 VDD.t3579 44.495
R2262 VDD.t891 VDD.n354 44.495
R2263 VDD.t883 VDD.n353 44.495
R2264 VDD.n351 VDD.t2815 44.495
R2265 VDD.n451 VDD.t1702 44.495
R2266 VDD.t567 VDD.n453 44.495
R2267 VDD.t571 VDD.n452 44.495
R2268 VDD.n450 VDD.t1640 44.495
R2269 VDD.n519 VDD.t95 44.495
R2270 VDD.t1501 VDD.n521 44.495
R2271 VDD.t4256 VDD.n520 44.495
R2272 VDD.n518 VDD.t85 44.495
R2273 VDD.n2803 VDD.t4156 44.495
R2274 VDD.t4428 VDD.n2805 44.495
R2275 VDD.t4432 VDD.n2804 44.495
R2276 VDD.n2802 VDD.t4170 44.495
R2277 VDD.n2740 VDD.t1951 44.495
R2278 VDD.t3660 VDD.n2742 44.495
R2279 VDD.t3664 VDD.n2741 44.495
R2280 VDD.n2739 VDD.t1945 44.495
R2281 VDD.t4338 VDD.t4283 44.494
R2282 VDD.t4346 VDD.t4281 44.494
R2283 VDD.t950 VDD.t4282 44.494
R2284 VDD.t3702 VDD.t2882 44.494
R2285 VDD.t3706 VDD.t3222 44.494
R2286 VDD.t3718 VDD.t3223 44.494
R2287 VDD.t512 VDD.t331 44.494
R2288 VDD.t3800 VDD.t332 44.494
R2289 VDD.t3591 VDD.t330 44.494
R2290 VDD.t160 VDD.t1861 44.494
R2291 VDD.t172 VDD.t1862 44.494
R2292 VDD.t156 VDD.t1860 44.494
R2293 VDD.t1620 VDD.t2669 44.494
R2294 VDD.t2268 VDD.t2518 44.494
R2295 VDD.t1616 VDD.t2519 44.494
R2296 VDD.t900 VDD.t3695 44.494
R2297 VDD.t910 VDD.t4422 44.494
R2298 VDD.t914 VDD.t4423 44.494
R2299 VDD.t1558 VDD.t227 44.494
R2300 VDD.t3412 VDD.t228 44.494
R2301 VDD.t3408 VDD.t229 44.494
R2302 VDD.t2402 VDD.t3653 44.494
R2303 VDD.t4528 VDD.t3654 44.494
R2304 VDD.t2398 VDD.t4151 44.494
R2305 VDD.t623 VDD.t30 44.494
R2306 VDD.t1020 VDD.t28 44.494
R2307 VDD.t1024 VDD.t29 44.494
R2308 VDD.t1314 VDD.t2073 44.494
R2309 VDD.t4467 VDD.t2497 44.494
R2310 VDD.t490 VDD.t2498 44.494
R2311 VDD.t778 VDD.t4472 44.494
R2312 VDD.t784 VDD.t4473 44.494
R2313 VDD.t973 VDD.t4471 44.494
R2314 VDD.t1236 VDD.t2138 44.494
R2315 VDD.t679 VDD.t2137 44.494
R2316 VDD.t1232 VDD.t2136 44.494
R2317 VDD.t1671 VDD.t1690 44.494
R2318 VDD.t1685 VDD.t3327 44.494
R2319 VDD.t1669 VDD.t1689 44.494
R2320 VDD.t4106 VDD.t1980 44.494
R2321 VDD.t4090 VDD.t1979 44.494
R2322 VDD.t4098 VDD.t1981 44.494
R2323 VDD.t181 VDD.t4517 44.494
R2324 VDD.t2705 VDD.t4503 44.494
R2325 VDD.t179 VDD.t146 44.494
R2326 VDD.t206 VDD.t2836 44.494
R2327 VDD.t212 VDD.t1968 44.494
R2328 VDD.t3560 VDD.t1969 44.494
R2329 VDD.n2173 VDD.t3877 44.17
R2330 VDD.n2174 VDD.t2036 44.17
R2331 VDD.t3724 VDD.n2177 44.17
R2332 VDD.t439 VDD.n2176 44.17
R2333 VDD.n2157 VDD.t1741 44.17
R2334 VDD.n2158 VDD.t2880 44.17
R2335 VDD.t2460 VDD.n2161 44.17
R2336 VDD.t4138 VDD.n2160 44.17
R2337 VDD.n1460 VDD.t3943 44.17
R2338 VDD.n1461 VDD.t1807 44.17
R2339 VDD.t2222 VDD.n1464 44.17
R2340 VDD.t2210 VDD.n1463 44.17
R2341 VDD.t3305 VDD.n2040 44.17
R2342 VDD.n2037 VDD.t1440 44.17
R2343 VDD.n2038 VDD.t1464 44.17
R2344 VDD.t3307 VDD.n2041 44.17
R2345 VDD.t1360 VDD.n1940 44.17
R2346 VDD.n1937 VDD.t3961 44.17
R2347 VDD.n1938 VDD.t3985 44.17
R2348 VDD.t437 VDD.n1941 44.17
R2349 VDD.t2216 VDD.n1890 44.17
R2350 VDD.n1887 VDD.t2316 44.17
R2351 VDD.n1888 VDD.t2326 44.17
R2352 VDD.t2208 VDD.n1891 44.17
R2353 VDD.t2466 VDD.n1915 44.17
R2354 VDD.n1912 VDD.t191 44.17
R2355 VDD.n1913 VDD.t1922 44.17
R2356 VDD.t2470 VDD.n1916 44.17
R2357 VDD.t4129 VDD.n1965 44.17
R2358 VDD.n1962 VDD.t3546 44.17
R2359 VDD.n1963 VDD.t4383 44.17
R2360 VDD.t2433 VDD.n1966 44.17
R2361 VDD.t922 VDD.n1990 44.17
R2362 VDD.n1987 VDD.t282 44.17
R2363 VDD.n1988 VDD.t2007 44.17
R2364 VDD.t936 VDD.n1991 44.17
R2365 VDD.t1819 VDD.n2015 44.17
R2366 VDD.n2012 VDD.t3430 44.17
R2367 VDD.n2013 VDD.t2095 44.17
R2368 VDD.t4110 VDD.n2016 44.17
R2369 VDD.t2617 VDD.n2065 44.17
R2370 VDD.n2062 VDD.t3744 44.17
R2371 VDD.n2063 VDD.t3757 44.17
R2372 VDD.t1550 VDD.n2066 44.17
R2373 VDD.n2625 VDD.t1739 44.17
R2374 VDD.n2626 VDD.t3853 44.17
R2375 VDD.t2599 VDD.n2629 44.17
R2376 VDD.t2613 VDD.n2628 44.17
R2377 VDD.n2432 VDD.t3268 44.17
R2378 VDD.n2433 VDD.t1731 44.17
R2379 VDD.t1399 VDD.n2436 44.17
R2380 VDD.t1409 VDD.n2435 44.17
R2381 VDD.n2407 VDD.t3252 44.17
R2382 VDD.n2408 VDD.t1777 44.17
R2383 VDD.t4112 VDD.n2411 44.17
R2384 VDD.t2412 VDD.n2410 44.17
R2385 VDD.n2223 VDD.t3855 44.17
R2386 VDD.n2224 VDD.t4005 44.17
R2387 VDD.t1863 VDD.n2227 44.17
R2388 VDD.t924 VDD.n2226 44.17
R2389 VDD.n2198 VDD.t1513 44.17
R2390 VDD.n2199 VDD.t1799 44.17
R2391 VDD.t2435 VDD.n2202 44.17
R2392 VDD.t2424 VDD.n2201 44.17
R2393 VDD.t1611 VDD.t4227 42.976
R2394 VDD.t4173 VDD.t4233 42.976
R2395 VDD.t4172 VDD.t4223 42.976
R2396 VDD.t3483 VDD.t1327 42.976
R2397 VDD.t3491 VDD.t1326 42.976
R2398 VDD.t1111 VDD.t3061 42.976
R2399 VDD.t516 VDD.t4568 42.976
R2400 VDD.t514 VDD.t4574 42.976
R2401 VDD.t515 VDD.t4582 42.976
R2402 VDD.t360 VDD.t4051 42.976
R2403 VDD.t4455 VDD.t376 42.976
R2404 VDD.t4457 VDD.t377 42.976
R2405 VDD.t2055 VDD.t1144 42.976
R2406 VDD.t2053 VDD.t1150 42.976
R2407 VDD.t2054 VDD.t1140 42.976
R2408 VDD.t468 VDD.t1332 42.976
R2409 VDD.t476 VDD.t1333 42.976
R2410 VDD.t1056 VDD.t1331 42.976
R2411 VDD.t16 VDD.t2564 42.976
R2412 VDD.t15 VDD.t2562 42.976
R2413 VDD.t2864 VDD.t2560 42.976
R2414 VDD.t3622 VDD.t19 42.976
R2415 VDD.t3618 VDD.t18 42.976
R2416 VDD.t3616 VDD.t17 42.976
R2417 VDD.t2036 VDD.n2173 41.273
R2418 VDD.t3802 VDD.n2174 41.273
R2419 VDD.n2177 VDD.t439 41.273
R2420 VDD.n2176 VDD.t433 41.273
R2421 VDD.t2880 VDD.n2157 41.273
R2422 VDD.t2384 VDD.n2158 41.273
R2423 VDD.n2161 VDD.t4138 41.273
R2424 VDD.n2160 VDD.t4142 41.273
R2425 VDD.t1807 VDD.n1460 41.273
R2426 VDD.t3922 VDD.n1461 41.273
R2427 VDD.n1464 VDD.t2210 41.273
R2428 VDD.n1463 VDD.t2196 41.273
R2429 VDD.t1464 VDD.n2037 41.273
R2430 VDD.t3035 VDD.n2038 41.273
R2431 VDD.n2041 VDD.t3305 41.273
R2432 VDD.n2040 VDD.t1395 41.273
R2433 VDD.t3985 VDD.n1937 41.273
R2434 VDD.t4025 VDD.n1938 41.273
R2435 VDD.n1941 VDD.t1360 41.273
R2436 VDD.n1940 VDD.t3726 41.273
R2437 VDD.t2326 VDD.n1887 41.273
R2438 VDD.t2305 VDD.n1888 41.273
R2439 VDD.n1891 VDD.t2216 41.273
R2440 VDD.n1890 VDD.t2204 41.273
R2441 VDD.t1922 VDD.n1912 41.273
R2442 VDD.t3391 VDD.n1913 41.273
R2443 VDD.n1916 VDD.t2466 41.273
R2444 VDD.n1915 VDD.t2474 41.273
R2445 VDD.t4383 VDD.n1962 41.273
R2446 VDD.t4375 VDD.n1963 41.273
R2447 VDD.n1966 VDD.t4129 41.273
R2448 VDD.n1965 VDD.t2651 41.273
R2449 VDD.t2007 VDD.n1987 41.273
R2450 VDD.t267 VDD.n1988 41.273
R2451 VDD.n1991 VDD.t922 41.273
R2452 VDD.n1990 VDD.t920 41.273
R2453 VDD.t2095 VDD.n2012 41.273
R2454 VDD.t3469 VDD.n2013 41.273
R2455 VDD.n2016 VDD.t1819 41.273
R2456 VDD.n2015 VDD.t2410 41.273
R2457 VDD.t3757 VDD.n2062 41.273
R2458 VDD.t3773 VDD.n2063 41.273
R2459 VDD.n2066 VDD.t2617 41.273
R2460 VDD.n2065 VDD.t1548 41.273
R2461 VDD.t3853 VDD.n2625 41.273
R2462 VDD.t3246 VDD.n2626 41.273
R2463 VDD.n2629 VDD.t2613 41.273
R2464 VDD.n2628 VDD.t1546 41.273
R2465 VDD.t1731 VDD.n2432 41.273
R2466 VDD.t3185 VDD.n2433 41.273
R2467 VDD.n2436 VDD.t1409 41.273
R2468 VDD.n2435 VDD.t3313 41.273
R2469 VDD.t1777 VDD.n2407 41.273
R2470 VDD.t3816 VDD.n2408 41.273
R2471 VDD.n2411 VDD.t2412 41.273
R2472 VDD.n2410 VDD.t1815 41.273
R2473 VDD.t4005 VDD.n2223 41.273
R2474 VDD.t1515 VDD.n2224 41.273
R2475 VDD.n2227 VDD.t924 41.273
R2476 VDD.n2226 VDD.t1871 41.273
R2477 VDD.t1799 VDD.n2198 41.273
R2478 VDD.t3248 VDD.n2199 41.273
R2479 VDD.n2202 VDD.t2424 41.273
R2480 VDD.n2201 VDD.t2659 41.273
R2481 VDD.n1168 VDD.n1167 41.219
R2482 VDD.n1213 VDD.n1212 41.219
R2483 VDD.n1198 VDD.n1197 39.256
R2484 VDD.n1183 VDD.n1182 39.256
R2485 VDD.n599 VDD.t3483 37.698
R2486 VDD.n585 VDD.t360 37.698
R2487 VDD.n263 VDD.t468 37.698
R2488 VDD.n729 VDD.t3622 37.698
R2489 VDD.n2145 VDD.t4055 30.726
R2490 VDD.n3258 VDD.t1999 30.238
R2491 VDD.n549 VDD.t1017 30.238
R2492 VDD.n409 VDD.t1382 30.238
R2493 VDD.n2926 VDD.t1830 30.238
R2494 VDD.n283 VDD.t4567 30.238
R2495 VDD.n272 VDD.t1149 30.238
R2496 VDD.n424 VDD.t620 30.238
R2497 VDD.n485 VDD.t781 30.238
R2498 VDD.n2775 VDD.t1678 30.238
R2499 VDD.n2708 VDD.t2704 30.238
R2500 VDD.n1077 VDD.t3969 30.238
R2501 VDD.n1085 VDD.t4403 30.238
R2502 VDD.n1118 VDD.t3753 30.238
R2503 VDD.n1110 VDD.t1452 30.238
R2504 VDD.n1101 VDD.t2081 30.238
R2505 VDD.n1093 VDD.t277 30.238
R2506 VDD.n1068 VDD.t2584 30.238
R2507 VDD.n1060 VDD.t2320 30.238
R2508 VDD.n3244 VDD.t4345 30.163
R2509 VDD.n2907 VDD.t2656 30.163
R2510 VDD.n2680 VDD.t3453 30.163
R2511 VDD.n2671 VDD.t2662 30.163
R2512 VDD.n2893 VDD.t184 30.163
R2513 VDD.n2858 VDD.t1666 30.163
R2514 VDD.n2827 VDD.t646 30.163
R2515 VDD.n2915 VDD.t1814 30.163
R2516 VDD.n310 VDD.t4401 30.163
R2517 VDD.n301 VDD.t2006 30.163
R2518 VDD.n392 VDD.t289 30.163
R2519 VDD.n401 VDD.t1402 30.163
R2520 VDD.n3110 VDD.t3411 30.163
R2521 VDD.n3134 VDD.t2267 30.163
R2522 VDD.n3222 VDD.t3594 30.163
R2523 VDD.n2982 VDD.t2173 30.163
R2524 VDD.n2973 VDD.t955 30.163
R2525 VDD.n3157 VDD.t253 30.163
R2526 VDD.n3145 VDD.t3793 30.163
R2527 VDD.n3051 VDD.t1073 30.163
R2528 VDD.n3039 VDD.t2261 30.163
R2529 VDD.n2661 VDD.t3435 30.163
R2530 VDD.n714 VDD.t3032 30.163
R2531 VDD.n2653 VDD.t1882 30.163
R2532 VDD.n706 VDD.t2427 30.163
R2533 VDD.n732 VDD.t4496 30.163
R2534 VDD.n608 VDD.t4232 30.163
R2535 VDD.n293 VDD.t927 30.163
R2536 VDD.n3270 VDD.t3740 30.163
R2537 VDD.n3327 VDD.t1444 30.163
R2538 VDD.n3384 VDD.t668 30.163
R2539 VDD.n193 VDD.t2016 30.163
R2540 VDD.n848 VDD.t2294 30.163
R2541 VDD.n828 VDD.t3261 30.163
R2542 VDD.n24 VDD.t3401 30.163
R2543 VDD.n823 VDD.t2307 30.163
R2544 VDD.n805 VDD.t3959 30.163
R2545 VDD.n134 VDD.t4394 30.163
R2546 VDD.n160 VDD.t1306 30.163
R2547 VDD.n152 VDD.t4399 30.163
R2548 VDD.n101 VDD.t995 30.163
R2549 VDD.n93 VDD.t3989 30.163
R2550 VDD.n50 VDD.t2573 30.163
R2551 VDD.n42 VDD.t3393 30.163
R2552 VDD.n3430 VDD.t3537 30.163
R2553 VDD.n3440 VDD.t3742 30.163
R2554 VDD.n3288 VDD.t3299 30.163
R2555 VDD.n3298 VDD.t3030 30.163
R2556 VDD.n3345 VDD.t2986 30.163
R2557 VDD.n3355 VDD.t3468 30.163
R2558 VDD.n221 VDD.t986 30.163
R2559 VDD.n231 VDD.t2002 30.163
R2560 VDD.n326 VDD.t2346 30.163
R2561 VDD.n314 VDD.t3500 30.163
R2562 VDD.n433 VDD.t1643 30.163
R2563 VDD.n493 VDD.t88 30.163
R2564 VDD.n2784 VDD.t4153 30.163
R2565 VDD.n2722 VDD.t1940 30.163
R2566 VDD.n2175 VDD.t1424 29.891
R2567 VDD.n2159 VDD.t2152 29.891
R2568 VDD.n1462 VDD.t3909 29.891
R2569 VDD.n2039 VDD.t135 29.891
R2570 VDD.n1939 VDD.t3386 29.891
R2571 VDD.n1889 VDD.t1480 29.891
R2572 VDD.n1914 VDD.t4447 29.891
R2573 VDD.n1964 VDD.t2121 29.891
R2574 VDD.n1989 VDD.t310 29.891
R2575 VDD.n2014 VDD.t2908 29.891
R2576 VDD.n2064 VDD.t3235 29.891
R2577 VDD.n2627 VDD.t4116 29.891
R2578 VDD.n2434 VDD.t42 29.891
R2579 VDD.n2409 VDD.t3670 29.891
R2580 VDD.n2225 VDD.t1133 29.891
R2581 VDD.n2200 VDD.t2516 29.891
R2582 VDD.n1155 VDD.t413 29.305
R2583 VDD.n1170 VDD.n1169 29.305
R2584 VDD.n1200 VDD.n1199 29.305
R2585 VDD.n1128 VDD.n1127 29.305
R2586 VDD.n1233 VDD.t2895 29.305
R2587 VDD.n1215 VDD.n1214 29.23
R2588 VDD.n1185 VDD.n1184 29.23
R2589 VDD.n1143 VDD.n1142 29.23
R2590 VDD.n2124 VDD.t3784 29.208
R2591 VDD.n2118 VDD.t1457 29.208
R2592 VDD.n2112 VDD.t2085 29.208
R2593 VDD.n2106 VDD.t262 29.208
R2594 VDD.n2100 VDD.t4391 29.208
R2595 VDD.n2082 VDD.t2324 29.208
R2596 VDD.n2094 VDD.t3992 29.202
R2597 VDD.n2088 VDD.t149 29.191
R2598 VDD.n3003 VDD.t972 28.957
R2599 VDD.n3191 VDD.t4024 28.957
R2600 VDD.n3073 VDD.t786 28.957
R2601 VDD.n355 VDD.t3140 28.957
R2602 VDD.n454 VDD.t1773 28.957
R2603 VDD.n522 VDD.t109 28.957
R2604 VDD.n2806 VDD.t2575 28.957
R2605 VDD.n2743 VDD.t2988 28.957
R2606 VDD.n2218 VDD.t1880 28.913
R2607 VDD.n2953 VDD.t3127 28.664
R2608 VDD.n2958 VDD.t1662 28.664
R2609 VDD.n2988 VDD.t3709 28.664
R2610 VDD.n2993 VDD.t4349 28.664
R2611 VDD.n3177 VDD.t2645 28.664
R2612 VDD.n3182 VDD.t245 28.664
R2613 VDD.n3164 VDD.t167 28.664
R2614 VDD.n3169 VDD.t3795 28.664
R2615 VDD.n3077 VDD.t1535 28.664
R2616 VDD.n3082 VDD.t4285 28.664
R2617 VDD.n3058 VDD.t903 28.664
R2618 VDD.n3063 VDD.t2273 28.664
R2619 VDD.n724 VDD.t2488 28.664
R2620 VDD.n719 VDD.t2559 28.664
R2621 VDD.n594 VDD.t3486 28.664
R2622 VDD.n589 VDD.t2874 28.664
R2623 VDD.n580 VDD.t363 28.664
R2624 VDD.n575 VDD.t4577 28.664
R2625 VDD.n258 VDD.t471 28.664
R2626 VDD.n253 VDD.t1155 28.664
R2627 VDD.n180 VDD.t3139 28.664
R2628 VDD.n185 VDD.t1309 28.664
R2629 VDD.n168 VDD.t759 28.664
R2630 VDD.n173 VDD.t4398 28.664
R2631 VDD.n121 VDD.t879 28.664
R2632 VDD.n126 VDD.t994 28.664
R2633 VDD.n109 VDD.t1916 28.664
R2634 VDD.n114 VDD.t3988 28.664
R2635 VDD.n835 VDD.t1492 28.664
R2636 VDD.n840 VDD.t2299 28.664
R2637 VDD.n11 VDD.t525 28.664
R2638 VDD.n16 VDD.t3804 28.664
R2639 VDD.n70 VDD.t4082 28.664
R2640 VDD.n75 VDD.t2571 28.664
R2641 VDD.n58 VDD.t2590 28.664
R2642 VDD.n63 VDD.t1925 28.664
R2643 VDD.n3423 VDD.t3813 28.664
R2644 VDD.n3418 VDD.t3769 28.664
R2645 VDD.n3412 VDD.t1265 28.664
R2646 VDD.n3407 VDD.t3541 28.664
R2647 VDD.n3281 VDD.t1461 28.664
R2648 VDD.n3276 VDD.t3106 28.664
R2649 VDD.n3309 VDD.t3293 28.664
R2650 VDD.n3304 VDD.t4509 28.664
R2651 VDD.n3338 VDD.t3445 28.664
R2652 VDD.n3333 VDD.t77 28.664
R2653 VDD.n3366 VDD.t2987 28.664
R2654 VDD.n3361 VDD.t1374 28.664
R2655 VDD.n214 VDD.t1996 28.664
R2656 VDD.n209 VDD.t2509 28.664
R2657 VDD.n242 VDD.t982 28.664
R2658 VDD.n237 VDD.t4560 28.664
R2659 VDD.n358 VDD.t886 28.664
R2660 VDD.n363 VDD.t2810 28.664
R2661 VDD.n340 VDD.t4531 28.664
R2662 VDD.n345 VDD.t2543 28.664
R2663 VDD.n458 VDD.t574 28.664
R2664 VDD.n463 VDD.t1707 28.664
R2665 VDD.n439 VDD.t4470 28.664
R2666 VDD.n444 VDD.t618 28.664
R2667 VDD.n470 VDD.t4262 28.664
R2668 VDD.n475 VDD.t92 28.664
R2669 VDD.n507 VDD.t1245 28.664
R2670 VDD.n512 VDD.t783 28.664
R2671 VDD.n2757 VDD.t4431 28.664
R2672 VDD.n2762 VDD.t2064 28.664
R2673 VDD.n2791 VDD.t4093 28.664
R2674 VDD.n2796 VDD.t1680 28.664
R2675 VDD.n2693 VDD.t3667 28.664
R2676 VDD.n2698 VDD.t552 28.664
R2677 VDD.n2728 VDD.t215 28.664
R2678 VDD.n2733 VDD.t2708 28.664
R2679 VDD.n2182 VDD.t2041 28.664
R2680 VDD.n2168 VDD.t430 28.664
R2681 VDD.n2150 VDD.t2459 28.664
R2682 VDD.n1469 VDD.t1512 28.664
R2683 VDD.n1455 VDD.t2221 28.664
R2684 VDD.n2030 VDD.t3310 28.664
R2685 VDD.n2045 VDD.t1463 28.664
R2686 VDD.n1930 VDD.t432 28.664
R2687 VDD.n1945 VDD.t3982 28.664
R2688 VDD.n1880 VDD.t2213 28.664
R2689 VDD.n1895 VDD.t2330 28.664
R2690 VDD.n1905 VDD.t2473 28.664
R2691 VDD.n1920 VDD.t1933 28.664
R2692 VDD.n1955 VDD.t2419 28.664
R2693 VDD.n1970 VDD.t4389 28.664
R2694 VDD.n1980 VDD.t941 28.664
R2695 VDD.n1995 VDD.t2004 28.664
R2696 VDD.n2005 VDD.t4115 28.664
R2697 VDD.n2020 VDD.t2077 28.664
R2698 VDD.n2055 VDD.t2608 28.664
R2699 VDD.n2070 VDD.t3756 28.664
R2700 VDD.n2618 VDD.t2612 28.664
R2701 VDD.n2613 VDD.t4010 28.664
R2702 VDD.n2441 VDD.t3819 28.664
R2703 VDD.n2427 VDD.t1388 28.664
R2704 VDD.n2416 VDD.t3209 28.664
R2705 VDD.n2402 VDD.t1824 28.664
R2706 VDD.n2232 VDD.t104 28.664
R2707 VDD.n2207 VDD.t1797 28.664
R2708 VDD.n2193 VDD.t2654 28.664
R2709 VDD.n2687 VDD.t3119 28.57
R2710 VDD.n2868 VDD.t4177 28.57
R2711 VDD.n2752 VDD.t3145 28.57
R2712 VDD.n2840 VDD.t2886 28.57
R2713 VDD.n2815 VDD.t3162 28.57
R2714 VDD.n529 VDD.t3638 28.57
R2715 VDD.n558 VDD.t2100 28.57
R2716 VDD.n565 VDD.t4590 28.57
R2717 VDD.n3093 VDD.t2549 28.57
R2718 VDD.n375 VDD.t3536 28.57
R2719 VDD.n3022 VDD.t1631 28.57
R2720 VDD.n3029 VDD.t4253 28.57
R2721 VDD.n3206 VDD.t1085 28.57
R2722 VDD.n2941 VDD.t426 28.57
R2723 VDD.n2947 VDD.t2630 28.57
R2724 VDD.n3012 VDD.t969 28.57
R2725 VDD.n3374 VDD.t396 28.57
R2726 VDD.n3379 VDD.t2742 28.57
R2727 VDD.n3322 VDD.t3632 28.57
R2728 VDD.n3317 VDD.t1106 28.57
R2729 VDD.n200 VDD.t1032 28.57
R2730 VDD.n205 VDD.t1747 28.57
R2731 VDD.n3265 VDD.t1920 28.57
R2732 VDD.n32 VDD.t418 28.57
R2733 VDD.n37 VDD.t2522 28.57
R2734 VDD.n2 VDD.t1435 28.57
R2735 VDD.n7 VDD.t346 28.57
R2736 VDD.n88 VDD.t1350 28.57
R2737 VDD.n83 VDD.t3051 28.57
R2738 VDD.n142 VDD.t959 28.57
R2739 VDD.n147 VDD.t1573 28.57
R2740 VDD.n3401 VDD.t614 28.57
R2741 VDD.n1163 VDD.t412 28.57
R2742 VDD.n1178 VDD.t10 28.57
R2743 VDD.n1223 VDD.t4299 28.57
R2744 VDD.n1208 VDD.t301 28.57
R2745 VDD.n1193 VDD.t3381 28.57
R2746 VDD.n1151 VDD.t3507 28.57
R2747 VDD.n1136 VDD.t640 28.57
R2748 VDD.n1241 VDD.t3239 28.57
R2749 VDD.n1043 VDD.t597 28.568
R2750 VDD.n918 VDD.t1264 28.568
R2751 VDD.n943 VDD.t2481 28.568
R2752 VDD.n1018 VDD.t2146 28.568
R2753 VDD.n993 VDD.t2154 28.568
R2754 VDD.n968 VDD.t676 28.568
R2755 VDD.n893 VDD.t79 28.568
R2756 VDD.n869 VDD.t947 28.568
R2757 VDD.n639 VDD.t2757 28.568
R2758 VDD.n657 VDD.t1900 28.568
R2759 VDD.n675 VDD.t2894 28.568
R2760 VDD.n692 VDD.t2342 28.568
R2761 VDD.n621 VDD.t3042 28.568
R2762 VDD.n752 VDD.t1038 28.568
R2763 VDD.n770 VDD.t3324 28.568
R2764 VDD.n788 VDD.t1761 28.568
R2765 VDD.n1744 VDD.t2803 28.568
R2766 VDD.n1769 VDD.t3571 28.568
R2767 VDD.n1862 VDD.t2844 28.568
R2768 VDD.n1837 VDD.t352 28.568
R2769 VDD.n1819 VDD.t1721 28.568
R2770 VDD.n1794 VDD.t2681 28.568
R2771 VDD.n1719 VDD.t1281 28.568
R2772 VDD.n1695 VDD.t2344 28.568
R2773 VDD.n1537 VDD.t3329 28.568
R2774 VDD.n1562 VDD.t2762 28.568
R2775 VDD.n1662 VDD.t1159 28.568
R2776 VDD.n1637 VDD.t4222 28.568
R2777 VDD.n1612 VDD.t399 28.568
R2778 VDD.n1587 VDD.t483 28.568
R2779 VDD.n1512 VDD.t2693 28.568
R2780 VDD.n1488 VDD.t1595 28.568
R2781 VDD.n1387 VDD.t2313 28.568
R2782 VDD.n1362 VDD.t519 28.568
R2783 VDD.n1263 VDD.t4244 28.568
R2784 VDD.n1287 VDD.t375 28.568
R2785 VDD.n1312 VDD.t638 28.568
R2786 VDD.n1337 VDD.t313 28.568
R2787 VDD.n1412 VDD.t3936 28.568
R2788 VDD.n1437 VDD.t2490 28.568
R2789 VDD.n2605 VDD.t4212 28.568
R2790 VDD.n2466 VDD.t1537 28.568
R2791 VDD.n2485 VDD.t1302 28.568
R2792 VDD.n2545 VDD.t4182 28.568
R2793 VDD.n2565 VDD.t1971 28.568
R2794 VDD.n2585 VDD.t2 28.568
R2795 VDD.n2525 VDD.t875 28.568
R2796 VDD.n2505 VDD.t3182 28.568
R2797 VDD.n2389 VDD.t2545 28.568
R2798 VDD.n2257 VDD.t1579 28.568
R2799 VDD.n2276 VDD.t2131 28.568
R2800 VDD.n2329 VDD.t1854 28.568
R2801 VDD.n2349 VDD.t1555 28.568
R2802 VDD.n2369 VDD.t3044 28.568
R2803 VDD.n2316 VDD.t2555 28.568
R2804 VDD.n2296 VDD.t2689 28.568
R2805 VDD.n1045 VDD.t2371 28.565
R2806 VDD.n1045 VDD.t3215 28.565
R2807 VDD.n1048 VDD.t3203 28.565
R2808 VDD.n1042 VDD.t595 28.565
R2809 VDD.n1042 VDD.t593 28.565
R2810 VDD.n920 VDD.t2049 28.565
R2811 VDD.n920 VDD.t3921 28.565
R2812 VDD.n923 VDD.t1806 28.565
R2813 VDD.n917 VDD.t1262 28.565
R2814 VDD.n917 VDD.t1260 28.565
R2815 VDD.n945 VDD.t4053 28.565
R2816 VDD.n945 VDD.t3180 28.565
R2817 VDD.n948 VDD.t3678 28.565
R2818 VDD.n942 VDD.t2485 28.565
R2819 VDD.n942 VDD.t2483 28.565
R2820 VDD.n1020 VDD.t3832 28.565
R2821 VDD.n1020 VDD.t3207 28.565
R2822 VDD.n1023 VDD.t3199 28.565
R2823 VDD.n1017 VDD.t2144 28.565
R2824 VDD.n1017 VDD.t2148 28.565
R2825 VDD.n995 VDD.t3263 28.565
R2826 VDD.n995 VDD.t2039 28.565
R2827 VDD.n998 VDD.t3946 28.565
R2828 VDD.n992 VDD.t2158 28.565
R2829 VDD.n992 VDD.t2156 28.565
R2830 VDD.n970 VDD.t3217 28.565
R2831 VDD.n970 VDD.t3205 28.565
R2832 VDD.n973 VDD.t4000 28.565
R2833 VDD.n967 VDD.t674 28.565
R2834 VDD.n967 VDD.t672 28.565
R2835 VDD.n895 VDD.t3938 28.565
R2836 VDD.n895 VDD.t1599 28.565
R2837 VDD.n898 VDD.t4535 28.565
R2838 VDD.n892 VDD.t3658 28.565
R2839 VDD.n892 VDD.t3656 28.565
R2840 VDD.n871 VDD.t1784 28.565
R2841 VDD.n871 VDD.t2879 28.565
R2842 VDD.n874 VDD.t1011 28.565
R2843 VDD.n868 VDD.t945 28.565
R2844 VDD.n868 VDD.t943 28.565
R2845 VDD.n3243 VDD.t953 28.565
R2846 VDD.n3243 VDD.t4337 28.565
R2847 VDD.n2936 VDD.t3342 28.565
R2848 VDD.n2936 VDD.t3344 28.565
R2849 VDD.n2937 VDD.t3340 28.565
R2850 VDD.n2937 VDD.t3713 28.565
R2851 VDD.n3242 VDD.t3723 28.565
R2852 VDD.n3242 VDD.t3711 28.565
R2853 VDD.n3257 VDD.t2013 28.565
R2854 VDD.n3257 VDD.t291 28.565
R2855 VDD.n3252 VDD.t1649 28.565
R2856 VDD.n3252 VDD.t1645 28.565
R2857 VDD.n3253 VDD.t4352 28.565
R2858 VDD.n3253 VDD.t1651 28.565
R2859 VDD.n3254 VDD.t4356 28.565
R2860 VDD.n3254 VDD.t4354 28.565
R2861 VDD.n2906 VDD.t2438 28.565
R2862 VDD.n2906 VDD.t1908 28.565
R2863 VDD.n2901 VDD.t2736 28.565
R2864 VDD.n2901 VDD.t1983 28.565
R2865 VDD.n2902 VDD.t1985 28.565
R2866 VDD.n2902 VDD.t3025 28.565
R2867 VDD.n2904 VDD.t1455 28.565
R2868 VDD.n2904 VDD.t3014 28.565
R2869 VDD.n2679 VDD.t2088 28.565
R2870 VDD.n2679 VDD.t3457 28.565
R2871 VDD.n2674 VDD.t1570 28.565
R2872 VDD.n2674 VDD.t1575 28.565
R2873 VDD.n2675 VDD.t1568 28.565
R2874 VDD.n2675 VDD.t1878 28.565
R2875 VDD.n2677 VDD.t935 28.565
R2876 VDD.n2677 VDD.t1874 28.565
R2877 VDD.n2670 VDD.t1910 28.565
R2878 VDD.n2670 VDD.t2421 28.565
R2879 VDD.n2665 VDD.t2796 28.565
R2880 VDD.n2665 VDD.t2798 28.565
R2881 VDD.n2666 VDD.t2794 28.565
R2882 VDD.n2666 VDD.t2093 28.565
R2883 VDD.n2668 VDD.t3466 28.565
R2884 VDD.n2668 VDD.t2083 28.565
R2885 VDD.n2686 VDD.t3121 28.565
R2886 VDD.n2686 VDD.t3117 28.565
R2887 VDD.n2867 VDD.t3369 28.565
R2888 VDD.n2867 VDD.t4175 28.565
R2889 VDD.n2892 VDD.t178 28.565
R2890 VDD.n2892 VDD.t2714 28.565
R2891 VDD.n2682 VDD.t4557 28.565
R2892 VDD.n2682 VDD.t4553 28.565
R2893 VDD.n2683 VDD.t4555 28.565
R2894 VDD.n2683 VDD.t209 28.565
R2895 VDD.n2891 VDD.t3559 28.565
R2896 VDD.n2891 VDD.t205 28.565
R2897 VDD.n2751 VDD.t3147 28.565
R2898 VDD.n2751 VDD.t3149 28.565
R2899 VDD.n2839 VDD.t2884 28.565
R2900 VDD.n2839 VDD.t2888 28.565
R2901 VDD.n2857 VDD.t1668 28.565
R2902 VDD.n2857 VDD.t1676 28.565
R2903 VDD.n2747 VDD.t2854 28.565
R2904 VDD.n2747 VDD.t2852 28.565
R2905 VDD.n2748 VDD.t2856 28.565
R2906 VDD.n2748 VDD.t4103 28.565
R2907 VDD.n2856 VDD.t4089 28.565
R2908 VDD.n2856 VDD.t4095 28.565
R2909 VDD.n2814 VDD.t14 28.565
R2910 VDD.n2814 VDD.t3164 28.565
R2911 VDD.n528 VDD.t3642 28.565
R2912 VDD.n528 VDD.t3640 28.565
R2913 VDD.n2826 VDD.t648 28.565
R2914 VDD.n2826 VDD.t771 28.565
R2915 VDD.n2810 VDD.t2190 28.565
R2916 VDD.n2810 VDD.t2192 28.565
R2917 VDD.n2811 VDD.t2188 28.565
R2918 VDD.n2811 VDD.t1243 28.565
R2919 VDD.n2825 VDD.t1249 28.565
R2920 VDD.n2825 VDD.t1239 28.565
R2921 VDD.n548 VDD.t1019 28.565
R2922 VDD.n548 VDD.t626 28.565
R2923 VDD.n547 VDD.t489 28.565
R2924 VDD.n547 VDD.t1313 28.565
R2925 VDD.n544 VDD.t1430 28.565
R2926 VDD.n544 VDD.t4464 28.565
R2927 VDD.n545 VDD.t1428 28.565
R2928 VDD.n545 VDD.t1426 28.565
R2929 VDD.n557 VDD.t4511 28.565
R2930 VDD.n557 VDD.t4513 28.565
R2931 VDD.n564 VDD.t32 28.565
R2932 VDD.n564 VDD.t4588 28.565
R2933 VDD.n2914 VDD.t1844 28.565
R2934 VDD.n2914 VDD.t1838 28.565
R2935 VDD.n2909 VDD.t2356 28.565
R2936 VDD.n2909 VDD.t2354 28.565
R2937 VDD.n2910 VDD.t2352 28.565
R2938 VDD.n2910 VDD.t2024 28.565
R2939 VDD.n2912 VDD.t2020 28.565
R2940 VDD.n2912 VDD.t2018 28.565
R2941 VDD.n405 VDD.t3006 28.565
R2942 VDD.n405 VDD.t3004 28.565
R2943 VDD.n404 VDD.t3002 28.565
R2944 VDD.n404 VDD.t3455 28.565
R2945 VDD.n403 VDD.t3451 28.565
R2946 VDD.n403 VDD.t3447 28.565
R2947 VDD.n408 VDD.t1378 28.565
R2948 VDD.n408 VDD.t1384 28.565
R2949 VDD.n2922 VDD.t422 28.565
R2950 VDD.n2922 VDD.t4441 28.565
R2951 VDD.n2921 VDD.t420 28.565
R2952 VDD.n2921 VDD.t1475 28.565
R2953 VDD.n2920 VDD.t1473 28.565
R2954 VDD.n2920 VDD.t1470 28.565
R2955 VDD.n2925 VDD.t1840 28.565
R2956 VDD.n2925 VDD.t1834 28.565
R2957 VDD.n309 VDD.t4397 28.565
R2958 VDD.n309 VDD.t4378 28.565
R2959 VDD.n304 VDD.t2072 28.565
R2960 VDD.n304 VDD.t2068 28.565
R2961 VDD.n305 VDD.t2070 28.565
R2962 VDD.n305 VDD.t2409 28.565
R2963 VDD.n307 VDD.t1852 28.565
R2964 VDD.n307 VDD.t1812 28.565
R2965 VDD.n300 VDD.t2011 28.565
R2966 VDD.n300 VDD.t275 28.565
R2967 VDD.n295 VDD.t1277 28.565
R2968 VDD.n295 VDD.t1273 28.565
R2969 VDD.n296 VDD.t1275 28.565
R2970 VDD.n296 VDD.t4122 28.565
R2971 VDD.n298 VDD.t4120 28.565
R2972 VDD.n298 VDD.t2423 28.565
R2973 VDD.n391 VDD.t2015 28.565
R2974 VDD.n391 VDD.t2027 28.565
R2975 VDD.n386 VDD.t1793 28.565
R2976 VDD.n386 VDD.t1795 28.565
R2977 VDD.n387 VDD.t1791 28.565
R2978 VDD.n387 VDD.t1408 28.565
R2979 VDD.n389 VDD.t3312 28.565
R2980 VDD.n389 VDD.t1380 28.565
R2981 VDD.n400 VDD.t1420 28.565
R2982 VDD.n400 VDD.t1404 28.565
R2983 VDD.n395 VDD.t124 28.565
R2984 VDD.n395 VDD.t4239 28.565
R2985 VDD.n396 VDD.t126 28.565
R2986 VDD.n396 VDD.t3549 28.565
R2987 VDD.n398 VDD.t3551 28.565
R2988 VDD.n398 VDD.t4410 28.565
R2989 VDD.n3092 VDD.t2551 28.565
R2990 VDD.n3092 VDD.t2547 28.565
R2991 VDD.n374 VDD.t2537 28.565
R2992 VDD.n374 VDD.t2539 28.565
R2993 VDD.n3109 VDD.t1561 28.565
R2994 VDD.n3109 VDD.t3496 28.565
R2995 VDD.n3088 VDD.t546 28.565
R2996 VDD.n3088 VDD.t542 28.565
R2997 VDD.n3089 VDD.t544 28.565
R2998 VDD.n3089 VDD.t4260 28.565
R2999 VDD.n3108 VDD.t4519 28.565
R3000 VDD.n3108 VDD.t4525 28.565
R3001 VDD.n3021 VDD.t1629 28.565
R3002 VDD.n3021 VDD.t1627 28.565
R3003 VDD.n3028 VDD.t4195 28.565
R3004 VDD.n3028 VDD.t4251 28.565
R3005 VDD.n3133 VDD.t2275 28.565
R3006 VDD.n3133 VDD.t1619 28.565
R3007 VDD.n3017 VDD.t1347 28.565
R3008 VDD.n3017 VDD.t1343 28.565
R3009 VDD.n3018 VDD.t1345 28.565
R3010 VDD.n3018 VDD.t2167 28.565
R3011 VDD.n3132 VDD.t907 28.565
R3012 VDD.n3132 VDD.t917 28.565
R3013 VDD.n3205 VDD.t1756 28.565
R3014 VDD.n3205 VDD.t1083 28.565
R3015 VDD.n3221 VDD.t3590 28.565
R3016 VDD.n3221 VDD.t511 28.565
R3017 VDD.n3007 VDD.t2823 28.565
R3018 VDD.n3007 VDD.t2866 28.565
R3019 VDD.n3008 VDD.t2821 28.565
R3020 VDD.n3008 VDD.t169 28.565
R3021 VDD.n3220 VDD.t153 28.565
R3022 VDD.n3220 VDD.t163 28.565
R3023 VDD.n2940 VDD.t428 28.565
R3024 VDD.n2940 VDD.t424 28.565
R3025 VDD.n2946 VDD.t2140 28.565
R3026 VDD.n2946 VDD.t2142 28.565
R3027 VDD.n2954 VDD.t3227 28.565
R3028 VDD.n2954 VDD.t3123 28.565
R3029 VDD.n2959 VDD.t2250 28.565
R3030 VDD.n2959 VDD.t2175 28.565
R3031 VDD.n2989 VDD.t3721 28.565
R3032 VDD.n2989 VDD.t3705 28.565
R3033 VDD.n2994 VDD.t949 28.565
R3034 VDD.n2994 VDD.t4335 28.565
R3035 VDD.n2981 VDD.t61 28.565
R3036 VDD.n2981 VDD.t59 28.565
R3037 VDD.n2963 VDD.t2906 28.565
R3038 VDD.n2963 VDD.t2902 28.565
R3039 VDD.n2964 VDD.t2904 28.565
R3040 VDD.n2964 VDD.t3717 28.565
R3041 VDD.n2980 VDD.t3701 28.565
R3042 VDD.n2980 VDD.t3715 28.565
R3043 VDD.n2972 VDD.t4343 28.565
R3044 VDD.n2972 VDD.t4341 28.565
R3045 VDD.n2967 VDD.t2165 28.565
R3046 VDD.n2967 VDD.t2108 28.565
R3047 VDD.n2968 VDD.t2163 28.565
R3048 VDD.n2968 VDD.t57 28.565
R3049 VDD.n2971 VDD.t2171 28.565
R3050 VDD.n2971 VDD.t2179 28.565
R3051 VDD.n3011 VDD.t971 28.565
R3052 VDD.n3011 VDD.t967 28.565
R3053 VDD.n3178 VDD.t2647 28.565
R3054 VDD.n3178 VDD.t4437 28.565
R3055 VDD.n3183 VDD.t247 28.565
R3056 VDD.n3183 VDD.t231 28.565
R3057 VDD.n3165 VDD.t72 28.565
R3058 VDD.n3165 VDD.t159 28.565
R3059 VDD.n3170 VDD.t509 28.565
R3060 VDD.n3170 VDD.t3799 28.565
R3061 VDD.n3156 VDD.t237 28.565
R3062 VDD.n3156 VDD.t243 28.565
R3063 VDD.n3139 VDD.t2835 28.565
R3064 VDD.n3139 VDD.t2831 28.565
R3065 VDD.n3140 VDD.t2833 28.565
R3066 VDD.n3140 VDD.t171 28.565
R3067 VDD.n3155 VDD.t155 28.565
R3068 VDD.n3155 VDD.t165 28.565
R3069 VDD.n3144 VDD.t3797 28.565
R3070 VDD.n3144 VDD.t3588 28.565
R3071 VDD.n3149 VDD.t1254 28.565
R3072 VDD.n3149 VDD.t1256 28.565
R3073 VDD.n3150 VDD.t1258 28.565
R3074 VDD.n3150 VDD.t239 28.565
R3075 VDD.n3143 VDD.t249 28.565
R3076 VDD.n3143 VDD.t233 28.565
R3077 VDD.n3078 VDD.t2596 28.565
R3078 VDD.n3078 VDD.t1531 28.565
R3079 VDD.n3083 VDD.t4287 28.565
R3080 VDD.n3083 VDD.t1075 28.565
R3081 VDD.n3059 VDD.t913 28.565
R3082 VDD.n3059 VDD.t2169 28.565
R3083 VDD.n3064 VDD.t2265 28.565
R3084 VDD.n3064 VDD.t2263 28.565
R3085 VDD.n3050 VDD.t1081 28.565
R3086 VDD.n3050 VDD.t1067 28.565
R3087 VDD.n3034 VDD.t1288 28.565
R3088 VDD.n3034 VDD.t1290 28.565
R3089 VDD.n3035 VDD.t1286 28.565
R3090 VDD.n3035 VDD.t909 28.565
R3091 VDD.n3049 VDD.t919 28.565
R3092 VDD.n3049 VDD.t905 28.565
R3093 VDD.n3038 VDD.t2271 28.565
R3094 VDD.n3038 VDD.t2277 28.565
R3095 VDD.n3043 VDD.t3502 28.565
R3096 VDD.n3043 VDD.t4547 28.565
R3097 VDD.n3044 VDD.t4549 28.565
R3098 VDD.n3044 VDD.t1079 28.565
R3099 VDD.n3037 VDD.t4291 28.565
R3100 VDD.n3037 VDD.t1071 28.565
R3101 VDD.n2660 VDD.t2090 28.565
R3102 VDD.n2660 VDD.t3439 28.565
R3103 VDD.n2655 VDD.t344 28.565
R3104 VDD.n2655 VDD.t4446 28.565
R3105 VDD.n2656 VDD.t4444 28.565
R3106 VDD.n2656 VDD.t1850 28.565
R3107 VDD.n2658 VDD.t1846 28.565
R3108 VDD.n2658 VDD.t1842 28.565
R3109 VDD.n713 VDD.t3027 28.565
R3110 VDD.n713 VDD.t3034 28.565
R3111 VDD.n708 VDD.t2098 28.565
R3112 VDD.n708 VDD.t2288 28.565
R3113 VDD.n709 VDD.t3160 28.565
R3114 VDD.n709 VDD.t3316 28.565
R3115 VDD.n711 VDD.t1398 28.565
R3116 VDD.n711 VDD.t1394 28.565
R3117 VDD.n2652 VDD.t1647 28.565
R3118 VDD.n2652 VDD.t1890 28.565
R3119 VDD.n2647 VDD.t8 28.565
R3120 VDD.n2647 VDD.t114 28.565
R3121 VDD.n2648 VDD.t112 28.565
R3122 VDD.n2648 VDD.t1443 28.565
R3123 VDD.n2650 VDD.t3012 28.565
R3124 VDD.n2650 VDD.t1477 28.565
R3125 VDD.n705 VDD.t3067 28.565
R3126 VDD.n705 VDD.t2429 28.565
R3127 VDD.n700 VDD.t2114 28.565
R3128 VDD.n700 VDD.t2112 28.565
R3129 VDD.n701 VDD.t2116 28.565
R3130 VDD.n701 VDD.t3545 28.565
R3131 VDD.n703 VDD.t1319 28.565
R3132 VDD.n703 VDD.t1323 28.565
R3133 VDD.n725 VDD.t3631 28.565
R3134 VDD.n725 VDD.t3621 28.565
R3135 VDD.n720 VDD.t4502 28.565
R3136 VDD.n720 VDD.t4500 28.565
R3137 VDD.n731 VDD.t2557 28.565
R3138 VDD.n731 VDD.t4498 28.565
R3139 VDD.n733 VDD.t535 28.565
R3140 VDD.n733 VDD.t4545 28.565
R3141 VDD.n734 VDD.t4543 28.565
R3142 VDD.n734 VDD.t3629 28.565
R3143 VDD.n736 VDD.t3627 28.565
R3144 VDD.n736 VDD.t3625 28.565
R3145 VDD.n638 VDD.t2755 28.565
R3146 VDD.n638 VDD.t2753 28.565
R3147 VDD.n630 VDD.t796 28.565
R3148 VDD.n629 VDD.t1179 28.565
R3149 VDD.n629 VDD.t830 28.565
R3150 VDD.n656 VDD.t1904 28.565
R3151 VDD.n656 VDD.t1902 28.565
R3152 VDD.n648 VDD.t1187 28.565
R3153 VDD.n647 VDD.t682 28.565
R3154 VDD.n647 VDD.t806 28.565
R3155 VDD.n674 VDD.t2892 28.565
R3156 VDD.n674 VDD.t2890 28.565
R3157 VDD.n666 VDD.t724 28.565
R3158 VDD.n665 VDD.t4364 28.565
R3159 VDD.n665 VDD.t1167 28.565
R3160 VDD.n691 VDD.t2338 28.565
R3161 VDD.n691 VDD.t2340 28.565
R3162 VDD.n683 VDD.t728 28.565
R3163 VDD.n682 VDD.t4368 28.565
R3164 VDD.n682 VDD.t1169 28.565
R3165 VDD.n595 VDD.t3480 28.565
R3166 VDD.n595 VDD.t3488 28.565
R3167 VDD.n590 VDD.t2876 28.565
R3168 VDD.n590 VDD.t4230 28.565
R3169 VDD.n607 VDD.t2872 28.565
R3170 VDD.n607 VDD.t4226 28.565
R3171 VDD.n602 VDD.t2998 28.565
R3172 VDD.n602 VDD.t3000 28.565
R3173 VDD.n603 VDD.t2996 28.565
R3174 VDD.n603 VDD.t3482 28.565
R3175 VDD.n605 VDD.t3490 28.565
R3176 VDD.n605 VDD.t1110 28.565
R3177 VDD.n581 VDD.t4462 28.565
R3178 VDD.n581 VDD.t365 28.565
R3179 VDD.n576 VDD.t4579 28.565
R3180 VDD.n576 VDD.t4573 28.565
R3181 VDD.n292 VDD.t1870 28.565
R3182 VDD.n292 VDD.t1886 28.565
R3183 VDD.n287 VDD.t4014 28.565
R3184 VDD.n287 VDD.t4016 28.565
R3185 VDD.n288 VDD.t2801 28.565
R3186 VDD.n288 VDD.t4393 28.565
R3187 VDD.n290 VDD.t1321 28.565
R3188 VDD.n290 VDD.t4382 28.565
R3189 VDD.n282 VDD.t4571 28.565
R3190 VDD.n282 VDD.t4581 28.565
R3191 VDD.n277 VDD.t359 28.565
R3192 VDD.n277 VDD.t367 28.565
R3193 VDD.n278 VDD.t4069 28.565
R3194 VDD.n278 VDD.t4460 28.565
R3195 VDD.n279 VDD.t4071 28.565
R3196 VDD.n279 VDD.t4073 28.565
R3197 VDD.n259 VDD.t1059 28.565
R3198 VDD.n259 VDD.t475 28.565
R3199 VDD.n254 VDD.t1139 28.565
R3200 VDD.n254 VDD.t1147 28.565
R3201 VDD.n271 VDD.t1153 28.565
R3202 VDD.n271 VDD.t1143 28.565
R3203 VDD.n266 VDD.t473 28.565
R3204 VDD.n266 VDD.t1055 28.565
R3205 VDD.n267 VDD.t600 28.565
R3206 VDD.n267 VDD.t1061 28.565
R3207 VDD.n268 VDD.t602 28.565
R3208 VDD.n268 VDD.t604 28.565
R3209 VDD.n620 VDD.t3038 28.565
R3210 VDD.n620 VDD.t3040 28.565
R3211 VDD.n612 VDD.t822 28.565
R3212 VDD.n611 VDD.t804 28.565
R3213 VDD.n611 VDD.t1219 28.565
R3214 VDD.n751 VDD.t1036 28.565
R3215 VDD.n751 VDD.t1040 28.565
R3216 VDD.n743 VDD.t684 28.565
R3217 VDD.n742 VDD.t1205 28.565
R3218 VDD.n742 VDD.t1173 28.565
R3219 VDD.n769 VDD.t3322 28.565
R3220 VDD.n769 VDD.t3326 28.565
R3221 VDD.n761 VDD.t802 28.565
R3222 VDD.n760 VDD.t1189 28.565
R3223 VDD.n760 VDD.t742 28.565
R3224 VDD.n787 VDD.t1765 28.565
R3225 VDD.n787 VDD.t1763 28.565
R3226 VDD.n779 VDD.t810 28.565
R3227 VDD.n778 VDD.t4360 28.565
R3228 VDD.n778 VDD.t744 28.565
R3229 VDD.n3373 VDD.t395 28.565
R3230 VDD.n3373 VDD.t397 28.565
R3231 VDD.n3378 VDD.t2741 28.565
R3232 VDD.n3378 VDD.t2740 28.565
R3233 VDD.n3321 VDD.t3634 28.565
R3234 VDD.n3321 VDD.t3633 28.565
R3235 VDD.n3316 VDD.t1108 28.565
R3236 VDD.n3316 VDD.t1107 28.565
R3237 VDD.n3272 VDD.t960 28.565
R3238 VDD.n3272 VDD.t962 28.565
R3239 VDD.n3273 VDD.t3869 28.565
R3240 VDD.n3273 VDD.t961 28.565
R3241 VDD.n3269 VDD.t3766 28.565
R3242 VDD.n3269 VDD.t3765 28.565
R3243 VDD.n3268 VDD.t3104 28.565
R3244 VDD.n3268 VDD.t3870 28.565
R3245 VDD.n3329 VDD.t4540 28.565
R3246 VDD.n3329 VDD.t4539 28.565
R3247 VDD.n3330 VDD.t3367 28.565
R3248 VDD.n3330 VDD.t4541 28.565
R3249 VDD.n3326 VDD.t1439 28.565
R3250 VDD.n3326 VDD.t1438 28.565
R3251 VDD.n3325 VDD.t3364 28.565
R3252 VDD.n3325 VDD.t3112 28.565
R3253 VDD.n3386 VDD.t2506 28.565
R3254 VDD.n3386 VDD.t2505 28.565
R3255 VDD.n3387 VDD.t2405 28.565
R3256 VDD.n3387 VDD.t2507 28.565
R3257 VDD.n3383 VDD.t3458 28.565
R3258 VDD.n3383 VDD.t2094 28.565
R3259 VDD.n3382 VDD.t2407 28.565
R3260 VDD.n3382 VDD.t2406 28.565
R3261 VDD.n195 VDD.t653 28.565
R3262 VDD.n195 VDD.t652 28.565
R3263 VDD.n196 VDD.t536 28.565
R3264 VDD.n196 VDD.t654 28.565
R3265 VDD.n192 VDD.t1995 28.565
R3266 VDD.n192 VDD.t263 28.565
R3267 VDD.n191 VDD.t538 28.565
R3268 VDD.n191 VDD.t537 28.565
R3269 VDD.n199 VDD.t1034 28.565
R3270 VDD.n199 VDD.t1033 28.565
R3271 VDD.n204 VDD.t3158 28.565
R3272 VDD.n204 VDD.t1748 28.565
R3273 VDD.n3264 VDD.t1029 28.565
R3274 VDD.n3264 VDD.t1028 28.565
R3275 VDD.n847 VDD.t2302 28.565
R3276 VDD.n847 VDD.t2298 28.565
R3277 VDD.n850 VDD.t3349 28.565
R3278 VDD.n850 VDD.t3351 28.565
R3279 VDD.n851 VDD.t3350 28.565
R3280 VDD.n851 VDD.t3258 28.565
R3281 VDD.n846 VDD.t3245 28.565
R3282 VDD.n846 VDD.t2388 28.565
R3283 VDD.n827 VDD.t1787 28.565
R3284 VDD.n827 VDD.t3822 28.565
R3285 VDD.n830 VDD.t3698 28.565
R3286 VDD.n830 VDD.t3697 28.565
R3287 VDD.n831 VDD.t3595 28.565
R3288 VDD.n831 VDD.t1499 28.565
R3289 VDD.n826 VDD.t1498 28.565
R3290 VDD.n826 VDD.t1496 28.565
R3291 VDD.n23 VDD.t188 28.565
R3292 VDD.n23 VDD.t187 28.565
R3293 VDD.n26 VDD.t2639 28.565
R3294 VDD.n26 VDD.t2638 28.565
R3295 VDD.n27 VDD.t2637 28.565
R3296 VDD.n27 VDD.t2587 28.565
R3297 VDD.n22 VDD.t2293 28.565
R3298 VDD.n22 VDD.t2292 28.565
R3299 VDD.n31 VDD.t416 28.565
R3300 VDD.n31 VDD.t417 28.565
R3301 VDD.n36 VDD.t2521 28.565
R3302 VDD.n36 VDD.t2520 28.565
R3303 VDD.n1 VDD.t1434 28.565
R3304 VDD.n1 VDD.t1088 28.565
R3305 VDD.n6 VDD.t345 28.565
R3306 VDD.n6 VDD.t2721 28.565
R3307 VDD.n822 VDD.t899 28.565
R3308 VDD.n822 VDD.t895 28.565
R3309 VDD.n818 VDD.t3680 28.565
R3310 VDD.n818 VDD.t3679 28.565
R3311 VDD.n819 VDD.t1543 28.565
R3312 VDD.n819 VDD.t1489 28.565
R3313 VDD.n821 VDD.t1500 28.565
R3314 VDD.n821 VDD.t1493 28.565
R3315 VDD.n804 VDD.t3995 28.565
R3316 VDD.n804 VDD.t3976 28.565
R3317 VDD.n807 VDD.t3652 28.565
R3318 VDD.n807 VDD.t3651 28.565
R3319 VDD.n808 VDD.t3650 28.565
R3320 VDD.n808 VDD.t339 28.565
R3321 VDD.n803 VDD.t338 28.565
R3322 VDD.n803 VDD.t337 28.565
R3323 VDD.n87 VDD.t1349 28.565
R3324 VDD.n87 VDD.t1348 28.565
R3325 VDD.n82 VDD.t3050 28.565
R3326 VDD.n82 VDD.t3049 28.565
R3327 VDD.n133 VDD.t4408 28.565
R3328 VDD.n133 VDD.t4413 28.565
R3329 VDD.n136 VDD.t1015 28.565
R3330 VDD.n136 VDD.t1014 28.565
R3331 VDD.n137 VDD.t1013 28.565
R3332 VDD.n137 VDD.t757 28.565
R3333 VDD.n132 VDD.t755 28.565
R3334 VDD.n132 VDD.t754 28.565
R3335 VDD.n141 VDD.t3233 28.565
R3336 VDD.n141 VDD.t3232 28.565
R3337 VDD.n146 VDD.t3231 28.565
R3338 VDD.n146 VDD.t3230 28.565
R3339 VDD.n181 VDD.t3138 28.565
R3340 VDD.n181 VDD.t3137 28.565
R3341 VDD.n186 VDD.t1307 28.565
R3342 VDD.n186 VDD.t1305 28.565
R3343 VDD.n169 VDD.t758 28.565
R3344 VDD.n169 VDD.t756 28.565
R3345 VDD.n174 VDD.t3552 28.565
R3346 VDD.n174 VDD.t4416 28.565
R3347 VDD.n159 VDD.t1311 28.565
R3348 VDD.n159 VDD.t1308 28.565
R3349 VDD.n162 VDD.t4200 28.565
R3350 VDD.n162 VDD.t4202 28.565
R3351 VDD.n163 VDD.t4201 28.565
R3352 VDD.n163 VDD.t762 28.565
R3353 VDD.n158 VDD.t761 28.565
R3354 VDD.n158 VDD.t760 28.565
R3355 VDD.n151 VDD.t4417 28.565
R3356 VDD.n151 VDD.t4419 28.565
R3357 VDD.n154 VDD.t2525 28.565
R3358 VDD.n154 VDD.t3525 28.565
R3359 VDD.n155 VDD.t3524 28.565
R3360 VDD.n155 VDD.t1963 28.565
R3361 VDD.n150 VDD.t1962 28.565
R3362 VDD.n150 VDD.t1961 28.565
R3363 VDD.n122 VDD.t750 28.565
R3364 VDD.n122 VDD.t749 28.565
R3365 VDD.n127 VDD.t993 28.565
R3366 VDD.n127 VDD.t1003 28.565
R3367 VDD.n110 VDD.t1915 28.565
R3368 VDD.n110 VDD.t340 28.565
R3369 VDD.n115 VDD.t3963 28.565
R3370 VDD.n115 VDD.t4032 28.565
R3371 VDD.n100 VDD.t997 28.565
R3372 VDD.n100 VDD.t996 28.565
R3373 VDD.n103 VDD.t3557 28.565
R3374 VDD.n103 VDD.t4135 28.565
R3375 VDD.n104 VDD.t4134 28.565
R3376 VDD.n104 VDD.t342 28.565
R3377 VDD.n99 VDD.t341 28.565
R3378 VDD.n99 VDD.t335 28.565
R3379 VDD.n92 VDD.t4029 28.565
R3380 VDD.n92 VDD.t3990 28.565
R3381 VDD.n95 VDD.t3103 28.565
R3382 VDD.n95 VDD.t3102 28.565
R3383 VDD.n96 VDD.t4532 28.565
R3384 VDD.n96 VDD.t992 28.565
R3385 VDD.n91 VDD.t1002 28.565
R3386 VDD.n91 VDD.t1001 28.565
R3387 VDD.n836 VDD.t1491 28.565
R3388 VDD.n836 VDD.t1490 28.565
R3389 VDD.n841 VDD.t2304 28.565
R3390 VDD.n841 VDD.t2303 28.565
R3391 VDD.n12 VDD.t524 28.565
R3392 VDD.n12 VDD.t523 28.565
R3393 VDD.n17 VDD.t2391 28.565
R3394 VDD.n17 VDD.t3848 28.565
R3395 VDD.n71 VDD.t4081 28.565
R3396 VDD.n71 VDD.t4080 28.565
R3397 VDD.n76 VDD.t2570 28.565
R3398 VDD.n76 VDD.t2572 28.565
R3399 VDD.n59 VDD.t2589 28.565
R3400 VDD.n59 VDD.t2588 28.565
R3401 VDD.n64 VDD.t1924 28.565
R3402 VDD.n64 VDD.t151 28.565
R3403 VDD.n49 VDD.t2566 28.565
R3404 VDD.n49 VDD.t2574 28.565
R3405 VDD.n52 VDD.t878 28.565
R3406 VDD.n52 VDD.t877 28.565
R3407 VDD.n53 VDD.t876 28.565
R3408 VDD.n53 VDD.t2586 28.565
R3409 VDD.n48 VDD.t2585 28.565
R3410 VDD.n48 VDD.t256 28.565
R3411 VDD.n41 VDD.t2578 28.565
R3412 VDD.n41 VDD.t3399 28.565
R3413 VDD.n44 VDD.t3174 28.565
R3414 VDD.n44 VDD.t3173 28.565
R3415 VDD.n45 VDD.t3172 28.565
R3416 VDD.n45 VDD.t2569 28.565
R3417 VDD.n40 VDD.t2783 28.565
R3418 VDD.n40 VDD.t2782 28.565
R3419 VDD.n3400 VDD.t3615 28.565
R3420 VDD.n3400 VDD.t3614 28.565
R3421 VDD.n3424 VDD.t3178 28.565
R3422 VDD.n3424 VDD.t3177 28.565
R3423 VDD.n3419 VDD.t3749 28.565
R3424 VDD.n3419 VDD.t3746 28.565
R3425 VDD.n3413 VDD.t2650 28.565
R3426 VDD.n3413 VDD.t1266 28.565
R3427 VDD.n3408 VDD.t3540 28.565
R3428 VDD.n3408 VDD.t1657 28.565
R3429 VDD.n3432 VDD.t3285 28.565
R3430 VDD.n3432 VDD.t3284 28.565
R3431 VDD.n3433 VDD.t3105 28.565
R3432 VDD.n3433 VDD.t1660 28.565
R3433 VDD.n3429 VDD.t1658 28.565
R3434 VDD.n3429 VDD.t1656 28.565
R3435 VDD.n3428 VDD.t1601 28.565
R3436 VDD.n3428 VDD.t1600 28.565
R3437 VDD.n3435 VDD.t677 28.565
R3438 VDD.n3435 VDD.t3136 28.565
R3439 VDD.n3436 VDD.t1654 28.565
R3440 VDD.n3436 VDD.t678 28.565
R3441 VDD.n3439 VDD.t3771 28.565
R3442 VDD.n3439 VDD.t3770 28.565
R3443 VDD.n3438 VDD.t1652 28.565
R3444 VDD.n3438 VDD.t1653 28.565
R3445 VDD.n3282 VDD.t1460 28.565
R3446 VDD.n3282 VDD.t1459 28.565
R3447 VDD.n3277 VDD.t3108 28.565
R3448 VDD.n3277 VDD.t3107 28.565
R3449 VDD.n3310 VDD.t3292 28.565
R3450 VDD.n3310 VDD.t3291 28.565
R3451 VDD.n3305 VDD.t4505 28.565
R3452 VDD.n3305 VDD.t4504 28.565
R3453 VDD.n3290 VDD.t4187 28.565
R3454 VDD.n3290 VDD.t3330 28.565
R3455 VDD.n3291 VDD.t3111 28.565
R3456 VDD.n3291 VDD.t4188 28.565
R3457 VDD.n3287 VDD.t3298 28.565
R3458 VDD.n3287 VDD.t3297 28.565
R3459 VDD.n3286 VDD.t3366 28.565
R3460 VDD.n3286 VDD.t3113 28.565
R3461 VDD.n3293 VDD.t224 28.565
R3462 VDD.n3293 VDD.t223 28.565
R3463 VDD.n3294 VDD.t3295 28.565
R3464 VDD.n3294 VDD.t225 28.565
R3465 VDD.n3297 VDD.t3023 28.565
R3466 VDD.n3297 VDD.t3016 28.565
R3467 VDD.n3296 VDD.t3300 28.565
R3468 VDD.n3296 VDD.t3296 28.565
R3469 VDD.n3339 VDD.t2091 28.565
R3470 VDD.n3339 VDD.t669 28.565
R3471 VDD.n3334 VDD.t3132 28.565
R3472 VDD.n3334 VDD.t2404 28.565
R3473 VDD.n3367 VDD.t2980 28.565
R3474 VDD.n3367 VDD.t2977 28.565
R3475 VDD.n3362 VDD.t1376 28.565
R3476 VDD.n3362 VDD.t1375 28.565
R3477 VDD.n3347 VDD.t2720 28.565
R3478 VDD.n3347 VDD.t2719 28.565
R3479 VDD.n3348 VDD.t3130 28.565
R3480 VDD.n3348 VDD.t2718 28.565
R3481 VDD.n3344 VDD.t2985 28.565
R3482 VDD.n3344 VDD.t2984 28.565
R3483 VDD.n3343 VDD.t3133 28.565
R3484 VDD.n3343 VDD.t3131 28.565
R3485 VDD.n3350 VDD.t3504 28.565
R3486 VDD.n3350 VDD.t3503 28.565
R3487 VDD.n3351 VDD.t2976 28.565
R3488 VDD.n3351 VDD.t612 28.565
R3489 VDD.n3354 VDD.t3467 28.565
R3490 VDD.n3354 VDD.t3442 28.565
R3491 VDD.n3353 VDD.t2981 28.565
R3492 VDD.n3353 VDD.t2978 28.565
R3493 VDD.n215 VDD.t1994 28.565
R3494 VDD.n215 VDD.t2031 28.565
R3495 VDD.n210 VDD.t2511 28.565
R3496 VDD.n210 VDD.t2510 28.565
R3497 VDD.n243 VDD.t981 28.565
R3498 VDD.n243 VDD.t988 28.565
R3499 VDD.n238 VDD.t4565 28.565
R3500 VDD.n238 VDD.t4561 28.565
R3501 VDD.n223 VDD.t2759 28.565
R3502 VDD.n223 VDD.t2758 28.565
R3503 VDD.n224 VDD.t539 28.565
R3504 VDD.n224 VDD.t2760 28.565
R3505 VDD.n220 VDD.t985 28.565
R3506 VDD.n220 VDD.t984 28.565
R3507 VDD.n219 VDD.t2508 28.565
R3508 VDD.n219 VDD.t540 28.565
R3509 VDD.n226 VDD.t3515 28.565
R3510 VDD.n226 VDD.t3514 28.565
R3511 VDD.n227 VDD.t987 28.565
R3512 VDD.n227 VDD.t3516 28.565
R3513 VDD.n230 VDD.t265 28.565
R3514 VDD.n230 VDD.t264 28.565
R3515 VDD.n229 VDD.t980 28.565
R3516 VDD.n229 VDD.t979 28.565
R3517 VDD.n359 VDD.t890 28.565
R3518 VDD.n359 VDD.t894 28.565
R3519 VDD.n364 VDD.t2814 28.565
R3520 VDD.n364 VDD.t2350 28.565
R3521 VDD.n341 VDD.t2401 28.565
R3522 VDD.n341 VDD.t4523 28.565
R3523 VDD.n346 VDD.t958 28.565
R3524 VDD.n346 VDD.t651 28.565
R3525 VDD.n325 VDD.t2348 28.565
R3526 VDD.n325 VDD.t3586 28.565
R3527 VDD.n329 VDD.t3155 28.565
R3528 VDD.n329 VDD.t2361 28.565
R3529 VDD.n330 VDD.t3157 28.565
R3530 VDD.n330 VDD.t2397 28.565
R3531 VDD.n324 VDD.t4521 28.565
R3532 VDD.n324 VDD.t4527 28.565
R3533 VDD.n313 VDD.t3498 28.565
R3534 VDD.n313 VDD.t1557 28.565
R3535 VDD.n318 VDD.t66 28.565
R3536 VDD.n318 VDD.t68 28.565
R3537 VDD.n319 VDD.t70 28.565
R3538 VDD.n319 VDD.t3584 28.565
R3539 VDD.n312 VDD.t2818 28.565
R3540 VDD.n312 VDD.t3582 28.565
R3541 VDD.n459 VDD.t566 28.565
R3542 VDD.n459 VDD.t570 28.565
R3543 VDD.n464 VDD.t1639 28.565
R3544 VDD.n464 VDD.t1701 28.565
R3545 VDD.n440 VDD.t493 28.565
R3546 VDD.n440 VDD.t4466 28.565
R3547 VDD.n445 VDD.t622 28.565
R3548 VDD.n445 VDD.t628 28.565
R3549 VDD.n432 VDD.t1699 28.565
R3550 VDD.n432 VDD.t3694 28.565
R3551 VDD.n416 VDD.t3071 28.565
R3552 VDD.n416 VDD.t3073 28.565
R3553 VDD.n417 VDD.t3069 28.565
R3554 VDD.n417 VDD.t487 28.565
R3555 VDD.n431 VDD.t495 28.565
R3556 VDD.n431 VDD.t485 28.565
R3557 VDD.n423 VDD.t616 28.565
R3558 VDD.n423 VDD.t1023 28.565
R3559 VDD.n422 VDD.t1711 28.565
R3560 VDD.n422 VDD.t1713 28.565
R3561 VDD.n419 VDD.t1065 28.565
R3562 VDD.n419 VDD.t1705 28.565
R3563 VDD.n420 VDD.t1063 28.565
R3564 VDD.n420 VDD.t2685 28.565
R3565 VDD.n471 VDD.t4266 28.565
R3566 VDD.n471 VDD.t4264 28.565
R3567 VDD.n476 VDD.t100 28.565
R3568 VDD.n476 VDD.t1488 28.565
R3569 VDD.n508 VDD.t1229 28.565
R3570 VDD.n508 VDD.t1235 28.565
R3571 VDD.n513 VDD.t777 28.565
R3572 VDD.n513 VDD.t775 28.565
R3573 VDD.n492 VDD.t98 28.565
R3574 VDD.n492 VDD.t1486 28.565
R3575 VDD.n497 VDD.t1047 28.565
R3576 VDD.n497 VDD.t3578 28.565
R3577 VDD.n498 VDD.t1045 28.565
R3578 VDD.n498 VDD.t1247 28.565
R3579 VDD.n491 VDD.t1231 28.565
R3580 VDD.n491 VDD.t1241 28.565
R3581 VDD.n484 VDD.t976 28.565
R3582 VDD.n484 VDD.t773 28.565
R3583 VDD.n483 VDD.t90 28.565
R3584 VDD.n483 VDD.t94 28.565
R3585 VDD.n480 VDD.t3361 28.565
R3586 VDD.n480 VDD.t84 28.565
R3587 VDD.n481 VDD.t3357 28.565
R3588 VDD.n481 VDD.t3359 28.565
R3589 VDD.n2758 VDD.t4435 28.565
R3590 VDD.n2758 VDD.t4427 28.565
R3591 VDD.n2763 VDD.t4167 28.565
R3592 VDD.n2763 VDD.t4161 28.565
R3593 VDD.n2792 VDD.t4097 28.565
R3594 VDD.n2792 VDD.t4105 28.565
R3595 VDD.n2797 VDD.t1684 28.565
R3596 VDD.n2797 VDD.t1688 28.565
R3597 VDD.n2783 VDD.t4159 28.565
R3598 VDD.n2783 VDD.t4163 28.565
R3599 VDD.n2767 VDD.t3529 28.565
R3600 VDD.n2767 VDD.t3531 28.565
R3601 VDD.n2768 VDD.t3143 28.565
R3602 VDD.n2768 VDD.t4087 28.565
R3603 VDD.n2782 VDD.t4101 28.565
R3604 VDD.n2782 VDD.t4085 28.565
R3605 VDD.n2774 VDD.t1674 28.565
R3606 VDD.n2774 VDD.t1682 28.565
R3607 VDD.n2773 VDD.t2066 28.565
R3608 VDD.n2773 VDD.t4155 28.565
R3609 VDD.n2770 VDD.t3332 28.565
R3610 VDD.n2770 VDD.t4169 28.565
R3611 VDD.n2771 VDD.t1585 28.565
R3612 VDD.n2771 VDD.t1587 28.565
R3613 VDD.n2694 VDD.t1752 28.565
R3614 VDD.n2694 VDD.t3663 28.565
R3615 VDD.n2699 VDD.t1936 28.565
R3616 VDD.n2699 VDD.t1944 28.565
R3617 VDD.n2729 VDD.t3563 28.565
R3618 VDD.n2729 VDD.t211 28.565
R3619 VDD.n2734 VDD.t2710 28.565
R3620 VDD.n2734 VDD.t2702 28.565
R3621 VDD.n2721 VDD.t550 28.565
R3622 VDD.n2721 VDD.t548 28.565
R3623 VDD.n2714 VDD.t1635 28.565
R3624 VDD.n2714 VDD.t1637 28.565
R3625 VDD.n2715 VDD.t1633 28.565
R3626 VDD.n2715 VDD.t219 28.565
R3627 VDD.n2720 VDD.t203 28.565
R3628 VDD.n2720 VDD.t217 28.565
R3629 VDD.n2707 VDD.t2712 28.565
R3630 VDD.n2707 VDD.t186 28.565
R3631 VDD.n2706 VDD.t1950 28.565
R3632 VDD.n2706 VDD.t1948 28.565
R3633 VDD.n2703 VDD.t392 28.565
R3634 VDD.n2703 VDD.t1942 28.565
R3635 VDD.n2704 VDD.t1119 28.565
R3636 VDD.n2704 VDD.t390 28.565
R3637 VDD.n2183 VDD.t4059 28.565
R3638 VDD.n2183 VDD.t3211 28.565
R3639 VDD.n2169 VDD.t3731 28.565
R3640 VDD.n2169 VDD.t1357 28.565
R3641 VDD.n2151 VDD.t2479 28.565
R3642 VDD.n2151 VDD.t2465 28.565
R3643 VDD.n2144 VDD.t3919 28.565
R3644 VDD.n2144 VDD.t3219 28.565
R3645 VDD.n1470 VDD.t3911 28.565
R3646 VDD.n1470 VDD.t1031 28.565
R3647 VDD.n1456 VDD.t2207 28.565
R3648 VDD.n1456 VDD.t2229 28.565
R3649 VDD.n2031 VDD.t1386 28.565
R3650 VDD.n2031 VDD.t1406 28.565
R3651 VDD.n2046 VDD.t1467 28.565
R3652 VDD.n2046 VDD.t1437 28.565
R3653 VDD.n1931 VDD.t1355 28.565
R3654 VDD.n1931 VDD.t3737 28.565
R3655 VDD.n1946 VDD.t4031 28.565
R3656 VDD.n1946 VDD.t3984 28.565
R3657 VDD.n1881 VDD.t2219 28.565
R3658 VDD.n1881 VDD.t2195 28.565
R3659 VDD.n1896 VDD.t2335 28.565
R3660 VDD.n1896 VDD.t2322 28.565
R3661 VDD.n1906 VDD.t4141 28.565
R3662 VDD.n1906 VDD.t2477 28.565
R3663 VDD.n1921 VDD.t3398 28.565
R3664 VDD.n1921 VDD.t194 28.565
R3665 VDD.n1956 VDD.t1906 28.565
R3666 VDD.n1956 VDD.t2658 28.565
R3667 VDD.n1971 VDD.t4415 28.565
R3668 VDD.n1971 VDD.t4372 28.565
R3669 VDD.n1981 VDD.t1876 28.565
R3670 VDD.n1981 VDD.t933 28.565
R3671 VDD.n1996 VDD.t279 28.565
R3672 VDD.n1996 VDD.t273 28.565
R3673 VDD.n2006 VDD.t1822 28.565
R3674 VDD.n2006 VDD.t2417 28.565
R3675 VDD.n2021 VDD.t3444 28.565
R3676 VDD.n2021 VDD.t3426 28.565
R3677 VDD.n2056 VDD.t2624 28.565
R3678 VDD.n2056 VDD.t2604 28.565
R3679 VDD.n2071 VDD.t3760 28.565
R3680 VDD.n2071 VDD.t3776 28.565
R3681 VDD.n2123 VDD.t3762 28.565
R3682 VDD.n2123 VDD.t3778 28.565
R3683 VDD.n2117 VDD.t3022 28.565
R3684 VDD.n2117 VDD.t3018 28.565
R3685 VDD.n2111 VDD.t3449 28.565
R3686 VDD.n2111 VDD.t2079 28.565
R3687 VDD.n2105 VDD.t1993 28.565
R3688 VDD.n2105 VDD.t2022 28.565
R3689 VDD.n2099 VDD.t4405 28.565
R3690 VDD.n2099 VDD.t4374 28.565
R3691 VDD.n2093 VDD.t4028 28.565
R3692 VDD.n2093 VDD.t3980 28.565
R3693 VDD.n2087 VDD.t3389 28.565
R3694 VDD.n2087 VDD.t190 28.565
R3695 VDD.n2081 VDD.t2332 28.565
R3696 VDD.n2081 VDD.t897 28.565
R3697 VDD.n1743 VDD.t2805 28.565
R3698 VDD.n1743 VDD.t1504 28.565
R3699 VDD.n1734 VDD.t3810 28.565
R3700 VDD.n1734 VDD.t3915 28.565
R3701 VDD.n1735 VDD.t2243 28.565
R3702 VDD.n1768 VDD.t3573 28.565
R3703 VDD.n1768 VDD.t3569 28.565
R3704 VDD.n1759 VDD.t1604 28.565
R3705 VDD.n1759 VDD.t4050 28.565
R3706 VDD.n1760 VDD.t3868 28.565
R3707 VDD.n1864 VDD.t1520 28.565
R3708 VDD.n1864 VDD.t1518 28.565
R3709 VDD.n1865 VDD.t1353 28.565
R3710 VDD.n1861 VDD.t2768 28.565
R3711 VDD.n1861 VDD.t2770 28.565
R3712 VDD.n1839 VDD.t2375 28.565
R3713 VDD.n1839 VDD.t1510 28.565
R3714 VDD.n1840 VDD.t3690 28.565
R3715 VDD.n1836 VDD.t348 28.565
R3716 VDD.n1836 VDD.t350 28.565
R3717 VDD.n1818 VDD.t1723 28.565
R3718 VDD.n1818 VDD.t3874 28.565
R3719 VDD.n1809 VDD.t3201 28.565
R3720 VDD.n1809 VDD.t3940 28.565
R3721 VDD.n1810 VDD.t1522 28.565
R3722 VDD.n1793 VDD.t2677 28.565
R3723 VDD.n1793 VDD.t2679 28.565
R3724 VDD.n1784 VDD.t1810 28.565
R3725 VDD.n1784 VDD.t2377 28.565
R3726 VDD.n1785 VDD.t4002 28.565
R3727 VDD.n1718 VDD.t2541 28.565
R3728 VDD.n1718 VDD.t1279 28.565
R3729 VDD.n1709 VDD.t1786 28.565
R3730 VDD.n1709 VDD.t2241 28.565
R3731 VDD.n1710 VDD.t2235 28.565
R3732 VDD.n1694 VDD.t1564 28.565
R3733 VDD.n1694 VDD.t1566 28.565
R3734 VDD.n1685 VDD.t3998 28.565
R3735 VDD.n1685 VDD.t4036 28.565
R3736 VDD.n1686 VDD.t3279 28.565
R3737 VDD.n1539 VDD.t704 28.565
R3738 VDD.n1539 VDD.t698 28.565
R3739 VDD.n1540 VDD.t4366 28.565
R3740 VDD.n1536 VDD.t2673 28.565
R3741 VDD.n1536 VDD.t2671 28.565
R3742 VDD.n1564 VDD.t694 28.565
R3743 VDD.n1564 VDD.t686 28.565
R3744 VDD.n1565 VDD.t4358 28.565
R3745 VDD.n1561 VDD.t2766 28.565
R3746 VDD.n1561 VDD.t2764 28.565
R3747 VDD.n1664 VDD.t1185 28.565
R3748 VDD.n1664 VDD.t1217 28.565
R3749 VDD.n1665 VDD.t1207 28.565
R3750 VDD.n1661 VDD.t1157 28.565
R3751 VDD.n1661 VDD.t531 28.565
R3752 VDD.n1639 VDD.t4370 28.565
R3753 VDD.n1639 VDD.t1213 28.565
R3754 VDD.n1640 VDD.t1203 28.565
R3755 VDD.n1636 VDD.t4493 28.565
R3756 VDD.n1636 VDD.t4491 28.565
R3757 VDD.n1614 VDD.t722 28.565
R3758 VDD.n1614 VDD.t718 28.565
R3759 VDD.n1615 VDD.t816 28.565
R3760 VDD.n1611 VDD.t403 28.565
R3761 VDD.n1611 VDD.t401 28.565
R3762 VDD.n1589 VDD.t1221 28.565
R3763 VDD.n1589 VDD.t1211 28.565
R3764 VDD.n1590 VDD.t716 28.565
R3765 VDD.n1586 VDD.t481 28.565
R3766 VDD.n1586 VDD.t479 28.565
R3767 VDD.n1514 VDD.t814 28.565
R3768 VDD.n1514 VDD.t798 28.565
R3769 VDD.n1515 VDD.t832 28.565
R3770 VDD.n1511 VDD.t2691 28.565
R3771 VDD.n1511 VDD.t1087 28.565
R3772 VDD.n1490 VDD.t734 28.565
R3773 VDD.n1490 VDD.t836 28.565
R3774 VDD.n1491 VDD.t828 28.565
R3775 VDD.n1487 VDD.t3556 28.565
R3776 VDD.n1487 VDD.t3554 28.565
R3777 VDD.n1389 VDD.t1782 28.565
R3778 VDD.n1389 VDD.t4034 28.565
R3779 VDD.n1390 VDD.t1789 28.565
R3780 VDD.n1386 VDD.t2311 28.565
R3781 VDD.n1386 VDD.t2309 28.565
R3782 VDD.n1364 VDD.t2237 28.565
R3783 VDD.n1364 VDD.t3275 28.565
R3784 VDD.n1365 VDD.t3841 28.565
R3785 VDD.n1361 VDD.t457 28.565
R3786 VDD.n1361 VDD.t455 28.565
R3787 VDD.n1265 VDD.t2051 28.565
R3788 VDD.n1265 VDD.t4063 28.565
R3789 VDD.n1266 VDD.t3835 28.565
R3790 VDD.n1262 VDD.t2730 28.565
R3791 VDD.n1262 VDD.t1283 28.565
R3792 VDD.n1289 VDD.t3828 28.565
R3793 VDD.n1289 VDD.t1744 28.565
R3794 VDD.n1290 VDD.t1482 28.565
R3795 VDD.n1286 VDD.t373 28.565
R3796 VDD.n1286 VDD.t371 28.565
R3797 VDD.n1314 VDD.t1776 28.565
R3798 VDD.n1314 VDD.t3837 28.565
R3799 VDD.n1315 VDD.t1005 28.565
R3800 VDD.n1311 VDD.t636 28.565
R3801 VDD.n1311 VDD.t634 28.565
R3802 VDD.n1339 VDD.t4046 28.565
R3803 VDD.n1339 VDD.t4038 28.565
R3804 VDD.n1340 VDD.t3830 28.565
R3805 VDD.n1336 VDD.t317 28.565
R3806 VDD.n1336 VDD.t315 28.565
R3807 VDD.n1414 VDD.t1780 28.565
R3808 VDD.n1414 VDD.t3281 28.565
R3809 VDD.n1415 VDD.t3267 28.565
R3810 VDD.n1411 VDD.t3934 28.565
R3811 VDD.n1411 VDD.t3932 28.565
R3812 VDD.n1439 VDD.t2390 28.565
R3813 VDD.n1439 VDD.t2233 28.565
R3814 VDD.n1440 VDD.t3273 28.565
R3815 VDD.n1436 VDD.t2494 28.565
R3816 VDD.n1436 VDD.t2492 28.565
R3817 VDD.n1080 VDD.t3353 28.565
R3818 VDD.n1080 VDD.t3599 28.565
R3819 VDD.n1079 VDD.t1359 28.565
R3820 VDD.n1079 VDD.t3355 28.565
R3821 VDD.n1078 VDD.t3735 28.565
R3822 VDD.n1078 VDD.t1363 28.565
R3823 VDD.n1076 VDD.t3967 28.565
R3824 VDD.n1076 VDD.t3975 28.565
R3825 VDD.n1088 VDD.t1369 28.565
R3826 VDD.n1088 VDD.t1371 28.565
R3827 VDD.n1087 VDD.t1912 28.565
R3828 VDD.n1087 VDD.t1373 28.565
R3829 VDD.n1086 VDD.t3065 28.565
R3830 VDD.n1086 VDD.t3063 28.565
R3831 VDD.n1084 VDD.t4380 28.565
R3832 VDD.n1084 VDD.t1325 28.565
R3833 VDD.n1121 VDD.t3676 28.565
R3834 VDD.n1121 VDD.t3674 28.565
R3835 VDD.n1120 VDD.t2622 28.565
R3836 VDD.n1120 VDD.t3672 28.565
R3837 VDD.n1119 VDD.t2598 28.565
R3838 VDD.n1119 VDD.t1545 28.565
R3839 VDD.n1117 VDD.t3751 28.565
R3840 VDD.n1117 VDD.t3748 28.565
R3841 VDD.n1113 VDD.t1365 28.565
R3842 VDD.n1113 VDD.t2451 28.565
R3843 VDD.n1112 VDD.t3318 28.565
R3844 VDD.n1112 VDD.t1367 28.565
R3845 VDD.n1111 VDD.t1392 28.565
R3846 VDD.n1111 VDD.t1390 28.565
R3847 VDD.n1109 VDD.t1450 28.565
R3848 VDD.n1109 VDD.t1447 28.565
R3849 VDD.n1104 VDD.t3956 28.565
R3850 VDD.n1104 VDD.t3952 28.565
R3851 VDD.n1103 VDD.t1828 28.565
R3852 VDD.n1103 VDD.t3954 28.565
R3853 VDD.n1102 VDD.t1836 28.565
R3854 VDD.n1102 VDD.t1832 28.565
R3855 VDD.n1100 VDD.t3441 28.565
R3856 VDD.n1100 VDD.t3437 28.565
R3857 VDD.n1096 VDD.t4303 28.565
R3858 VDD.n1096 VDD.t4301 28.565
R3859 VDD.n1095 VDD.t1868 28.565
R3860 VDD.n1095 VDD.t4305 28.565
R3861 VDD.n1094 VDD.t1892 28.565
R3862 VDD.n1094 VDD.t1888 28.565
R3863 VDD.n1092 VDD.t270 28.565
R3864 VDD.n1092 VDD.t2030 28.565
R3865 VDD.n1071 VDD.t2446 28.565
R3866 VDD.n1071 VDD.t2444 28.565
R3867 VDD.n1070 VDD.t4145 28.565
R3868 VDD.n1070 VDD.t2448 28.565
R3869 VDD.n1069 VDD.t2463 28.565
R3870 VDD.n1069 VDD.t2455 28.565
R3871 VDD.n1067 VDD.t2582 28.565
R3872 VDD.n1067 VDD.t2580 28.565
R3873 VDD.n1063 VDD.t3608 28.565
R3874 VDD.n1063 VDD.t3606 28.565
R3875 VDD.n1062 VDD.t2215 28.565
R3876 VDD.n1062 VDD.t3610 28.565
R3877 VDD.n1061 VDD.t2227 28.565
R3878 VDD.n1061 VDD.t2225 28.565
R3879 VDD.n1059 VDD.t2301 28.565
R3880 VDD.n1059 VDD.t2297 28.565
R3881 VDD.n1162 VDD.t221 28.565
R3882 VDD.n1162 VDD.t414 28.565
R3883 VDD.n1177 VDD.t2181 28.565
R3884 VDD.n1177 VDD.t12 28.565
R3885 VDD.n1222 VDD.t4297 28.565
R3886 VDD.n1222 VDD.t4204 28.565
R3887 VDD.n1207 VDD.t305 28.565
R3888 VDD.n1207 VDD.t303 28.565
R3889 VDD.n1192 VDD.t3379 28.565
R3890 VDD.n1192 VDD.t3383 28.565
R3891 VDD.n1150 VDD.t3511 28.565
R3892 VDD.n1150 VDD.t3509 28.565
R3893 VDD.n1135 VDD.t644 28.565
R3894 VDD.n1135 VDD.t642 28.565
R3895 VDD.n1240 VDD.t3237 28.565
R3896 VDD.n1240 VDD.t2896 28.565
R3897 VDD.n2619 VDD.t2620 28.565
R3898 VDD.n2619 VDD.t2602 28.565
R3899 VDD.n2614 VDD.t3191 28.565
R3900 VDD.n2614 VDD.t1597 28.565
R3901 VDD.n2442 VDD.t3494 28.565
R3902 VDD.n2442 VDD.t1529 28.565
R3903 VDD.n2428 VDD.t1418 28.565
R3904 VDD.n2428 VDD.t3304 28.565
R3905 VDD.n2417 VDD.t1746 28.565
R3906 VDD.n2417 VDD.t2239 28.565
R3907 VDD.n2403 VDD.t1818 28.565
R3908 VDD.n2403 VDD.t4109 28.565
R3909 VDD.n2233 VDD.t2043 28.565
R3910 VDD.n2233 VDD.t3925 28.565
R3911 VDD.n2219 VDD.t939 28.565
R3912 VDD.n2219 VDD.t931 28.565
R3913 VDD.n2208 VDD.t2381 28.565
R3914 VDD.n2208 VDD.t4048 28.565
R3915 VDD.n2194 VDD.t4128 28.565
R3916 VDD.n2194 VDD.t2440 28.565
R3917 VDD.n2604 VDD.t4216 28.565
R3918 VDD.n2604 VDD.t4214 28.565
R3919 VDD.n2595 VDD.t3888 28.565
R3920 VDD.n2595 VDD.t4270 28.565
R3921 VDD.n2596 VDD.t4325 28.565
R3922 VDD.n2465 VDD.t1541 28.565
R3923 VDD.n2465 VDD.t1539 28.565
R3924 VDD.n2456 VDD.t4311 28.565
R3925 VDD.n2456 VDD.t4309 28.565
R3926 VDD.n2457 VDD.t4315 28.565
R3927 VDD.n2484 VDD.t1300 28.565
R3928 VDD.n2484 VDD.t1298 28.565
R3929 VDD.n2475 VDD.t4551 28.565
R3930 VDD.n2475 VDD.t3086 28.565
R3931 VDD.n2476 VDD.t3906 28.565
R3932 VDD.n2544 VDD.t4186 28.565
R3933 VDD.n2544 VDD.t4184 28.565
R3934 VDD.n2535 VDD.t4321 28.565
R3935 VDD.n2535 VDD.t3904 28.565
R3936 VDD.n2536 VDD.t4323 28.565
R3937 VDD.n2564 VDD.t1975 28.565
R3938 VDD.n2564 VDD.t1973 28.565
R3939 VDD.n2555 VDD.t3892 28.565
R3940 VDD.n2555 VDD.t3890 28.565
R3941 VDD.n2556 VDD.t3896 28.565
R3942 VDD.n2584 VDD.t4220 28.565
R3943 VDD.n2584 VDD.t4218 28.565
R3944 VDD.n2575 VDD.t3882 28.565
R3945 VDD.n2575 VDD.t3880 28.565
R3946 VDD.n2576 VDD.t3886 28.565
R3947 VDD.n2524 VDD.t746 28.565
R3948 VDD.n2524 VDD.t748 28.565
R3949 VDD.n2515 VDD.t4331 28.565
R3950 VDD.n2515 VDD.t4327 28.565
R3951 VDD.n2516 VDD.t3078 28.565
R3952 VDD.n2504 VDD.t1009 28.565
R3953 VDD.n2504 VDD.t1007 28.565
R3954 VDD.n2495 VDD.t4268 28.565
R3955 VDD.n2495 VDD.t3098 28.565
R3956 VDD.n2496 VDD.t4272 28.565
R3957 VDD.n2391 VDD.t2958 28.565
R3958 VDD.n2391 VDD.t850 28.565
R3959 VDD.n2392 VDD.t2922 28.565
R3960 VDD.n2388 VDD.t3789 28.565
R3961 VDD.n2388 VDD.t3791 28.565
R3962 VDD.n2256 VDD.t2126 28.565
R3963 VDD.n2256 VDD.t1577 28.565
R3964 VDD.n2247 VDD.t2962 28.565
R3965 VDD.n2247 VDD.t852 28.565
R3966 VDD.n2248 VDD.t2926 28.565
R3967 VDD.n2275 VDD.t2133 28.565
R3968 VDD.n2275 VDD.t2135 28.565
R3969 VDD.n2266 VDD.t2950 28.565
R3970 VDD.n2266 VDD.t866 28.565
R3971 VDD.n2267 VDD.t2914 28.565
R3972 VDD.n2331 VDD.t2970 28.565
R3973 VDD.n2331 VDD.t2968 28.565
R3974 VDD.n2332 VDD.t2934 28.565
R3975 VDD.n2328 VDD.t1856 28.565
R3976 VDD.n2328 VDD.t1117 28.565
R3977 VDD.n2351 VDD.t2920 28.565
R3978 VDD.n2351 VDD.t2956 28.565
R3979 VDD.n2352 VDD.t2936 28.565
R3980 VDD.n2348 VDD.t108 28.565
R3981 VDD.n2348 VDD.t106 28.565
R3982 VDD.n2371 VDD.t2940 28.565
R3983 VDD.n2371 VDD.t2972 28.565
R3984 VDD.n2372 VDD.t868 28.565
R3985 VDD.n2368 VDD.t3046 28.565
R3986 VDD.n2368 VDD.t3048 28.565
R3987 VDD.n2315 VDD.t2553 28.565
R3988 VDD.n2315 VDD.t3534 28.565
R3989 VDD.n2306 VDD.t2916 28.565
R3990 VDD.n2306 VDD.t2954 28.565
R3991 VDD.n2307 VDD.t846 28.565
R3992 VDD.n2295 VDD.t3055 28.565
R3993 VDD.n2295 VDD.t3053 28.565
R3994 VDD.n2286 VDD.t854 28.565
R3995 VDD.n2286 VDD.t2952 28.565
R3996 VDD.n2287 VDD.t2928 28.565
R3997 VDD.n3003 VDD.t3228 23.418
R3998 VDD.n3191 VDD.t4438 23.418
R3999 VDD.n3073 VDD.t1532 23.418
R4000 VDD.n355 VDD.t891 23.418
R4001 VDD.n454 VDD.t567 23.418
R4002 VDD.n522 VDD.t1501 23.418
R4003 VDD.n2806 VDD.t4428 23.418
R4004 VDD.n2743 VDD.t3660 23.418
R4005 VDD.n3251 VDD.t2012 23.317
R4006 VDD.n2900 VDD.t2437 23.317
R4007 VDD.n2673 VDD.t2087 23.317
R4008 VDD.n2664 VDD.t1909 23.317
R4009 VDD.n411 VDD.t1377 23.317
R4010 VDD.n2928 VDD.t1839 23.317
R4011 VDD.n303 VDD.t4396 23.317
R4012 VDD.n294 VDD.t2010 23.317
R4013 VDD.n385 VDD.t2014 23.317
R4014 VDD.n394 VDD.t1419 23.317
R4015 VDD.n2654 VDD.t2089 23.317
R4016 VDD.n707 VDD.t3026 23.317
R4017 VDD.n2646 VDD.t1646 23.317
R4018 VDD.n699 VDD.t3066 23.317
R4019 VDD.n286 VDD.t1869 23.317
R4020 VDD.n276 VDD.t4570 23.317
R4021 VDD.n265 VDD.t1152 23.317
R4022 VDD.n1075 VDD.t3974 23.317
R4023 VDD.n1108 VDD.t1446 23.317
R4024 VDD.n1058 VDD.t2296 23.317
R4025 VDD.n601 VDD.t2871 23.316
R4026 VDD.n738 VDD.t2556 23.316
R4027 VDD.n2881 VDD.t3120 22.813
R4028 VDD.n2851 VDD.t3146 22.813
R4029 VDD.n2820 VDD.t13 22.813
R4030 VDD.n554 VDD.t4510 22.813
R4031 VDD.n3100 VDD.t2550 22.813
R4032 VDD.n3124 VDD.t1628 22.813
R4033 VDD.n3213 VDD.t1755 22.813
R4034 VDD.n3237 VDD.t427 22.813
R4035 VDD.n2175 VDD.t3802 20.998
R4036 VDD.n2159 VDD.t2384 20.998
R4037 VDD.n1462 VDD.t3922 20.998
R4038 VDD.n2039 VDD.t3035 20.998
R4039 VDD.n1939 VDD.t4025 20.998
R4040 VDD.n1889 VDD.t2305 20.998
R4041 VDD.n1914 VDD.t3391 20.998
R4042 VDD.n1964 VDD.t4375 20.998
R4043 VDD.n1989 VDD.t267 20.998
R4044 VDD.n2014 VDD.t3469 20.998
R4045 VDD.n2064 VDD.t3773 20.998
R4046 VDD.n2627 VDD.t3246 20.998
R4047 VDD.n2434 VDD.t3185 20.998
R4048 VDD.n2409 VDD.t3816 20.998
R4049 VDD.n2225 VDD.t1515 20.998
R4050 VDD.n2200 VDD.t3248 20.998
R4051 VDD.n601 VDD.t1109 20.186
R4052 VDD.n738 VDD.t3624 20.186
R4053 VDD.n3251 VDD.t1644 20.183
R4054 VDD.n2900 VDD.t3013 20.183
R4055 VDD.n2673 VDD.t1873 20.183
R4056 VDD.n2664 VDD.t2082 20.183
R4057 VDD.n411 VDD.t3446 20.183
R4058 VDD.n2928 VDD.t1469 20.183
R4059 VDD.n303 VDD.t1811 20.183
R4060 VDD.n294 VDD.t2422 20.183
R4061 VDD.n385 VDD.t1379 20.183
R4062 VDD.n394 VDD.t4409 20.183
R4063 VDD.n2654 VDD.t1841 20.183
R4064 VDD.n707 VDD.t1393 20.183
R4065 VDD.n2646 VDD.t1476 20.183
R4066 VDD.n699 VDD.t1322 20.183
R4067 VDD.n286 VDD.t4381 20.183
R4068 VDD.n276 VDD.t366 20.183
R4069 VDD.n265 VDD.t1054 20.183
R4070 VDD.n1075 VDD.t3734 20.183
R4071 VDD.n1108 VDD.t1391 20.183
R4072 VDD.n1058 VDD.t2226 20.183
R4073 VDD.t3194 VDD.n1036 17.506
R4074 VDD.t3264 VDD.n911 17.506
R4075 VDD.t3820 VDD.n936 17.506
R4076 VDD.t3825 VDD.n1011 17.506
R4077 VDD.t3865 VDD.n986 17.506
R4078 VDD.t2378 VDD.n961 17.506
R4079 VDD.t1735 VDD.n886 17.506
R4080 VDD.t3926 VDD.n862 17.506
R4081 VDD.n1730 VDD.t3276 17.506
R4082 VDD.n1755 VDD.t4011 17.506
R4083 VDD.n1855 VDD.t3947 17.506
R4084 VDD.n1830 VDD.t2244 17.506
R4085 VDD.n1805 VDD.t1505 17.506
R4086 VDD.n1780 VDD.t2046 17.506
R4087 VDD.n1705 VDD.t4039 17.506
R4088 VDD.n1681 VDD.t3259 17.506
R4089 VDD.n1530 VDD.t1162 17.506
R4090 VDD.n1555 VDD.t719 17.506
R4091 VDD.n1655 VDD.t1198 17.506
R4092 VDD.n1630 VDD.t699 17.506
R4093 VDD.n1605 VDD.t1196 17.506
R4094 VDD.n1580 VDD.t1192 17.506
R4095 VDD.n1505 VDD.t825 17.506
R4096 VDD.n1481 VDD.t1214 17.506
R4097 VDD.n1380 VDD.t3250 17.506
R4098 VDD.n1355 VDD.t2394 17.506
R4099 VDD.n1256 VDD.t2230 17.506
R4100 VDD.n1280 VDD.t4060 17.506
R4101 VDD.n1305 VDD.t3192 17.506
R4102 VDD.n1330 VDD.t3941 17.506
R4103 VDD.n1405 VDD.t3838 17.506
R4104 VDD.n1430 VDD.t3256 17.506
R4105 VDD.n2593 VDD.t4277 17.506
R4106 VDD.n2454 VDD.t3883 17.506
R4107 VDD.n2473 VDD.t3091 17.506
R4108 VDD.n2533 VDD.t3897 17.506
R4109 VDD.n2553 VDD.t4273 17.506
R4110 VDD.n2573 VDD.t3893 17.506
R4111 VDD.n2513 VDD.t4318 17.506
R4112 VDD.n2493 VDD.t3081 17.506
R4113 VDD.n2384 VDD.t859 17.506
R4114 VDD.n2245 VDD.t2965 17.506
R4115 VDD.n2264 VDD.t855 17.506
R4116 VDD.n2324 VDD.t2937 17.506
R4117 VDD.n2344 VDD.t2943 17.506
R4118 VDD.n2364 VDD.t837 17.506
R4119 VDD.n2304 VDD.t2947 17.506
R4120 VDD.n2284 VDD.t2931 17.506
R4121 VDD.n2688 VDD.t4020 14.284
R4122 VDD.n2869 VDD.t4199 14.284
R4123 VDD.n2753 VDD.t2636 14.284
R4124 VDD.n2841 VDD.t2780 14.284
R4125 VDD.n2816 VDD.t2668 14.284
R4126 VDD.n530 VDD.t1128 14.284
R4127 VDD.n559 VDD.t3476 14.284
R4128 VDD.n566 VDD.t1896 14.284
R4129 VDD.n3094 VDD.t2994 14.284
R4130 VDD.n376 VDD.t325 14.284
R4131 VDD.n3023 VDD.t2734 14.284
R4132 VDD.n3030 VDD.t309 14.284
R4133 VDD.n3207 VDD.t965 14.284
R4134 VDD.n2942 VDD.t410 14.284
R4135 VDD.n2948 VDD.t307 14.284
R4136 VDD.n2953 VDD.t3225 14.284
R4137 VDD.n2958 VDD.t2177 14.284
R4138 VDD.n2988 VDD.t3719 14.284
R4139 VDD.n2993 VDD.t4339 14.284
R4140 VDD.n3013 VDD.t3417 14.284
R4141 VDD.n3177 VDD.t2649 14.284
R4142 VDD.n3182 VDD.t251 14.284
R4143 VDD.n3164 VDD.t157 14.284
R4144 VDD.n3169 VDD.t513 14.284
R4145 VDD.n3077 VDD.t2592 14.284
R4146 VDD.n3082 VDD.t1069 14.284
R4147 VDD.n3058 VDD.t915 14.284
R4148 VDD.n3063 VDD.t1621 14.284
R4149 VDD.n724 VDD.t3617 14.284
R4150 VDD.n719 VDD.t2565 14.284
R4151 VDD.n594 VDD.t1112 14.284
R4152 VDD.n589 VDD.t4228 14.284
R4153 VDD.n580 VDD.t4458 14.284
R4154 VDD.n575 VDD.t4569 14.284
R4155 VDD.n258 VDD.t1057 14.284
R4156 VDD.n253 VDD.t1145 14.284
R4157 VDD.n3375 VDD.t1250 14.284
R4158 VDD.n3380 VDD.t259 14.284
R4159 VDD.n3323 VDD.t1757 14.284
R4160 VDD.n3318 VDD.t607 14.284
R4161 VDD.n201 VDD.t3187 14.284
R4162 VDD.n206 VDD.t990 14.284
R4163 VDD.n3266 VDD.t4197 14.284
R4164 VDD.n33 VDD.t1913 14.284
R4165 VDD.n38 VDD.t3600 14.284
R4166 VDD.n3 VDD.t1967 14.284
R4167 VDD.n8 VDD.t3691 14.284
R4168 VDD.n89 VDD.t64 14.284
R4169 VDD.n84 VDD.t2973 14.284
R4170 VDD.n143 VDD.t2715 14.284
R4171 VDD.n148 VDD.t3738 14.284
R4172 VDD.n180 VDD.t527 14.284
R4173 VDD.n185 VDD.t1310 14.284
R4174 VDD.n168 VDD.t763 14.284
R4175 VDD.n173 VDD.t4386 14.284
R4176 VDD.n121 VDD.t880 14.284
R4177 VDD.n126 VDD.t999 14.284
R4178 VDD.n109 VDD.t333 14.284
R4179 VDD.n114 VDD.t3960 14.284
R4180 VDD.n835 VDD.t1494 14.284
R4181 VDD.n840 VDD.t2318 14.284
R4182 VDD.n11 VDD.t520 14.284
R4183 VDD.n16 VDD.t1527 14.284
R4184 VDD.n70 VDD.t4077 14.284
R4185 VDD.n75 VDD.t2781 14.284
R4186 VDD.n58 VDD.t2291 14.284
R4187 VDD.n63 VDD.t3390 14.284
R4188 VDD.n3402 VDD.t2862 14.284
R4189 VDD.n3423 VDD.t1804 14.284
R4190 VDD.n3418 VDD.t3741 14.284
R4191 VDD.n3412 VDD.t3518 14.284
R4192 VDD.n3407 VDD.t3539 14.284
R4193 VDD.n3281 VDD.t1453 14.284
R4194 VDD.n3276 VDD.t3365 14.284
R4195 VDD.n3309 VDD.t3301 14.284
R4196 VDD.n3304 VDD.t4508 14.284
R4197 VDD.n3338 VDD.t670 14.284
R4198 VDD.n3333 VDD.t76 14.284
R4199 VDD.n3366 VDD.t2979 14.284
R4200 VDD.n3361 VDD.t1131 14.284
R4201 VDD.n214 VDD.t266 14.284
R4202 VDD.n209 VDD.t2514 14.284
R4203 VDD.n242 VDD.t977 14.284
R4204 VDD.n237 VDD.t4562 14.284
R4205 VDD.n358 VDD.t888 14.284
R4206 VDD.n363 VDD.t2816 14.284
R4207 VDD.n340 VDD.t2399 14.284
R4208 VDD.n345 VDD.t1559 14.284
R4209 VDD.n458 VDD.t564 14.284
R4210 VDD.n463 VDD.t1641 14.284
R4211 VDD.n439 VDD.t491 14.284
R4212 VDD.n444 VDD.t624 14.284
R4213 VDD.n470 VDD.t4255 14.284
R4214 VDD.n475 VDD.t86 14.284
R4215 VDD.n507 VDD.t1233 14.284
R4216 VDD.n512 VDD.t779 14.284
R4217 VDD.n2757 VDD.t4425 14.284
R4218 VDD.n2762 VDD.t4171 14.284
R4219 VDD.n2791 VDD.t4099 14.284
R4220 VDD.n2796 VDD.t1672 14.284
R4221 VDD.n2693 VDD.t1754 14.284
R4222 VDD.n2698 VDD.t1946 14.284
R4223 VDD.n2728 VDD.t3561 14.284
R4224 VDD.n2733 VDD.t182 14.284
R4225 VDD.n2182 VDD.t3878 14.284
R4226 VDD.n2168 VDD.t434 14.284
R4227 VDD.n2150 VDD.t4143 14.284
R4228 VDD.n2145 VDD.t1742 14.284
R4229 VDD.n1469 VDD.t3944 14.284
R4230 VDD.n1455 VDD.t2197 14.284
R4231 VDD.n2030 VDD.t1396 14.284
R4232 VDD.n2045 VDD.t1441 14.284
R4233 VDD.n1930 VDD.t3727 14.284
R4234 VDD.n1945 VDD.t3962 14.284
R4235 VDD.n1880 VDD.t2205 14.284
R4236 VDD.n1895 VDD.t2317 14.284
R4237 VDD.n1905 VDD.t2475 14.284
R4238 VDD.n1920 VDD.t192 14.284
R4239 VDD.n1955 VDD.t2652 14.284
R4240 VDD.n1970 VDD.t3547 14.284
R4241 VDD.n1980 VDD.t921 14.284
R4242 VDD.n1995 VDD.t283 14.284
R4243 VDD.n2005 VDD.t2411 14.284
R4244 VDD.n2020 VDD.t3431 14.284
R4245 VDD.n2055 VDD.t1549 14.284
R4246 VDD.n2070 VDD.t3745 14.284
R4247 VDD.n1164 VDD.t2442 14.284
R4248 VDD.n1179 VDD.t929 14.284
R4249 VDD.n1224 VDD.t2606 14.284
R4250 VDD.n1209 VDD.t1412 14.284
R4251 VDD.n1194 VDD.t1848 14.284
R4252 VDD.n1152 VDD.t3729 14.284
R4253 VDD.n1137 VDD.t2469 14.284
R4254 VDD.n1242 VDD.t2199 14.284
R4255 VDD.n2618 VDD.t1547 14.284
R4256 VDD.n2613 VDD.t1740 14.284
R4257 VDD.n2441 VDD.t3269 14.284
R4258 VDD.n2427 VDD.t3314 14.284
R4259 VDD.n2416 VDD.t3253 14.284
R4260 VDD.n2402 VDD.t1816 14.284
R4261 VDD.n2232 VDD.t3856 14.284
R4262 VDD.n2218 VDD.t1872 14.284
R4263 VDD.n2207 VDD.t1514 14.284
R4264 VDD.n2193 VDD.t2660 14.284
R4265 VDD.n1041 VDD.t1524 14.283
R4266 VDD.n916 VDD.t1802 14.283
R4267 VDD.n941 VDD.t1340 14.283
R4268 VDD.n1016 VDD.t3812 14.283
R4269 VDD.n991 VDD.t1768 14.283
R4270 VDD.n966 VDD.t3213 14.283
R4271 VDD.n891 VDD.t3338 14.283
R4272 VDD.n867 VDD.t1738 14.283
R4273 VDD.n637 VDD.t712 14.283
R4274 VDD.n655 VDD.t834 14.283
R4275 VDD.n673 VDD.t1195 14.283
R4276 VDD.n690 VDD.t726 14.283
R4277 VDD.n619 VDD.t1175 14.283
R4278 VDD.n750 VDD.t732 14.283
R4279 VDD.n768 VDD.t800 14.283
R4280 VDD.n786 VDD.t714 14.283
R4281 VDD.n1742 VDD.t1725 14.283
R4282 VDD.n1767 VDD.t3808 14.283
R4283 VDD.n1860 VDD.t3876 14.283
R4284 VDD.n1835 VDD.t3255 14.283
R4285 VDD.n1817 VDD.t3806 14.283
R4286 VDD.n1792 VDD.t3815 14.283
R4287 VDD.n1717 VDD.t1338 14.283
R4288 VDD.n1693 VDD.t3221 14.283
R4289 VDD.n1535 VDD.t702 14.283
R4290 VDD.n1560 VDD.t690 14.283
R4291 VDD.n1660 VDD.t1181 14.283
R4292 VDD.n1635 VDD.t4362 14.283
R4293 VDD.n1610 VDD.t708 14.283
R4294 VDD.n1585 VDD.t1177 14.283
R4295 VDD.n1510 VDD.t808 14.283
R4296 VDD.n1486 VDD.t730 14.283
R4297 VDD.n1385 VDD.t1727 14.283
R4298 VDD.n1360 VDD.t2373 14.283
R4299 VDD.n1261 VDD.t2045 14.283
R4300 VDD.n1285 VDD.t3847 14.283
R4301 VDD.n1310 VDD.t3852 14.283
R4302 VDD.n1335 VDD.t4004 14.283
R4303 VDD.n1410 VDD.t3824 14.283
R4304 VDD.n1435 VDD.t2383 14.283
R4305 VDD.n2603 VDD.t3900 14.283
R4306 VDD.n2464 VDD.t4317 14.283
R4307 VDD.n2483 VDD.t3096 14.283
R4308 VDD.n2543 VDD.t4329 14.283
R4309 VDD.n2563 VDD.t4307 14.283
R4310 VDD.n2583 VDD.t3080 14.283
R4311 VDD.n2523 VDD.t3090 14.283
R4312 VDD.n2503 VDD.t3100 14.283
R4313 VDD.n2387 VDD.t872 14.283
R4314 VDD.n2255 VDD.t840 14.283
R4315 VDD.n2274 VDD.t858 14.283
R4316 VDD.n2327 VDD.t2924 14.283
R4317 VDD.n2347 VDD.t842 14.283
R4318 VDD.n2367 VDD.t844 14.283
R4319 VDD.n2314 VDD.t848 14.283
R4320 VDD.n2294 VDD.t864 14.283
R4321 VDD.n1049 VDD.t3396 14.283
R4322 VDD.n924 VDD.t3029 14.283
R4323 VDD.n949 VDD.t3464 14.283
R4324 VDD.n1024 VDD.t3994 14.283
R4325 VDD.n999 VDD.t4407 14.283
R4326 VDD.n974 VDD.t287 14.283
R4327 VDD.n899 VDD.t3780 14.283
R4328 VDD.n875 VDD.t4600 14.283
R4329 VDD.n633 VDD.t3858 14.283
R4330 VDD.n651 VDD.t1610 14.283
R4331 VDD.n669 VDD.t2700 14.283
R4332 VDD.n686 VDD.t3862 14.283
R4333 VDD.n615 VDD.t561 14.283
R4334 VDD.n746 VDD.t453 14.283
R4335 VDD.n764 VDD.t2785 14.283
R4336 VDD.n782 VDD.t2848 14.283
R4337 VDD.n1738 VDD.t2110 14.283
R4338 VDD.n1763 VDD.t1098 14.283
R4339 VDD.n1868 VDD.t2732 14.283
R4340 VDD.n1843 VDD.t4594 14.283
R4341 VDD.n1813 VDD.t1695 14.283
R4342 VDD.n1788 VDD.t4450 14.283
R4343 VDD.n1713 VDD.t49 14.283
R4344 VDD.n1689 VDD.t1719 14.283
R4345 VDD.n1543 VDD.t4488 14.283
R4346 VDD.n1568 VDD.t1296 14.283
R4347 VDD.n1668 VDD.t4206 14.283
R4348 VDD.n1643 VDD.t38 14.283
R4349 VDD.n1618 VDD.t3684 14.283
R4350 VDD.n1593 VDD.t1090 14.283
R4351 VDD.n1518 VDD.t2256 14.283
R4352 VDD.n1494 VDD.t2500 14.283
R4353 VDD.n1393 VDD.t445 14.283
R4354 VDD.n1368 VDD.t3422 14.283
R4355 VDD.n1269 VDD.t383 14.283
R4356 VDD.n1293 VDD.t2102 14.283
R4357 VDD.n1318 VDD.t3375 14.283
R4358 VDD.n1343 VDD.t3334 14.283
R4359 VDD.n1418 VDD.t2751 14.283
R4360 VDD.n1443 VDD.t4479 14.283
R4361 VDD.n2599 VDD.t3320 14.283
R4362 VDD.n2460 VDD.t2723 14.283
R4363 VDD.n2479 VDD.t297 14.283
R4364 VDD.n2539 VDD.t133 14.283
R4365 VDD.n2559 VDD.t3527 14.283
R4366 VDD.n2579 VDD.t2825 14.283
R4367 VDD.n2519 VDD.t1593 14.283
R4368 VDD.n2499 VDD.t2772 14.283
R4369 VDD.n2395 VDD.t3167 14.283
R4370 VDD.n2251 VDD.t587 14.283
R4371 VDD.n2270 VDD.t1051 14.283
R4372 VDD.n2335 VDD.t2281 14.283
R4373 VDD.n2355 VDD.t464 14.283
R4374 VDD.n2375 VDD.t1269 14.283
R4375 VDD.n2310 VDD.t319 14.283
R4376 VDD.n2290 VDD.t2058 14.283
R4377 VDD.n1047 VDD.t1929 14.282
R4378 VDD.n1047 VDD.t1927 14.282
R4379 VDD.n1040 VDD.t3195 14.282
R4380 VDD.n1040 VDD.t1526 14.282
R4381 VDD.n922 VDD.t3020 14.282
R4382 VDD.n922 VDD.t3008 14.282
R4383 VDD.n915 VDD.t3265 14.282
R4384 VDD.n915 VDD.t1730 14.282
R4385 VDD.n947 VDD.t3462 14.282
R4386 VDD.n947 VDD.t3460 14.282
R4387 VDD.n940 VDD.t3821 14.282
R4388 VDD.n940 VDD.t3872 14.282
R4389 VDD.n1022 VDD.t3973 14.282
R4390 VDD.n1022 VDD.t3971 14.282
R4391 VDD.n1015 VDD.t3826 14.282
R4392 VDD.n1015 VDD.t3682 14.282
R4393 VDD.n997 VDD.t4412 14.282
R4394 VDD.n997 VDD.t1317 14.282
R4395 VDD.n990 VDD.t3866 14.282
R4396 VDD.n990 VDD.t3950 14.282
R4397 VDD.n972 VDD.t285 14.282
R4398 VDD.n972 VDD.t281 14.282
R4399 VDD.n965 VDD.t2379 14.282
R4400 VDD.n965 VDD.t2369 14.282
R4401 VDD.n897 VDD.t3764 14.282
R4402 VDD.n897 VDD.t3768 14.282
R4403 VDD.n890 VDD.t1736 14.282
R4404 VDD.n890 VDD.t4044 14.282
R4405 VDD.n873 VDD.t4605 14.282
R4406 VDD.n873 VDD.t4607 14.282
R4407 VDD.n866 VDD.t3927 14.282
R4408 VDD.n866 VDD.t4008 14.282
R4409 VDD.n2685 VDD.t4022 14.282
R4410 VDD.n2685 VDD.t4018 14.282
R4411 VDD.n2866 VDD.t4 14.282
R4412 VDD.n2866 VDD.t6 14.282
R4413 VDD.n2750 VDD.t2632 14.282
R4414 VDD.n2750 VDD.t2634 14.282
R4415 VDD.n2838 VDD.t2776 14.282
R4416 VDD.n2838 VDD.t2778 14.282
R4417 VDD.n2813 VDD.t2664 14.282
R4418 VDD.n2813 VDD.t2666 14.282
R4419 VDD.n527 VDD.t2860 14.282
R4420 VDD.n527 VDD.t2858 14.282
R4421 VDD.n560 VDD.t3478 14.282
R4422 VDD.n560 VDD.t3474 14.282
R4423 VDD.n567 VDD.t1894 14.282
R4424 VDD.n567 VDD.t1898 14.282
R4425 VDD.n3091 VDD.t2990 14.282
R4426 VDD.n3091 VDD.t2992 14.282
R4427 VDD.n373 VDD.t329 14.282
R4428 VDD.n373 VDD.t327 14.282
R4429 VDD.n3020 VDD.t580 14.282
R4430 VDD.n3020 VDD.t582 14.282
R4431 VDD.n3027 VDD.t2626 14.282
R4432 VDD.n3027 VDD.t2628 14.282
R4433 VDD.n3204 VDD.t660 14.282
R4434 VDD.n3204 VDD.t658 14.282
R4435 VDD.n2939 VDD.t40 14.282
R4436 VDD.n2939 VDD.t408 14.282
R4437 VDD.n2945 VDD.t1123 14.282
R4438 VDD.n2945 VDD.t1125 14.282
R4439 VDD.n2952 VDD.t3229 14.282
R4440 VDD.n2952 VDD.t3125 14.282
R4441 VDD.n2957 VDD.t1664 14.282
R4442 VDD.n2957 VDD.t2252 14.282
R4443 VDD.n2987 VDD.t3703 14.282
R4444 VDD.n2987 VDD.t3707 14.282
R4445 VDD.n2992 VDD.t4347 14.282
R4446 VDD.n2992 VDD.t951 14.282
R4447 VDD.n3010 VDD.t2120 14.282
R4448 VDD.n3010 VDD.t3415 14.282
R4449 VDD.n3176 VDD.t4439 14.282
R4450 VDD.n3176 VDD.t2643 14.282
R4451 VDD.n3181 VDD.t235 14.282
R4452 VDD.n3181 VDD.t241 14.282
R4453 VDD.n3163 VDD.t161 14.282
R4454 VDD.n3163 VDD.t173 14.282
R4455 VDD.n3168 VDD.t3801 14.282
R4456 VDD.n3168 VDD.t3592 14.282
R4457 VDD.n3076 VDD.t1533 14.282
R4458 VDD.n3076 VDD.t2594 14.282
R4459 VDD.n3081 VDD.t1077 14.282
R4460 VDD.n3081 VDD.t4289 14.282
R4461 VDD.n3057 VDD.t901 14.282
R4462 VDD.n3057 VDD.t911 14.282
R4463 VDD.n3062 VDD.t2269 14.282
R4464 VDD.n3062 VDD.t1617 14.282
R4465 VDD.n723 VDD.t3623 14.282
R4466 VDD.n723 VDD.t3619 14.282
R4467 VDD.n718 VDD.t2563 14.282
R4468 VDD.n718 VDD.t2561 14.282
R4469 VDD.n636 VDD.t812 14.282
R4470 VDD.n636 VDD.t1209 14.282
R4471 VDD.n632 VDD.t556 14.282
R4472 VDD.n632 VDD.t554 14.282
R4473 VDD.n654 VDD.t736 14.282
R4474 VDD.n654 VDD.t792 14.282
R4475 VDD.n650 VDD.t1608 14.282
R4476 VDD.n650 VDD.t1606 14.282
R4477 VDD.n672 VDD.t1161 14.282
R4478 VDD.n672 VDD.t794 14.282
R4479 VDD.n668 VDD.t2698 14.282
R4480 VDD.n668 VDD.t606 14.282
R4481 VDD.n689 VDD.t692 14.282
R4482 VDD.n689 VDD.t1227 14.282
R4483 VDD.n685 VDD.t3860 14.282
R4484 VDD.n685 VDD.t3864 14.282
R4485 VDD.n593 VDD.t3484 14.282
R4486 VDD.n593 VDD.t3492 14.282
R4487 VDD.n588 VDD.t4234 14.282
R4488 VDD.n588 VDD.t4224 14.282
R4489 VDD.n579 VDD.t361 14.282
R4490 VDD.n579 VDD.t4456 14.282
R4491 VDD.n574 VDD.t4575 14.282
R4492 VDD.n574 VDD.t4583 14.282
R4493 VDD.n257 VDD.t469 14.282
R4494 VDD.n257 VDD.t477 14.282
R4495 VDD.n252 VDD.t1151 14.282
R4496 VDD.n252 VDD.t1141 14.282
R4497 VDD.n618 VDD.t1225 14.282
R4498 VDD.n618 VDD.t688 14.282
R4499 VDD.n614 VDD.t357 14.282
R4500 VDD.n614 VDD.t3523 14.282
R4501 VDD.n749 VDD.t1201 14.282
R4502 VDD.n749 VDD.t1165 14.282
R4503 VDD.n745 VDD.t451 14.282
R4504 VDD.n745 VDD.t449 14.282
R4505 VDD.n767 VDD.t1171 14.282
R4506 VDD.n767 VDD.t740 14.282
R4507 VDD.n763 VDD.t2789 14.282
R4508 VDD.n763 VDD.t2787 14.282
R4509 VDD.n785 VDD.t824 14.282
R4510 VDD.n785 VDD.t1223 14.282
R4511 VDD.n781 VDD.t2846 14.282
R4512 VDD.n781 VDD.t2850 14.282
R4513 VDD.n3372 VDD.t1252 14.282
R4514 VDD.n3372 VDD.t1251 14.282
R4515 VDD.n3377 VDD.t258 14.282
R4516 VDD.n3377 VDD.t257 14.282
R4517 VDD.n3320 VDD.t1759 14.282
R4518 VDD.n3320 VDD.t1758 14.282
R4519 VDD.n3315 VDD.t609 14.282
R4520 VDD.n3315 VDD.t608 14.282
R4521 VDD.n198 VDD.t3189 14.282
R4522 VDD.n198 VDD.t3188 14.282
R4523 VDD.n203 VDD.t989 14.282
R4524 VDD.n203 VDD.t991 14.282
R4525 VDD.n3263 VDD.t1351 14.282
R4526 VDD.n3263 VDD.t4196 14.282
R4527 VDD.n30 VDD.t2640 14.282
R4528 VDD.n30 VDD.t1914 14.282
R4529 VDD.n35 VDD.t3601 14.282
R4530 VDD.n35 VDD.t3602 14.282
R4531 VDD.n0 VDD.t1966 14.282
R4532 VDD.n0 VDD.t1965 14.282
R4533 VDD.n5 VDD.t2799 14.282
R4534 VDD.n5 VDD.t3692 14.282
R4535 VDD.n86 VDD.t63 14.282
R4536 VDD.n86 VDD.t62 14.282
R4537 VDD.n81 VDD.t2975 14.282
R4538 VDD.n81 VDD.t2974 14.282
R4539 VDD.n140 VDD.t497 14.282
R4540 VDD.n140 VDD.t496 14.282
R4541 VDD.n145 VDD.t2363 14.282
R4542 VDD.n145 VDD.t3739 14.282
R4543 VDD.n179 VDD.t529 14.282
R4544 VDD.n179 VDD.t528 14.282
R4545 VDD.n184 VDD.t1304 14.282
R4546 VDD.n184 VDD.t1303 14.282
R4547 VDD.n167 VDD.t765 14.282
R4548 VDD.n167 VDD.t764 14.282
R4549 VDD.n172 VDD.t4418 14.282
R4550 VDD.n172 VDD.t3542 14.282
R4551 VDD.n120 VDD.t882 14.282
R4552 VDD.n120 VDD.t881 14.282
R4553 VDD.n125 VDD.t998 14.282
R4554 VDD.n125 VDD.t1000 14.282
R4555 VDD.n108 VDD.t336 14.282
R4556 VDD.n108 VDD.t334 14.282
R4557 VDD.n113 VDD.t3958 14.282
R4558 VDD.n113 VDD.t3957 14.282
R4559 VDD.n834 VDD.t1497 14.282
R4560 VDD.n834 VDD.t1495 14.282
R4561 VDD.n839 VDD.t2336 14.282
R4562 VDD.n839 VDD.t2295 14.282
R4563 VDD.n10 VDD.t522 14.282
R4564 VDD.n10 VDD.t521 14.282
R4565 VDD.n15 VDD.t2365 14.282
R4566 VDD.n15 VDD.t1728 14.282
R4567 VDD.n69 VDD.t4079 14.282
R4568 VDD.n69 VDD.t4078 14.282
R4569 VDD.n74 VDD.t2568 14.282
R4570 VDD.n74 VDD.t2567 14.282
R4571 VDD.n57 VDD.t255 14.282
R4572 VDD.n57 VDD.t254 14.282
R4573 VDD.n62 VDD.t150 14.282
R4574 VDD.n62 VDD.t147 14.282
R4575 VDD.n3399 VDD.t3234 14.282
R4576 VDD.n3399 VDD.t2863 14.282
R4577 VDD.n3422 VDD.t1803 14.282
R4578 VDD.n3422 VDD.t1602 14.282
R4579 VDD.n3417 VDD.t3754 14.282
R4580 VDD.n3417 VDD.t3743 14.282
R4581 VDD.n3411 VDD.t3517 14.282
R4582 VDD.n3411 VDD.t1267 14.282
R4583 VDD.n3406 VDD.t1655 14.282
R4584 VDD.n3406 VDD.t3538 14.282
R4585 VDD.n3280 VDD.t1471 14.282
R4586 VDD.n3280 VDD.t1468 14.282
R4587 VDD.n3275 VDD.t3110 14.282
R4588 VDD.n3275 VDD.t3109 14.282
R4589 VDD.n3308 VDD.t3294 14.282
R4590 VDD.n3308 VDD.t3302 14.282
R4591 VDD.n3303 VDD.t4507 14.282
R4592 VDD.n3303 VDD.t4506 14.282
R4593 VDD.n3337 VDD.t2075 14.282
R4594 VDD.n3337 VDD.t2074 14.282
R4595 VDD.n3332 VDD.t3135 14.282
R4596 VDD.n3332 VDD.t3134 14.282
R4597 VDD.n3365 VDD.t2983 14.282
R4598 VDD.n3365 VDD.t2982 14.282
R4599 VDD.n3360 VDD.t1130 14.282
R4600 VDD.n3360 VDD.t1129 14.282
R4601 VDD.n213 VDD.t1997 14.282
R4602 VDD.n213 VDD.t271 14.282
R4603 VDD.n208 VDD.t2513 14.282
R4604 VDD.n208 VDD.t2512 14.282
R4605 VDD.n241 VDD.t983 14.282
R4606 VDD.n241 VDD.t978 14.282
R4607 VDD.n236 VDD.t4563 14.282
R4608 VDD.n236 VDD.t4564 14.282
R4609 VDD.n357 VDD.t892 14.282
R4610 VDD.n357 VDD.t884 14.282
R4611 VDD.n362 VDD.t3580 14.282
R4612 VDD.n362 VDD.t2812 14.282
R4613 VDD.n339 VDD.t2403 14.282
R4614 VDD.n339 VDD.t4529 14.282
R4615 VDD.n344 VDD.t3413 14.282
R4616 VDD.n344 VDD.t3409 14.282
R4617 VDD.n457 VDD.t568 14.282
R4618 VDD.n457 VDD.t572 14.282
R4619 VDD.n462 VDD.t1703 14.282
R4620 VDD.n462 VDD.t1709 14.282
R4621 VDD.n438 VDD.t1315 14.282
R4622 VDD.n438 VDD.t4468 14.282
R4623 VDD.n443 VDD.t1021 14.282
R4624 VDD.n443 VDD.t1025 14.282
R4625 VDD.n469 VDD.t1502 14.282
R4626 VDD.n469 VDD.t4257 14.282
R4627 VDD.n474 VDD.t96 14.282
R4628 VDD.n474 VDD.t102 14.282
R4629 VDD.n506 VDD.t1237 14.282
R4630 VDD.n506 VDD.t680 14.282
R4631 VDD.n511 VDD.t785 14.282
R4632 VDD.n511 VDD.t974 14.282
R4633 VDD.n2756 VDD.t4429 14.282
R4634 VDD.n2756 VDD.t4433 14.282
R4635 VDD.n2761 VDD.t4157 14.282
R4636 VDD.n2761 VDD.t4165 14.282
R4637 VDD.n2790 VDD.t4107 14.282
R4638 VDD.n2790 VDD.t4091 14.282
R4639 VDD.n2795 VDD.t1686 14.282
R4640 VDD.n2795 VDD.t1670 14.282
R4641 VDD.n2692 VDD.t3661 14.282
R4642 VDD.n2692 VDD.t3665 14.282
R4643 VDD.n2697 VDD.t1952 14.282
R4644 VDD.n2697 VDD.t1938 14.282
R4645 VDD.n2727 VDD.t207 14.282
R4646 VDD.n2727 VDD.t213 14.282
R4647 VDD.n2732 VDD.t2706 14.282
R4648 VDD.n2732 VDD.t180 14.282
R4649 VDD.n2181 VDD.t2037 14.282
R4650 VDD.n2181 VDD.t3803 14.282
R4651 VDD.n2167 VDD.t3725 14.282
R4652 VDD.n2167 VDD.t440 14.282
R4653 VDD.n2149 VDD.t2461 14.282
R4654 VDD.n2149 VDD.t4139 14.282
R4655 VDD.n2147 VDD.t2881 14.282
R4656 VDD.n2147 VDD.t2385 14.282
R4657 VDD.n1468 VDD.t1808 14.282
R4658 VDD.n1468 VDD.t3923 14.282
R4659 VDD.n1454 VDD.t2223 14.282
R4660 VDD.n1454 VDD.t2211 14.282
R4661 VDD.n2029 VDD.t3308 14.282
R4662 VDD.n2029 VDD.t3306 14.282
R4663 VDD.n2044 VDD.t1465 14.282
R4664 VDD.n2044 VDD.t3036 14.282
R4665 VDD.n1929 VDD.t438 14.282
R4666 VDD.n1929 VDD.t1361 14.282
R4667 VDD.n1944 VDD.t3986 14.282
R4668 VDD.n1944 VDD.t4026 14.282
R4669 VDD.n1879 VDD.t2209 14.282
R4670 VDD.n1879 VDD.t2217 14.282
R4671 VDD.n1894 VDD.t2327 14.282
R4672 VDD.n1894 VDD.t2306 14.282
R4673 VDD.n1904 VDD.t2471 14.282
R4674 VDD.n1904 VDD.t2467 14.282
R4675 VDD.n1919 VDD.t1923 14.282
R4676 VDD.n1919 VDD.t3392 14.282
R4677 VDD.n1954 VDD.t2434 14.282
R4678 VDD.n1954 VDD.t4130 14.282
R4679 VDD.n1969 VDD.t4384 14.282
R4680 VDD.n1969 VDD.t4376 14.282
R4681 VDD.n1979 VDD.t937 14.282
R4682 VDD.n1979 VDD.t923 14.282
R4683 VDD.n1994 VDD.t2008 14.282
R4684 VDD.n1994 VDD.t268 14.282
R4685 VDD.n2004 VDD.t4111 14.282
R4686 VDD.n2004 VDD.t1820 14.282
R4687 VDD.n2019 VDD.t2096 14.282
R4688 VDD.n2019 VDD.t3470 14.282
R4689 VDD.n2054 VDD.t1551 14.282
R4690 VDD.n2054 VDD.t2618 14.282
R4691 VDD.n2069 VDD.t3758 14.282
R4692 VDD.n2069 VDD.t3774 14.282
R4693 VDD.n1741 VDD.t3277 14.282
R4694 VDD.n1741 VDD.t3271 14.282
R4695 VDD.n1737 VDD.t1613 14.282
R4696 VDD.n1737 VDD.t1615 14.282
R4697 VDD.n1766 VDD.t4012 14.282
R4698 VDD.n1766 VDD.t3850 14.282
R4699 VDD.n1762 VDD.t1100 14.282
R4700 VDD.n1762 VDD.t1096 14.282
R4701 VDD.n1867 VDD.t4065 14.282
R4702 VDD.n1867 VDD.t4067 14.282
R4703 VDD.n1859 VDD.t3948 14.282
R4704 VDD.n1859 VDD.t2367 14.282
R4705 VDD.n1842 VDD.t4596 14.282
R4706 VDD.n1842 VDD.t4592 14.282
R4707 VDD.n1834 VDD.t2245 14.282
R4708 VDD.n1834 VDD.t4042 14.282
R4709 VDD.n1816 VDD.t1506 14.282
R4710 VDD.n1816 VDD.t1734 14.282
R4711 VDD.n1812 VDD.t1697 14.282
R4712 VDD.n1812 VDD.t1693 14.282
R4713 VDD.n1791 VDD.t2047 14.282
R4714 VDD.n1791 VDD.t2247 14.282
R4715 VDD.n1787 VDD.t4454 14.282
R4716 VDD.n1787 VDD.t4452 14.282
R4717 VDD.n1716 VDD.t4040 14.282
R4718 VDD.n1716 VDD.t3197 14.282
R4719 VDD.n1712 VDD.t45 14.282
R4720 VDD.n1712 VDD.t47 14.282
R4721 VDD.n1692 VDD.t3260 14.282
R4722 VDD.n1692 VDD.t3184 14.282
R4723 VDD.n1688 VDD.t1715 14.282
R4724 VDD.n1688 VDD.t1717 14.282
R4725 VDD.n1542 VDD.t4486 14.282
R4726 VDD.n1542 VDD.t4484 14.282
R4727 VDD.n1534 VDD.t1163 14.282
R4728 VDD.n1534 VDD.t706 14.282
R4729 VDD.n1567 VDD.t1294 14.282
R4730 VDD.n1567 VDD.t1292 14.282
R4731 VDD.n1559 VDD.t720 14.282
R4732 VDD.n1559 VDD.t820 14.282
R4733 VDD.n1667 VDD.t4210 14.282
R4734 VDD.n1667 VDD.t4208 14.282
R4735 VDD.n1659 VDD.t1199 14.282
R4736 VDD.n1659 VDD.t1191 14.282
R4737 VDD.n1642 VDD.t36 14.282
R4738 VDD.n1642 VDD.t34 14.282
R4739 VDD.n1634 VDD.t700 14.282
R4740 VDD.n1634 VDD.t696 14.282
R4741 VDD.n1617 VDD.t3688 14.282
R4742 VDD.n1617 VDD.t3686 14.282
R4743 VDD.n1609 VDD.t1197 14.282
R4744 VDD.n1609 VDD.t710 14.282
R4745 VDD.n1592 VDD.t1094 14.282
R4746 VDD.n1592 VDD.t1092 14.282
R4747 VDD.n1584 VDD.t1193 14.282
R4748 VDD.n1584 VDD.t1183 14.282
R4749 VDD.n1517 VDD.t2254 14.282
R4750 VDD.n1517 VDD.t1102 14.282
R4751 VDD.n1509 VDD.t826 14.282
R4752 VDD.n1509 VDD.t818 14.282
R4753 VDD.n1493 VDD.t2504 14.282
R4754 VDD.n1493 VDD.t2502 14.282
R4755 VDD.n1485 VDD.t1215 14.282
R4756 VDD.n1485 VDD.t738 14.282
R4757 VDD.n1392 VDD.t443 14.282
R4758 VDD.n1392 VDD.t447 14.282
R4759 VDD.n1384 VDD.t3251 14.282
R4760 VDD.n1384 VDD.t3913 14.282
R4761 VDD.n1367 VDD.t3420 14.282
R4762 VDD.n1367 VDD.t3424 14.282
R4763 VDD.n1359 VDD.t2395 14.282
R4764 VDD.n1359 VDD.t2387 14.282
R4765 VDD.n1268 VDD.t381 14.282
R4766 VDD.n1268 VDD.t379 14.282
R4767 VDD.n1260 VDD.t2231 14.282
R4768 VDD.n1260 VDD.t1508 14.282
R4769 VDD.n1292 VDD.t2106 14.282
R4770 VDD.n1292 VDD.t2104 14.282
R4771 VDD.n1284 VDD.t4061 14.282
R4772 VDD.n1284 VDD.t3843 14.282
R4773 VDD.n1317 VDD.t3373 14.282
R4774 VDD.n1317 VDD.t3377 14.282
R4775 VDD.n1309 VDD.t3193 14.282
R4776 VDD.n1309 VDD.t3917 14.282
R4777 VDD.n1342 VDD.t4190 14.282
R4778 VDD.n1342 VDD.t3336 14.282
R4779 VDD.n1334 VDD.t3942 14.282
R4780 VDD.n1334 VDD.t3845 14.282
R4781 VDD.n1417 VDD.t2749 14.282
R4782 VDD.n1417 VDD.t2747 14.282
R4783 VDD.n1409 VDD.t3839 14.282
R4784 VDD.n1409 VDD.t4057 14.282
R4785 VDD.n1442 VDD.t4477 14.282
R4786 VDD.n1442 VDD.t4475 14.282
R4787 VDD.n1434 VDD.t3257 14.282
R4788 VDD.n1434 VDD.t2393 14.282
R4789 VDD.n1161 VDD.t4126 14.282
R4790 VDD.n1161 VDD.t4124 14.282
R4791 VDD.n1176 VDD.t1884 14.282
R4792 VDD.n1176 VDD.t1866 14.282
R4793 VDD.n1221 VDD.t2616 14.282
R4794 VDD.n1221 VDD.t2610 14.282
R4795 VDD.n1206 VDD.t1416 14.282
R4796 VDD.n1206 VDD.t1414 14.282
R4797 VDD.n1191 VDD.t2415 14.282
R4798 VDD.n1191 VDD.t1826 14.282
R4799 VDD.n1149 VDD.t436 14.282
R4800 VDD.n1149 VDD.t3733 14.282
R4801 VDD.n1134 VDD.t2457 14.282
R4802 VDD.n1134 VDD.t4137 14.282
R4803 VDD.n1239 VDD.t2203 14.282
R4804 VDD.n1239 VDD.t2201 14.282
R4805 VDD.n2617 VDD.t2600 14.282
R4806 VDD.n2617 VDD.t2614 14.282
R4807 VDD.n2612 VDD.t3854 14.282
R4808 VDD.n2612 VDD.t3247 14.282
R4809 VDD.n2440 VDD.t1732 14.282
R4810 VDD.n2440 VDD.t3186 14.282
R4811 VDD.n2426 VDD.t1400 14.282
R4812 VDD.n2426 VDD.t1410 14.282
R4813 VDD.n2415 VDD.t1778 14.282
R4814 VDD.n2415 VDD.t3817 14.282
R4815 VDD.n2401 VDD.t4113 14.282
R4816 VDD.n2401 VDD.t2413 14.282
R4817 VDD.n2231 VDD.t4006 14.282
R4818 VDD.n2231 VDD.t1516 14.282
R4819 VDD.n2217 VDD.t1864 14.282
R4820 VDD.n2217 VDD.t925 14.282
R4821 VDD.n2206 VDD.t1800 14.282
R4822 VDD.n2206 VDD.t3249 14.282
R4823 VDD.n2192 VDD.t2436 14.282
R4824 VDD.n2192 VDD.t2425 14.282
R4825 VDD.n2602 VDD.t4280 14.282
R4826 VDD.n2602 VDD.t4278 14.282
R4827 VDD.n2598 VDD.t2910 14.282
R4828 VDD.n2598 VDD.t2912 14.282
R4829 VDD.n2463 VDD.t4313 14.282
R4830 VDD.n2463 VDD.t3884 14.282
R4831 VDD.n2459 VDD.t2727 14.282
R4832 VDD.n2459 VDD.t2725 14.282
R4833 VDD.n2482 VDD.t3094 14.282
R4834 VDD.n2482 VDD.t3092 14.282
R4835 VDD.n2478 VDD.t299 14.282
R4836 VDD.n2478 VDD.t295 14.282
R4837 VDD.n2542 VDD.t3902 14.282
R4838 VDD.n2542 VDD.t3898 14.282
R4839 VDD.n2538 VDD.t131 14.282
R4840 VDD.n2538 VDD.t2453 14.282
R4841 VDD.n2562 VDD.t4276 14.282
R4842 VDD.n2562 VDD.t4274 14.282
R4843 VDD.n2558 VDD.t2532 14.282
R4844 VDD.n2558 VDD.t2530 14.282
R4845 VDD.n2582 VDD.t4333 14.282
R4846 VDD.n2582 VDD.t3894 14.282
R4847 VDD.n2578 VDD.t2829 14.282
R4848 VDD.n2578 VDD.t2827 14.282
R4849 VDD.n2522 VDD.t3088 14.282
R4850 VDD.n2522 VDD.t4319 14.282
R4851 VDD.n2518 VDD.t1591 14.282
R4852 VDD.n2518 VDD.t1589 14.282
R4853 VDD.n2502 VDD.t3084 14.282
R4854 VDD.n2502 VDD.t3082 14.282
R4855 VDD.n2498 VDD.t2118 14.282
R4856 VDD.n2498 VDD.t2774 14.282
R4857 VDD.n2394 VDD.t3171 14.282
R4858 VDD.n2394 VDD.t3169 14.282
R4859 VDD.n2386 VDD.t2946 14.282
R4860 VDD.n2386 VDD.t860 14.282
R4861 VDD.n2254 VDD.t2930 14.282
R4862 VDD.n2254 VDD.t2966 14.282
R4863 VDD.n2250 VDD.t589 14.282
R4864 VDD.n2250 VDD.t585 14.282
R4865 VDD.n2273 VDD.t2964 14.282
R4866 VDD.n2273 VDD.t856 14.282
R4867 VDD.n2269 VDD.t1049 14.282
R4868 VDD.n2269 VDD.t1053 14.282
R4869 VDD.n2334 VDD.t2283 14.282
R4870 VDD.n2334 VDD.t2279 14.282
R4871 VDD.n2326 VDD.t2960 14.282
R4872 VDD.n2326 VDD.t2938 14.282
R4873 VDD.n2354 VDD.t466 14.282
R4874 VDD.n2354 VDD.t462 14.282
R4875 VDD.n2346 VDD.t870 14.282
R4876 VDD.n2346 VDD.t2944 14.282
R4877 VDD.n2374 VDD.t3346 14.282
R4878 VDD.n2374 VDD.t3348 14.282
R4879 VDD.n2366 VDD.t2942 14.282
R4880 VDD.n2366 VDD.t838 14.282
R4881 VDD.n2313 VDD.t2918 14.282
R4882 VDD.n2313 VDD.t2948 14.282
R4883 VDD.n2309 VDD.t321 14.282
R4884 VDD.n2309 VDD.t323 14.282
R4885 VDD.n2293 VDD.t862 14.282
R4886 VDD.n2293 VDD.t2932 14.282
R4887 VDD.n2289 VDD.t2060 14.282
R4888 VDD.n2289 VDD.t2062 14.282
R4889 VDD.n1156 VDD.t2441 13.431
R4890 VDD.n1171 VDD.t928 13.431
R4891 VDD.n1201 VDD.t1411 13.431
R4892 VDD.n1129 VDD.t2468 13.431
R4893 VDD.n1234 VDD.t2198 13.431
R4894 VDD.n1216 VDD.t2605 13.397
R4895 VDD.n1186 VDD.t1847 13.397
R4896 VDD.n1144 VDD.t3728 13.397
R4897 VDD.n643 VDD.t811 12.385
R4898 VDD.n661 VDD.t735 12.385
R4899 VDD.n679 VDD.t1160 12.385
R4900 VDD.n696 VDD.t691 12.385
R4901 VDD.n625 VDD.t1224 12.385
R4902 VDD.n756 VDD.t1200 12.385
R4903 VDD.n774 VDD.t1170 12.385
R4904 VDD.n792 VDD.t823 12.385
R4905 VDD.n1054 VDD.n1053 9
R4906 VDD.n929 VDD.n928 9
R4907 VDD.n954 VDD.n953 9
R4908 VDD.n1029 VDD.n1028 9
R4909 VDD.n1004 VDD.n1003 9
R4910 VDD.n979 VDD.n978 9
R4911 VDD.n904 VDD.n903 9
R4912 VDD.n880 VDD.n879 9
R4913 VDD.n599 VDD.t4172 8.293
R4914 VDD.n585 VDD.t515 8.293
R4915 VDD.n263 VDD.t2054 8.293
R4916 VDD.n729 VDD.t2864 8.293
R4917 VDD.n1036 VDD.n1035 6.626
R4918 VDD.n911 VDD.n910 6.626
R4919 VDD.n936 VDD.n935 6.626
R4920 VDD.n1011 VDD.n1010 6.626
R4921 VDD.n986 VDD.n985 6.626
R4922 VDD.n961 VDD.n960 6.626
R4923 VDD.n886 VDD.n885 6.626
R4924 VDD.n862 VDD.n861 6.626
R4925 VDD.n1731 VDD.n1730 6.626
R4926 VDD.n1756 VDD.n1755 6.626
R4927 VDD.n1856 VDD.n1855 6.626
R4928 VDD.n1831 VDD.n1830 6.626
R4929 VDD.n1806 VDD.n1805 6.626
R4930 VDD.n1781 VDD.n1780 6.626
R4931 VDD.n1706 VDD.n1705 6.626
R4932 VDD.n1682 VDD.n1681 6.626
R4933 VDD.n1531 VDD.n1530 6.626
R4934 VDD.n1556 VDD.n1555 6.626
R4935 VDD.n1656 VDD.n1655 6.626
R4936 VDD.n1631 VDD.n1630 6.626
R4937 VDD.n1606 VDD.n1605 6.626
R4938 VDD.n1581 VDD.n1580 6.626
R4939 VDD.n1506 VDD.n1505 6.626
R4940 VDD.n1482 VDD.n1481 6.626
R4941 VDD.n1381 VDD.n1380 6.626
R4942 VDD.n1356 VDD.n1355 6.626
R4943 VDD.n1257 VDD.n1256 6.626
R4944 VDD.n1281 VDD.n1280 6.626
R4945 VDD.n1306 VDD.n1305 6.626
R4946 VDD.n1331 VDD.n1330 6.626
R4947 VDD.n1406 VDD.n1405 6.626
R4948 VDD.n1431 VDD.n1430 6.626
R4949 VDD.n2594 VDD.n2593 6.626
R4950 VDD.n2455 VDD.n2454 6.626
R4951 VDD.n2474 VDD.n2473 6.626
R4952 VDD.n2534 VDD.n2533 6.626
R4953 VDD.n2554 VDD.n2553 6.626
R4954 VDD.n2574 VDD.n2573 6.626
R4955 VDD.n2514 VDD.n2513 6.626
R4956 VDD.n2494 VDD.n2493 6.626
R4957 VDD.n2385 VDD.n2384 6.626
R4958 VDD.n2246 VDD.n2245 6.626
R4959 VDD.n2265 VDD.n2264 6.626
R4960 VDD.n2325 VDD.n2324 6.626
R4961 VDD.n2345 VDD.n2344 6.626
R4962 VDD.n2365 VDD.n2364 6.626
R4963 VDD.n2305 VDD.n2304 6.626
R4964 VDD.n2285 VDD.n2284 6.626
R4965 VDD.n644 VDD.n642 6.376
R4966 VDD.n662 VDD.n660 6.376
R4967 VDD.n680 VDD.n678 6.376
R4968 VDD.n697 VDD.n695 6.376
R4969 VDD.n626 VDD.n624 6.376
R4970 VDD.n757 VDD.n755 6.376
R4971 VDD.n775 VDD.n773 6.376
R4972 VDD.n793 VDD.n791 6.376
R4973 VDD.n2173 VDD.t4294 6.189
R4974 VDD.n2174 VDD.t3643 6.189
R4975 VDD.n2177 VDD.t1423 6.189
R4976 VDD.n2176 VDD.t1422 6.189
R4977 VDD.n2157 VDD.t2364 6.189
R4978 VDD.n2158 VDD.t766 6.189
R4979 VDD.n2161 VDD.t2151 6.189
R4980 VDD.n2160 VDD.t2150 6.189
R4981 VDD.n1460 VDD.t199 6.189
R4982 VDD.n1461 VDD.t201 6.189
R4983 VDD.n1464 VDD.t3908 6.189
R4984 VDD.n1463 VDD.t3907 6.189
R4985 VDD.n2037 VDD.t2257 6.189
R4986 VDD.n2038 VDD.t2258 6.189
R4987 VDD.n2041 VDD.t136 6.189
R4988 VDD.n2040 VDD.t137 6.189
R4989 VDD.n1937 VDD.t1041 6.189
R4990 VDD.n1938 VDD.t1042 6.189
R4991 VDD.n1941 VDD.t3387 6.189
R4992 VDD.n1940 VDD.t3385 6.189
R4993 VDD.n1887 VDD.t2576 6.189
R4994 VDD.n1888 VDD.t2577 6.189
R4995 VDD.n1891 VDD.t1478 6.189
R4996 VDD.n1890 VDD.t1479 6.189
R4997 VDD.n1912 VDD.t3176 6.189
R4998 VDD.n1913 VDD.t3150 6.189
R4999 VDD.n1916 VDD.t4448 6.189
R5000 VDD.n1915 VDD.t1126 6.189
R5001 VDD.n1962 VDD.t1623 6.189
R5002 VDD.n1963 VDD.t1624 6.189
R5003 VDD.n1966 VDD.t198 6.189
R5004 VDD.n1965 VDD.t2122 6.189
R5005 VDD.n1987 VDD.t1953 6.189
R5006 VDD.n1988 VDD.t1954 6.189
R5007 VDD.n1991 VDD.t311 6.189
R5008 VDD.n1990 VDD.t2743 6.189
R5009 VDD.n2012 VDD.t3060 6.189
R5010 VDD.n2013 VDD.t3058 6.189
R5011 VDD.n2016 VDD.t3636 6.189
R5012 VDD.n2015 VDD.t3635 6.189
R5013 VDD.n2062 VDD.t50 6.189
R5014 VDD.n2063 VDD.t52 6.189
R5015 VDD.n2066 VDD.t3362 6.189
R5016 VDD.n2065 VDD.t3363 6.189
R5017 VDD.n2625 VDD.t4350 6.189
R5018 VDD.n2626 VDD.t1750 6.189
R5019 VDD.n2629 VDD.t4117 6.189
R5020 VDD.n2628 VDD.t4118 6.189
R5021 VDD.n2432 VDD.t3370 6.189
R5022 VDD.n2433 VDD.t532 6.189
R5023 VDD.n2436 VDD.t43 6.189
R5024 VDD.n2435 VDD.t41 6.189
R5025 VDD.n2407 VDD.t526 6.189
R5026 VDD.n2408 VDD.t517 6.189
R5027 VDD.n2411 VDD.t3669 6.189
R5028 VDD.n2410 VDD.t3668 6.189
R5029 VDD.n2223 VDD.t1431 6.189
R5030 VDD.n2224 VDD.t1433 6.189
R5031 VDD.n2227 VDD.t1132 6.189
R5032 VDD.n2226 VDD.t1134 6.189
R5033 VDD.n2198 VDD.t3287 6.189
R5034 VDD.n2199 VDD.t3286 6.189
R5035 VDD.n2202 VDD.t2515 6.189
R5036 VDD.n2201 VDD.t441 6.189
R5037 VDD.t4123 VDD.n1158 6.105
R5038 VDD.t1865 VDD.n1173 6.105
R5039 VDD.t1413 VDD.n1203 6.105
R5040 VDD.t4136 VDD.n1131 6.105
R5041 VDD.t2200 VDD.n1236 6.105
R5042 VDD.t2609 VDD.n1218 6.089
R5043 VDD.t1825 VDD.n1188 6.089
R5044 VDD.t3732 VDD.n1146 6.089
R5045 VDD.n1039 VDD.n1038 6
R5046 VDD.n914 VDD.n913 6
R5047 VDD.n939 VDD.n938 6
R5048 VDD.n1014 VDD.n1013 6
R5049 VDD.n989 VDD.n988 6
R5050 VDD.n964 VDD.n963 6
R5051 VDD.n889 VDD.n888 6
R5052 VDD.n865 VDD.n864 6
R5053 VDD.n1733 VDD.n1732 6
R5054 VDD.n1758 VDD.n1757 6
R5055 VDD.n1858 VDD.n1857 6
R5056 VDD.n1833 VDD.n1832 6
R5057 VDD.n1808 VDD.n1807 6
R5058 VDD.n1783 VDD.n1782 6
R5059 VDD.n1708 VDD.n1707 6
R5060 VDD.n1684 VDD.n1683 6
R5061 VDD.n1533 VDD.n1532 6
R5062 VDD.n1558 VDD.n1557 6
R5063 VDD.n1658 VDD.n1657 6
R5064 VDD.n1633 VDD.n1632 6
R5065 VDD.n1608 VDD.n1607 6
R5066 VDD.n1583 VDD.n1582 6
R5067 VDD.n1508 VDD.n1507 6
R5068 VDD.n1484 VDD.n1483 6
R5069 VDD.n1383 VDD.n1382 6
R5070 VDD.n1358 VDD.n1357 6
R5071 VDD.n1259 VDD.n1258 6
R5072 VDD.n1283 VDD.n1282 6
R5073 VDD.n1308 VDD.n1307 6
R5074 VDD.n1333 VDD.n1332 6
R5075 VDD.n1408 VDD.n1407 6
R5076 VDD.n1433 VDD.n1432 6
R5077 VDD.n2591 VDD.n2590 6
R5078 VDD.n2452 VDD.n2451 6
R5079 VDD.n2471 VDD.n2470 6
R5080 VDD.n2531 VDD.n2530 6
R5081 VDD.n2551 VDD.n2550 6
R5082 VDD.n2571 VDD.n2570 6
R5083 VDD.n2511 VDD.n2510 6
R5084 VDD.n2491 VDD.n2490 6
R5085 VDD.n2382 VDD.n2381 6
R5086 VDD.n2243 VDD.n2242 6
R5087 VDD.n2262 VDD.n2261 6
R5088 VDD.n2322 VDD.n2321 6
R5089 VDD.n2342 VDD.n2341 6
R5090 VDD.n2362 VDD.n2361 6
R5091 VDD.n2302 VDD.n2301 6
R5092 VDD.n2282 VDD.n2281 6
R5093 VDD.n1157 VDD.n1156 5.506
R5094 VDD.n1172 VDD.n1171 5.506
R5095 VDD.n1217 VDD.n1216 5.506
R5096 VDD.n1202 VDD.n1201 5.506
R5097 VDD.n1187 VDD.n1186 5.506
R5098 VDD.n1145 VDD.n1144 5.506
R5099 VDD.n1130 VDD.n1129 5.506
R5100 VDD.n1235 VDD.n1234 5.506
R5101 VDD.n644 VDD.n643 4.688
R5102 VDD.n662 VDD.n661 4.688
R5103 VDD.n680 VDD.n679 4.688
R5104 VDD.n697 VDD.n696 4.688
R5105 VDD.n626 VDD.n625 4.688
R5106 VDD.n757 VDD.n756 4.688
R5107 VDD.n775 VDD.n774 4.688
R5108 VDD.n793 VDD.n792 4.688
R5109 VDD.n628 VDD.n627 4.623
R5110 VDD.n2999 VDD.t4147 4.524
R5111 VDD.n3000 VDD.t4146 4.524
R5112 VDD.n3002 VDD.t3612 4.524
R5113 VDD.n3001 VDD.t3613 4.524
R5114 VDD.n3187 VDD.t4083 4.524
R5115 VDD.n3188 VDD.t4023 4.524
R5116 VDD.n3190 VDD.t2159 4.524
R5117 VDD.n3189 VDD.t2160 4.524
R5118 VDD.n3069 VDD.t787 4.524
R5119 VDD.n3070 VDD.t2056 4.524
R5120 VDD.n3072 VDD.t460 4.524
R5121 VDD.n3071 VDD.t459 4.524
R5122 VDD.n351 VDD.t2877 4.524
R5123 VDD.n352 VDD.t3141 4.524
R5124 VDD.n354 VDD.t1858 4.524
R5125 VDD.n353 VDD.t1857 4.524
R5126 VDD.n450 VDD.t1772 4.524
R5127 VDD.n451 VDD.t1771 4.524
R5128 VDD.n453 VDD.t2841 4.524
R5129 VDD.n452 VDD.t2842 4.524
R5130 VDD.n518 VDD.t110 4.524
R5131 VDD.n519 VDD.t0 4.524
R5132 VDD.n521 VDD.t1552 4.524
R5133 VDD.n520 VDD.t1553 4.524
R5134 VDD.n2802 VDD.t2907 4.524
R5135 VDD.n2803 VDD.t1542 4.524
R5136 VDD.n2805 VDD.t3406 4.524
R5137 VDD.n2804 VDD.t3407 4.524
R5138 VDD.n2739 VDD.t393 4.524
R5139 VDD.n2740 VDD.t769 4.524
R5140 VDD.n2742 VDD.t1580 4.524
R5141 VDD.n2741 VDD.t1581 4.524
R5142 VDD.n728 VDD.n727 4.331
R5143 VDD.n598 VDD.n597 4.331
R5144 VDD.n262 VDD.n261 4.331
R5145 VDD.n2962 VDD.n2956 4.276
R5146 VDD.n2997 VDD.n2991 4.276
R5147 VDD.n3186 VDD.n3180 4.276
R5148 VDD.n3173 VDD.n3167 4.276
R5149 VDD.n3086 VDD.n3080 4.276
R5150 VDD.n3067 VDD.n3061 4.276
R5151 VDD.n189 VDD.n183 4.276
R5152 VDD.n177 VDD.n171 4.276
R5153 VDD.n130 VDD.n124 4.276
R5154 VDD.n118 VDD.n112 4.276
R5155 VDD.n844 VDD.n838 4.276
R5156 VDD.n20 VDD.n14 4.276
R5157 VDD.n79 VDD.n73 4.276
R5158 VDD.n67 VDD.n61 4.276
R5159 VDD.n367 VDD.n361 4.276
R5160 VDD.n349 VDD.n343 4.276
R5161 VDD.n467 VDD.n461 4.276
R5162 VDD.n448 VDD.n442 4.276
R5163 VDD.n479 VDD.n473 4.276
R5164 VDD.n516 VDD.n510 4.276
R5165 VDD.n2766 VDD.n2760 4.276
R5166 VDD.n2800 VDD.n2794 4.276
R5167 VDD.n2702 VDD.n2696 4.276
R5168 VDD.n2737 VDD.n2731 4.276
R5169 VDD VDD.n3450 3.655
R5170 VDD.n1140 VDD.t3508 3.442
R5171 VDD.n1125 VDD.t641 3.442
R5172 VDD.n1055 VDD.n1054 3.418
R5173 VDD.n930 VDD.n929 3.418
R5174 VDD.n955 VDD.n954 3.418
R5175 VDD.n1030 VDD.n1029 3.418
R5176 VDD.n1005 VDD.n1004 3.418
R5177 VDD.n980 VDD.n979 3.418
R5178 VDD.n905 VDD.n904 3.418
R5179 VDD.n881 VDD.n880 3.418
R5180 VDD.n1167 VDD.t11 3.368
R5181 VDD.n1212 VDD.t4203 3.368
R5182 VDD.n1197 VDD.t302 3.356
R5183 VDD.n1182 VDD.t3382 3.356
R5184 VDD.n2917 VDD.t2019 2.932
R5185 VDD.n1746 VDD.n1740 2.682
R5186 VDD.n1771 VDD.n1765 2.682
R5187 VDD.n1821 VDD.n1815 2.682
R5188 VDD.n1796 VDD.n1790 2.682
R5189 VDD.n1721 VDD.n1715 2.682
R5190 VDD.n1697 VDD.n1691 2.682
R5191 VDD.n2398 VDD.n2397 2.682
R5192 VDD.n2338 VDD.n2337 2.682
R5193 VDD.n2358 VDD.n2357 2.682
R5194 VDD.n2378 VDD.n2377 2.682
R5195 VDD.n1052 VDD.n1051 2.572
R5196 VDD.n927 VDD.n926 2.572
R5197 VDD.n952 VDD.n951 2.572
R5198 VDD.n1027 VDD.n1026 2.572
R5199 VDD.n1002 VDD.n1001 2.572
R5200 VDD.n977 VDD.n976 2.572
R5201 VDD.n902 VDD.n901 2.572
R5202 VDD.n878 VDD.n877 2.572
R5203 VDD.n641 VDD.n635 2.572
R5204 VDD.n659 VDD.n653 2.572
R5205 VDD.n677 VDD.n671 2.572
R5206 VDD.n694 VDD.n688 2.572
R5207 VDD.n623 VDD.n617 2.572
R5208 VDD.n754 VDD.n748 2.572
R5209 VDD.n772 VDD.n766 2.572
R5210 VDD.n790 VDD.n784 2.572
R5211 VDD.n1871 VDD.n1870 2.572
R5212 VDD.n1846 VDD.n1845 2.572
R5213 VDD.n1546 VDD.n1545 2.572
R5214 VDD.n1571 VDD.n1570 2.572
R5215 VDD.n1671 VDD.n1670 2.572
R5216 VDD.n1646 VDD.n1645 2.572
R5217 VDD.n1621 VDD.n1620 2.572
R5218 VDD.n1596 VDD.n1595 2.572
R5219 VDD.n1521 VDD.n1520 2.572
R5220 VDD.n1497 VDD.n1496 2.572
R5221 VDD.n1396 VDD.n1395 2.572
R5222 VDD.n1371 VDD.n1370 2.572
R5223 VDD.n1272 VDD.n1271 2.572
R5224 VDD.n1296 VDD.n1295 2.572
R5225 VDD.n1321 VDD.n1320 2.572
R5226 VDD.n1346 VDD.n1345 2.572
R5227 VDD.n1421 VDD.n1420 2.572
R5228 VDD.n1446 VDD.n1445 2.572
R5229 VDD.n2607 VDD.n2601 2.572
R5230 VDD.n2468 VDD.n2462 2.572
R5231 VDD.n2487 VDD.n2481 2.572
R5232 VDD.n2547 VDD.n2541 2.572
R5233 VDD.n2567 VDD.n2561 2.572
R5234 VDD.n2587 VDD.n2581 2.572
R5235 VDD.n2527 VDD.n2521 2.572
R5236 VDD.n2507 VDD.n2501 2.572
R5237 VDD.n2259 VDD.n2253 2.572
R5238 VDD.n2278 VDD.n2272 2.572
R5239 VDD.n2318 VDD.n2312 2.572
R5240 VDD.n2298 VDD.n2292 2.572
R5241 VDD.n2404 VDD.n2403 2.546
R5242 VDD.n2220 VDD.n2219 2.546
R5243 VDD.n1044 VDD.n1043 2.542
R5244 VDD.n919 VDD.n918 2.542
R5245 VDD.n944 VDD.n943 2.542
R5246 VDD.n1019 VDD.n1018 2.542
R5247 VDD.n994 VDD.n993 2.542
R5248 VDD.n969 VDD.n968 2.542
R5249 VDD.n894 VDD.n893 2.542
R5250 VDD.n870 VDD.n869 2.542
R5251 VDD.n640 VDD.n639 2.542
R5252 VDD.n658 VDD.n657 2.542
R5253 VDD.n676 VDD.n675 2.542
R5254 VDD.n693 VDD.n692 2.542
R5255 VDD.n622 VDD.n621 2.542
R5256 VDD.n753 VDD.n752 2.542
R5257 VDD.n771 VDD.n770 2.542
R5258 VDD.n789 VDD.n788 2.542
R5259 VDD.n1745 VDD.n1744 2.542
R5260 VDD.n1770 VDD.n1769 2.542
R5261 VDD.n1863 VDD.n1862 2.542
R5262 VDD.n1838 VDD.n1837 2.542
R5263 VDD.n1820 VDD.n1819 2.542
R5264 VDD.n1795 VDD.n1794 2.542
R5265 VDD.n1720 VDD.n1719 2.542
R5266 VDD.n1696 VDD.n1695 2.542
R5267 VDD.n1538 VDD.n1537 2.542
R5268 VDD.n1563 VDD.n1562 2.542
R5269 VDD.n1663 VDD.n1662 2.542
R5270 VDD.n1638 VDD.n1637 2.542
R5271 VDD.n1613 VDD.n1612 2.542
R5272 VDD.n1588 VDD.n1587 2.542
R5273 VDD.n1513 VDD.n1512 2.542
R5274 VDD.n1489 VDD.n1488 2.542
R5275 VDD.n1388 VDD.n1387 2.542
R5276 VDD.n1363 VDD.n1362 2.542
R5277 VDD.n1264 VDD.n1263 2.542
R5278 VDD.n1288 VDD.n1287 2.542
R5279 VDD.n1313 VDD.n1312 2.542
R5280 VDD.n1338 VDD.n1337 2.542
R5281 VDD.n1413 VDD.n1412 2.542
R5282 VDD.n1438 VDD.n1437 2.542
R5283 VDD.n2606 VDD.n2605 2.54
R5284 VDD.n2467 VDD.n2466 2.54
R5285 VDD.n2486 VDD.n2485 2.54
R5286 VDD.n2546 VDD.n2545 2.54
R5287 VDD.n2566 VDD.n2565 2.54
R5288 VDD.n2586 VDD.n2585 2.54
R5289 VDD.n2526 VDD.n2525 2.54
R5290 VDD.n2506 VDD.n2505 2.54
R5291 VDD.n2390 VDD.n2389 2.54
R5292 VDD.n2258 VDD.n2257 2.54
R5293 VDD.n2277 VDD.n2276 2.54
R5294 VDD.n2330 VDD.n2329 2.54
R5295 VDD.n2350 VDD.n2349 2.54
R5296 VDD.n2370 VDD.n2369 2.54
R5297 VDD.n2317 VDD.n2316 2.54
R5298 VDD.n2297 VDD.n2296 2.54
R5299 VDD.n2146 VDD.n2144 2.531
R5300 VDD.n1224 VDD.n1223 2.521
R5301 VDD.n2955 VDD.n2954 2.451
R5302 VDD.n2990 VDD.n2989 2.451
R5303 VDD.n3179 VDD.n3178 2.451
R5304 VDD.n3166 VDD.n3165 2.451
R5305 VDD.n3079 VDD.n3078 2.451
R5306 VDD.n3060 VDD.n3059 2.451
R5307 VDD.n726 VDD.n725 2.451
R5308 VDD.n596 VDD.n595 2.451
R5309 VDD.n582 VDD.n581 2.451
R5310 VDD.n260 VDD.n259 2.451
R5311 VDD.n182 VDD.n181 2.451
R5312 VDD.n170 VDD.n169 2.451
R5313 VDD.n123 VDD.n122 2.451
R5314 VDD.n111 VDD.n110 2.451
R5315 VDD.n837 VDD.n836 2.451
R5316 VDD.n13 VDD.n12 2.451
R5317 VDD.n72 VDD.n71 2.451
R5318 VDD.n60 VDD.n59 2.451
R5319 VDD.n3425 VDD.n3424 2.451
R5320 VDD.n3414 VDD.n3413 2.451
R5321 VDD.n3278 VDD.n3277 2.451
R5322 VDD.n3306 VDD.n3305 2.451
R5323 VDD.n3335 VDD.n3334 2.451
R5324 VDD.n3363 VDD.n3362 2.451
R5325 VDD.n211 VDD.n210 2.451
R5326 VDD.n239 VDD.n238 2.451
R5327 VDD.n360 VDD.n359 2.451
R5328 VDD.n342 VDD.n341 2.451
R5329 VDD.n460 VDD.n459 2.451
R5330 VDD.n441 VDD.n440 2.451
R5331 VDD.n472 VDD.n471 2.451
R5332 VDD.n509 VDD.n508 2.451
R5333 VDD.n2759 VDD.n2758 2.451
R5334 VDD.n2793 VDD.n2792 2.451
R5335 VDD.n2695 VDD.n2694 2.451
R5336 VDD.n2730 VDD.n2729 2.451
R5337 VDD.n2184 VDD.n2183 2.451
R5338 VDD.n1471 VDD.n1470 2.451
R5339 VDD.n2047 VDD.n2046 2.451
R5340 VDD.n1947 VDD.n1946 2.451
R5341 VDD.n1897 VDD.n1896 2.451
R5342 VDD.n1922 VDD.n1921 2.451
R5343 VDD.n1972 VDD.n1971 2.451
R5344 VDD.n1997 VDD.n1996 2.451
R5345 VDD.n2022 VDD.n2021 2.451
R5346 VDD.n2072 VDD.n2071 2.451
R5347 VDD.n2615 VDD.n2614 2.451
R5348 VDD.n2443 VDD.n2442 2.451
R5349 VDD.n2418 VDD.n2417 2.451
R5350 VDD.n2234 VDD.n2233 2.451
R5351 VDD.n2209 VDD.n2208 2.451
R5352 VDD.n2960 VDD.n2959 2.449
R5353 VDD.n2995 VDD.n2994 2.449
R5354 VDD.n3184 VDD.n3183 2.449
R5355 VDD.n3171 VDD.n3170 2.449
R5356 VDD.n3084 VDD.n3083 2.449
R5357 VDD.n3065 VDD.n3064 2.449
R5358 VDD.n721 VDD.n720 2.449
R5359 VDD.n591 VDD.n590 2.449
R5360 VDD.n577 VDD.n576 2.449
R5361 VDD.n255 VDD.n254 2.449
R5362 VDD.n187 VDD.n186 2.449
R5363 VDD.n175 VDD.n174 2.449
R5364 VDD.n128 VDD.n127 2.449
R5365 VDD.n116 VDD.n115 2.449
R5366 VDD.n842 VDD.n841 2.449
R5367 VDD.n18 VDD.n17 2.449
R5368 VDD.n77 VDD.n76 2.449
R5369 VDD.n65 VDD.n64 2.449
R5370 VDD.n3420 VDD.n3419 2.449
R5371 VDD.n3409 VDD.n3408 2.449
R5372 VDD.n3283 VDD.n3282 2.449
R5373 VDD.n3311 VDD.n3310 2.449
R5374 VDD.n3340 VDD.n3339 2.449
R5375 VDD.n3368 VDD.n3367 2.449
R5376 VDD.n216 VDD.n215 2.449
R5377 VDD.n244 VDD.n243 2.449
R5378 VDD.n365 VDD.n364 2.449
R5379 VDD.n347 VDD.n346 2.449
R5380 VDD.n465 VDD.n464 2.449
R5381 VDD.n446 VDD.n445 2.449
R5382 VDD.n477 VDD.n476 2.449
R5383 VDD.n514 VDD.n513 2.449
R5384 VDD.n2764 VDD.n2763 2.449
R5385 VDD.n2798 VDD.n2797 2.449
R5386 VDD.n2700 VDD.n2699 2.449
R5387 VDD.n2735 VDD.n2734 2.449
R5388 VDD.n2170 VDD.n2169 2.449
R5389 VDD.n2152 VDD.n2151 2.449
R5390 VDD.n1457 VDD.n1456 2.449
R5391 VDD.n2032 VDD.n2031 2.449
R5392 VDD.n1932 VDD.n1931 2.449
R5393 VDD.n1882 VDD.n1881 2.449
R5394 VDD.n1907 VDD.n1906 2.449
R5395 VDD.n1957 VDD.n1956 2.449
R5396 VDD.n1982 VDD.n1981 2.449
R5397 VDD.n2007 VDD.n2006 2.449
R5398 VDD.n2057 VDD.n2056 2.449
R5399 VDD.n2620 VDD.n2619 2.449
R5400 VDD.n2429 VDD.n2428 2.449
R5401 VDD.n2195 VDD.n2194 2.449
R5402 VDD.n1209 VDD.n1208 2.225
R5403 VDD.n1179 VDD.n1178 2.221
R5404 VDD.n1242 VDD.n1241 2.221
R5405 VDD.n1194 VDD.n1193 2.218
R5406 VDD.n1164 VDD.n1163 2.199
R5407 VDD.n1137 VDD.n1136 2.199
R5408 VDD.n2688 VDD.n2687 2.195
R5409 VDD.n2869 VDD.n2868 2.195
R5410 VDD.n2753 VDD.n2752 2.195
R5411 VDD.n2841 VDD.n2840 2.195
R5412 VDD.n2816 VDD.n2815 2.195
R5413 VDD.n530 VDD.n529 2.195
R5414 VDD.n559 VDD.n558 2.195
R5415 VDD.n566 VDD.n565 2.195
R5416 VDD.n3094 VDD.n3093 2.195
R5417 VDD.n376 VDD.n375 2.195
R5418 VDD.n3023 VDD.n3022 2.195
R5419 VDD.n3030 VDD.n3029 2.195
R5420 VDD.n3207 VDD.n3206 2.195
R5421 VDD.n2942 VDD.n2941 2.195
R5422 VDD.n2948 VDD.n2947 2.195
R5423 VDD.n3013 VDD.n3012 2.195
R5424 VDD.n3375 VDD.n3374 2.195
R5425 VDD.n3380 VDD.n3379 2.195
R5426 VDD.n3323 VDD.n3322 2.195
R5427 VDD.n3318 VDD.n3317 2.195
R5428 VDD.n201 VDD.n200 2.195
R5429 VDD.n206 VDD.n205 2.195
R5430 VDD.n3266 VDD.n3265 2.195
R5431 VDD.n33 VDD.n32 2.195
R5432 VDD.n38 VDD.n37 2.195
R5433 VDD.n3 VDD.n2 2.195
R5434 VDD.n8 VDD.n7 2.195
R5435 VDD.n89 VDD.n88 2.195
R5436 VDD.n84 VDD.n83 2.195
R5437 VDD.n143 VDD.n142 2.195
R5438 VDD.n148 VDD.n147 2.195
R5439 VDD.n3402 VDD.n3401 2.195
R5440 VDD.n1152 VDD.n1151 2.192
R5441 VDD.n1039 VDD.n1037 1.929
R5442 VDD.n914 VDD.n912 1.929
R5443 VDD.n939 VDD.n937 1.929
R5444 VDD.n1014 VDD.n1012 1.929
R5445 VDD.n989 VDD.n987 1.929
R5446 VDD.n964 VDD.n962 1.929
R5447 VDD.n889 VDD.n887 1.929
R5448 VDD.n865 VDD.n863 1.929
R5449 VDD.n568 VDD.n567 1.833
R5450 VDD.n561 VDD.n560 1.811
R5451 VDD.n2870 VDD.n2866 1.72
R5452 VDD.n2842 VDD.n2838 1.72
R5453 VDD.n531 VDD.n527 1.72
R5454 VDD.n377 VDD.n373 1.72
R5455 VDD.n3031 VDD.n3027 1.72
R5456 VDD.n2949 VDD.n2945 1.72
R5457 VDD.n3014 VDD.n3010 1.72
R5458 VDD.n3376 VDD.n3372 1.72
R5459 VDD.n3319 VDD.n3315 1.72
R5460 VDD.n207 VDD.n203 1.72
R5461 VDD.n39 VDD.n35 1.72
R5462 VDD.n9 VDD.n5 1.72
R5463 VDD.n90 VDD.n86 1.72
R5464 VDD.n149 VDD.n145 1.72
R5465 VDD.n3403 VDD.n3399 1.72
R5466 VDD.n2689 VDD.n2685 1.698
R5467 VDD.n2754 VDD.n2750 1.698
R5468 VDD.n2817 VDD.n2813 1.698
R5469 VDD.n3095 VDD.n3091 1.698
R5470 VDD.n3024 VDD.n3020 1.698
R5471 VDD.n3208 VDD.n3204 1.698
R5472 VDD.n2943 VDD.n2939 1.698
R5473 VDD.n3381 VDD.n3377 1.698
R5474 VDD.n3324 VDD.n3320 1.698
R5475 VDD.n202 VDD.n198 1.698
R5476 VDD.n3267 VDD.n3263 1.698
R5477 VDD.n34 VDD.n30 1.698
R5478 VDD.n4 VDD.n0 1.698
R5479 VDD.n85 VDD.n81 1.698
R5480 VDD.n144 VDD.n140 1.698
R5481 VDD.n2687 VDD.n2686 1.651
R5482 VDD.n2868 VDD.n2867 1.651
R5483 VDD.n2752 VDD.n2751 1.651
R5484 VDD.n2840 VDD.n2839 1.651
R5485 VDD.n2815 VDD.n2814 1.651
R5486 VDD.n529 VDD.n528 1.651
R5487 VDD.n558 VDD.n557 1.651
R5488 VDD.n565 VDD.n564 1.651
R5489 VDD.n3093 VDD.n3092 1.651
R5490 VDD.n375 VDD.n374 1.651
R5491 VDD.n3022 VDD.n3021 1.651
R5492 VDD.n3029 VDD.n3028 1.651
R5493 VDD.n3206 VDD.n3205 1.651
R5494 VDD.n2941 VDD.n2940 1.651
R5495 VDD.n2947 VDD.n2946 1.651
R5496 VDD.n3012 VDD.n3011 1.651
R5497 VDD.n3374 VDD.n3373 1.651
R5498 VDD.n3379 VDD.n3378 1.651
R5499 VDD.n3322 VDD.n3321 1.651
R5500 VDD.n3317 VDD.n3316 1.651
R5501 VDD.n200 VDD.n199 1.651
R5502 VDD.n205 VDD.n204 1.651
R5503 VDD.n3265 VDD.n3264 1.651
R5504 VDD.n32 VDD.n31 1.651
R5505 VDD.n37 VDD.n36 1.651
R5506 VDD.n2 VDD.n1 1.651
R5507 VDD.n7 VDD.n6 1.651
R5508 VDD.n88 VDD.n87 1.651
R5509 VDD.n83 VDD.n82 1.651
R5510 VDD.n142 VDD.n141 1.651
R5511 VDD.n147 VDD.n146 1.651
R5512 VDD.n3401 VDD.n3400 1.651
R5513 VDD.n1163 VDD.n1162 1.651
R5514 VDD.n1151 VDD.n1150 1.651
R5515 VDD.n1136 VDD.n1135 1.651
R5516 VDD.n3255 VDD.n3254 1.647
R5517 VDD.n546 VDD.n545 1.647
R5518 VDD.n406 VDD.n405 1.647
R5519 VDD.n2923 VDD.n2922 1.647
R5520 VDD.n280 VDD.n279 1.647
R5521 VDD.n269 VDD.n268 1.647
R5522 VDD.n421 VDD.n420 1.647
R5523 VDD.n482 VDD.n481 1.647
R5524 VDD.n2772 VDD.n2771 1.647
R5525 VDD.n2705 VDD.n2704 1.647
R5526 VDD.n1081 VDD.n1080 1.647
R5527 VDD.n1089 VDD.n1088 1.647
R5528 VDD.n1122 VDD.n1121 1.647
R5529 VDD.n1114 VDD.n1113 1.647
R5530 VDD.n1105 VDD.n1104 1.647
R5531 VDD.n1097 VDD.n1096 1.647
R5532 VDD.n1072 VDD.n1071 1.647
R5533 VDD.n1064 VDD.n1063 1.647
R5534 VDD.n1178 VDD.n1177 1.607
R5535 VDD.n1223 VDD.n1222 1.607
R5536 VDD.n1241 VDD.n1240 1.607
R5537 VDD.n1208 VDD.n1207 1.599
R5538 VDD.n1193 VDD.n1192 1.599
R5539 VDD.n2938 VDD.n2936 1.564
R5540 VDD.n2903 VDD.n2901 1.564
R5541 VDD.n2676 VDD.n2674 1.564
R5542 VDD.n2667 VDD.n2665 1.564
R5543 VDD.n2684 VDD.n2682 1.564
R5544 VDD.n2749 VDD.n2747 1.564
R5545 VDD.n2812 VDD.n2810 1.564
R5546 VDD.n2911 VDD.n2909 1.564
R5547 VDD.n306 VDD.n304 1.564
R5548 VDD.n297 VDD.n295 1.564
R5549 VDD.n388 VDD.n386 1.564
R5550 VDD.n397 VDD.n395 1.564
R5551 VDD.n3090 VDD.n3088 1.564
R5552 VDD.n3019 VDD.n3017 1.564
R5553 VDD.n3009 VDD.n3007 1.564
R5554 VDD.n2965 VDD.n2963 1.564
R5555 VDD.n2969 VDD.n2967 1.564
R5556 VDD.n3141 VDD.n3139 1.564
R5557 VDD.n3151 VDD.n3149 1.564
R5558 VDD.n3036 VDD.n3034 1.564
R5559 VDD.n3045 VDD.n3043 1.564
R5560 VDD.n2657 VDD.n2655 1.564
R5561 VDD.n710 VDD.n708 1.564
R5562 VDD.n2649 VDD.n2647 1.564
R5563 VDD.n702 VDD.n700 1.564
R5564 VDD.n735 VDD.n733 1.564
R5565 VDD.n604 VDD.n602 1.564
R5566 VDD.n289 VDD.n287 1.564
R5567 VDD.n3274 VDD.n3272 1.564
R5568 VDD.n3331 VDD.n3329 1.564
R5569 VDD.n3388 VDD.n3386 1.564
R5570 VDD.n197 VDD.n195 1.564
R5571 VDD.n852 VDD.n850 1.564
R5572 VDD.n832 VDD.n830 1.564
R5573 VDD.n28 VDD.n26 1.564
R5574 VDD.n820 VDD.n818 1.564
R5575 VDD.n809 VDD.n807 1.564
R5576 VDD.n138 VDD.n136 1.564
R5577 VDD.n164 VDD.n162 1.564
R5578 VDD.n156 VDD.n154 1.564
R5579 VDD.n105 VDD.n103 1.564
R5580 VDD.n97 VDD.n95 1.564
R5581 VDD.n54 VDD.n52 1.564
R5582 VDD.n46 VDD.n44 1.564
R5583 VDD.n3434 VDD.n3432 1.564
R5584 VDD.n3437 VDD.n3435 1.564
R5585 VDD.n3292 VDD.n3290 1.564
R5586 VDD.n3295 VDD.n3293 1.564
R5587 VDD.n3349 VDD.n3347 1.564
R5588 VDD.n3352 VDD.n3350 1.564
R5589 VDD.n225 VDD.n223 1.564
R5590 VDD.n228 VDD.n226 1.564
R5591 VDD.n331 VDD.n329 1.564
R5592 VDD.n320 VDD.n318 1.564
R5593 VDD.n418 VDD.n416 1.564
R5594 VDD.n499 VDD.n497 1.564
R5595 VDD.n2769 VDD.n2767 1.564
R5596 VDD.n2716 VDD.n2714 1.564
R5597 VDD.n414 VDD.n413 1.496
R5598 VDD.n2932 VDD.n2931 1.224
R5599 VDD.n2931 VDD.n2930 1.214
R5600 VDD.n716 VDD.n715 1.212
R5601 VDD.n2148 VDD.n2147 1.195
R5602 VDD.n2146 VDD.n2145 1.194
R5603 VDD.n1453 VDD.n1452 1.187
R5604 VDD.n1225 VDD.n1224 1.158
R5605 VDD.n1195 VDD.n1194 1.158
R5606 VDD.n1153 VDD.n1152 1.158
R5607 VDD.n1165 VDD.n1164 1.151
R5608 VDD.n1180 VDD.n1179 1.151
R5609 VDD.n1210 VDD.n1209 1.151
R5610 VDD.n1138 VDD.n1137 1.151
R5611 VDD.n1243 VDD.n1242 1.151
R5612 VDD.n2616 VDD.n2612 1.114
R5613 VDD.n1225 VDD.n1221 1.11
R5614 VDD.n1195 VDD.n1191 1.11
R5615 VDD.n1153 VDD.n1149 1.11
R5616 VDD.n1165 VDD.n1161 1.103
R5617 VDD.n1180 VDD.n1176 1.103
R5618 VDD.n1210 VDD.n1206 1.103
R5619 VDD.n1138 VDD.n1134 1.103
R5620 VDD.n1243 VDD.n1239 1.103
R5621 VDD.n1038 VDD.t2182 1.057
R5622 VDD.n913 VDD.t2867 1.057
R5623 VDD.n938 VDD.t2033 1.057
R5624 VDD.n1013 VDD.t2806 1.057
R5625 VDD.n988 VDD.t353 1.057
R5626 VDD.n963 VDD.t3057 1.057
R5627 VDD.n888 VDD.t4148 1.057
R5628 VDD.n864 VDD.t4191 1.057
R5629 VDD.n1732 VDD.t2745 1.057
R5630 VDD.n1757 VDD.t2717 1.057
R5631 VDD.n1857 VDD.t2123 1.057
R5632 VDD.n1832 VDD.t4533 1.057
R5633 VDD.n1807 VDD.t415 1.057
R5634 VDD.n1782 VDD.t963 1.057
R5635 VDD.n1707 VDD.t3647 1.057
R5636 VDD.n1683 VDD.t1562 1.057
R5637 VDD.n1532 VDD.t2523 1.057
R5638 VDD.n1557 VDD.t4074 1.057
R5639 VDD.n1657 VDD.t3699 1.057
R5640 VDD.n1632 VDD.t127 1.057
R5641 VDD.n1607 VDD.t1026 1.057
R5642 VDD.n1582 VDD.t2675 1.057
R5643 VDD.n1507 VDD.t53 1.057
R5644 VDD.n1483 VDD.t4442 1.057
R5645 VDD.n1382 VDD.t1990 1.057
R5646 VDD.n1357 VDD.t387 1.057
R5647 VDD.n1258 VDD.t2527 1.057
R5648 VDD.n1282 VDD.t139 1.057
R5649 VDD.n1307 VDD.t1329 1.057
R5650 VDD.n1332 VDD.t3565 1.057
R5651 VDD.n1407 VDD.t1955 1.057
R5652 VDD.n1432 VDD.t2868 1.057
R5653 VDD.n2590 VDD.t1919 1.057
R5654 VDD.n2451 VDD.t75 1.057
R5655 VDD.n2470 VDD.t4559 1.057
R5656 VDD.n2530 VDD.t4489 1.057
R5657 VDD.n2550 VDD.t467 1.057
R5658 VDD.n2570 VDD.t2286 1.057
R5659 VDD.n2510 VDD.t4494 1.057
R5660 VDD.n2490 VDD.t4180 1.057
R5661 VDD.n2381 VDD.t3115 1.057
R5662 VDD.n2242 VDD.t80 1.057
R5663 VDD.n2261 VDD.t2289 1.057
R5664 VDD.n2321 VDD.t24 1.057
R5665 VDD.n2341 VDD.t3521 1.057
R5666 VDD.n2361 VDD.t2535 1.057
R5667 VDD.n2301 VDD.t1691 1.057
R5668 VDD.n2281 VDD.t3603 1.057
R5669 VDD.n642 VDD.t611 1.057
R5670 VDD.n660 VDD.t1960 1.057
R5671 VDD.n678 VDD.t3243 1.057
R5672 VDD.n695 VDD.t2838 1.057
R5673 VDD.n624 VDD.t4133 1.057
R5674 VDD.n755 VDD.t2248 1.057
R5675 VDD.n773 VDD.t3371 1.057
R5676 VDD.n791 VDD.t655 1.057
R5677 VDD.n1453 VDD.n1253 1.052
R5678 VDD.n2663 VDD.n2662 1.031
R5679 VDD.n3256 VDD.n3255 0.983
R5680 VDD.n550 VDD.n549 0.983
R5681 VDD.n407 VDD.n406 0.983
R5682 VDD.n2924 VDD.n2923 0.983
R5683 VDD.n281 VDD.n280 0.983
R5684 VDD.n270 VDD.n269 0.983
R5685 VDD.n425 VDD.n424 0.983
R5686 VDD.n486 VDD.n485 0.983
R5687 VDD.n2776 VDD.n2775 0.983
R5688 VDD.n2709 VDD.n2708 0.983
R5689 VDD.n1082 VDD.n1081 0.983
R5690 VDD.n1090 VDD.n1089 0.983
R5691 VDD.n1123 VDD.n1122 0.983
R5692 VDD.n1115 VDD.n1114 0.983
R5693 VDD.n1106 VDD.n1105 0.983
R5694 VDD.n1098 VDD.n1097 0.983
R5695 VDD.n1073 VDD.n1072 0.983
R5696 VDD.n1065 VDD.n1064 0.983
R5697 VDD.n2956 VDD.n2952 0.922
R5698 VDD.n2961 VDD.n2957 0.922
R5699 VDD.n2991 VDD.n2987 0.922
R5700 VDD.n2996 VDD.n2992 0.922
R5701 VDD.n3180 VDD.n3176 0.922
R5702 VDD.n3185 VDD.n3181 0.922
R5703 VDD.n3167 VDD.n3163 0.922
R5704 VDD.n3172 VDD.n3168 0.922
R5705 VDD.n3080 VDD.n3076 0.922
R5706 VDD.n3085 VDD.n3081 0.922
R5707 VDD.n3061 VDD.n3057 0.922
R5708 VDD.n3066 VDD.n3062 0.922
R5709 VDD.n727 VDD.n723 0.922
R5710 VDD.n722 VDD.n718 0.922
R5711 VDD.n597 VDD.n593 0.922
R5712 VDD.n592 VDD.n588 0.922
R5713 VDD.n583 VDD.n579 0.922
R5714 VDD.n578 VDD.n574 0.922
R5715 VDD.n261 VDD.n257 0.922
R5716 VDD.n256 VDD.n252 0.922
R5717 VDD.n183 VDD.n179 0.922
R5718 VDD.n188 VDD.n184 0.922
R5719 VDD.n171 VDD.n167 0.922
R5720 VDD.n176 VDD.n172 0.922
R5721 VDD.n124 VDD.n120 0.922
R5722 VDD.n129 VDD.n125 0.922
R5723 VDD.n112 VDD.n108 0.922
R5724 VDD.n117 VDD.n113 0.922
R5725 VDD.n838 VDD.n834 0.922
R5726 VDD.n843 VDD.n839 0.922
R5727 VDD.n14 VDD.n10 0.922
R5728 VDD.n19 VDD.n15 0.922
R5729 VDD.n73 VDD.n69 0.922
R5730 VDD.n78 VDD.n74 0.922
R5731 VDD.n61 VDD.n57 0.922
R5732 VDD.n66 VDD.n62 0.922
R5733 VDD.n3426 VDD.n3422 0.922
R5734 VDD.n3421 VDD.n3417 0.922
R5735 VDD.n3415 VDD.n3411 0.922
R5736 VDD.n3410 VDD.n3406 0.922
R5737 VDD.n3284 VDD.n3280 0.922
R5738 VDD.n3279 VDD.n3275 0.922
R5739 VDD.n3312 VDD.n3308 0.922
R5740 VDD.n3307 VDD.n3303 0.922
R5741 VDD.n3341 VDD.n3337 0.922
R5742 VDD.n3336 VDD.n3332 0.922
R5743 VDD.n3369 VDD.n3365 0.922
R5744 VDD.n3364 VDD.n3360 0.922
R5745 VDD.n217 VDD.n213 0.922
R5746 VDD.n212 VDD.n208 0.922
R5747 VDD.n245 VDD.n241 0.922
R5748 VDD.n240 VDD.n236 0.922
R5749 VDD.n361 VDD.n357 0.922
R5750 VDD.n366 VDD.n362 0.922
R5751 VDD.n343 VDD.n339 0.922
R5752 VDD.n348 VDD.n344 0.922
R5753 VDD.n461 VDD.n457 0.922
R5754 VDD.n466 VDD.n462 0.922
R5755 VDD.n442 VDD.n438 0.922
R5756 VDD.n447 VDD.n443 0.922
R5757 VDD.n473 VDD.n469 0.922
R5758 VDD.n478 VDD.n474 0.922
R5759 VDD.n510 VDD.n506 0.922
R5760 VDD.n515 VDD.n511 0.922
R5761 VDD.n2760 VDD.n2756 0.922
R5762 VDD.n2765 VDD.n2761 0.922
R5763 VDD.n2794 VDD.n2790 0.922
R5764 VDD.n2799 VDD.n2795 0.922
R5765 VDD.n2696 VDD.n2692 0.922
R5766 VDD.n2701 VDD.n2697 0.922
R5767 VDD.n2731 VDD.n2727 0.922
R5768 VDD.n2736 VDD.n2732 0.922
R5769 VDD.n2185 VDD.n2181 0.922
R5770 VDD.n2171 VDD.n2167 0.922
R5771 VDD.n2153 VDD.n2149 0.922
R5772 VDD.n1472 VDD.n1468 0.922
R5773 VDD.n1458 VDD.n1454 0.922
R5774 VDD.n2033 VDD.n2029 0.922
R5775 VDD.n2048 VDD.n2044 0.922
R5776 VDD.n1933 VDD.n1929 0.922
R5777 VDD.n1948 VDD.n1944 0.922
R5778 VDD.n1883 VDD.n1879 0.922
R5779 VDD.n1898 VDD.n1894 0.922
R5780 VDD.n1908 VDD.n1904 0.922
R5781 VDD.n1923 VDD.n1919 0.922
R5782 VDD.n1958 VDD.n1954 0.922
R5783 VDD.n1973 VDD.n1969 0.922
R5784 VDD.n1983 VDD.n1979 0.922
R5785 VDD.n1998 VDD.n1994 0.922
R5786 VDD.n2008 VDD.n2004 0.922
R5787 VDD.n2023 VDD.n2019 0.922
R5788 VDD.n2058 VDD.n2054 0.922
R5789 VDD.n2073 VDD.n2069 0.922
R5790 VDD.n2621 VDD.n2617 0.922
R5791 VDD.n2444 VDD.n2440 0.922
R5792 VDD.n2430 VDD.n2426 0.922
R5793 VDD.n2419 VDD.n2415 0.922
R5794 VDD.n2405 VDD.n2401 0.922
R5795 VDD.n2235 VDD.n2231 0.922
R5796 VDD.n2221 VDD.n2217 0.922
R5797 VDD.n2210 VDD.n2206 0.922
R5798 VDD.n2196 VDD.n2192 0.922
R5799 VDD.n2955 VDD.n2953 0.921
R5800 VDD.n2960 VDD.n2958 0.921
R5801 VDD.n2990 VDD.n2988 0.921
R5802 VDD.n2995 VDD.n2993 0.921
R5803 VDD.n3179 VDD.n3177 0.921
R5804 VDD.n3184 VDD.n3182 0.921
R5805 VDD.n3166 VDD.n3164 0.921
R5806 VDD.n3171 VDD.n3169 0.921
R5807 VDD.n3079 VDD.n3077 0.921
R5808 VDD.n3084 VDD.n3082 0.921
R5809 VDD.n3060 VDD.n3058 0.921
R5810 VDD.n3065 VDD.n3063 0.921
R5811 VDD.n726 VDD.n724 0.921
R5812 VDD.n721 VDD.n719 0.921
R5813 VDD.n596 VDD.n594 0.921
R5814 VDD.n591 VDD.n589 0.921
R5815 VDD.n582 VDD.n580 0.921
R5816 VDD.n577 VDD.n575 0.921
R5817 VDD.n260 VDD.n258 0.921
R5818 VDD.n255 VDD.n253 0.921
R5819 VDD.n182 VDD.n180 0.921
R5820 VDD.n187 VDD.n185 0.921
R5821 VDD.n170 VDD.n168 0.921
R5822 VDD.n175 VDD.n173 0.921
R5823 VDD.n123 VDD.n121 0.921
R5824 VDD.n128 VDD.n126 0.921
R5825 VDD.n111 VDD.n109 0.921
R5826 VDD.n116 VDD.n114 0.921
R5827 VDD.n837 VDD.n835 0.921
R5828 VDD.n842 VDD.n840 0.921
R5829 VDD.n13 VDD.n11 0.921
R5830 VDD.n18 VDD.n16 0.921
R5831 VDD.n72 VDD.n70 0.921
R5832 VDD.n77 VDD.n75 0.921
R5833 VDD.n60 VDD.n58 0.921
R5834 VDD.n65 VDD.n63 0.921
R5835 VDD.n3425 VDD.n3423 0.921
R5836 VDD.n3420 VDD.n3418 0.921
R5837 VDD.n3414 VDD.n3412 0.921
R5838 VDD.n3409 VDD.n3407 0.921
R5839 VDD.n3283 VDD.n3281 0.921
R5840 VDD.n3278 VDD.n3276 0.921
R5841 VDD.n3311 VDD.n3309 0.921
R5842 VDD.n3306 VDD.n3304 0.921
R5843 VDD.n3340 VDD.n3338 0.921
R5844 VDD.n3335 VDD.n3333 0.921
R5845 VDD.n3368 VDD.n3366 0.921
R5846 VDD.n3363 VDD.n3361 0.921
R5847 VDD.n216 VDD.n214 0.921
R5848 VDD.n211 VDD.n209 0.921
R5849 VDD.n244 VDD.n242 0.921
R5850 VDD.n239 VDD.n237 0.921
R5851 VDD.n360 VDD.n358 0.921
R5852 VDD.n365 VDD.n363 0.921
R5853 VDD.n342 VDD.n340 0.921
R5854 VDD.n347 VDD.n345 0.921
R5855 VDD.n460 VDD.n458 0.921
R5856 VDD.n465 VDD.n463 0.921
R5857 VDD.n441 VDD.n439 0.921
R5858 VDD.n446 VDD.n444 0.921
R5859 VDD.n472 VDD.n470 0.921
R5860 VDD.n477 VDD.n475 0.921
R5861 VDD.n509 VDD.n507 0.921
R5862 VDD.n514 VDD.n512 0.921
R5863 VDD.n2759 VDD.n2757 0.921
R5864 VDD.n2764 VDD.n2762 0.921
R5865 VDD.n2793 VDD.n2791 0.921
R5866 VDD.n2798 VDD.n2796 0.921
R5867 VDD.n2695 VDD.n2693 0.921
R5868 VDD.n2700 VDD.n2698 0.921
R5869 VDD.n2730 VDD.n2728 0.921
R5870 VDD.n2735 VDD.n2733 0.921
R5871 VDD.n2184 VDD.n2182 0.921
R5872 VDD.n2170 VDD.n2168 0.921
R5873 VDD.n2152 VDD.n2150 0.921
R5874 VDD.n1471 VDD.n1469 0.921
R5875 VDD.n1457 VDD.n1455 0.921
R5876 VDD.n2032 VDD.n2030 0.921
R5877 VDD.n2047 VDD.n2045 0.921
R5878 VDD.n1932 VDD.n1930 0.921
R5879 VDD.n1947 VDD.n1945 0.921
R5880 VDD.n1882 VDD.n1880 0.921
R5881 VDD.n1897 VDD.n1895 0.921
R5882 VDD.n1907 VDD.n1905 0.921
R5883 VDD.n1922 VDD.n1920 0.921
R5884 VDD.n1957 VDD.n1955 0.921
R5885 VDD.n1972 VDD.n1970 0.921
R5886 VDD.n1982 VDD.n1980 0.921
R5887 VDD.n1997 VDD.n1995 0.921
R5888 VDD.n2007 VDD.n2005 0.921
R5889 VDD.n2022 VDD.n2020 0.921
R5890 VDD.n2057 VDD.n2055 0.921
R5891 VDD.n2072 VDD.n2070 0.921
R5892 VDD.n2620 VDD.n2618 0.921
R5893 VDD.n2615 VDD.n2613 0.921
R5894 VDD.n2443 VDD.n2441 0.921
R5895 VDD.n2429 VDD.n2427 0.921
R5896 VDD.n2418 VDD.n2416 0.921
R5897 VDD.n2404 VDD.n2402 0.921
R5898 VDD.n2234 VDD.n2232 0.921
R5899 VDD.n2220 VDD.n2218 0.921
R5900 VDD.n2209 VDD.n2207 0.921
R5901 VDD.n2195 VDD.n2193 0.921
R5902 VDD.n551 VDD.n546 0.908
R5903 VDD.n426 VDD.n421 0.908
R5904 VDD.n487 VDD.n482 0.908
R5905 VDD.n2777 VDD.n2772 0.908
R5906 VDD.n2710 VDD.n2705 0.908
R5907 VDD.n1044 VDD.n1041 0.863
R5908 VDD.n919 VDD.n916 0.863
R5909 VDD.n944 VDD.n941 0.863
R5910 VDD.n1019 VDD.n1016 0.863
R5911 VDD.n994 VDD.n991 0.863
R5912 VDD.n969 VDD.n966 0.863
R5913 VDD.n894 VDD.n891 0.863
R5914 VDD.n870 VDD.n867 0.863
R5915 VDD.n640 VDD.n637 0.863
R5916 VDD.n658 VDD.n655 0.863
R5917 VDD.n676 VDD.n673 0.863
R5918 VDD.n693 VDD.n690 0.863
R5919 VDD.n622 VDD.n619 0.863
R5920 VDD.n753 VDD.n750 0.863
R5921 VDD.n771 VDD.n768 0.863
R5922 VDD.n789 VDD.n786 0.863
R5923 VDD.n1745 VDD.n1742 0.863
R5924 VDD.n1770 VDD.n1767 0.863
R5925 VDD.n1863 VDD.n1860 0.863
R5926 VDD.n1838 VDD.n1835 0.863
R5927 VDD.n1820 VDD.n1817 0.863
R5928 VDD.n1795 VDD.n1792 0.863
R5929 VDD.n1720 VDD.n1717 0.863
R5930 VDD.n1696 VDD.n1693 0.863
R5931 VDD.n1538 VDD.n1535 0.863
R5932 VDD.n1563 VDD.n1560 0.863
R5933 VDD.n1663 VDD.n1660 0.863
R5934 VDD.n1638 VDD.n1635 0.863
R5935 VDD.n1613 VDD.n1610 0.863
R5936 VDD.n1588 VDD.n1585 0.863
R5937 VDD.n1513 VDD.n1510 0.863
R5938 VDD.n1489 VDD.n1486 0.863
R5939 VDD.n1388 VDD.n1385 0.863
R5940 VDD.n1363 VDD.n1360 0.863
R5941 VDD.n1264 VDD.n1261 0.863
R5942 VDD.n1288 VDD.n1285 0.863
R5943 VDD.n1313 VDD.n1310 0.863
R5944 VDD.n1338 VDD.n1335 0.863
R5945 VDD.n1413 VDD.n1410 0.863
R5946 VDD.n1438 VDD.n1435 0.863
R5947 VDD.n2606 VDD.n2603 0.863
R5948 VDD.n2467 VDD.n2464 0.863
R5949 VDD.n2486 VDD.n2483 0.863
R5950 VDD.n2546 VDD.n2543 0.863
R5951 VDD.n2566 VDD.n2563 0.863
R5952 VDD.n2586 VDD.n2583 0.863
R5953 VDD.n2526 VDD.n2523 0.863
R5954 VDD.n2506 VDD.n2503 0.863
R5955 VDD.n2390 VDD.n2387 0.863
R5956 VDD.n2258 VDD.n2255 0.863
R5957 VDD.n2277 VDD.n2274 0.863
R5958 VDD.n2330 VDD.n2327 0.863
R5959 VDD.n2350 VDD.n2347 0.863
R5960 VDD.n2370 VDD.n2367 0.863
R5961 VDD.n2317 VDD.n2314 0.863
R5962 VDD.n2297 VDD.n2294 0.863
R5963 VDD.n2905 VDD.n2903 0.85
R5964 VDD.n2678 VDD.n2676 0.85
R5965 VDD.n2669 VDD.n2667 0.85
R5966 VDD.n2913 VDD.n2911 0.85
R5967 VDD.n308 VDD.n306 0.85
R5968 VDD.n299 VDD.n297 0.85
R5969 VDD.n390 VDD.n388 0.85
R5970 VDD.n399 VDD.n397 0.85
R5971 VDD.n2659 VDD.n2657 0.85
R5972 VDD.n712 VDD.n710 0.85
R5973 VDD.n2651 VDD.n2649 0.85
R5974 VDD.n704 VDD.n702 0.85
R5975 VDD.n737 VDD.n735 0.85
R5976 VDD.n606 VDD.n604 0.85
R5977 VDD.n291 VDD.n289 0.85
R5978 VDD.n2689 VDD.n2688 0.806
R5979 VDD.n2754 VDD.n2753 0.806
R5980 VDD.n2817 VDD.n2816 0.806
R5981 VDD.n3095 VDD.n3094 0.806
R5982 VDD.n3024 VDD.n3023 0.806
R5983 VDD.n3208 VDD.n3207 0.806
R5984 VDD.n2943 VDD.n2942 0.806
R5985 VDD.n3381 VDD.n3380 0.806
R5986 VDD.n3324 VDD.n3323 0.806
R5987 VDD.n202 VDD.n201 0.806
R5988 VDD.n3267 VDD.n3266 0.806
R5989 VDD.n34 VDD.n33 0.806
R5990 VDD.n4 VDD.n3 0.806
R5991 VDD.n85 VDD.n84 0.806
R5992 VDD.n144 VDD.n143 0.806
R5993 VDD.n3262 VDD.n2663 0.793
R5994 VDD.n2870 VDD.n2869 0.778
R5995 VDD.n2842 VDD.n2841 0.778
R5996 VDD.n531 VDD.n530 0.778
R5997 VDD.n377 VDD.n376 0.778
R5998 VDD.n3031 VDD.n3030 0.778
R5999 VDD.n2949 VDD.n2948 0.778
R6000 VDD.n3014 VDD.n3013 0.778
R6001 VDD.n3376 VDD.n3375 0.778
R6002 VDD.n3319 VDD.n3318 0.778
R6003 VDD.n207 VDD.n206 0.778
R6004 VDD.n39 VDD.n38 0.778
R6005 VDD.n9 VDD.n8 0.778
R6006 VDD.n90 VDD.n89 0.778
R6007 VDD.n149 VDD.n148 0.778
R6008 VDD.n3403 VDD.n3402 0.778
R6009 VDD.n561 VDD.n559 0.777
R6010 VDD.n1746 VDD.n1745 0.756
R6011 VDD.n1771 VDD.n1770 0.756
R6012 VDD.n1821 VDD.n1820 0.756
R6013 VDD.n1796 VDD.n1795 0.756
R6014 VDD.n1721 VDD.n1720 0.756
R6015 VDD.n1697 VDD.n1696 0.756
R6016 VDD.n2398 VDD.n2390 0.756
R6017 VDD.n2338 VDD.n2330 0.756
R6018 VDD.n2358 VDD.n2350 0.756
R6019 VDD.n2378 VDD.n2370 0.756
R6020 VDD.n3244 VDD.n3243 0.747
R6021 VDD.n2938 VDD.n2937 0.747
R6022 VDD.n2907 VDD.n2906 0.747
R6023 VDD.n2903 VDD.n2902 0.747
R6024 VDD.n2905 VDD.n2904 0.747
R6025 VDD.n2680 VDD.n2679 0.747
R6026 VDD.n2676 VDD.n2675 0.747
R6027 VDD.n2678 VDD.n2677 0.747
R6028 VDD.n2671 VDD.n2670 0.747
R6029 VDD.n2667 VDD.n2666 0.747
R6030 VDD.n2669 VDD.n2668 0.747
R6031 VDD.n2893 VDD.n2892 0.747
R6032 VDD.n2684 VDD.n2683 0.747
R6033 VDD.n2858 VDD.n2857 0.747
R6034 VDD.n2749 VDD.n2748 0.747
R6035 VDD.n2827 VDD.n2826 0.747
R6036 VDD.n2812 VDD.n2811 0.747
R6037 VDD.n2915 VDD.n2914 0.747
R6038 VDD.n2911 VDD.n2910 0.747
R6039 VDD.n2913 VDD.n2912 0.747
R6040 VDD.n310 VDD.n309 0.747
R6041 VDD.n306 VDD.n305 0.747
R6042 VDD.n308 VDD.n307 0.747
R6043 VDD.n301 VDD.n300 0.747
R6044 VDD.n297 VDD.n296 0.747
R6045 VDD.n299 VDD.n298 0.747
R6046 VDD.n392 VDD.n391 0.747
R6047 VDD.n388 VDD.n387 0.747
R6048 VDD.n390 VDD.n389 0.747
R6049 VDD.n401 VDD.n400 0.747
R6050 VDD.n397 VDD.n396 0.747
R6051 VDD.n399 VDD.n398 0.747
R6052 VDD.n3110 VDD.n3109 0.747
R6053 VDD.n3090 VDD.n3089 0.747
R6054 VDD.n3134 VDD.n3133 0.747
R6055 VDD.n3019 VDD.n3018 0.747
R6056 VDD.n3222 VDD.n3221 0.747
R6057 VDD.n3009 VDD.n3008 0.747
R6058 VDD.n2982 VDD.n2981 0.747
R6059 VDD.n2965 VDD.n2964 0.747
R6060 VDD.n2973 VDD.n2972 0.747
R6061 VDD.n2969 VDD.n2968 0.747
R6062 VDD.n3157 VDD.n3156 0.747
R6063 VDD.n3141 VDD.n3140 0.747
R6064 VDD.n3145 VDD.n3144 0.747
R6065 VDD.n3151 VDD.n3150 0.747
R6066 VDD.n3051 VDD.n3050 0.747
R6067 VDD.n3036 VDD.n3035 0.747
R6068 VDD.n3039 VDD.n3038 0.747
R6069 VDD.n3045 VDD.n3044 0.747
R6070 VDD.n2661 VDD.n2660 0.747
R6071 VDD.n2657 VDD.n2656 0.747
R6072 VDD.n2659 VDD.n2658 0.747
R6073 VDD.n714 VDD.n713 0.747
R6074 VDD.n710 VDD.n709 0.747
R6075 VDD.n712 VDD.n711 0.747
R6076 VDD.n2653 VDD.n2652 0.747
R6077 VDD.n2649 VDD.n2648 0.747
R6078 VDD.n2651 VDD.n2650 0.747
R6079 VDD.n706 VDD.n705 0.747
R6080 VDD.n702 VDD.n701 0.747
R6081 VDD.n704 VDD.n703 0.747
R6082 VDD.n732 VDD.n731 0.747
R6083 VDD.n735 VDD.n734 0.747
R6084 VDD.n737 VDD.n736 0.747
R6085 VDD.n608 VDD.n607 0.747
R6086 VDD.n604 VDD.n603 0.747
R6087 VDD.n606 VDD.n605 0.747
R6088 VDD.n293 VDD.n292 0.747
R6089 VDD.n289 VDD.n288 0.747
R6090 VDD.n291 VDD.n290 0.747
R6091 VDD.n3274 VDD.n3273 0.747
R6092 VDD.n3270 VDD.n3269 0.747
R6093 VDD.n3331 VDD.n3330 0.747
R6094 VDD.n3327 VDD.n3326 0.747
R6095 VDD.n3388 VDD.n3387 0.747
R6096 VDD.n3384 VDD.n3383 0.747
R6097 VDD.n197 VDD.n196 0.747
R6098 VDD.n193 VDD.n192 0.747
R6099 VDD.n848 VDD.n847 0.747
R6100 VDD.n852 VDD.n851 0.747
R6101 VDD.n828 VDD.n827 0.747
R6102 VDD.n832 VDD.n831 0.747
R6103 VDD.n24 VDD.n23 0.747
R6104 VDD.n28 VDD.n27 0.747
R6105 VDD.n823 VDD.n822 0.747
R6106 VDD.n820 VDD.n819 0.747
R6107 VDD.n805 VDD.n804 0.747
R6108 VDD.n809 VDD.n808 0.747
R6109 VDD.n134 VDD.n133 0.747
R6110 VDD.n138 VDD.n137 0.747
R6111 VDD.n160 VDD.n159 0.747
R6112 VDD.n164 VDD.n163 0.747
R6113 VDD.n152 VDD.n151 0.747
R6114 VDD.n156 VDD.n155 0.747
R6115 VDD.n101 VDD.n100 0.747
R6116 VDD.n105 VDD.n104 0.747
R6117 VDD.n93 VDD.n92 0.747
R6118 VDD.n97 VDD.n96 0.747
R6119 VDD.n50 VDD.n49 0.747
R6120 VDD.n54 VDD.n53 0.747
R6121 VDD.n42 VDD.n41 0.747
R6122 VDD.n46 VDD.n45 0.747
R6123 VDD.n3434 VDD.n3433 0.747
R6124 VDD.n3430 VDD.n3429 0.747
R6125 VDD.n3437 VDD.n3436 0.747
R6126 VDD.n3440 VDD.n3439 0.747
R6127 VDD.n3292 VDD.n3291 0.747
R6128 VDD.n3288 VDD.n3287 0.747
R6129 VDD.n3295 VDD.n3294 0.747
R6130 VDD.n3298 VDD.n3297 0.747
R6131 VDD.n3349 VDD.n3348 0.747
R6132 VDD.n3345 VDD.n3344 0.747
R6133 VDD.n3352 VDD.n3351 0.747
R6134 VDD.n3355 VDD.n3354 0.747
R6135 VDD.n225 VDD.n224 0.747
R6136 VDD.n221 VDD.n220 0.747
R6137 VDD.n228 VDD.n227 0.747
R6138 VDD.n231 VDD.n230 0.747
R6139 VDD.n326 VDD.n325 0.747
R6140 VDD.n331 VDD.n330 0.747
R6141 VDD.n314 VDD.n313 0.747
R6142 VDD.n320 VDD.n319 0.747
R6143 VDD.n433 VDD.n432 0.747
R6144 VDD.n418 VDD.n417 0.747
R6145 VDD.n493 VDD.n492 0.747
R6146 VDD.n499 VDD.n498 0.747
R6147 VDD.n2784 VDD.n2783 0.747
R6148 VDD.n2769 VDD.n2768 0.747
R6149 VDD.n2722 VDD.n2721 0.747
R6150 VDD.n2716 VDD.n2715 0.747
R6151 VDD.n568 VDD.n566 0.74
R6152 VDD.n3246 VDD.n3242 0.689
R6153 VDD.n3258 VDD.n3257 0.689
R6154 VDD.n3256 VDD.n3252 0.689
R6155 VDD.n3255 VDD.n3253 0.689
R6156 VDD.n2895 VDD.n2891 0.689
R6157 VDD.n2860 VDD.n2856 0.689
R6158 VDD.n2829 VDD.n2825 0.689
R6159 VDD.n549 VDD.n548 0.689
R6160 VDD.n550 VDD.n547 0.689
R6161 VDD.n546 VDD.n544 0.689
R6162 VDD.n406 VDD.n404 0.689
R6163 VDD.n407 VDD.n403 0.689
R6164 VDD.n409 VDD.n408 0.689
R6165 VDD.n2923 VDD.n2921 0.689
R6166 VDD.n2924 VDD.n2920 0.689
R6167 VDD.n2926 VDD.n2925 0.689
R6168 VDD.n3112 VDD.n3108 0.689
R6169 VDD.n3136 VDD.n3132 0.689
R6170 VDD.n3224 VDD.n3220 0.689
R6171 VDD.n2984 VDD.n2980 0.689
R6172 VDD.n2975 VDD.n2971 0.689
R6173 VDD.n3159 VDD.n3155 0.689
R6174 VDD.n3147 VDD.n3143 0.689
R6175 VDD.n3053 VDD.n3049 0.689
R6176 VDD.n3041 VDD.n3037 0.689
R6177 VDD.n283 VDD.n282 0.689
R6178 VDD.n281 VDD.n277 0.689
R6179 VDD.n280 VDD.n278 0.689
R6180 VDD.n272 VDD.n271 0.689
R6181 VDD.n270 VDD.n266 0.689
R6182 VDD.n269 VDD.n267 0.689
R6183 VDD.n3271 VDD.n3268 0.689
R6184 VDD.n3328 VDD.n3325 0.689
R6185 VDD.n3385 VDD.n3382 0.689
R6186 VDD.n194 VDD.n191 0.689
R6187 VDD.n849 VDD.n846 0.689
R6188 VDD.n829 VDD.n826 0.689
R6189 VDD.n25 VDD.n22 0.689
R6190 VDD.n824 VDD.n821 0.689
R6191 VDD.n806 VDD.n803 0.689
R6192 VDD.n135 VDD.n132 0.689
R6193 VDD.n161 VDD.n158 0.689
R6194 VDD.n153 VDD.n150 0.689
R6195 VDD.n102 VDD.n99 0.689
R6196 VDD.n94 VDD.n91 0.689
R6197 VDD.n51 VDD.n48 0.689
R6198 VDD.n43 VDD.n40 0.689
R6199 VDD.n3431 VDD.n3428 0.689
R6200 VDD.n3441 VDD.n3438 0.689
R6201 VDD.n3289 VDD.n3286 0.689
R6202 VDD.n3299 VDD.n3296 0.689
R6203 VDD.n3346 VDD.n3343 0.689
R6204 VDD.n3356 VDD.n3353 0.689
R6205 VDD.n222 VDD.n219 0.689
R6206 VDD.n232 VDD.n229 0.689
R6207 VDD.n328 VDD.n324 0.689
R6208 VDD.n316 VDD.n312 0.689
R6209 VDD.n435 VDD.n431 0.689
R6210 VDD.n424 VDD.n423 0.689
R6211 VDD.n425 VDD.n422 0.689
R6212 VDD.n421 VDD.n419 0.689
R6213 VDD.n495 VDD.n491 0.689
R6214 VDD.n485 VDD.n484 0.689
R6215 VDD.n486 VDD.n483 0.689
R6216 VDD.n482 VDD.n480 0.689
R6217 VDD.n2786 VDD.n2782 0.689
R6218 VDD.n2775 VDD.n2774 0.689
R6219 VDD.n2776 VDD.n2773 0.689
R6220 VDD.n2772 VDD.n2770 0.689
R6221 VDD.n2724 VDD.n2720 0.689
R6222 VDD.n2708 VDD.n2707 0.689
R6223 VDD.n2709 VDD.n2706 0.689
R6224 VDD.n2705 VDD.n2703 0.689
R6225 VDD.n1081 VDD.n1079 0.689
R6226 VDD.n1082 VDD.n1078 0.689
R6227 VDD.n1077 VDD.n1076 0.689
R6228 VDD.n1089 VDD.n1087 0.689
R6229 VDD.n1090 VDD.n1086 0.689
R6230 VDD.n1085 VDD.n1084 0.689
R6231 VDD.n1122 VDD.n1120 0.689
R6232 VDD.n1123 VDD.n1119 0.689
R6233 VDD.n1118 VDD.n1117 0.689
R6234 VDD.n1114 VDD.n1112 0.689
R6235 VDD.n1115 VDD.n1111 0.689
R6236 VDD.n1110 VDD.n1109 0.689
R6237 VDD.n1105 VDD.n1103 0.689
R6238 VDD.n1106 VDD.n1102 0.689
R6239 VDD.n1101 VDD.n1100 0.689
R6240 VDD.n1097 VDD.n1095 0.689
R6241 VDD.n1098 VDD.n1094 0.689
R6242 VDD.n1093 VDD.n1092 0.689
R6243 VDD.n1072 VDD.n1070 0.689
R6244 VDD.n1073 VDD.n1069 0.689
R6245 VDD.n1068 VDD.n1067 0.689
R6246 VDD.n1064 VDD.n1062 0.689
R6247 VDD.n1065 VDD.n1061 0.689
R6248 VDD.n1060 VDD.n1059 0.689
R6249 VDD.n2956 VDD.n2955 0.686
R6250 VDD.n2961 VDD.n2960 0.686
R6251 VDD.n2991 VDD.n2990 0.686
R6252 VDD.n2996 VDD.n2995 0.686
R6253 VDD.n3180 VDD.n3179 0.686
R6254 VDD.n3185 VDD.n3184 0.686
R6255 VDD.n3167 VDD.n3166 0.686
R6256 VDD.n3172 VDD.n3171 0.686
R6257 VDD.n3080 VDD.n3079 0.686
R6258 VDD.n3085 VDD.n3084 0.686
R6259 VDD.n3061 VDD.n3060 0.686
R6260 VDD.n3066 VDD.n3065 0.686
R6261 VDD.n727 VDD.n726 0.686
R6262 VDD.n722 VDD.n721 0.686
R6263 VDD.n597 VDD.n596 0.686
R6264 VDD.n592 VDD.n591 0.686
R6265 VDD.n578 VDD.n577 0.686
R6266 VDD.n583 VDD.n582 0.686
R6267 VDD.n261 VDD.n260 0.686
R6268 VDD.n256 VDD.n255 0.686
R6269 VDD.n183 VDD.n182 0.686
R6270 VDD.n188 VDD.n187 0.686
R6271 VDD.n171 VDD.n170 0.686
R6272 VDD.n176 VDD.n175 0.686
R6273 VDD.n124 VDD.n123 0.686
R6274 VDD.n129 VDD.n128 0.686
R6275 VDD.n112 VDD.n111 0.686
R6276 VDD.n117 VDD.n116 0.686
R6277 VDD.n838 VDD.n837 0.686
R6278 VDD.n843 VDD.n842 0.686
R6279 VDD.n14 VDD.n13 0.686
R6280 VDD.n19 VDD.n18 0.686
R6281 VDD.n73 VDD.n72 0.686
R6282 VDD.n78 VDD.n77 0.686
R6283 VDD.n61 VDD.n60 0.686
R6284 VDD.n66 VDD.n65 0.686
R6285 VDD.n3426 VDD.n3425 0.686
R6286 VDD.n3421 VDD.n3420 0.686
R6287 VDD.n3415 VDD.n3414 0.686
R6288 VDD.n3410 VDD.n3409 0.686
R6289 VDD.n3279 VDD.n3278 0.686
R6290 VDD.n3284 VDD.n3283 0.686
R6291 VDD.n3307 VDD.n3306 0.686
R6292 VDD.n3312 VDD.n3311 0.686
R6293 VDD.n3336 VDD.n3335 0.686
R6294 VDD.n3341 VDD.n3340 0.686
R6295 VDD.n3364 VDD.n3363 0.686
R6296 VDD.n3369 VDD.n3368 0.686
R6297 VDD.n212 VDD.n211 0.686
R6298 VDD.n217 VDD.n216 0.686
R6299 VDD.n240 VDD.n239 0.686
R6300 VDD.n245 VDD.n244 0.686
R6301 VDD.n361 VDD.n360 0.686
R6302 VDD.n366 VDD.n365 0.686
R6303 VDD.n343 VDD.n342 0.686
R6304 VDD.n348 VDD.n347 0.686
R6305 VDD.n461 VDD.n460 0.686
R6306 VDD.n466 VDD.n465 0.686
R6307 VDD.n442 VDD.n441 0.686
R6308 VDD.n447 VDD.n446 0.686
R6309 VDD.n473 VDD.n472 0.686
R6310 VDD.n478 VDD.n477 0.686
R6311 VDD.n510 VDD.n509 0.686
R6312 VDD.n515 VDD.n514 0.686
R6313 VDD.n2760 VDD.n2759 0.686
R6314 VDD.n2765 VDD.n2764 0.686
R6315 VDD.n2794 VDD.n2793 0.686
R6316 VDD.n2799 VDD.n2798 0.686
R6317 VDD.n2696 VDD.n2695 0.686
R6318 VDD.n2701 VDD.n2700 0.686
R6319 VDD.n2731 VDD.n2730 0.686
R6320 VDD.n2736 VDD.n2735 0.686
R6321 VDD.n2185 VDD.n2184 0.686
R6322 VDD.n2171 VDD.n2170 0.686
R6323 VDD.n2153 VDD.n2152 0.686
R6324 VDD.n1472 VDD.n1471 0.686
R6325 VDD.n1458 VDD.n1457 0.686
R6326 VDD.n2033 VDD.n2032 0.686
R6327 VDD.n2048 VDD.n2047 0.686
R6328 VDD.n1933 VDD.n1932 0.686
R6329 VDD.n1948 VDD.n1947 0.686
R6330 VDD.n1883 VDD.n1882 0.686
R6331 VDD.n1898 VDD.n1897 0.686
R6332 VDD.n1908 VDD.n1907 0.686
R6333 VDD.n1923 VDD.n1922 0.686
R6334 VDD.n1958 VDD.n1957 0.686
R6335 VDD.n1973 VDD.n1972 0.686
R6336 VDD.n1983 VDD.n1982 0.686
R6337 VDD.n1998 VDD.n1997 0.686
R6338 VDD.n2008 VDD.n2007 0.686
R6339 VDD.n2023 VDD.n2022 0.686
R6340 VDD.n2058 VDD.n2057 0.686
R6341 VDD.n2073 VDD.n2072 0.686
R6342 VDD.n2621 VDD.n2620 0.686
R6343 VDD.n2616 VDD.n2615 0.686
R6344 VDD.n2444 VDD.n2443 0.686
R6345 VDD.n2430 VDD.n2429 0.686
R6346 VDD.n2419 VDD.n2418 0.686
R6347 VDD.n2405 VDD.n2404 0.686
R6348 VDD.n2235 VDD.n2234 0.686
R6349 VDD.n2221 VDD.n2220 0.686
R6350 VDD.n2210 VDD.n2209 0.686
R6351 VDD.n2196 VDD.n2195 0.686
R6352 VDD.n1052 VDD.n1044 0.646
R6353 VDD.n927 VDD.n919 0.646
R6354 VDD.n952 VDD.n944 0.646
R6355 VDD.n1027 VDD.n1019 0.646
R6356 VDD.n1002 VDD.n994 0.646
R6357 VDD.n977 VDD.n969 0.646
R6358 VDD.n902 VDD.n894 0.646
R6359 VDD.n878 VDD.n870 0.646
R6360 VDD.n641 VDD.n640 0.646
R6361 VDD.n659 VDD.n658 0.646
R6362 VDD.n677 VDD.n676 0.646
R6363 VDD.n694 VDD.n693 0.646
R6364 VDD.n623 VDD.n622 0.646
R6365 VDD.n754 VDD.n753 0.646
R6366 VDD.n772 VDD.n771 0.646
R6367 VDD.n790 VDD.n789 0.646
R6368 VDD.n1871 VDD.n1863 0.646
R6369 VDD.n1846 VDD.n1838 0.646
R6370 VDD.n1546 VDD.n1538 0.646
R6371 VDD.n1571 VDD.n1563 0.646
R6372 VDD.n1671 VDD.n1663 0.646
R6373 VDD.n1646 VDD.n1638 0.646
R6374 VDD.n1621 VDD.n1613 0.646
R6375 VDD.n1596 VDD.n1588 0.646
R6376 VDD.n1521 VDD.n1513 0.646
R6377 VDD.n1497 VDD.n1489 0.646
R6378 VDD.n1396 VDD.n1388 0.646
R6379 VDD.n1371 VDD.n1363 0.646
R6380 VDD.n1272 VDD.n1264 0.646
R6381 VDD.n1296 VDD.n1288 0.646
R6382 VDD.n1321 VDD.n1313 0.646
R6383 VDD.n1346 VDD.n1338 0.646
R6384 VDD.n1421 VDD.n1413 0.646
R6385 VDD.n1446 VDD.n1438 0.646
R6386 VDD.n2607 VDD.n2606 0.646
R6387 VDD.n2468 VDD.n2467 0.646
R6388 VDD.n2487 VDD.n2486 0.646
R6389 VDD.n2547 VDD.n2546 0.646
R6390 VDD.n2567 VDD.n2566 0.646
R6391 VDD.n2587 VDD.n2586 0.646
R6392 VDD.n2527 VDD.n2526 0.646
R6393 VDD.n2507 VDD.n2506 0.646
R6394 VDD.n2259 VDD.n2258 0.646
R6395 VDD.n2278 VDD.n2277 0.646
R6396 VDD.n2318 VDD.n2317 0.646
R6397 VDD.n2298 VDD.n2297 0.646
R6398 VDD.n982 VDD.n957 0.643
R6399 VDD.n1802 VDD.n1777 0.643
R6400 VDD.n1602 VDD.n1577 0.643
R6401 VDD.n1377 VDD.n1352 0.643
R6402 VDD.n907 VDD.n882 0.632
R6403 VDD.n1727 VDD.n1702 0.632
R6404 VDD.n1527 VDD.n1502 0.632
R6405 VDD.n1302 VDD.n1277 0.632
R6406 VDD.n1007 VDD.n982 0.631
R6407 VDD.n957 VDD.n932 0.631
R6408 VDD.n1877 VDD.n1852 0.631
R6409 VDD.n1827 VDD.n1802 0.631
R6410 VDD.n1777 VDD.n1752 0.631
R6411 VDD.n1677 VDD.n1652 0.631
R6412 VDD.n1627 VDD.n1602 0.631
R6413 VDD.n1577 VDD.n1552 0.631
R6414 VDD.n1452 VDD.n1427 0.631
R6415 VDD.n1402 VDD.n1377 0.631
R6416 VDD.n1352 VDD.n1327 0.631
R6417 VDD.n1032 VDD.n1007 0.629
R6418 VDD.n932 VDD.n907 0.629
R6419 VDD.n1852 VDD.n1827 0.629
R6420 VDD.n1752 VDD.n1727 0.629
R6421 VDD.n1652 VDD.n1627 0.629
R6422 VDD.n1552 VDD.n1527 0.629
R6423 VDD.n1427 VDD.n1402 0.629
R6424 VDD.n1327 VDD.n1302 0.629
R6425 VDD.n3271 VDD.n3270 0.59
R6426 VDD.n3328 VDD.n3327 0.59
R6427 VDD.n3385 VDD.n3384 0.59
R6428 VDD.n194 VDD.n193 0.59
R6429 VDD.n849 VDD.n848 0.59
R6430 VDD.n829 VDD.n828 0.59
R6431 VDD.n25 VDD.n24 0.59
R6432 VDD.n824 VDD.n823 0.59
R6433 VDD.n806 VDD.n805 0.59
R6434 VDD.n135 VDD.n134 0.59
R6435 VDD.n161 VDD.n160 0.59
R6436 VDD.n153 VDD.n152 0.59
R6437 VDD.n102 VDD.n101 0.59
R6438 VDD.n94 VDD.n93 0.59
R6439 VDD.n51 VDD.n50 0.59
R6440 VDD.n43 VDD.n42 0.59
R6441 VDD.n3431 VDD.n3430 0.59
R6442 VDD.n3441 VDD.n3440 0.59
R6443 VDD.n3289 VDD.n3288 0.59
R6444 VDD.n3299 VDD.n3298 0.59
R6445 VDD.n3346 VDD.n3345 0.59
R6446 VDD.n3356 VDD.n3355 0.59
R6447 VDD.n222 VDD.n221 0.59
R6448 VDD.n232 VDD.n231 0.59
R6449 VDD.n2148 VDD.n2146 0.587
R6450 VDD.n3245 VDD.n3244 0.571
R6451 VDD.n2859 VDD.n2858 0.571
R6452 VDD.n3223 VDD.n3222 0.571
R6453 VDD.n2974 VDD.n2973 0.571
R6454 VDD.n3158 VDD.n3157 0.571
R6455 VDD.n3052 VDD.n3051 0.571
R6456 VDD.n3040 VDD.n3039 0.571
R6457 VDD.n327 VDD.n326 0.571
R6458 VDD.n315 VDD.n314 0.571
R6459 VDD.n494 VDD.n493 0.571
R6460 VDD.n2723 VDD.n2722 0.571
R6461 VDD.n3135 VDD.n3134 0.57
R6462 VDD.n2983 VDD.n2982 0.57
R6463 VDD.n434 VDD.n433 0.57
R6464 VDD.n2894 VDD.n2893 0.569
R6465 VDD.n2828 VDD.n2827 0.569
R6466 VDD.n3111 VDD.n3110 0.569
R6467 VDD.n3146 VDD.n3145 0.569
R6468 VDD.n2785 VDD.n2784 0.569
R6469 VDD.n3259 VDD.n3258 0.5
R6470 VDD.n410 VDD.n409 0.5
R6471 VDD.n2927 VDD.n2926 0.5
R6472 VDD.n284 VDD.n283 0.5
R6473 VDD.n273 VDD.n272 0.5
R6474 VDD.n1083 VDD.n1077 0.5
R6475 VDD.n1091 VDD.n1085 0.5
R6476 VDD.n1124 VDD.n1118 0.5
R6477 VDD.n1116 VDD.n1110 0.5
R6478 VDD.n1107 VDD.n1101 0.5
R6479 VDD.n1099 VDD.n1093 0.5
R6480 VDD.n1074 VDD.n1068 0.5
R6481 VDD.n1066 VDD.n1060 0.5
R6482 VDD.n3259 VDD.n3256 0.483
R6483 VDD.n410 VDD.n407 0.483
R6484 VDD.n2927 VDD.n2924 0.483
R6485 VDD.n284 VDD.n281 0.483
R6486 VDD.n273 VDD.n270 0.483
R6487 VDD.n1083 VDD.n1082 0.483
R6488 VDD.n1091 VDD.n1090 0.483
R6489 VDD.n1124 VDD.n1123 0.483
R6490 VDD.n1116 VDD.n1115 0.483
R6491 VDD.n1107 VDD.n1106 0.483
R6492 VDD.n1099 VDD.n1098 0.483
R6493 VDD.n1074 VDD.n1073 0.483
R6494 VDD.n1066 VDD.n1065 0.483
R6495 VDD.n1053 VDD.n1039 0.465
R6496 VDD.n928 VDD.n914 0.465
R6497 VDD.n953 VDD.n939 0.465
R6498 VDD.n1028 VDD.n1014 0.465
R6499 VDD.n1003 VDD.n989 0.465
R6500 VDD.n978 VDD.n964 0.465
R6501 VDD.n903 VDD.n889 0.465
R6502 VDD.n879 VDD.n865 0.465
R6503 VDD.n1747 VDD.n1733 0.465
R6504 VDD.n1772 VDD.n1758 0.465
R6505 VDD.n1872 VDD.n1858 0.465
R6506 VDD.n1847 VDD.n1833 0.465
R6507 VDD.n1822 VDD.n1808 0.465
R6508 VDD.n1797 VDD.n1783 0.465
R6509 VDD.n1722 VDD.n1708 0.465
R6510 VDD.n1698 VDD.n1684 0.465
R6511 VDD.n1547 VDD.n1533 0.465
R6512 VDD.n1572 VDD.n1558 0.465
R6513 VDD.n1672 VDD.n1658 0.465
R6514 VDD.n1647 VDD.n1633 0.465
R6515 VDD.n1622 VDD.n1608 0.465
R6516 VDD.n1597 VDD.n1583 0.465
R6517 VDD.n1522 VDD.n1508 0.465
R6518 VDD.n1498 VDD.n1484 0.465
R6519 VDD.n1397 VDD.n1383 0.465
R6520 VDD.n1372 VDD.n1358 0.465
R6521 VDD.n1273 VDD.n1259 0.465
R6522 VDD.n1297 VDD.n1283 0.465
R6523 VDD.n1322 VDD.n1308 0.465
R6524 VDD.n1347 VDD.n1333 0.465
R6525 VDD.n1422 VDD.n1408 0.465
R6526 VDD.n1447 VDD.n1433 0.465
R6527 VDD.n2608 VDD.n2591 0.465
R6528 VDD.n2469 VDD.n2452 0.465
R6529 VDD.n2488 VDD.n2471 0.465
R6530 VDD.n2548 VDD.n2531 0.465
R6531 VDD.n2568 VDD.n2551 0.465
R6532 VDD.n2588 VDD.n2571 0.465
R6533 VDD.n2528 VDD.n2511 0.465
R6534 VDD.n2508 VDD.n2491 0.465
R6535 VDD.n2399 VDD.n2382 0.465
R6536 VDD.n2260 VDD.n2243 0.465
R6537 VDD.n2279 VDD.n2262 0.465
R6538 VDD.n2339 VDD.n2322 0.465
R6539 VDD.n2359 VDD.n2342 0.465
R6540 VDD.n2379 VDD.n2362 0.465
R6541 VDD.n2319 VDD.n2302 0.465
R6542 VDD.n2299 VDD.n2282 0.465
R6543 VDD.n3105 VDD.n3090 0.452
R6544 VDD.n2986 VDD.n2965 0.452
R6545 VDD.n2789 VDD.n2769 0.452
R6546 VDD.n2888 VDD.n2684 0.452
R6547 VDD.n2824 VDD.n2812 0.452
R6548 VDD.n3130 VDD.n3019 0.452
R6549 VDD.n437 VDD.n418 0.452
R6550 VDD.n3152 VDD.n3151 0.452
R6551 VDD.n3241 VDD.n2938 0.451
R6552 VDD.n2855 VDD.n2749 0.451
R6553 VDD.n3219 VDD.n3009 0.451
R6554 VDD.n3162 VDD.n3141 0.451
R6555 VDD.n3056 VDD.n3036 0.451
R6556 VDD.n3397 VDD.n3274 0.451
R6557 VDD.n3393 VDD.n3331 0.451
R6558 VDD.n3389 VDD.n3388 0.451
R6559 VDD.n251 VDD.n197 0.451
R6560 VDD.n853 VDD.n852 0.451
R6561 VDD.n833 VDD.n832 0.451
R6562 VDD.n29 VDD.n28 0.451
R6563 VDD.n825 VDD.n820 0.451
R6564 VDD.n810 VDD.n809 0.451
R6565 VDD.n139 VDD.n138 0.451
R6566 VDD.n165 VDD.n164 0.451
R6567 VDD.n157 VDD.n156 0.451
R6568 VDD.n106 VDD.n105 0.451
R6569 VDD.n98 VDD.n97 0.451
R6570 VDD.n55 VDD.n54 0.451
R6571 VDD.n47 VDD.n46 0.451
R6572 VDD.n3443 VDD.n3434 0.451
R6573 VDD.n3442 VDD.n3437 0.451
R6574 VDD.n3301 VDD.n3292 0.451
R6575 VDD.n3300 VDD.n3295 0.451
R6576 VDD.n3358 VDD.n3349 0.451
R6577 VDD.n3357 VDD.n3352 0.451
R6578 VDD.n234 VDD.n225 0.451
R6579 VDD.n233 VDD.n228 0.451
R6580 VDD.n3046 VDD.n3045 0.451
R6581 VDD.n321 VDD.n320 0.451
R6582 VDD.n2970 VDD.n2969 0.45
R6583 VDD.n1250 VDD.n1249 0.45
R6584 VDD.n2717 VDD.n2716 0.449
R6585 VDD.n2141 VDD.n2140 0.446
R6586 VDD.n1252 VDD.n1251 0.444
R6587 VDD.n1248 VDD.n1247 0.444
R6588 VDD.n2916 VDD.n2915 0.433
R6589 VDD.n1253 VDD.n1252 0.429
R6590 VDD.n1251 VDD.n1250 0.429
R6591 VDD.n1249 VDD.n1248 0.429
R6592 VDD.n1247 VDD.n1246 0.429
R6593 VDD.n332 VDD.n331 0.419
R6594 VDD.n500 VDD.n499 0.419
R6595 VDD.n2916 VDD.n2913 0.416
R6596 VDD.n2691 VDD.n2690 0.4
R6597 VDD.n2844 VDD.n2843 0.4
R6598 VDD.n3097 VDD.n3096 0.4
R6599 VDD.n379 VDD.n378 0.4
R6600 VDD.n3026 VDD.n3025 0.4
R6601 VDD.n3033 VDD.n3032 0.4
R6602 VDD.n3210 VDD.n3209 0.4
R6603 VDD.n2951 VDD.n2950 0.4
R6604 VDD.n3016 VDD.n3015 0.4
R6605 VDD.n2140 VDD.n2139 0.398
R6606 VDD.n2139 VDD.n2138 0.398
R6607 VDD.n2138 VDD.n2137 0.398
R6608 VDD.n2137 VDD.n2136 0.398
R6609 VDD.n2136 VDD.n2135 0.398
R6610 VDD.n2135 VDD.n2134 0.398
R6611 VDD.n2134 VDD.n2133 0.398
R6612 VDD.n2124 VDD.n2123 0.386
R6613 VDD.n2118 VDD.n2117 0.386
R6614 VDD.n2112 VDD.n2111 0.386
R6615 VDD.n2106 VDD.n2105 0.386
R6616 VDD.n2100 VDD.n2099 0.386
R6617 VDD.n2082 VDD.n2081 0.386
R6618 VDD.n2094 VDD.n2093 0.38
R6619 VDD.n2088 VDD.n2087 0.369
R6620 VDD.n2639 VDD.n2400 0.347
R6621 VDD.n3285 VDD.n3279 0.345
R6622 VDD.n3313 VDD.n3307 0.345
R6623 VDD.n3342 VDD.n3336 0.345
R6624 VDD.n3370 VDD.n3364 0.345
R6625 VDD.n218 VDD.n212 0.345
R6626 VDD.n246 VDD.n240 0.345
R6627 VDD.n584 VDD.n578 0.343
R6628 VDD.n584 VDD.n583 0.343
R6629 VDD.n3427 VDD.n3421 0.342
R6630 VDD.n3416 VDD.n3410 0.342
R6631 VDD.n3285 VDD.n3284 0.34
R6632 VDD.n3313 VDD.n3312 0.34
R6633 VDD.n3342 VDD.n3341 0.34
R6634 VDD.n3370 VDD.n3369 0.34
R6635 VDD.n218 VDD.n217 0.34
R6636 VDD.n246 VDD.n245 0.34
R6637 VDD.n3427 VDD.n3426 0.336
R6638 VDD.n3416 VDD.n3415 0.336
R6639 VDD.n2622 VDD.n2616 0.334
R6640 VDD.n777 VDD.n251 0.326
R6641 VDD.n1246 VDD.n1245 0.315
R6642 VDD.n2133 VDD.n2132 0.309
R6643 VDD.n2154 VDD.n2153 0.305
R6644 VDD.n2622 VDD.n2621 0.305
R6645 VDD.n384 VDD.n383 0.303
R6646 VDD.n2636 VDD.n2609 0.297
R6647 VDD.n562 VDD.n561 0.295
R6648 VDD.n569 VDD.n568 0.286
R6649 VDD.n571 VDD.n415 0.286
R6650 VDD.n2154 VDD.n2148 0.284
R6651 VDD.n415 VDD.n414 0.283
R6652 VDD.n1227 VDD.n1226 0.283
R6653 VDD.n1230 VDD.n1229 0.281
R6654 VDD.n1245 VDD.n1232 0.28
R6655 VDD.n1232 VDD.n1231 0.28
R6656 VDD.n1231 VDD.n1230 0.28
R6657 VDD.n1229 VDD.n1228 0.28
R6658 VDD.n1228 VDD.n1227 0.28
R6659 VDD.n166 VDD.n157 0.276
R6660 VDD.n107 VDD.n98 0.276
R6661 VDD.n56 VDD.n47 0.276
R6662 VDD.n3262 VDD.n3261 0.275
R6663 VDD.n490 VDD.n489 0.272
R6664 VDD.n429 VDD.n428 0.272
R6665 VDD.n3443 VDD.n3442 0.272
R6666 VDD.n3301 VDD.n3300 0.272
R6667 VDD.n3358 VDD.n3357 0.272
R6668 VDD.n234 VDD.n233 0.272
R6669 VDD.n2780 VDD.n2779 0.271
R6670 VDD.n2713 VDD.n2712 0.271
R6671 VDD.n627 VDD.n626 0.271
R6672 VDD.n3048 VDD.n3047 0.271
R6673 VDD.n323 VDD.n322 0.271
R6674 VDD.n2978 VDD.n2977 0.271
R6675 VDD.n3154 VDD.n3153 0.271
R6676 VDD.n3450 VDD.n1453 0.255
R6677 VDD.n3390 VDD.n3381 0.254
R6678 VDD.n3394 VDD.n3324 0.254
R6679 VDD.n250 VDD.n202 0.254
R6680 VDD.n3398 VDD.n3267 0.254
R6681 VDD.n813 VDD.n34 0.253
R6682 VDD.n817 VDD.n4 0.253
R6683 VDD.n802 VDD.n85 0.253
R6684 VDD.n798 VDD.n144 0.253
R6685 VDD.n610 VDD.n600 0.252
R6686 VDD.n3196 VDD.n3195 0.244
R6687 VDD.n2085 VDD.t3388 0.243
R6688 VDD.n2091 VDD.t4027 0.243
R6689 VDD.n2121 VDD.t3761 0.243
R6690 VDD.n2115 VDD.t3021 0.243
R6691 VDD.n2109 VDD.t3448 0.243
R6692 VDD.n2103 VDD.t1992 0.243
R6693 VDD.n2097 VDD.t4404 0.243
R6694 VDD.n2079 VDD.t2331 0.243
R6695 VDD.n3404 VDD.n3403 0.242
R6696 VDD.n3391 VDD.n3376 0.242
R6697 VDD.n3395 VDD.n3319 0.242
R6698 VDD.n249 VDD.n207 0.242
R6699 VDD.n1166 VDD.n1165 0.241
R6700 VDD.n1181 VDD.n1180 0.241
R6701 VDD.n1226 VDD.n1225 0.241
R6702 VDD.n1211 VDD.n1210 0.241
R6703 VDD.n1196 VDD.n1195 0.241
R6704 VDD.n1154 VDD.n1153 0.241
R6705 VDD.n1139 VDD.n1138 0.241
R6706 VDD.n1244 VDD.n1243 0.241
R6707 VDD.n812 VDD.n39 0.241
R6708 VDD.n816 VDD.n9 0.241
R6709 VDD.n801 VDD.n90 0.241
R6710 VDD.n797 VDD.n149 0.241
R6711 VDD.n1678 VDD.n1677 0.238
R6712 VDD.n2141 VDD.n1877 0.236
R6713 VDD.n730 VDD.n717 0.233
R6714 VDD.n2280 VDD.n2260 0.231
R6715 VDD.n2691 VDD.n2689 0.23
R6716 VDD.n2755 VDD.n2754 0.23
R6717 VDD.n2818 VDD.n2817 0.23
R6718 VDD.n3097 VDD.n3095 0.23
R6719 VDD.n3026 VDD.n3024 0.23
R6720 VDD.n3210 VDD.n3208 0.23
R6721 VDD.n2944 VDD.n2943 0.23
R6722 VDD.n2935 VDD.n2934 0.228
R6723 VDD.n2340 VDD.n2320 0.228
R6724 VDD.n2360 VDD.n2340 0.224
R6725 VDD.n2320 VDD.n2300 0.224
R6726 VDD.n2380 VDD.n2360 0.223
R6727 VDD.n2300 VDD.n2280 0.223
R6728 VDD.n2644 VDD.n2141 0.221
R6729 VDD.n2871 VDD.n2870 0.218
R6730 VDD.n2844 VDD.n2842 0.218
R6731 VDD.n532 VDD.n531 0.218
R6732 VDD.n379 VDD.n377 0.218
R6733 VDD.n3033 VDD.n3031 0.218
R6734 VDD.n2951 VDD.n2949 0.218
R6735 VDD.n3016 VDD.n3014 0.218
R6736 VDD.n3449 VDD.n3448 0.217
R6737 VDD.n2400 VDD.n2380 0.211
R6738 VDD.n2908 VDD.n2907 0.208
R6739 VDD.n2681 VDD.n2680 0.208
R6740 VDD.n2672 VDD.n2671 0.208
R6741 VDD.n311 VDD.n310 0.208
R6742 VDD.n302 VDD.n301 0.208
R6743 VDD.n393 VDD.n392 0.208
R6744 VDD.n402 VDD.n401 0.208
R6745 VDD.n2662 VDD.n2661 0.208
R6746 VDD.n715 VDD.n714 0.208
R6747 VDD.n2663 VDD.n2653 0.208
R6748 VDD.n717 VDD.n706 0.208
R6749 VDD.n739 VDD.n732 0.208
R6750 VDD.n609 VDD.n608 0.208
R6751 VDD.n573 VDD.n293 0.208
R6752 VDD.n728 VDD.n722 0.203
R6753 VDD.n598 VDD.n592 0.203
R6754 VDD.n262 VDD.n256 0.203
R6755 VDD.n2908 VDD.n2905 0.195
R6756 VDD.n2681 VDD.n2678 0.195
R6757 VDD.n2672 VDD.n2669 0.195
R6758 VDD.n311 VDD.n308 0.195
R6759 VDD.n302 VDD.n299 0.195
R6760 VDD.n393 VDD.n390 0.195
R6761 VDD.n402 VDD.n399 0.195
R6762 VDD.n2662 VDD.n2659 0.195
R6763 VDD.n715 VDD.n712 0.195
R6764 VDD.n2663 VDD.n2651 0.195
R6765 VDD.n717 VDD.n704 0.195
R6766 VDD.n739 VDD.n737 0.195
R6767 VDD.n609 VDD.n606 0.195
R6768 VDD.n573 VDD.n291 0.195
R6769 VDD.n2489 VDD.n2469 0.195
R6770 VDD.n275 VDD.n264 0.195
R6771 VDD.n586 VDD.n573 0.194
R6772 VDD.n2186 VDD.n2185 0.193
R6773 VDD.n1473 VDD.n1472 0.193
R6774 VDD.n2049 VDD.n2048 0.193
R6775 VDD.n1949 VDD.n1948 0.193
R6776 VDD.n1899 VDD.n1898 0.193
R6777 VDD.n1924 VDD.n1923 0.193
R6778 VDD.n1974 VDD.n1973 0.193
R6779 VDD.n1999 VDD.n1998 0.193
R6780 VDD.n2024 VDD.n2023 0.193
R6781 VDD.n2074 VDD.n2073 0.193
R6782 VDD.n2445 VDD.n2444 0.193
R6783 VDD.n2420 VDD.n2419 0.193
R6784 VDD.n2236 VDD.n2235 0.193
R6785 VDD.n2211 VDD.n2210 0.193
R6786 VDD.n2549 VDD.n2529 0.192
R6787 VDD.n2172 VDD.n2171 0.189
R6788 VDD.n1459 VDD.n1458 0.189
R6789 VDD.n2034 VDD.n2033 0.189
R6790 VDD.n1934 VDD.n1933 0.189
R6791 VDD.n1884 VDD.n1883 0.189
R6792 VDD.n1909 VDD.n1908 0.189
R6793 VDD.n1959 VDD.n1958 0.189
R6794 VDD.n1984 VDD.n1983 0.189
R6795 VDD.n2009 VDD.n2008 0.189
R6796 VDD.n2059 VDD.n2058 0.189
R6797 VDD.n2431 VDD.n2430 0.189
R6798 VDD.n2406 VDD.n2405 0.189
R6799 VDD.n2222 VDD.n2221 0.189
R6800 VDD.n2197 VDD.n2196 0.189
R6801 VDD.n2589 VDD.n2569 0.188
R6802 VDD.n2569 VDD.n2549 0.188
R6803 VDD.n2529 VDD.n2509 0.188
R6804 VDD.n2509 VDD.n2489 0.188
R6805 VDD.n3228 VDD.n3227 0.186
R6806 VDD.n2835 VDD.n2834 0.186
R6807 VDD.n572 VDD.n384 0.185
R6808 VDD.n3196 VDD.n3138 0.185
R6809 VDD.n543 VDD.n540 0.184
R6810 VDD.n2609 VDD.n2589 0.184
R6811 VDD.n2130 VDD.n2129 0.183
R6812 VDD.n2126 VDD.n2125 0.182
R6813 VDD.n3117 VDD.n3116 0.182
R6814 VDD.n3219 VDD.n3218 0.182
R6815 VDD.n3105 VDD.n3104 0.182
R6816 VDD.n2132 VDD.n2131 0.182
R6817 VDD.n2131 VDD.n2130 0.182
R6818 VDD.n2129 VDD.n2128 0.182
R6819 VDD.n2128 VDD.n2127 0.182
R6820 VDD.n2127 VDD.n2126 0.182
R6821 VDD.n1166 VDD.n1157 0.182
R6822 VDD.n1181 VDD.n1172 0.182
R6823 VDD.n1226 VDD.n1217 0.182
R6824 VDD.n1211 VDD.n1202 0.182
R6825 VDD.n1196 VDD.n1187 0.182
R6826 VDD.n1154 VDD.n1145 0.182
R6827 VDD.n1139 VDD.n1130 0.182
R6828 VDD.n1244 VDD.n1235 0.182
R6829 VDD.n2864 VDD.n2863 0.18
R6830 VDD.n2962 VDD.n2961 0.179
R6831 VDD.n2997 VDD.n2996 0.179
R6832 VDD.n3186 VDD.n3185 0.179
R6833 VDD.n3173 VDD.n3172 0.179
R6834 VDD.n3086 VDD.n3085 0.179
R6835 VDD.n3067 VDD.n3066 0.179
R6836 VDD.n189 VDD.n188 0.179
R6837 VDD.n177 VDD.n176 0.179
R6838 VDD.n130 VDD.n129 0.179
R6839 VDD.n118 VDD.n117 0.179
R6840 VDD.n844 VDD.n843 0.179
R6841 VDD.n20 VDD.n19 0.179
R6842 VDD.n79 VDD.n78 0.179
R6843 VDD.n67 VDD.n66 0.179
R6844 VDD.n367 VDD.n366 0.179
R6845 VDD.n349 VDD.n348 0.179
R6846 VDD.n467 VDD.n466 0.179
R6847 VDD.n448 VDD.n447 0.179
R6848 VDD.n479 VDD.n478 0.179
R6849 VDD.n516 VDD.n515 0.179
R6850 VDD.n2766 VDD.n2765 0.179
R6851 VDD.n2800 VDD.n2799 0.179
R6852 VDD.n2702 VDD.n2701 0.179
R6853 VDD.n2737 VDD.n2736 0.179
R6854 VDD.n2933 VDD.n2932 0.179
R6855 VDD.n3445 VDD.n3444 0.177
R6856 VDD.n2888 VDD.n2887 0.177
R6857 VDD.n2855 VDD.n2854 0.176
R6858 VDD.n456 VDD.n449 0.175
R6859 VDD.n524 VDD.n517 0.175
R6860 VDD.n2808 VDD.n2801 0.175
R6861 VDD.n3005 VDD.n2998 0.175
R6862 VDD.n2745 VDD.n2738 0.175
R6863 VDD.n368 VDD.n350 0.175
R6864 VDD.n3075 VDD.n3068 0.174
R6865 VDD.n2824 VDD.n2823 0.174
R6866 VDD.n3314 VDD.n3302 0.174
R6867 VDD.n3371 VDD.n3359 0.174
R6868 VDD.n247 VDD.n235 0.174
R6869 VDD.n190 VDD.n178 0.174
R6870 VDD.n131 VDD.n119 0.174
R6871 VDD.n80 VDD.n68 0.174
R6872 VDD.n556 VDD.n553 0.173
R6873 VDD.n2934 VDD.n2681 0.17
R6874 VDD.n3117 VDD.n3087 0.168
R6875 VDD.n3175 VDD.n3174 0.168
R6876 VDD.n3261 VDD.n3260 0.167
R6877 VDD.n2932 VDD.n2908 0.167
R6878 VDD.n2935 VDD.n2672 0.166
R6879 VDD.n3130 VDD.n3129 0.164
R6880 VDD.n1057 VDD.n1032 0.162
R6881 VDD.n3447 VDD.n858 0.162
R6882 VDD.n3397 VDD.n3396 0.162
R6883 VDD.n2998 VDD.n2986 0.162
R6884 VDD.n3174 VDD.n3162 0.162
R6885 VDD.n3068 VDD.n3056 0.162
R6886 VDD.n449 VDD.n437 0.162
R6887 VDD.n2801 VDD.n2789 0.162
R6888 VDD.n178 VDD.n166 0.161
R6889 VDD.n119 VDD.n107 0.161
R6890 VDD.n68 VDD.n56 0.161
R6891 VDD.n3393 VDD.n3392 0.161
R6892 VDD.n3398 VDD.n3397 0.161
R6893 VDD.n350 VDD.n338 0.161
R6894 VDD.n517 VDD.n505 0.161
R6895 VDD.n2738 VDD.n2726 0.161
R6896 VDD.n3241 VDD.n3240 0.16
R6897 VDD.n3444 VDD.n3443 0.159
R6898 VDD.n3302 VDD.n3301 0.159
R6899 VDD.n3359 VDD.n3358 0.159
R6900 VDD.n235 VDD.n234 0.159
R6901 VDD.n251 VDD.n250 0.158
R6902 VDD.n3390 VDD.n3389 0.158
R6903 VDD.n3394 VDD.n3393 0.158
R6904 VDD.n3446 VDD.n3445 0.158
R6905 VDD.n3228 VDD.n3006 0.155
R6906 VDD.n3444 VDD.n3427 0.15
R6907 VDD.n3445 VDD.n3416 0.15
R6908 VDD.n855 VDD.n845 0.148
R6909 VDD.n796 VDD.n190 0.146
R6910 VDD.n2998 VDD.n2997 0.142
R6911 VDD.n3174 VDD.n3173 0.142
R6912 VDD.n3068 VDD.n3067 0.142
R6913 VDD.n178 VDD.n177 0.142
R6914 VDD.n119 VDD.n118 0.142
R6915 VDD.n845 VDD.n844 0.142
R6916 VDD.n68 VDD.n67 0.142
R6917 VDD.n350 VDD.n349 0.142
R6918 VDD.n449 VDD.n448 0.142
R6919 VDD.n517 VDD.n516 0.142
R6920 VDD.n2801 VDD.n2800 0.142
R6921 VDD.n2738 VDD.n2737 0.142
R6922 VDD.n190 VDD.n189 0.141
R6923 VDD.n131 VDD.n130 0.141
R6924 VDD.n21 VDD.n20 0.141
R6925 VDD.n80 VDD.n79 0.141
R6926 VDD.n3250 VDD.n2935 0.137
R6927 VDD.n740 VDD.n730 0.131
R6928 VDD.n586 VDD.n584 0.129
R6929 VDD.n800 VDD.n131 0.129
R6930 VDD.n815 VDD.n21 0.129
R6931 VDD.n811 VDD.n80 0.129
R6932 VDD.n3396 VDD.n3314 0.129
R6933 VDD.n3392 VDD.n3371 0.128
R6934 VDD.n248 VDD.n247 0.128
R6935 VDD.n381 VDD.n368 0.128
R6936 VDD.n570 VDD.n468 0.128
R6937 VDD.n540 VDD.n525 0.128
R6938 VDD.n2835 VDD.n2809 0.128
R6939 VDD.n2864 VDD.n2746 0.128
R6940 VDD.n3006 VDD.n2962 0.125
R6941 VDD.n3194 VDD.n3186 0.125
R6942 VDD.n468 VDD.n467 0.125
R6943 VDD.n525 VDD.n479 0.125
R6944 VDD.n2809 VDD.n2766 0.125
R6945 VDD.n2746 VDD.n2702 0.125
R6946 VDD.n368 VDD.n367 0.124
R6947 VDD.n3087 VDD.n3086 0.123
R6948 VDD.n1053 VDD.n1052 0.12
R6949 VDD.n928 VDD.n927 0.12
R6950 VDD.n953 VDD.n952 0.12
R6951 VDD.n1028 VDD.n1027 0.12
R6952 VDD.n1003 VDD.n1002 0.12
R6953 VDD.n978 VDD.n977 0.12
R6954 VDD.n903 VDD.n902 0.12
R6955 VDD.n879 VDD.n878 0.12
R6956 VDD.n1872 VDD.n1871 0.12
R6957 VDD.n1847 VDD.n1846 0.12
R6958 VDD.n1547 VDD.n1546 0.12
R6959 VDD.n1572 VDD.n1571 0.12
R6960 VDD.n1672 VDD.n1671 0.12
R6961 VDD.n1647 VDD.n1646 0.12
R6962 VDD.n1622 VDD.n1621 0.12
R6963 VDD.n1597 VDD.n1596 0.12
R6964 VDD.n1522 VDD.n1521 0.12
R6965 VDD.n1498 VDD.n1497 0.12
R6966 VDD.n1397 VDD.n1396 0.12
R6967 VDD.n1372 VDD.n1371 0.12
R6968 VDD.n1273 VDD.n1272 0.12
R6969 VDD.n1297 VDD.n1296 0.12
R6970 VDD.n1322 VDD.n1321 0.12
R6971 VDD.n1347 VDD.n1346 0.12
R6972 VDD.n1422 VDD.n1421 0.12
R6973 VDD.n1447 VDD.n1446 0.12
R6974 VDD.n2608 VDD.n2607 0.12
R6975 VDD.n2469 VDD.n2468 0.12
R6976 VDD.n2488 VDD.n2487 0.12
R6977 VDD.n2548 VDD.n2547 0.12
R6978 VDD.n2568 VDD.n2567 0.12
R6979 VDD.n2588 VDD.n2587 0.12
R6980 VDD.n2528 VDD.n2527 0.12
R6981 VDD.n2508 VDD.n2507 0.12
R6982 VDD.n2260 VDD.n2259 0.12
R6983 VDD.n2279 VDD.n2278 0.12
R6984 VDD.n2319 VDD.n2318 0.12
R6985 VDD.n2299 VDD.n2298 0.12
R6986 VDD.n644 VDD.n641 0.118
R6987 VDD.n662 VDD.n659 0.118
R6988 VDD.n680 VDD.n677 0.118
R6989 VDD.n697 VDD.n694 0.118
R6990 VDD.n626 VDD.n623 0.118
R6991 VDD.n757 VDD.n754 0.118
R6992 VDD.n775 VDD.n772 0.118
R6993 VDD.n793 VDD.n790 0.118
R6994 VDD.n3250 VDD.n3249 0.117
R6995 VDD.n414 VDD.n402 0.114
R6996 VDD.n587 VDD.n586 0.113
R6997 VDD.n415 VDD.n393 0.113
R6998 VDD VDD.n858 0.107
R6999 VDD.n2933 VDD.n2899 0.105
R7000 VDD.n628 VDD.n610 0.104
R7001 VDD.n2644 VDD.n1678 0.104
R7002 VDD.n796 VDD.n795 0.103
R7003 VDD.n2641 VDD.n2640 0.102
R7004 VDD.n2638 VDD.n2637 0.102
R7005 VDD.n383 VDD.n311 0.1
R7006 VDD.n384 VDD.n302 0.1
R7007 VDD.n3447 VDD.n3446 0.098
R7008 VDD.n2847 VDD.n2837 0.098
R7009 VDD.n3216 VDD.n3203 0.098
R7010 VDD.n371 VDD.n370 0.097
R7011 VDD.n3127 VDD.n3126 0.097
R7012 VDD.n3120 VDD.n3119 0.097
R7013 VDD.n3199 VDD.n3198 0.097
R7014 VDD.n3232 VDD.n3231 0.095
R7015 VDD.n1051 VDD.n1046 0.095
R7016 VDD.n926 VDD.n921 0.095
R7017 VDD.n951 VDD.n946 0.095
R7018 VDD.n1026 VDD.n1021 0.095
R7019 VDD.n1001 VDD.n996 0.095
R7020 VDD.n976 VDD.n971 0.095
R7021 VDD.n901 VDD.n896 0.095
R7022 VDD.n877 VDD.n872 0.095
R7023 VDD.n635 VDD.n631 0.095
R7024 VDD.n653 VDD.n649 0.095
R7025 VDD.n671 VDD.n667 0.095
R7026 VDD.n688 VDD.n684 0.095
R7027 VDD.n617 VDD.n613 0.095
R7028 VDD.n748 VDD.n744 0.095
R7029 VDD.n766 VDD.n762 0.095
R7030 VDD.n784 VDD.n780 0.095
R7031 VDD.n1740 VDD.n1736 0.095
R7032 VDD.n1765 VDD.n1761 0.095
R7033 VDD.n1870 VDD.n1866 0.095
R7034 VDD.n1845 VDD.n1841 0.095
R7035 VDD.n1815 VDD.n1811 0.095
R7036 VDD.n1790 VDD.n1786 0.095
R7037 VDD.n1715 VDD.n1711 0.095
R7038 VDD.n1691 VDD.n1687 0.095
R7039 VDD.n1545 VDD.n1541 0.095
R7040 VDD.n1570 VDD.n1566 0.095
R7041 VDD.n1670 VDD.n1666 0.095
R7042 VDD.n1645 VDD.n1641 0.095
R7043 VDD.n1620 VDD.n1616 0.095
R7044 VDD.n1595 VDD.n1591 0.095
R7045 VDD.n1520 VDD.n1516 0.095
R7046 VDD.n1496 VDD.n1492 0.095
R7047 VDD.n1395 VDD.n1391 0.095
R7048 VDD.n1370 VDD.n1366 0.095
R7049 VDD.n1271 VDD.n1267 0.095
R7050 VDD.n1295 VDD.n1291 0.095
R7051 VDD.n1320 VDD.n1316 0.095
R7052 VDD.n1345 VDD.n1341 0.095
R7053 VDD.n1420 VDD.n1416 0.095
R7054 VDD.n1445 VDD.n1441 0.095
R7055 VDD.n2601 VDD.n2597 0.095
R7056 VDD.n2462 VDD.n2458 0.095
R7057 VDD.n2481 VDD.n2477 0.095
R7058 VDD.n2541 VDD.n2537 0.095
R7059 VDD.n2561 VDD.n2557 0.095
R7060 VDD.n2581 VDD.n2577 0.095
R7061 VDD.n2521 VDD.n2517 0.095
R7062 VDD.n2501 VDD.n2497 0.095
R7063 VDD.n2397 VDD.n2393 0.095
R7064 VDD.n2253 VDD.n2249 0.095
R7065 VDD.n2272 VDD.n2268 0.095
R7066 VDD.n2337 VDD.n2333 0.095
R7067 VDD.n2357 VDD.n2353 0.095
R7068 VDD.n2377 VDD.n2373 0.095
R7069 VDD.n2312 VDD.n2308 0.095
R7070 VDD.n2292 VDD.n2288 0.095
R7071 VDD.n2884 VDD.n2883 0.093
R7072 VDD.n3448 VDD.n3447 0.088
R7073 VDD.n3202 VDD.n3201 0.085
R7074 VDD VDD.n1057 0.084
R7075 VDD.n1747 VDD.n1746 0.083
R7076 VDD.n1772 VDD.n1771 0.083
R7077 VDD.n1822 VDD.n1821 0.083
R7078 VDD.n1797 VDD.n1796 0.083
R7079 VDD.n1722 VDD.n1721 0.083
R7080 VDD.n1698 VDD.n1697 0.083
R7081 VDD.n2399 VDD.n2398 0.083
R7082 VDD.n2339 VDD.n2338 0.083
R7083 VDD.n2359 VDD.n2358 0.083
R7084 VDD.n2379 VDD.n2378 0.083
R7085 VDD.n2879 VDD.n2878 0.082
R7086 VDD.n2850 VDD.n2849 0.082
R7087 VDD.n563 VDD.n562 0.081
R7088 VDD.n2125 VDD.n2124 0.079
R7089 VDD.n2119 VDD.n2118 0.079
R7090 VDD.n2113 VDD.n2112 0.079
R7091 VDD.n2107 VDD.n2106 0.079
R7092 VDD.n2101 VDD.n2100 0.079
R7093 VDD.n2095 VDD.n2094 0.079
R7094 VDD.n2089 VDD.n2088 0.079
R7095 VDD.n2083 VDD.n2082 0.079
R7096 VDD.n3123 VDD.n3122 0.077
R7097 VDD.n3236 VDD.n3235 0.076
R7098 VDD.n3404 VDD.n3398 0.075
R7099 VDD.n551 VDD.n550 0.075
R7100 VDD.n426 VDD.n425 0.075
R7101 VDD.n487 VDD.n486 0.075
R7102 VDD.n2777 VDD.n2776 0.075
R7103 VDD.n2710 VDD.n2709 0.075
R7104 VDD.n250 VDD.n249 0.073
R7105 VDD.n3391 VDD.n3390 0.073
R7106 VDD.n3395 VDD.n3394 0.073
R7107 VDD.n2640 VDD.n2639 0.072
R7108 VDD.n857 VDD.n856 0.07
R7109 VDD.n855 VDD.n854 0.067
R7110 VDD.n1157 VDD.n1155 0.065
R7111 VDD.n1172 VDD.n1170 0.065
R7112 VDD.n1217 VDD.n1215 0.065
R7113 VDD.n1202 VDD.n1200 0.065
R7114 VDD.n1187 VDD.n1185 0.065
R7115 VDD.n1145 VDD.n1143 0.065
R7116 VDD.n1130 VDD.n1128 0.065
R7117 VDD.n1235 VDD.n1233 0.065
R7118 VDD.n800 VDD.n799 0.064
R7119 VDD.n825 VDD.n817 0.064
R7120 VDD.n815 VDD.n814 0.063
R7121 VDD.n810 VDD.n802 0.063
R7122 VDD.n814 VDD.n813 0.063
R7123 VDD.n799 VDD.n798 0.063
R7124 VDD.n858 VDD.n857 0.062
R7125 VDD.n3302 VDD.n3285 0.062
R7126 VDD.n3314 VDD.n3313 0.062
R7127 VDD.n3359 VDD.n3342 0.062
R7128 VDD.n3371 VDD.n3370 0.062
R7129 VDD.n235 VDD.n218 0.062
R7130 VDD.n247 VDD.n246 0.062
R7131 VDD.n698 VDD.n681 0.062
R7132 VDD.n681 VDD.n275 0.061
R7133 VDD.n811 VDD.n810 0.061
R7134 VDD.n759 VDD.n758 0.06
R7135 VDD.n2155 VDD.n2154 0.059
R7136 VDD.n2623 VDD.n2622 0.059
R7137 VDD.n797 VDD.n796 0.058
R7138 VDD.n383 VDD.n382 0.057
R7139 VDD.n2637 VDD.n2636 0.057
R7140 VDD.n646 VDD.n645 0.056
R7141 VDD.n275 VDD.n274 0.055
R7142 VDD.n3260 VDD.n3259 0.054
R7143 VDD.n2919 VDD.n2916 0.054
R7144 VDD.n412 VDD.n410 0.054
R7145 VDD.n2929 VDD.n2927 0.054
R7146 VDD.n285 VDD.n284 0.054
R7147 VDD.n274 VDD.n273 0.054
R7148 VDD.n741 VDD.n740 0.054
R7149 VDD.n1251 VDD.n1083 0.054
R7150 VDD.n1250 VDD.n1091 0.054
R7151 VDD.n1246 VDD.n1124 0.054
R7152 VDD.n1247 VDD.n1116 0.054
R7153 VDD.n1248 VDD.n1107 0.054
R7154 VDD.n1249 VDD.n1099 0.054
R7155 VDD.n1252 VDD.n1074 0.054
R7156 VDD.n1253 VDD.n1066 0.054
R7157 VDD.n717 VDD.n716 0.053
R7158 VDD.n610 VDD.n609 0.053
R7159 VDD.n573 VDD.n572 0.051
R7160 VDD.n758 VDD.n741 0.049
R7161 VDD.n571 VDD.n570 0.048
R7162 VDD.n2712 VDD.n2710 0.047
R7163 VDD.n646 VDD.n587 0.046
R7164 VDD.n489 VDD.n487 0.045
R7165 VDD.n552 VDD.n551 0.045
R7166 VDD.n2779 VDD.n2777 0.045
R7167 VDD.n428 VDD.n426 0.044
R7168 VDD.n382 VDD.n381 0.044
R7169 VDD.n2636 VDD.n2635 0.044
R7170 VDD.n336 VDD.n335 0.043
R7171 VDD.n503 VDD.n502 0.042
R7172 VDD.n3114 VDD.n3106 0.042
R7173 VDD.n2885 VDD.n2880 0.042
R7174 VDD.n2642 VDD.n2641 0.042
R7175 VDD.n3233 VDD.n3230 0.042
R7176 VDD.n2897 VDD.n2889 0.041
R7177 VDD.n537 VDD.n536 0.041
R7178 VDD.n3448 VDD.n3262 0.041
R7179 VDD.n1054 VDD.n1033 0.04
R7180 VDD.n929 VDD.n908 0.04
R7181 VDD.n954 VDD.n933 0.04
R7182 VDD.n1029 VDD.n1008 0.04
R7183 VDD.n1004 VDD.n983 0.04
R7184 VDD.n979 VDD.n958 0.04
R7185 VDD.n904 VDD.n883 0.04
R7186 VDD.n880 VDD.n859 0.04
R7187 VDD.n2876 VDD.n2875 0.04
R7188 VDD.n2832 VDD.n2830 0.04
R7189 VDD.n1749 VDD.n1728 0.04
R7190 VDD.n1774 VDD.n1753 0.04
R7191 VDD.n1874 VDD.n1853 0.04
R7192 VDD.n1849 VDD.n1828 0.04
R7193 VDD.n1824 VDD.n1803 0.04
R7194 VDD.n1799 VDD.n1778 0.04
R7195 VDD.n1724 VDD.n1703 0.04
R7196 VDD.n1700 VDD.n1679 0.04
R7197 VDD.n1549 VDD.n1528 0.04
R7198 VDD.n1574 VDD.n1553 0.04
R7199 VDD.n1674 VDD.n1653 0.04
R7200 VDD.n1649 VDD.n1628 0.04
R7201 VDD.n1624 VDD.n1603 0.04
R7202 VDD.n1599 VDD.n1578 0.04
R7203 VDD.n1524 VDD.n1503 0.04
R7204 VDD.n1500 VDD.n1479 0.04
R7205 VDD.n1399 VDD.n1378 0.04
R7206 VDD.n1374 VDD.n1353 0.04
R7207 VDD.n1275 VDD.n1254 0.04
R7208 VDD.n1299 VDD.n1278 0.04
R7209 VDD.n1324 VDD.n1303 0.04
R7210 VDD.n1349 VDD.n1328 0.04
R7211 VDD.n1424 VDD.n1403 0.04
R7212 VDD.n1449 VDD.n1428 0.04
R7213 VDD.n740 VDD.n739 0.039
R7214 VDD.n777 VDD.n776 0.037
R7215 VDD.n587 VDD.n285 0.037
R7216 VDD.n794 VDD.n777 0.036
R7217 VDD.n681 VDD.n664 0.034
R7218 VDD.n572 VDD.n571 0.032
R7219 VDD.n798 VDD.n797 0.031
R7220 VDD.n813 VDD.n812 0.031
R7221 VDD.n817 VDD.n816 0.031
R7222 VDD.n802 VDD.n801 0.031
R7223 VDD.n730 VDD.n728 0.03
R7224 VDD.n600 VDD.n598 0.03
R7225 VDD.n264 VDD.n262 0.03
R7226 VDD.n645 VDD.n628 0.03
R7227 VDD.n334 VDD.n332 0.03
R7228 VDD.n501 VDD.n500 0.03
R7229 VDD.n2189 VDD.n2188 0.03
R7230 VDD.n2143 VDD.n2142 0.03
R7231 VDD.n1476 VDD.n1475 0.03
R7232 VDD.n2036 VDD.n2028 0.03
R7233 VDD.n1936 VDD.n1928 0.03
R7234 VDD.n1886 VDD.n1878 0.03
R7235 VDD.n1911 VDD.n1903 0.03
R7236 VDD.n1961 VDD.n1953 0.03
R7237 VDD.n1986 VDD.n1978 0.03
R7238 VDD.n2011 VDD.n2003 0.03
R7239 VDD.n2061 VDD.n2053 0.03
R7240 VDD.n2611 VDD.n2610 0.03
R7241 VDD.n2448 VDD.n2447 0.03
R7242 VDD.n2423 VDD.n2422 0.03
R7243 VDD.n2239 VDD.n2238 0.03
R7244 VDD.n2214 VDD.n2213 0.03
R7245 VDD.n2639 VDD.n2638 0.03
R7246 VDD.n570 VDD.n569 0.027
R7247 VDD.n2836 VDD.n2835 0.026
R7248 VDD.n2865 VDD.n2864 0.026
R7249 VDD.n664 VDD.n663 0.026
R7250 VDD.n381 VDD.n380 0.025
R7251 VDD.n540 VDD.n539 0.025
R7252 VDD.n3449 VDD.n2645 0.025
R7253 VDD.n543 VDD.n542 0.023
R7254 VDD.n2165 VDD.n2156 0.023
R7255 VDD.n2633 VDD.n2624 0.023
R7256 VDD.n249 VDD.n248 0.023
R7257 VDD.n3392 VDD.n3391 0.023
R7258 VDD.n3396 VDD.n3395 0.023
R7259 VDD.n3229 VDD.n3228 0.022
R7260 VDD.n2643 VDD.n2642 0.022
R7261 VDD.n3118 VDD.n3117 0.022
R7262 VDD.n380 VDD.n379 0.021
R7263 VDD.n3112 VDD.n3111 0.021
R7264 VDD.n2187 VDD.n2186 0.021
R7265 VDD.n2179 VDD.n2172 0.021
R7266 VDD.n1474 VDD.n1473 0.021
R7267 VDD.n1466 VDD.n1459 0.021
R7268 VDD.n2050 VDD.n2049 0.021
R7269 VDD.n2035 VDD.n2034 0.021
R7270 VDD.n1950 VDD.n1949 0.021
R7271 VDD.n1935 VDD.n1934 0.021
R7272 VDD.n1900 VDD.n1899 0.021
R7273 VDD.n1885 VDD.n1884 0.021
R7274 VDD.n1925 VDD.n1924 0.021
R7275 VDD.n1910 VDD.n1909 0.021
R7276 VDD.n1975 VDD.n1974 0.021
R7277 VDD.n1960 VDD.n1959 0.021
R7278 VDD.n2000 VDD.n1999 0.021
R7279 VDD.n1985 VDD.n1984 0.021
R7280 VDD.n2025 VDD.n2024 0.021
R7281 VDD.n2010 VDD.n2009 0.021
R7282 VDD.n2075 VDD.n2074 0.021
R7283 VDD.n2060 VDD.n2059 0.021
R7284 VDD.n2446 VDD.n2445 0.021
R7285 VDD.n2438 VDD.n2431 0.021
R7286 VDD.n2421 VDD.n2420 0.021
R7287 VDD.n2413 VDD.n2406 0.021
R7288 VDD.n2237 VDD.n2236 0.021
R7289 VDD.n2229 VDD.n2222 0.021
R7290 VDD.n2212 VDD.n2211 0.021
R7291 VDD.n2204 VDD.n2197 0.021
R7292 VDD.t3388 VDD.n2084 0.021
R7293 VDD.t4027 VDD.n2090 0.021
R7294 VDD.t3761 VDD.n2120 0.021
R7295 VDD.t3021 VDD.n2114 0.021
R7296 VDD.t3448 VDD.n2108 0.021
R7297 VDD.t1992 VDD.n2102 0.021
R7298 VDD.t4404 VDD.n2096 0.021
R7299 VDD.t2331 VDD.n2078 0.021
R7300 VDD.n2850 VDD.n2755 0.02
R7301 VDD.n2819 VDD.n2818 0.02
R7302 VDD.n3197 VDD.n3016 0.02
R7303 VDD.n3123 VDD.n3026 0.02
R7304 VDD.n3118 VDD.n3033 0.02
R7305 VDD.n3098 VDD.n3097 0.02
R7306 VDD.n3229 VDD.n2951 0.02
R7307 VDD.n2879 VDD.n2691 0.02
R7308 VDD.n2895 VDD.n2894 0.02
R7309 VDD.n2829 VDD.n2828 0.02
R7310 VDD.n3136 VDD.n3135 0.02
R7311 VDD.n2984 VDD.n2983 0.02
R7312 VDD.n3147 VDD.n3146 0.02
R7313 VDD.n435 VDD.n434 0.02
R7314 VDD.n2786 VDD.n2785 0.02
R7315 VDD.n3246 VDD.n3245 0.019
R7316 VDD.n2860 VDD.n2859 0.019
R7317 VDD.n3224 VDD.n3223 0.019
R7318 VDD.n2975 VDD.n2974 0.019
R7319 VDD.n3159 VDD.n3158 0.019
R7320 VDD.n3053 VDD.n3052 0.019
R7321 VDD.n3041 VDD.n3040 0.019
R7322 VDD.n795 VDD.n794 0.019
R7323 VDD.n741 VDD.n698 0.019
R7324 VDD.n316 VDD.n315 0.019
R7325 VDD.n3236 VDD.n2944 0.019
R7326 VDD.n328 VDD.n327 0.018
R7327 VDD.n495 VDD.n494 0.018
R7328 VDD.n2724 VDD.n2723 0.018
R7329 VDD.n3450 VDD.n3449 0.017
R7330 VDD.n3197 VDD.n3196 0.016
R7331 VDD.n2156 VDD.n2155 0.015
R7332 VDD.n2624 VDD.n2623 0.015
R7333 VDD.n776 VDD.n759 0.013
R7334 VDD.n2644 VDD.n2643 0.013
R7335 VDD.n856 VDD.n855 0.013
R7336 VDD.n857 VDD.n825 0.013
R7337 VDD.n3446 VDD.n3405 0.012
R7338 VDD.n3248 VDD.n3246 0.011
R7339 VDD.n2872 VDD.n2871 0.011
R7340 VDD.n2845 VDD.n2844 0.011
R7341 VDD.n2862 VDD.n2860 0.011
R7342 VDD.n533 VDD.n532 0.011
R7343 VDD.n3137 VDD.n3136 0.011
R7344 VDD.n3211 VDD.n3210 0.011
R7345 VDD.n3226 VDD.n3224 0.011
R7346 VDD.n2976 VDD.n2975 0.011
R7347 VDD.n3161 VDD.n3159 0.011
R7348 VDD.n3055 VDD.n3053 0.011
R7349 VDD.n3046 VDD.n3041 0.011
R7350 VDD.n3397 VDD.n3271 0.011
R7351 VDD.n3393 VDD.n3328 0.011
R7352 VDD.n3389 VDD.n3385 0.011
R7353 VDD.n251 VDD.n194 0.011
R7354 VDD.n853 VDD.n849 0.011
R7355 VDD.n833 VDD.n829 0.011
R7356 VDD.n29 VDD.n25 0.011
R7357 VDD.n825 VDD.n824 0.011
R7358 VDD.n810 VDD.n806 0.011
R7359 VDD.n139 VDD.n135 0.011
R7360 VDD.n165 VDD.n161 0.011
R7361 VDD.n157 VDD.n153 0.011
R7362 VDD.n106 VDD.n102 0.011
R7363 VDD.n98 VDD.n94 0.011
R7364 VDD.n55 VDD.n51 0.011
R7365 VDD.n47 VDD.n43 0.011
R7366 VDD.n3443 VDD.n3431 0.011
R7367 VDD.n3442 VDD.n3441 0.011
R7368 VDD.n3301 VDD.n3289 0.011
R7369 VDD.n3300 VDD.n3299 0.011
R7370 VDD.n3358 VDD.n3346 0.011
R7371 VDD.n3357 VDD.n3356 0.011
R7372 VDD.n234 VDD.n222 0.011
R7373 VDD.n233 VDD.n232 0.011
R7374 VDD.n337 VDD.n328 0.011
R7375 VDD.n321 VDD.n316 0.011
R7376 VDD.n436 VDD.n435 0.011
R7377 VDD.n504 VDD.n495 0.011
R7378 VDD.n2725 VDD.n2724 0.011
R7379 VDD.n2934 VDD.n2933 0.011
R7380 VDD.n854 VDD.n853 0.011
R7381 VDD.n2985 VDD.n2984 0.01
R7382 VDD.n3148 VDD.n3147 0.01
R7383 VDD.n2787 VDD.n2786 0.01
R7384 VDD.n2885 VDD.n2884 0.009
R7385 VDD.n2896 VDD.n2895 0.009
R7386 VDD.n2832 VDD.n2829 0.009
R7387 VDD.n801 VDD.n800 0.009
R7388 VDD.n812 VDD.n811 0.009
R7389 VDD.n816 VDD.n815 0.009
R7390 VDD.n3261 VDD.n3250 0.009
R7391 VDD.n3113 VDD.n3112 0.008
R7392 VDD.n2645 VDD.n2644 0.008
R7393 VDD.n3405 VDD.n3404 0.007
R7394 VDD.n2846 VDD.n2845 0.007
R7395 VDD.n2877 VDD.n2874 0.007
R7396 VDD.n2609 VDD.n2608 0.007
R7397 VDD.n2489 VDD.n2488 0.007
R7398 VDD.n2549 VDD.n2548 0.007
R7399 VDD.n2569 VDD.n2568 0.007
R7400 VDD.n2589 VDD.n2588 0.007
R7401 VDD.n2529 VDD.n2528 0.007
R7402 VDD.n2509 VDD.n2508 0.007
R7403 VDD.n2400 VDD.n2399 0.007
R7404 VDD.n2280 VDD.n2279 0.007
R7405 VDD.n2340 VDD.n2339 0.007
R7406 VDD.n2360 VDD.n2359 0.007
R7407 VDD.n2380 VDD.n2379 0.007
R7408 VDD.n2320 VDD.n2319 0.007
R7409 VDD.n2300 VDD.n2299 0.007
R7410 VDD.n1230 VDD.n1166 0.006
R7411 VDD.n3195 VDD.n3175 0.006
R7412 VDD.n3212 VDD.n3211 0.005
R7413 VDD.n535 VDD.n533 0.005
R7414 VDD.n3233 VDD.n3232 0.005
R7415 VDD.n2643 VDD.n2166 0.005
R7416 VDD.n2635 VDD.n2634 0.005
R7417 VDD.n1245 VDD.n1244 0.004
R7418 VDD.n663 VDD.n646 0.004
R7419 VDD.n3114 VDD.n3113 0.003
R7420 VDD.n1056 VDD.n1055 0.003
R7421 VDD.n931 VDD.n930 0.003
R7422 VDD.n956 VDD.n955 0.003
R7423 VDD.n1031 VDD.n1030 0.003
R7424 VDD.n1006 VDD.n1005 0.003
R7425 VDD.n981 VDD.n980 0.003
R7426 VDD.n906 VDD.n905 0.003
R7427 VDD.n882 VDD.n881 0.003
R7428 VDD.n1751 VDD.n1750 0.003
R7429 VDD.n1776 VDD.n1775 0.003
R7430 VDD.n1876 VDD.n1875 0.003
R7431 VDD.n1851 VDD.n1850 0.003
R7432 VDD.n1826 VDD.n1825 0.003
R7433 VDD.n1801 VDD.n1800 0.003
R7434 VDD.n1726 VDD.n1725 0.003
R7435 VDD.n1702 VDD.n1701 0.003
R7436 VDD.n1551 VDD.n1550 0.003
R7437 VDD.n1576 VDD.n1575 0.003
R7438 VDD.n1676 VDD.n1675 0.003
R7439 VDD.n1651 VDD.n1650 0.003
R7440 VDD.n1626 VDD.n1625 0.003
R7441 VDD.n1601 VDD.n1600 0.003
R7442 VDD.n1526 VDD.n1525 0.003
R7443 VDD.n1502 VDD.n1501 0.003
R7444 VDD.n1401 VDD.n1400 0.003
R7445 VDD.n1376 VDD.n1375 0.003
R7446 VDD.n1277 VDD.n1276 0.003
R7447 VDD.n1301 VDD.n1300 0.003
R7448 VDD.n1326 VDD.n1325 0.003
R7449 VDD.n1351 VDD.n1350 0.003
R7450 VDD.n1426 VDD.n1425 0.003
R7451 VDD.n1451 VDD.n1450 0.003
R7452 VDD.n645 VDD.n644 0.003
R7453 VDD.n663 VDD.n662 0.003
R7454 VDD.n681 VDD.n680 0.003
R7455 VDD.n698 VDD.n697 0.003
R7456 VDD.n758 VDD.n757 0.003
R7457 VDD.n776 VDD.n775 0.003
R7458 VDD.n794 VDD.n793 0.003
R7459 VDD.n538 VDD.n535 0.003
R7460 VDD.n2877 VDD.n2876 0.003
R7461 VDD.n1229 VDD.n1181 0.003
R7462 VDD.n1227 VDD.n1211 0.003
R7463 VDD.n1231 VDD.n1154 0.003
R7464 VDD.n1232 VDD.n1139 0.003
R7465 VDD.n1048 VDD.n1046 0.003
R7466 VDD.n923 VDD.n921 0.003
R7467 VDD.n948 VDD.n946 0.003
R7468 VDD.n1023 VDD.n1021 0.003
R7469 VDD.n998 VDD.n996 0.003
R7470 VDD.n973 VDD.n971 0.003
R7471 VDD.n898 VDD.n896 0.003
R7472 VDD.n874 VDD.n872 0.003
R7473 VDD.n631 VDD.n630 0.003
R7474 VDD.n649 VDD.n648 0.003
R7475 VDD.n667 VDD.n666 0.003
R7476 VDD.n684 VDD.n683 0.003
R7477 VDD.n613 VDD.n612 0.003
R7478 VDD.n744 VDD.n743 0.003
R7479 VDD.n762 VDD.n761 0.003
R7480 VDD.n780 VDD.n779 0.003
R7481 VDD.n1736 VDD.n1735 0.003
R7482 VDD.n1761 VDD.n1760 0.003
R7483 VDD.n1866 VDD.n1865 0.003
R7484 VDD.n1841 VDD.n1840 0.003
R7485 VDD.n1811 VDD.n1810 0.003
R7486 VDD.n1786 VDD.n1785 0.003
R7487 VDD.n1711 VDD.n1710 0.003
R7488 VDD.n1687 VDD.n1686 0.003
R7489 VDD.n1541 VDD.n1540 0.003
R7490 VDD.n1566 VDD.n1565 0.003
R7491 VDD.n1666 VDD.n1665 0.003
R7492 VDD.n1641 VDD.n1640 0.003
R7493 VDD.n1616 VDD.n1615 0.003
R7494 VDD.n1591 VDD.n1590 0.003
R7495 VDD.n1516 VDD.n1515 0.003
R7496 VDD.n1492 VDD.n1491 0.003
R7497 VDD.n1391 VDD.n1390 0.003
R7498 VDD.n1366 VDD.n1365 0.003
R7499 VDD.n1267 VDD.n1266 0.003
R7500 VDD.n1291 VDD.n1290 0.003
R7501 VDD.n1316 VDD.n1315 0.003
R7502 VDD.n1341 VDD.n1340 0.003
R7503 VDD.n1416 VDD.n1415 0.003
R7504 VDD.n1441 VDD.n1440 0.003
R7505 VDD.n2597 VDD.n2596 0.003
R7506 VDD.n2458 VDD.n2457 0.003
R7507 VDD.n2477 VDD.n2476 0.003
R7508 VDD.n2537 VDD.n2536 0.003
R7509 VDD.n2557 VDD.n2556 0.003
R7510 VDD.n2577 VDD.n2576 0.003
R7511 VDD.n2517 VDD.n2516 0.003
R7512 VDD.n2497 VDD.n2496 0.003
R7513 VDD.n2393 VDD.n2392 0.003
R7514 VDD.n2249 VDD.n2248 0.003
R7515 VDD.n2268 VDD.n2267 0.003
R7516 VDD.n2333 VDD.n2332 0.003
R7517 VDD.n2353 VDD.n2352 0.003
R7518 VDD.n2373 VDD.n2372 0.003
R7519 VDD.n2308 VDD.n2307 0.003
R7520 VDD.n2288 VDD.n2287 0.003
R7521 VDD.n1034 VDD.n1033 0.003
R7522 VDD.n909 VDD.n908 0.003
R7523 VDD.n934 VDD.n933 0.003
R7524 VDD.n1009 VDD.n1008 0.003
R7525 VDD.n984 VDD.n983 0.003
R7526 VDD.n959 VDD.n958 0.003
R7527 VDD.n884 VDD.n883 0.003
R7528 VDD.n860 VDD.n859 0.003
R7529 VDD.n1749 VDD.n1748 0.003
R7530 VDD.n1774 VDD.n1773 0.003
R7531 VDD.n1874 VDD.n1873 0.003
R7532 VDD.n1849 VDD.n1848 0.003
R7533 VDD.n1824 VDD.n1823 0.003
R7534 VDD.n1799 VDD.n1798 0.003
R7535 VDD.n1724 VDD.n1723 0.003
R7536 VDD.n1700 VDD.n1699 0.003
R7537 VDD.n1549 VDD.n1548 0.003
R7538 VDD.n1574 VDD.n1573 0.003
R7539 VDD.n1674 VDD.n1673 0.003
R7540 VDD.n1649 VDD.n1648 0.003
R7541 VDD.n1624 VDD.n1623 0.003
R7542 VDD.n1599 VDD.n1598 0.003
R7543 VDD.n1524 VDD.n1523 0.003
R7544 VDD.n1500 VDD.n1499 0.003
R7545 VDD.n1399 VDD.n1398 0.003
R7546 VDD.n1374 VDD.n1373 0.003
R7547 VDD.n1275 VDD.n1274 0.003
R7548 VDD.n1299 VDD.n1298 0.003
R7549 VDD.n1324 VDD.n1323 0.003
R7550 VDD.n1349 VDD.n1348 0.003
R7551 VDD.n1424 VDD.n1423 0.003
R7552 VDD.n1449 VDD.n1448 0.003
R7553 VDD.n2050 VDD.n2043 0.002
R7554 VDD.n1950 VDD.n1943 0.002
R7555 VDD.n1900 VDD.n1893 0.002
R7556 VDD.n1925 VDD.n1918 0.002
R7557 VDD.n1975 VDD.n1968 0.002
R7558 VDD.n2000 VDD.n1993 0.002
R7559 VDD.n2025 VDD.n2018 0.002
R7560 VDD.n2075 VDD.n2068 0.002
R7561 VDD.n1056 VDD.n1033 0.002
R7562 VDD.n931 VDD.n908 0.002
R7563 VDD.n956 VDD.n933 0.002
R7564 VDD.n1031 VDD.n1008 0.002
R7565 VDD.n1006 VDD.n983 0.002
R7566 VDD.n981 VDD.n958 0.002
R7567 VDD.n906 VDD.n883 0.002
R7568 VDD.n882 VDD.n859 0.002
R7569 VDD.n1751 VDD.n1749 0.002
R7570 VDD.n1776 VDD.n1774 0.002
R7571 VDD.n1876 VDD.n1874 0.002
R7572 VDD.n1851 VDD.n1849 0.002
R7573 VDD.n1826 VDD.n1824 0.002
R7574 VDD.n1801 VDD.n1799 0.002
R7575 VDD.n1726 VDD.n1724 0.002
R7576 VDD.n1702 VDD.n1700 0.002
R7577 VDD.n1551 VDD.n1549 0.002
R7578 VDD.n1576 VDD.n1574 0.002
R7579 VDD.n1676 VDD.n1674 0.002
R7580 VDD.n1651 VDD.n1649 0.002
R7581 VDD.n1626 VDD.n1624 0.002
R7582 VDD.n1601 VDD.n1599 0.002
R7583 VDD.n1526 VDD.n1524 0.002
R7584 VDD.n1502 VDD.n1500 0.002
R7585 VDD.n1401 VDD.n1399 0.002
R7586 VDD.n1376 VDD.n1374 0.002
R7587 VDD.n1277 VDD.n1275 0.002
R7588 VDD.n1301 VDD.n1299 0.002
R7589 VDD.n1326 VDD.n1324 0.002
R7590 VDD.n1351 VDD.n1349 0.002
R7591 VDD.n1426 VDD.n1424 0.002
R7592 VDD.n1451 VDD.n1449 0.002
R7593 VDD.n1055 VDD.n1034 0.002
R7594 VDD.n930 VDD.n909 0.002
R7595 VDD.n955 VDD.n934 0.002
R7596 VDD.n1030 VDD.n1009 0.002
R7597 VDD.n1005 VDD.n984 0.002
R7598 VDD.n980 VDD.n959 0.002
R7599 VDD.n905 VDD.n884 0.002
R7600 VDD.n881 VDD.n860 0.002
R7601 VDD.n2190 VDD.n2189 0.002
R7602 VDD.n1477 VDD.n1476 0.002
R7603 VDD.n2051 VDD.n2036 0.002
R7604 VDD.n1951 VDD.n1936 0.002
R7605 VDD.n1901 VDD.n1886 0.002
R7606 VDD.n1926 VDD.n1911 0.002
R7607 VDD.n1976 VDD.n1961 0.002
R7608 VDD.n2001 VDD.n1986 0.002
R7609 VDD.n2026 VDD.n2011 0.002
R7610 VDD.n2076 VDD.n2061 0.002
R7611 VDD.n2449 VDD.n2448 0.002
R7612 VDD.n2424 VDD.n2423 0.002
R7613 VDD.n2240 VDD.n2239 0.002
R7614 VDD.n2215 VDD.n2214 0.002
R7615 VDD.n2051 VDD.n2050 0.002
R7616 VDD.n1951 VDD.n1950 0.002
R7617 VDD.n1901 VDD.n1900 0.002
R7618 VDD.n1926 VDD.n1925 0.002
R7619 VDD.n1976 VDD.n1975 0.002
R7620 VDD.n2001 VDD.n2000 0.002
R7621 VDD.n2026 VDD.n2025 0.002
R7622 VDD.n2076 VDD.n2075 0.002
R7623 VDD.n1228 VDD.n1196 0.002
R7624 VDD.n336 VDD.n334 0.002
R7625 VDD.n2725 VDD.n2719 0.002
R7626 VDD.n2191 VDD.n2190 0.002
R7627 VDD.n1478 VDD.n1477 0.002
R7628 VDD.n2450 VDD.n2449 0.002
R7629 VDD.n2425 VDD.n2424 0.002
R7630 VDD.n2241 VDD.n2240 0.002
R7631 VDD.n2216 VDD.n2215 0.002
R7632 VDD.n2976 VDD.n2970 0.002
R7633 VDD.n2166 VDD.n2143 0.002
R7634 VDD.n2634 VDD.n2611 0.002
R7635 VDD.n2847 VDD.n2846 0.001
R7636 VDD.n2187 VDD.n2180 0.001
R7637 VDD.n1474 VDD.n1467 0.001
R7638 VDD.n2446 VDD.n2439 0.001
R7639 VDD.n2421 VDD.n2414 0.001
R7640 VDD.n2237 VDD.n2230 0.001
R7641 VDD.n2212 VDD.n2205 0.001
R7642 VDD.n2897 VDD.n2896 0.001
R7643 VDD.n503 VDD.n501 0.001
R7644 VDD.n2164 VDD.n2163 0.001
R7645 VDD.n2632 VDD.n2631 0.001
R7646 VDD.n3195 VDD.n3194 0.001
R7647 VDD.n2874 VDD.n2872 0.001
R7648 VDD.n3216 VDD.n3215 0.001
R7649 VDD.n2166 VDD.n2165 0.001
R7650 VDD.n2634 VDD.n2633 0.001
R7651 VDD.n3234 VDD.n3233 0.001
R7652 VDD.n1037 VDD.n1035 0.001
R7653 VDD.n912 VDD.n910 0.001
R7654 VDD.n937 VDD.n935 0.001
R7655 VDD.n1012 VDD.n1010 0.001
R7656 VDD.n987 VDD.n985 0.001
R7657 VDD.n962 VDD.n960 0.001
R7658 VDD.n887 VDD.n885 0.001
R7659 VDD.n863 VDD.n861 0.001
R7660 VDD.n538 VDD.n537 0.001
R7661 VDD.n2190 VDD.n2187 0.001
R7662 VDD.n1477 VDD.n1474 0.001
R7663 VDD.n2036 VDD.n2035 0.001
R7664 VDD.n1936 VDD.n1935 0.001
R7665 VDD.n1886 VDD.n1885 0.001
R7666 VDD.n1911 VDD.n1910 0.001
R7667 VDD.n1961 VDD.n1960 0.001
R7668 VDD.n1986 VDD.n1985 0.001
R7669 VDD.n2011 VDD.n2010 0.001
R7670 VDD.n2061 VDD.n2060 0.001
R7671 VDD.n1731 VDD.n1729 0.001
R7672 VDD.n1756 VDD.n1754 0.001
R7673 VDD.n1856 VDD.n1854 0.001
R7674 VDD.n1831 VDD.n1829 0.001
R7675 VDD.n1806 VDD.n1804 0.001
R7676 VDD.n1781 VDD.n1779 0.001
R7677 VDD.n1706 VDD.n1704 0.001
R7678 VDD.n1682 VDD.n1680 0.001
R7679 VDD.n1531 VDD.n1529 0.001
R7680 VDD.n1556 VDD.n1554 0.001
R7681 VDD.n1656 VDD.n1654 0.001
R7682 VDD.n1631 VDD.n1629 0.001
R7683 VDD.n1606 VDD.n1604 0.001
R7684 VDD.n1581 VDD.n1579 0.001
R7685 VDD.n1506 VDD.n1504 0.001
R7686 VDD.n1482 VDD.n1480 0.001
R7687 VDD.n1381 VDD.n1379 0.001
R7688 VDD.n1356 VDD.n1354 0.001
R7689 VDD.n1257 VDD.n1255 0.001
R7690 VDD.n1281 VDD.n1279 0.001
R7691 VDD.n1306 VDD.n1304 0.001
R7692 VDD.n1331 VDD.n1329 0.001
R7693 VDD.n1406 VDD.n1404 0.001
R7694 VDD.n1431 VDD.n1429 0.001
R7695 VDD.n1160 VDD.n1159 0.001
R7696 VDD.n1175 VDD.n1174 0.001
R7697 VDD.n1220 VDD.n1219 0.001
R7698 VDD.n1205 VDD.n1204 0.001
R7699 VDD.n1190 VDD.n1189 0.001
R7700 VDD.n1148 VDD.n1147 0.001
R7701 VDD.n1133 VDD.n1132 0.001
R7702 VDD.n1238 VDD.n1237 0.001
R7703 VDD.n2449 VDD.n2446 0.001
R7704 VDD.n2424 VDD.n2421 0.001
R7705 VDD.n2240 VDD.n2237 0.001
R7706 VDD.n2215 VDD.n2212 0.001
R7707 VDD.n2594 VDD.n2592 0.001
R7708 VDD.n2455 VDD.n2453 0.001
R7709 VDD.n2474 VDD.n2472 0.001
R7710 VDD.n2534 VDD.n2532 0.001
R7711 VDD.n2554 VDD.n2552 0.001
R7712 VDD.n2574 VDD.n2572 0.001
R7713 VDD.n2514 VDD.n2512 0.001
R7714 VDD.n2494 VDD.n2492 0.001
R7715 VDD.n2385 VDD.n2383 0.001
R7716 VDD.n2246 VDD.n2244 0.001
R7717 VDD.n2265 VDD.n2263 0.001
R7718 VDD.n2325 VDD.n2323 0.001
R7719 VDD.n2345 VDD.n2343 0.001
R7720 VDD.n2365 VDD.n2363 0.001
R7721 VDD.n2305 VDD.n2303 0.001
R7722 VDD.n2285 VDD.n2283 0.001
R7723 VDD.n372 VDD.n371 0.001
R7724 VDD.n3128 VDD.n3127 0.001
R7725 VDD.n3121 VDD.n3120 0.001
R7726 VDD.n3200 VDD.n3199 0.001
R7727 VDD.n3152 VDD.n3148 0.001
R7728 VDD.n2788 VDD.n2787 0.001
R7729 VDD.n2052 VDD.n2051 0.001
R7730 VDD.n1952 VDD.n1951 0.001
R7731 VDD.n1902 VDD.n1901 0.001
R7732 VDD.n1927 VDD.n1926 0.001
R7733 VDD.n1977 VDD.n1976 0.001
R7734 VDD.n2002 VDD.n2001 0.001
R7735 VDD.n2027 VDD.n2026 0.001
R7736 VDD.n2077 VDD.n2076 0.001
R7737 VDD.n814 VDD.n29 0.001
R7738 VDD.n799 VDD.n139 0.001
R7739 VDD.n166 VDD.n165 0.001
R7740 VDD.n107 VDD.n106 0.001
R7741 VDD.n56 VDD.n55 0.001
R7742 VDD.n3194 VDD.n3193 0.001
R7743 VDD.n856 VDD.n833 0.001
R7744 VDD.n2930 VDD.n2929 0.001
R7745 VDD.n413 VDD.n412 0.001
R7746 VDD.n2931 VDD.n2919 0.001
R7747 VDD.n2746 VDD.n2745 0.001
R7748 VDD.n3006 VDD.n3005 0.001
R7749 VDD.n2809 VDD.n2808 0.001
R7750 VDD.n525 VDD.n524 0.001
R7751 VDD.n1050 VDD.n1049 0.001
R7752 VDD.n925 VDD.n924 0.001
R7753 VDD.n950 VDD.n949 0.001
R7754 VDD.n1025 VDD.n1024 0.001
R7755 VDD.n1000 VDD.n999 0.001
R7756 VDD.n975 VDD.n974 0.001
R7757 VDD.n900 VDD.n899 0.001
R7758 VDD.n876 VDD.n875 0.001
R7759 VDD.n634 VDD.n633 0.001
R7760 VDD.n652 VDD.n651 0.001
R7761 VDD.n670 VDD.n669 0.001
R7762 VDD.n687 VDD.n686 0.001
R7763 VDD.n616 VDD.n615 0.001
R7764 VDD.n747 VDD.n746 0.001
R7765 VDD.n765 VDD.n764 0.001
R7766 VDD.n783 VDD.n782 0.001
R7767 VDD.n1739 VDD.n1738 0.001
R7768 VDD.n1764 VDD.n1763 0.001
R7769 VDD.n1869 VDD.n1868 0.001
R7770 VDD.n1844 VDD.n1843 0.001
R7771 VDD.n1814 VDD.n1813 0.001
R7772 VDD.n1789 VDD.n1788 0.001
R7773 VDD.n1714 VDD.n1713 0.001
R7774 VDD.n1690 VDD.n1689 0.001
R7775 VDD.n1544 VDD.n1543 0.001
R7776 VDD.n1569 VDD.n1568 0.001
R7777 VDD.n1669 VDD.n1668 0.001
R7778 VDD.n1644 VDD.n1643 0.001
R7779 VDD.n1619 VDD.n1618 0.001
R7780 VDD.n1594 VDD.n1593 0.001
R7781 VDD.n1519 VDD.n1518 0.001
R7782 VDD.n1495 VDD.n1494 0.001
R7783 VDD.n1394 VDD.n1393 0.001
R7784 VDD.n1369 VDD.n1368 0.001
R7785 VDD.n1270 VDD.n1269 0.001
R7786 VDD.n1294 VDD.n1293 0.001
R7787 VDD.n1319 VDD.n1318 0.001
R7788 VDD.n1344 VDD.n1343 0.001
R7789 VDD.n1419 VDD.n1418 0.001
R7790 VDD.n1444 VDD.n1443 0.001
R7791 VDD.n2600 VDD.n2599 0.001
R7792 VDD.n2461 VDD.n2460 0.001
R7793 VDD.n2480 VDD.n2479 0.001
R7794 VDD.n2540 VDD.n2539 0.001
R7795 VDD.n2560 VDD.n2559 0.001
R7796 VDD.n2580 VDD.n2579 0.001
R7797 VDD.n2520 VDD.n2519 0.001
R7798 VDD.n2500 VDD.n2499 0.001
R7799 VDD.n2396 VDD.n2395 0.001
R7800 VDD.n2252 VDD.n2251 0.001
R7801 VDD.n2271 VDD.n2270 0.001
R7802 VDD.n2336 VDD.n2335 0.001
R7803 VDD.n2356 VDD.n2355 0.001
R7804 VDD.n2376 VDD.n2375 0.001
R7805 VDD.n2311 VDD.n2310 0.001
R7806 VDD.n2291 VDD.n2290 0.001
R7807 VDD.n2122 VDD.n2121 0.001
R7808 VDD.n2116 VDD.n2115 0.001
R7809 VDD.n2110 VDD.n2109 0.001
R7810 VDD.n2104 VDD.n2103 0.001
R7811 VDD.n2098 VDD.n2097 0.001
R7812 VDD.n2080 VDD.n2079 0.001
R7813 VDD.n2092 VDD.n2091 0.001
R7814 VDD.n3102 VDD.n3099 0.001
R7815 VDD.n2086 VDD.n2085 0.001
R7816 VDD.n1053 VDD.n1034 0.001
R7817 VDD.n928 VDD.n909 0.001
R7818 VDD.n953 VDD.n934 0.001
R7819 VDD.n1028 VDD.n1009 0.001
R7820 VDD.n1003 VDD.n984 0.001
R7821 VDD.n978 VDD.n959 0.001
R7822 VDD.n903 VDD.n884 0.001
R7823 VDD.n879 VDD.n860 0.001
R7824 VDD.n1748 VDD.n1747 0.001
R7825 VDD.n1773 VDD.n1772 0.001
R7826 VDD.n1873 VDD.n1872 0.001
R7827 VDD.n1848 VDD.n1847 0.001
R7828 VDD.n1823 VDD.n1822 0.001
R7829 VDD.n1798 VDD.n1797 0.001
R7830 VDD.n1723 VDD.n1722 0.001
R7831 VDD.n1699 VDD.n1698 0.001
R7832 VDD.n1548 VDD.n1547 0.001
R7833 VDD.n1573 VDD.n1572 0.001
R7834 VDD.n1673 VDD.n1672 0.001
R7835 VDD.n1648 VDD.n1647 0.001
R7836 VDD.n1623 VDD.n1622 0.001
R7837 VDD.n1598 VDD.n1597 0.001
R7838 VDD.n1523 VDD.n1522 0.001
R7839 VDD.n1499 VDD.n1498 0.001
R7840 VDD.n1398 VDD.n1397 0.001
R7841 VDD.n1373 VDD.n1372 0.001
R7842 VDD.n1274 VDD.n1273 0.001
R7843 VDD.n1298 VDD.n1297 0.001
R7844 VDD.n1323 VDD.n1322 0.001
R7845 VDD.n1348 VDD.n1347 0.001
R7846 VDD.n1423 VDD.n1422 0.001
R7847 VDD.n1448 VDD.n1447 0.001
R7848 VDD.n3103 VDD.n3102 0.001
R7849 VDD.n337 VDD.n336 0.001
R7850 VDD.n535 VDD.n534 0.001
R7851 VDD.n2642 VDD.n2191 0.001
R7852 VDD.n2645 VDD.n1478 0.001
R7853 VDD.n2637 VDD.n2450 0.001
R7854 VDD.n2638 VDD.n2425 0.001
R7855 VDD.n2640 VDD.n2241 0.001
R7856 VDD.n2641 VDD.n2216 0.001
R7857 VDD.n3260 VDD.n3251 0.001
R7858 VDD.n2908 VDD.n2900 0.001
R7859 VDD.n2681 VDD.n2673 0.001
R7860 VDD.n2672 VDD.n2664 0.001
R7861 VDD.n412 VDD.n411 0.001
R7862 VDD.n2929 VDD.n2928 0.001
R7863 VDD.n311 VDD.n303 0.001
R7864 VDD.n302 VDD.n294 0.001
R7865 VDD.n393 VDD.n385 0.001
R7866 VDD.n402 VDD.n394 0.001
R7867 VDD.n2662 VDD.n2654 0.001
R7868 VDD.n715 VDD.n707 0.001
R7869 VDD.n2663 VDD.n2646 0.001
R7870 VDD.n717 VDD.n699 0.001
R7871 VDD.n573 VDD.n286 0.001
R7872 VDD.n285 VDD.n276 0.001
R7873 VDD.n274 VDD.n265 0.001
R7874 VDD.n1251 VDD.n1075 0.001
R7875 VDD.n1247 VDD.n1108 0.001
R7876 VDD.n1253 VDD.n1058 0.001
R7877 VDD.n609 VDD.n601 0.001
R7878 VDD.n739 VDD.n738 0.001
R7879 VDD.n2134 VDD.n2052 0.001
R7880 VDD.n2138 VDD.n1952 0.001
R7881 VDD.n2140 VDD.n1902 0.001
R7882 VDD.n2139 VDD.n1927 0.001
R7883 VDD.n2137 VDD.n1977 0.001
R7884 VDD.n2136 VDD.n2002 0.001
R7885 VDD.n2135 VDD.n2027 0.001
R7886 VDD.n2133 VDD.n2077 0.001
R7887 VDD.n2919 VDD.n2918 0.001
R7888 VDD.n2719 VDD.n2717 0.001
R7889 VDD.n2874 VDD.n2873 0.001
R7890 VDD.n3217 VDD.n3202 0.001
R7891 VDD.n3116 VDD.n3115 0.001
R7892 VDD.n3104 VDD.n3103 0.001
R7893 VDD.n539 VDD.n538 0.001
R7894 VDD.n2834 VDD.n2833 0.001
R7895 VDD.n2877 VDD.n2865 0.001
R7896 VDD.n2887 VDD.n2886 0.001
R7897 VDD.n2899 VDD.n2898 0.001
R7898 VDD.n3235 VDD.n3234 0.001
R7899 VDD.n3215 VDD.n3212 0.001
R7900 VDD.n338 VDD.n337 0.001
R7901 VDD.n505 VDD.n504 0.001
R7902 VDD.n2726 VDD.n2725 0.001
R7903 VDD.n553 VDD.n552 0.001
R7904 VDD.n2886 VDD.n2885 0.001
R7905 VDD.n1057 VDD.n1056 0.001
R7906 VDD.n932 VDD.n931 0.001
R7907 VDD.n957 VDD.n956 0.001
R7908 VDD.n1032 VDD.n1031 0.001
R7909 VDD.n1007 VDD.n1006 0.001
R7910 VDD.n982 VDD.n981 0.001
R7911 VDD.n907 VDD.n906 0.001
R7912 VDD.n1752 VDD.n1751 0.001
R7913 VDD.n1777 VDD.n1776 0.001
R7914 VDD.n1877 VDD.n1876 0.001
R7915 VDD.n1852 VDD.n1851 0.001
R7916 VDD.n1827 VDD.n1826 0.001
R7917 VDD.n1802 VDD.n1801 0.001
R7918 VDD.n1727 VDD.n1726 0.001
R7919 VDD.n1552 VDD.n1551 0.001
R7920 VDD.n1577 VDD.n1576 0.001
R7921 VDD.n1677 VDD.n1676 0.001
R7922 VDD.n1652 VDD.n1651 0.001
R7923 VDD.n1627 VDD.n1626 0.001
R7924 VDD.n1602 VDD.n1601 0.001
R7925 VDD.n1527 VDD.n1526 0.001
R7926 VDD.n1402 VDD.n1401 0.001
R7927 VDD.n1377 VDD.n1376 0.001
R7928 VDD.n1302 VDD.n1301 0.001
R7929 VDD.n1327 VDD.n1326 0.001
R7930 VDD.n1352 VDD.n1351 0.001
R7931 VDD.n1427 VDD.n1426 0.001
R7932 VDD.n1452 VDD.n1451 0.001
R7933 VDD.n3153 VDD.n3152 0.001
R7934 VDD.n3201 VDD.n3200 0.001
R7935 VDD.n372 VDD.n369 0.001
R7936 VDD.n2977 VDD.n2976 0.001
R7937 VDD.n3227 VDD.n3226 0.001
R7938 VDD.n3218 VDD.n3217 0.001
R7939 VDD.n3047 VDD.n3046 0.001
R7940 VDD.n322 VDD.n321 0.001
R7941 VDD.n2849 VDD.n2848 0.001
R7942 VDD.n2863 VDD.n2862 0.001
R7943 VDD.n3138 VDD.n3137 0.001
R7944 VDD.n3122 VDD.n3121 0.001
R7945 VDD.n3129 VDD.n3128 0.001
R7946 VDD.n3249 VDD.n3248 0.001
R7947 VDD.n3115 VDD.n3114 0.001
R7948 VDD.n562 VDD.n556 0.001
R7949 VDD.n2823 VDD.n2822 0.001
R7950 VDD.n2854 VDD.n2853 0.001
R7951 VDD.n538 VDD.n526 0.001
R7952 VDD.n2878 VDD.n2877 0.001
R7953 VDD.n552 VDD.n543 0.001
R7954 VDD.n569 VDD.n563 0.001
R7955 VDD.n2165 VDD.n2164 0.001
R7956 VDD.n2633 VDD.n2632 0.001
R7957 VDD.n2788 VDD.n2780 0.001
R7958 VDD.n2985 VDD.n2978 0.001
R7959 VDD.n436 VDD.n429 0.001
R7960 VDD.n3161 VDD.n3154 0.001
R7961 VDD.n3055 VDD.n3048 0.001
R7962 VDD.n337 VDD.n323 0.001
R7963 VDD.n504 VDD.n490 0.001
R7964 VDD.n2725 VDD.n2713 0.001
R7965 VDD.n3240 VDD.n3239 0.001
R7966 VDD.n380 VDD.n372 0.001
R7967 VDD.n468 VDD.n456 0.001
R7968 VDD.n3087 VDD.n3075 0.001
R7969 VDD.n504 VDD.n503 0.001
R7970 VDD.n2848 VDD.n2836 0.001
R7971 VDD.n2898 VDD.n2897 0.001
R7972 VDD.n2180 VDD.n2179 0.001
R7973 VDD.n1467 VDD.n1466 0.001
R7974 VDD.n2439 VDD.n2438 0.001
R7975 VDD.n2414 VDD.n2413 0.001
R7976 VDD.n2230 VDD.n2229 0.001
R7977 VDD.n2205 VDD.n2204 0.001
R7978 VDD.n3226 VDD.n3219 0.001
R7979 VDD.n2862 VDD.n2855 0.001
R7980 VDD.n3137 VDD.n3130 0.001
R7981 VDD.n2833 VDD.n2824 0.001
R7982 VDD.n2898 VDD.n2888 0.001
R7983 VDD.n3248 VDD.n3241 0.001
R7984 VDD.n437 VDD.n436 0.001
R7985 VDD.n3115 VDD.n3105 0.001
R7986 VDD.n3162 VDD.n3161 0.001
R7987 VDD.n3056 VDD.n3055 0.001
R7988 VDD.n2986 VDD.n2985 0.001
R7989 VDD.n2789 VDD.n2788 0.001
R7990 VDD.n2822 VDD.n2819 0.001
R7991 VDD.n2853 VDD.n2850 0.001
R7992 VDD.n3103 VDD.n3098 0.001
R7993 VDD.n2886 VDD.n2879 0.001
R7994 VDD.n3121 VDD.n3118 0.001
R7995 VDD.n3128 VDD.n3123 0.001
R7996 VDD.n3234 VDD.n3229 0.001
R7997 VDD.n3200 VDD.n3197 0.001
R7998 VDD.n3239 VDD.n3236 0.001
R7999 VDD.n1053 VDD.n1035 0.001
R8000 VDD.n1051 VDD.n1050 0.001
R8001 VDD.n928 VDD.n910 0.001
R8002 VDD.n926 VDD.n925 0.001
R8003 VDD.n953 VDD.n935 0.001
R8004 VDD.n951 VDD.n950 0.001
R8005 VDD.n1028 VDD.n1010 0.001
R8006 VDD.n1026 VDD.n1025 0.001
R8007 VDD.n1003 VDD.n985 0.001
R8008 VDD.n1001 VDD.n1000 0.001
R8009 VDD.n978 VDD.n960 0.001
R8010 VDD.n976 VDD.n975 0.001
R8011 VDD.n903 VDD.n885 0.001
R8012 VDD.n901 VDD.n900 0.001
R8013 VDD.n879 VDD.n861 0.001
R8014 VDD.n877 VDD.n876 0.001
R8015 VDD.n2848 VDD.n2847 0.001
R8016 VDD.n2833 VDD.n2832 0.001
R8017 VDD.n3217 VDD.n3216 0.001
R8018 VDD.n635 VDD.n634 0.001
R8019 VDD.n653 VDD.n652 0.001
R8020 VDD.n671 VDD.n670 0.001
R8021 VDD.n688 VDD.n687 0.001
R8022 VDD.n617 VDD.n616 0.001
R8023 VDD.n748 VDD.n747 0.001
R8024 VDD.n766 VDD.n765 0.001
R8025 VDD.n784 VDD.n783 0.001
R8026 VDD.n2125 VDD.n2122 0.001
R8027 VDD.n2126 VDD.n2119 0.001
R8028 VDD.n2119 VDD.n2116 0.001
R8029 VDD.n2127 VDD.n2113 0.001
R8030 VDD.n2113 VDD.n2110 0.001
R8031 VDD.n2128 VDD.n2107 0.001
R8032 VDD.n2107 VDD.n2104 0.001
R8033 VDD.n2129 VDD.n2101 0.001
R8034 VDD.n2101 VDD.n2098 0.001
R8035 VDD.n2130 VDD.n2095 0.001
R8036 VDD.n2095 VDD.n2092 0.001
R8037 VDD.n2131 VDD.n2089 0.001
R8038 VDD.n2089 VDD.n2086 0.001
R8039 VDD.n2132 VDD.n2083 0.001
R8040 VDD.n2083 VDD.n2080 0.001
R8041 VDD.n1747 VDD.n1731 0.001
R8042 VDD.n1740 VDD.n1739 0.001
R8043 VDD.n1772 VDD.n1756 0.001
R8044 VDD.n1765 VDD.n1764 0.001
R8045 VDD.n1872 VDD.n1856 0.001
R8046 VDD.n1870 VDD.n1869 0.001
R8047 VDD.n1847 VDD.n1831 0.001
R8048 VDD.n1845 VDD.n1844 0.001
R8049 VDD.n1822 VDD.n1806 0.001
R8050 VDD.n1815 VDD.n1814 0.001
R8051 VDD.n1797 VDD.n1781 0.001
R8052 VDD.n1790 VDD.n1789 0.001
R8053 VDD.n1722 VDD.n1706 0.001
R8054 VDD.n1715 VDD.n1714 0.001
R8055 VDD.n1698 VDD.n1682 0.001
R8056 VDD.n1691 VDD.n1690 0.001
R8057 VDD.n1547 VDD.n1531 0.001
R8058 VDD.n1545 VDD.n1544 0.001
R8059 VDD.n1572 VDD.n1556 0.001
R8060 VDD.n1570 VDD.n1569 0.001
R8061 VDD.n1672 VDD.n1656 0.001
R8062 VDD.n1670 VDD.n1669 0.001
R8063 VDD.n1647 VDD.n1631 0.001
R8064 VDD.n1645 VDD.n1644 0.001
R8065 VDD.n1622 VDD.n1606 0.001
R8066 VDD.n1620 VDD.n1619 0.001
R8067 VDD.n1597 VDD.n1581 0.001
R8068 VDD.n1595 VDD.n1594 0.001
R8069 VDD.n1522 VDD.n1506 0.001
R8070 VDD.n1520 VDD.n1519 0.001
R8071 VDD.n1498 VDD.n1482 0.001
R8072 VDD.n1496 VDD.n1495 0.001
R8073 VDD.n1397 VDD.n1381 0.001
R8074 VDD.n1395 VDD.n1394 0.001
R8075 VDD.n1372 VDD.n1356 0.001
R8076 VDD.n1370 VDD.n1369 0.001
R8077 VDD.n1273 VDD.n1257 0.001
R8078 VDD.n1271 VDD.n1270 0.001
R8079 VDD.n1297 VDD.n1281 0.001
R8080 VDD.n1295 VDD.n1294 0.001
R8081 VDD.n1322 VDD.n1306 0.001
R8082 VDD.n1320 VDD.n1319 0.001
R8083 VDD.n1347 VDD.n1331 0.001
R8084 VDD.n1345 VDD.n1344 0.001
R8085 VDD.n1422 VDD.n1406 0.001
R8086 VDD.n1420 VDD.n1419 0.001
R8087 VDD.n1447 VDD.n1431 0.001
R8088 VDD.n1445 VDD.n1444 0.001
R8089 VDD.n1166 VDD.n1160 0.001
R8090 VDD.n1181 VDD.n1175 0.001
R8091 VDD.n1226 VDD.n1220 0.001
R8092 VDD.n1211 VDD.n1205 0.001
R8093 VDD.n1196 VDD.n1190 0.001
R8094 VDD.n1154 VDD.n1148 0.001
R8095 VDD.n1139 VDD.n1133 0.001
R8096 VDD.n1244 VDD.n1238 0.001
R8097 VDD.n2608 VDD.n2594 0.001
R8098 VDD.n2601 VDD.n2600 0.001
R8099 VDD.n2469 VDD.n2455 0.001
R8100 VDD.n2462 VDD.n2461 0.001
R8101 VDD.n2488 VDD.n2474 0.001
R8102 VDD.n2481 VDD.n2480 0.001
R8103 VDD.n2548 VDD.n2534 0.001
R8104 VDD.n2541 VDD.n2540 0.001
R8105 VDD.n2568 VDD.n2554 0.001
R8106 VDD.n2561 VDD.n2560 0.001
R8107 VDD.n2588 VDD.n2574 0.001
R8108 VDD.n2581 VDD.n2580 0.001
R8109 VDD.n2528 VDD.n2514 0.001
R8110 VDD.n2521 VDD.n2520 0.001
R8111 VDD.n2508 VDD.n2494 0.001
R8112 VDD.n2501 VDD.n2500 0.001
R8113 VDD.n2399 VDD.n2385 0.001
R8114 VDD.n2397 VDD.n2396 0.001
R8115 VDD.n2260 VDD.n2246 0.001
R8116 VDD.n2253 VDD.n2252 0.001
R8117 VDD.n2279 VDD.n2265 0.001
R8118 VDD.n2272 VDD.n2271 0.001
R8119 VDD.n2339 VDD.n2325 0.001
R8120 VDD.n2337 VDD.n2336 0.001
R8121 VDD.n2359 VDD.n2345 0.001
R8122 VDD.n2357 VDD.n2356 0.001
R8123 VDD.n2379 VDD.n2365 0.001
R8124 VDD.n2377 VDD.n2376 0.001
R8125 VDD.n2319 VDD.n2305 0.001
R8126 VDD.n2312 VDD.n2311 0.001
R8127 VDD.n2299 VDD.n2285 0.001
R8128 VDD.n2292 VDD.n2291 0.001
R8129 a_3642_11724.n2 a_3642_11724.t4 990.34
R8130 a_3642_11724.n2 a_3642_11724.t5 408.211
R8131 a_3642_11724.n1 a_3642_11724.t6 286.438
R8132 a_3642_11724.n1 a_3642_11724.t7 286.438
R8133 a_3642_11724.n4 a_3642_11724.n0 185.55
R8134 a_3642_11724.t4 a_3642_11724.n1 160.666
R8135 a_3642_11724.t1 a_3642_11724.n4 28.568
R8136 a_3642_11724.n0 a_3642_11724.t3 28.565
R8137 a_3642_11724.n0 a_3642_11724.t2 28.565
R8138 a_3642_11724.n3 a_3642_11724.n2 21.382
R8139 a_3642_11724.n3 a_3642_11724.t0 21.376
R8140 a_3642_11724.n4 a_3642_11724.n3 1.637
R8141 a_3951_1740.n0 a_3951_1740.t6 14.282
R8142 a_3951_1740.t0 a_3951_1740.n0 14.282
R8143 a_3951_1740.n0 a_3951_1740.n9 89.977
R8144 a_3951_1740.n6 a_3951_1740.n7 75.815
R8145 a_3951_1740.n9 a_3951_1740.n6 77.456
R8146 a_3951_1740.n9 a_3951_1740.n4 77.456
R8147 a_3951_1740.n4 a_3951_1740.n2 77.784
R8148 a_3951_1740.n7 a_3951_1740.n8 167.433
R8149 a_3951_1740.n8 a_3951_1740.t4 14.282
R8150 a_3951_1740.n8 a_3951_1740.t5 14.282
R8151 a_3951_1740.n7 a_3951_1740.t3 104.259
R8152 a_3951_1740.n6 a_3951_1740.n5 89.977
R8153 a_3951_1740.n5 a_3951_1740.t7 14.282
R8154 a_3951_1740.n5 a_3951_1740.t2 14.282
R8155 a_3951_1740.n4 a_3951_1740.n3 89.977
R8156 a_3951_1740.n3 a_3951_1740.t8 14.282
R8157 a_3951_1740.n3 a_3951_1740.t1 14.282
R8158 a_3951_1740.n2 a_3951_1740.t9 104.259
R8159 a_3951_1740.n2 a_3951_1740.n1 167.433
R8160 a_3951_1740.n1 a_3951_1740.t11 14.282
R8161 a_3951_1740.n1 a_3951_1740.t10 14.282
R8162 a_38721_16161.n6 a_38721_16161.n5 501.28
R8163 a_38721_16161.t9 a_38721_16161.t16 437.233
R8164 a_38721_16161.t18 a_38721_16161.t13 415.315
R8165 a_38721_16161.t15 a_38721_16161.n3 313.873
R8166 a_38721_16161.n5 a_38721_16161.t14 294.986
R8167 a_38721_16161.n2 a_38721_16161.t10 272.288
R8168 a_38721_16161.n6 a_38721_16161.t8 236.009
R8169 a_38721_16161.n9 a_38721_16161.t9 216.627
R8170 a_38721_16161.n7 a_38721_16161.t18 216.111
R8171 a_38721_16161.n8 a_38721_16161.t7 214.686
R8172 a_38721_16161.t16 a_38721_16161.n8 214.686
R8173 a_38721_16161.n1 a_38721_16161.t11 214.335
R8174 a_38721_16161.t13 a_38721_16161.n1 214.335
R8175 a_38721_16161.n4 a_38721_16161.t19 190.152
R8176 a_38721_16161.n4 a_38721_16161.t15 190.152
R8177 a_38721_16161.n2 a_38721_16161.t5 160.666
R8178 a_38721_16161.n3 a_38721_16161.t4 160.666
R8179 a_38721_16161.n7 a_38721_16161.n6 148.428
R8180 a_38721_16161.n5 a_38721_16161.t6 110.859
R8181 a_38721_16161.n3 a_38721_16161.n2 96.129
R8182 a_38721_16161.n8 a_38721_16161.t17 80.333
R8183 a_38721_16161.n1 a_38721_16161.t12 80.333
R8184 a_38721_16161.t8 a_38721_16161.n4 80.333
R8185 a_38721_16161.n0 a_38721_16161.t2 28.57
R8186 a_38721_16161.n11 a_38721_16161.t1 28.565
R8187 a_38721_16161.t0 a_38721_16161.n11 28.565
R8188 a_38721_16161.n0 a_38721_16161.t3 17.638
R8189 a_38721_16161.n10 a_38721_16161.n9 5.638
R8190 a_38721_16161.n9 a_38721_16161.n7 2.923
R8191 a_38721_16161.n11 a_38721_16161.n10 0.693
R8192 a_38721_16161.n10 a_38721_16161.n0 0.597
R8193 a_39263_15765.n0 a_39263_15765.n1 0.001
R8194 a_39263_15765.n0 a_39263_15765.t1 14.282
R8195 a_39263_15765.t0 a_39263_15765.n0 14.282
R8196 a_39263_15765.n1 a_39263_15765.n9 267.767
R8197 a_39263_15765.n9 a_39263_15765.t3 14.282
R8198 a_39263_15765.n9 a_39263_15765.t2 14.282
R8199 a_39263_15765.n1 a_39263_15765.n7 0.669
R8200 a_39263_15765.n7 a_39263_15765.n8 1.511
R8201 a_39263_15765.n8 a_39263_15765.t10 14.282
R8202 a_39263_15765.n8 a_39263_15765.t11 14.282
R8203 a_39263_15765.n7 a_39263_15765.n6 0.227
R8204 a_39263_15765.n6 a_39263_15765.n3 0.2
R8205 a_39263_15765.n6 a_39263_15765.n5 0.575
R8206 a_39263_15765.n5 a_39263_15765.t5 16.058
R8207 a_39263_15765.n5 a_39263_15765.n4 0.999
R8208 a_39263_15765.n4 a_39263_15765.t6 14.282
R8209 a_39263_15765.n4 a_39263_15765.t4 14.282
R8210 a_39263_15765.n3 a_39263_15765.n2 0.999
R8211 a_39263_15765.n2 a_39263_15765.t8 14.282
R8212 a_39263_15765.n2 a_39263_15765.t9 14.282
R8213 a_39263_15765.n3 a_39263_15765.t7 16.058
R8214 a_13130_8992.n1 a_13130_8992.t7 990.34
R8215 a_13130_8992.n1 a_13130_8992.t6 408.211
R8216 a_13130_8992.n0 a_13130_8992.t5 286.438
R8217 a_13130_8992.n0 a_13130_8992.t4 286.438
R8218 a_13130_8992.n4 a_13130_8992.n3 185.55
R8219 a_13130_8992.t7 a_13130_8992.n0 160.666
R8220 a_13130_8992.n3 a_13130_8992.t2 28.568
R8221 a_13130_8992.n4 a_13130_8992.t3 28.565
R8222 a_13130_8992.t0 a_13130_8992.n4 28.565
R8223 a_13130_8992.n2 a_13130_8992.t1 21.476
R8224 a_13130_8992.n2 a_13130_8992.n1 12.305
R8225 a_13130_8992.n3 a_13130_8992.n2 1.537
R8226 a_13711_11724.t0 a_13711_11724.n0 14.282
R8227 a_13711_11724.n0 a_13711_11724.t1 14.282
R8228 a_13711_11724.n0 a_13711_11724.n9 89.977
R8229 a_13711_11724.n9 a_13711_11724.n7 77.784
R8230 a_13711_11724.n9 a_13711_11724.n6 77.456
R8231 a_13711_11724.n6 a_13711_11724.n4 77.456
R8232 a_13711_11724.n4 a_13711_11724.n2 75.815
R8233 a_13711_11724.n7 a_13711_11724.n8 167.433
R8234 a_13711_11724.n8 a_13711_11724.t9 14.282
R8235 a_13711_11724.n8 a_13711_11724.t10 14.282
R8236 a_13711_11724.n7 a_13711_11724.t11 104.259
R8237 a_13711_11724.n6 a_13711_11724.n5 89.977
R8238 a_13711_11724.n5 a_13711_11724.t2 14.282
R8239 a_13711_11724.n5 a_13711_11724.t7 14.282
R8240 a_13711_11724.n4 a_13711_11724.n3 89.977
R8241 a_13711_11724.n3 a_13711_11724.t8 14.282
R8242 a_13711_11724.n3 a_13711_11724.t6 14.282
R8243 a_13711_11724.n2 a_13711_11724.t4 104.259
R8244 a_13711_11724.n2 a_13711_11724.n1 167.433
R8245 a_13711_11724.n1 a_13711_11724.t3 14.282
R8246 a_13711_11724.n1 a_13711_11724.t5 14.282
R8247 A[3].n8 A[3].n7 3150.11
R8248 A[3].n36 A[3].n26 2170.52
R8249 A[3].n15 A[3].t39 990.34
R8250 A[3].n17 A[3].t12 867.497
R8251 A[3].n37 A[3].n19 647.392
R8252 A[3].n17 A[3].t6 591.811
R8253 A[3].t23 A[3].t31 575.234
R8254 A[3].n31 A[3].n30 535.449
R8255 A[3].t44 A[3].t0 437.233
R8256 A[3].t48 A[3].t36 437.233
R8257 A[3].t10 A[3].t41 437.233
R8258 A[3].t45 A[3].t50 437.233
R8259 A[3].t16 A[3].t1 415.315
R8260 A[3].t33 A[3].t18 415.315
R8261 A[3].t30 A[3].t40 415.315
R8262 A[3].n5 A[3].n4 412.11
R8263 A[3].n15 A[3].t20 408.211
R8264 A[3].n2 A[3].t57 394.151
R8265 A[3].t35 A[3].n28 313.873
R8266 A[3].n30 A[3].t11 294.986
R8267 A[3].n4 A[3].t53 294.653
R8268 A[3].n14 A[3].t4 286.438
R8269 A[3].n14 A[3].t42 286.438
R8270 A[3].n16 A[3].t5 286.438
R8271 A[3].n16 A[3].t15 286.438
R8272 A[3].n10 A[3].t59 284.688
R8273 A[3].n27 A[3].t46 272.288
R8274 A[3].n1 A[3].t7 269.523
R8275 A[3].t57 A[3].n1 269.523
R8276 A[3].n31 A[3].t51 245.184
R8277 A[3].n5 A[3].n3 224.13
R8278 A[3].n25 A[3].t33 221.468
R8279 A[3].n12 A[3].t44 221.268
R8280 A[3].n22 A[3].t48 219.798
R8281 A[3].n33 A[3].t45 218.628
R8282 A[3].n22 A[3].t16 217.276
R8283 A[3].n25 A[3].t30 217.129
R8284 A[3].n35 A[3].t10 217.024
R8285 A[3].n9 A[3].t37 214.686
R8286 A[3].t0 A[3].n9 214.686
R8287 A[3].n21 A[3].t32 214.686
R8288 A[3].t36 A[3].n21 214.686
R8289 A[3].n34 A[3].t24 214.686
R8290 A[3].t41 A[3].n34 214.686
R8291 A[3].n32 A[3].t34 214.686
R8292 A[3].t50 A[3].n32 214.686
R8293 A[3].n20 A[3].t58 214.335
R8294 A[3].t1 A[3].n20 214.335
R8295 A[3].n23 A[3].t26 214.335
R8296 A[3].t18 A[3].n23 214.335
R8297 A[3].n24 A[3].t56 214.335
R8298 A[3].t40 A[3].n24 214.335
R8299 A[3].n0 A[3].t52 198.043
R8300 A[3].n29 A[3].t35 190.152
R8301 A[3].n29 A[3].t54 190.152
R8302 A[3].n6 A[3].t27 185.301
R8303 A[3].n6 A[3].t8 185.301
R8304 A[3].n12 A[3].n11 182.757
R8305 A[3].n10 A[3].t21 160.666
R8306 A[3].n11 A[3].t23 160.666
R8307 A[3].n1 A[3].t17 160.666
R8308 A[3].t39 A[3].n14 160.666
R8309 A[3].t12 A[3].n16 160.666
R8310 A[3].n27 A[3].t49 160.666
R8311 A[3].n28 A[3].t14 160.666
R8312 A[3].n8 A[3].n5 141.789
R8313 A[3].n7 A[3].t29 140.583
R8314 A[3].n11 A[3].n10 115.593
R8315 A[3].n4 A[3].t25 111.663
R8316 A[3].n30 A[3].t22 110.859
R8317 A[3].n6 A[3].t43 107.646
R8318 A[3].n3 A[3].n2 97.816
R8319 A[3].n28 A[3].n27 96.129
R8320 A[3].n0 A[3].t9 93.989
R8321 A[3].n9 A[3].t19 80.333
R8322 A[3].n2 A[3].t28 80.333
R8323 A[3].n21 A[3].t13 80.333
R8324 A[3].n20 A[3].t3 80.333
R8325 A[3].n23 A[3].t2 80.333
R8326 A[3].n24 A[3].t55 80.333
R8327 A[3].n34 A[3].t38 80.333
R8328 A[3].t51 A[3].n29 80.333
R8329 A[3].n32 A[3].t47 80.333
R8330 A[3].n7 A[3].n6 61.856
R8331 A[3].n26 A[3].n25 54.612
R8332 A[3].n26 A[3].n22 49.781
R8333 A[3] A[3].n37 45.547
R8334 A[3].n13 A[3].n12 30.336
R8335 A[3].n36 A[3].n35 28.756
R8336 A[3].n18 A[3].n17 25.077
R8337 A[3].n19 A[3].n18 14.913
R8338 A[3].n33 A[3].n31 14.9
R8339 A[3].n13 A[3].n8 13.792
R8340 A[3].n19 A[3].n13 12.49
R8341 A[3].n3 A[3].n0 6.615
R8342 A[3].n37 A[3].n36 4.815
R8343 A[3].n35 A[3].n33 2.599
R8344 A[3].n18 A[3].n15 0.004
R8345 a_19763_16387.n0 a_19763_16387.t9 214.335
R8346 a_19763_16387.t7 a_19763_16387.n0 214.335
R8347 a_19763_16387.n1 a_19763_16387.t7 143.851
R8348 a_19763_16387.n1 a_19763_16387.t8 135.658
R8349 a_19763_16387.n0 a_19763_16387.t10 80.333
R8350 a_19763_16387.n2 a_19763_16387.t0 28.565
R8351 a_19763_16387.n2 a_19763_16387.t1 28.565
R8352 a_19763_16387.n4 a_19763_16387.t2 28.565
R8353 a_19763_16387.n4 a_19763_16387.t6 28.565
R8354 a_19763_16387.n7 a_19763_16387.t5 28.565
R8355 a_19763_16387.t4 a_19763_16387.n7 28.565
R8356 a_19763_16387.n3 a_19763_16387.t3 9.714
R8357 a_19763_16387.n3 a_19763_16387.n2 1.003
R8358 a_19763_16387.n6 a_19763_16387.n5 0.833
R8359 a_19763_16387.n5 a_19763_16387.n4 0.653
R8360 a_19763_16387.n7 a_19763_16387.n6 0.653
R8361 a_19763_16387.n5 a_19763_16387.n3 0.341
R8362 a_19763_16387.n6 a_19763_16387.n1 0.032
R8363 a_59223_16436.n0 a_59223_16436.t5 14.282
R8364 a_59223_16436.t1 a_59223_16436.n0 14.282
R8365 a_59223_16436.n0 a_59223_16436.n12 90.416
R8366 a_59223_16436.n12 a_59223_16436.n9 74.302
R8367 a_59223_16436.n12 a_59223_16436.n11 50.575
R8368 a_59223_16436.n11 a_59223_16436.n10 157.665
R8369 a_59223_16436.n10 a_59223_16436.t4 8.7
R8370 a_59223_16436.n10 a_59223_16436.t0 8.7
R8371 a_59223_16436.n9 a_59223_16436.n8 90.436
R8372 a_59223_16436.n8 a_59223_16436.t6 14.282
R8373 a_59223_16436.n8 a_59223_16436.t7 14.282
R8374 a_59223_16436.n11 a_59223_16436.n7 122.746
R8375 a_59223_16436.n7 a_59223_16436.t2 14.282
R8376 a_59223_16436.n7 a_59223_16436.t3 14.282
R8377 a_59223_16436.n9 a_59223_16436.n1 342.688
R8378 a_59223_16436.n1 a_59223_16436.n6 126.566
R8379 a_59223_16436.n6 a_59223_16436.t15 294.653
R8380 a_59223_16436.n6 a_59223_16436.t8 111.663
R8381 a_59223_16436.n1 a_59223_16436.n5 552.333
R8382 a_59223_16436.n5 a_59223_16436.n4 6.615
R8383 a_59223_16436.n4 a_59223_16436.t10 93.989
R8384 a_59223_16436.n4 a_59223_16436.t11 198.043
R8385 a_59223_16436.n5 a_59223_16436.n3 97.816
R8386 a_59223_16436.n3 a_59223_16436.t9 80.333
R8387 a_59223_16436.n3 a_59223_16436.t14 394.151
R8388 a_59223_16436.t14 a_59223_16436.n2 269.523
R8389 a_59223_16436.n2 a_59223_16436.t13 160.666
R8390 a_59223_16436.n2 a_59223_16436.t12 269.523
R8391 VSS.n637 VSS.t715 990.34
R8392 VSS.n495 VSS.t718 867.497
R8393 VSS.n495 VSS.t403 591.811
R8394 VSS.n637 VSS.t401 408.211
R8395 VSS.n636 VSS.t714 286.438
R8396 VSS.n636 VSS.t719 286.438
R8397 VSS.n494 VSS.t717 286.438
R8398 VSS.n494 VSS.t716 286.438
R8399 VSS.t715 VSS.n636 160.666
R8400 VSS.t718 VSS.n494 160.666
R8401 VSS.n453 VSS.t30 20.763
R8402 VSS.n31 VSS.t308 20.763
R8403 VSS.n389 VSS.t271 20.763
R8404 VSS.n67 VSS.t654 20.763
R8405 VSS.n344 VSS.t134 20.763
R8406 VSS.n305 VSS.t16 20.763
R8407 VSS.n175 VSS.t276 20.763
R8408 VSS.n160 VSS.t111 20.763
R8409 VSS.n667 VSS.t650 20.763
R8410 VSS.n534 VSS.t216 20.763
R8411 VSS.n545 VSS.t293 20.763
R8412 VSS.n521 VSS.t296 20.763
R8413 VSS.n711 VSS.t355 20.763
R8414 VSS.n694 VSS.t388 20.763
R8415 VSS.n679 VSS.t78 20.763
R8416 VSS.n572 VSS.t419 20.763
R8417 VSS.n347 VSS.t363 20.763
R8418 VSS.n302 VSS.t674 20.763
R8419 VSS.n57 VSS.t604 20.763
R8420 VSS.n75 VSS.t41 20.763
R8421 VSS.n34 VSS.t360 20.763
R8422 VSS.n23 VSS.t154 20.763
R8423 VSS.n172 VSS.t568 20.763
R8424 VSS.n296 VSS.t245 20.763
R8425 VSS.n317 VSS.t328 20.763
R8426 VSS.n341 VSS.t481 20.763
R8427 VSS.n456 VSS.t249 20.763
R8428 VSS.n429 VSS.t596 20.763
R8429 VSS.n392 VSS.t527 20.763
R8430 VSS.n369 VSS.t229 20.763
R8431 VSS.n129 VSS.t160 20.763
R8432 VSS.n271 VSS.t322 20.763
R8433 VSS.n418 VSS.t613 20.763
R8434 VSS.n415 VSS.t366 20.763
R8435 VSS.n352 VSS.t450 20.763
R8436 VSS.n355 VSS.t546 20.763
R8437 VSS.n126 VSS.t165 20.763
R8438 VSS.n123 VSS.t630 20.763
R8439 VSS.n182 VSS.t208 20.763
R8440 VSS.n266 VSS.t255 20.763
R8441 VSS.n5 VSS.t382 20.763
R8442 VSS.n3 VSS.t151 20.763
R8443 VSS.n481 VSS.t218 20.763
R8444 VSS.n1 VSS.t212 20.763
R8445 VSS.n488 VSS.t392 20.763
R8446 VSS.n484 VSS.t353 20.763
R8447 VSS.n721 VSS.t420 20.763
R8448 VSS.n7 VSS.t385 20.763
R8449 VSS.n672 VSS.t254 20.676
R8450 VSS.n651 VSS.t227 20.676
R8451 VSS.n651 VSS.t121 20.676
R8452 VSS.n672 VSS.t321 20.676
R8453 VSS.n718 VSS.t370 20.676
R8454 VSS.n695 VSS.t307 20.676
R8455 VSS.n683 VSS.t628 20.676
R8456 VSS.n651 VSS.t597 20.676
R8457 VSS VSS.t555 20.675
R8458 VSS VSS.t636 20.675
R8459 VSS VSS.t516 20.675
R8460 VSS VSS.t608 20.675
R8461 VSS VSS.t518 20.675
R8462 VSS VSS.t517 20.675
R8463 VSS.n486 VSS.t633 20.675
R8464 VSS.n482 VSS.t638 20.675
R8465 VSS.n454 VSS.t565 20.606
R8466 VSS.n32 VSS.t583 20.606
R8467 VSS.n390 VSS.t647 20.606
R8468 VSS.n68 VSS.t687 20.606
R8469 VSS.n345 VSS.t197 20.606
R8470 VSS.n306 VSS.t671 20.606
R8471 VSS.n176 VSS.t99 20.606
R8472 VSS.n161 VSS.t694 20.606
R8473 VSS.n348 VSS.t149 20.606
R8474 VSS.n303 VSS.t415 20.606
R8475 VSS.n58 VSS.t27 20.606
R8476 VSS.n76 VSS.t424 20.606
R8477 VSS.n35 VSS.t502 20.606
R8478 VSS.n24 VSS.t591 20.606
R8479 VSS.n173 VSS.t146 20.606
R8480 VSS.n297 VSS.t703 20.606
R8481 VSS.n318 VSS.t381 20.606
R8482 VSS.n342 VSS.t214 20.606
R8483 VSS.n457 VSS.t558 20.606
R8484 VSS.n430 VSS.t617 20.606
R8485 VSS.n393 VSS.t701 20.606
R8486 VSS.n370 VSS.t541 20.606
R8487 VSS.n130 VSS.t319 20.606
R8488 VSS.n272 VSS.t95 20.606
R8489 VSS.n419 VSS.t713 20.606
R8490 VSS.n416 VSS.t236 20.606
R8491 VSS.n353 VSS.t42 20.606
R8492 VSS.n356 VSS.t414 20.606
R8493 VSS.n127 VSS.t145 20.606
R8494 VSS.n124 VSS.t303 20.606
R8495 VSS.n183 VSS.t504 20.606
R8496 VSS.n267 VSS.t129 20.606
R8497 VSS.n185 VSS.t663 20.5
R8498 VSS.n192 VSS.t708 20.5
R8499 VSS.n190 VSS.t193 20.5
R8500 VSS.n188 VSS.t412 20.5
R8501 VSS.n186 VSS.t185 20.224
R8502 VSS.n256 VSS.t692 20.223
R8503 VSS.n256 VSS.t175 20.223
R8504 VSS.n256 VSS.t575 20.223
R8505 VSS.n599 VSS.t230 18.459
R8506 VSS.n601 VSS.t601 18.459
R8507 VSS.n563 VSS.t627 18.459
R8508 VSS.n532 VSS.t545 18.459
R8509 VSS.n650 VSS.t251 18.459
R8510 VSS.n596 VSS.t120 18.452
R8511 VSS.n577 VSS.t48 18.452
R8512 VSS.n536 VSS.t368 18.452
R8513 VSS.n496 VSS.n495 18.448
R8514 VSS.n546 VSS.t585 18.304
R8515 VSS.n652 VSS.t213 18.304
R8516 VSS.n665 VSS.t676 18.291
R8517 VSS.n674 VSS.t246 18.291
R8518 VSS.n503 VSS.t539 18.291
R8519 VSS.n668 VSS.t625 18.291
R8520 VSS.n696 VSS.t467 18.291
R8521 VSS.n709 VSS.t573 18.291
R8522 VSS.n284 VSS.t169 18.185
R8523 VSS.n332 VSS.t581 18.185
R8524 VSS.n379 VSS.t423 18.185
R8525 VSS.n464 VSS.t68 18.185
R8526 VSS.n396 VSS.t262 18.185
R8527 VSS.n95 VSS.t540 18.185
R8528 VSS.n153 VSS.t176 18.185
R8529 VSS.n17 VSS.t266 18.185
R8530 VSS.n50 VSS.t506 18.185
R8531 VSS.n90 VSS.t174 18.185
R8532 VSS.n132 VSS.t493 18.185
R8533 VSS.n407 VSS.t463 18.185
R8534 VSS.n108 VSS.t351 18.185
R8535 VSS.n131 VSS.t223 18.185
R8536 VSS.n471 VSS.t707 18.185
R8537 VSS.n11 VSS.t336 18.185
R8538 VSS.n44 VSS.t200 18.185
R8539 VSS.n84 VSS.t556 18.185
R8540 VSS.n142 VSS.t13 18.185
R8541 VSS.n460 VSS.t470 18.185
R8542 VSS.n78 VSS.t205 18.185
R8543 VSS.n148 VSS.t509 18.185
R8544 VSS.n38 VSS.t461 18.185
R8545 VSS.n102 VSS.t210 18.185
R8546 VSS.n469 VSS.t537 18.185
R8547 VSS.n136 VSS.t96 18.185
R8548 VSS.n402 VSS.t459 18.185
R8549 VSS.n423 VSS.t123 18.185
R8550 VSS.n361 VSS.t38 18.185
R8551 VSS.n120 VSS.t614 18.185
R8552 VSS.n179 VSS.t557 18.185
R8553 VSS.n358 VSS.t533 18.185
R8554 VSS.n121 VSS.t374 18.185
R8555 VSS.n180 VSS.t444 18.185
R8556 VSS.n420 VSS.t158 18.185
R8557 VSS.n357 VSS.t677 18.185
R8558 VSS.n299 VSS.t398 18.185
R8559 VSS.n178 VSS.t116 18.185
R8560 VSS.n25 VSS.t538 18.185
R8561 VSS.n60 VSS.t512 18.185
R8562 VSS.n328 VSS.t498 18.185
R8563 VSS.n283 VSS.t559 18.185
R8564 VSS.n327 VSS.t564 18.185
R8565 VSS.n282 VSS.t659 18.185
R8566 VSS.n59 VSS.t2 18.185
R8567 VSS.n26 VSS.t590 18.185
R8568 VSS.n444 VSS.t586 18.185
R8569 VSS.n262 VSS.t22 18.178
R8570 VSS.n193 VSS.t485 18.178
R8571 VSS.n260 VSS.t287 18.178
R8572 VSS.n478 VSS.t317 18.178
R8573 VSS.n477 VSS.t260 18.178
R8574 VSS.n194 VSS.t642 18.178
R8575 VSS.n261 VSS.t455 18.178
R8576 VSS.n257 VSS.t204 18.178
R8577 VSS.n195 VSS.t105 18.178
R8578 VSS.n9 VSS.t452 18.178
R8579 VSS.n258 VSS.t397 18.178
R8580 VSS.n8 VSS.t681 18.178
R8581 VSS.n196 VSS.t93 18.178
R8582 VSS.n424 VSS.t18 18.178
R8583 VSS.n362 VSS.t689 18.178
R8584 VSS.n259 VSS.t338 18.178
R8585 VSS.n300 VSS.t333 18.178
R8586 VSS.n119 VSS.t486 18.176
R8587 VSS.n363 VSS.t75 18.176
R8588 VSS.n425 VSS.t373 18.176
R8589 VSS.n36 VSS.t523 18.089
R8590 VSS.n639 VSS.t489 17.97
R8591 VSS.n648 VSS.t305 17.97
R8592 VSS.n631 VSS.t599 17.97
R8593 VSS.n62 VSS.t690 17.959
R8594 VSS.n330 VSS.t69 17.959
R8595 VSS.n315 VSS.t107 17.959
R8596 VSS.n163 VSS.t483 17.959
R8597 VSS.n367 VSS.t432 17.959
R8598 VSS.n281 VSS.t453 17.959
R8599 VSS.n648 VSS.t331 17.959
R8600 VSS.n648 VSS.t635 17.959
R8601 VSS.n648 VSS.t369 17.959
R8602 VSS.n648 VSS.t46 17.959
R8603 VSS.n648 VSS.t253 17.959
R8604 VSS.n170 VSS.t405 17.929
R8605 VSS.n118 VSS.t184 17.929
R8606 VSS.n435 VSS.t119 17.929
R8607 VSS.n64 VSS.t667 17.929
R8608 VSS.n115 VSS.t580 17.929
R8609 VSS.n276 VSS.t494 17.929
R8610 VSS.n375 VSS.t706 17.929
R8611 VSS.n440 VSS.t132 17.929
R8612 VSS.n323 VSS.t267 17.929
R8613 VSS.n269 VSS.t87 17.929
R8614 VSS.n360 VSS.t492 17.929
R8615 VSS.n422 VSS.t668 17.929
R8616 VSS.n427 VSS.t67 17.925
R8617 VSS.n365 VSS.t14 17.925
R8618 VSS.n313 VSS.t643 17.925
R8619 VSS.n264 VSS.t70 17.925
R8620 VSS.n339 VSS.t20 17.925
R8621 VSS.n292 VSS.t233 17.925
R8622 VSS.n451 VSS.t128 17.925
R8623 VSS.n387 VSS.t234 17.925
R8624 VSS.n383 VSS.t5 17.925
R8625 VSS.n447 VSS.t182 17.925
R8626 VSS.n335 VSS.t522 17.925
R8627 VSS.n287 VSS.t29 17.925
R8628 VSS.n28 VSS.t641 17.888
R8629 VSS.n432 VSS.t503 17.884
R8630 VSS.n614 VSS.t618 17.509
R8631 VSS.n644 VSS.t619 17.509
R8632 VSS.n564 VSS.t672 17.509
R8633 VSS.n703 VSS.t496 17.509
R8634 VSS.n675 VSS.t495 17.509
R8635 VSS.n653 VSS.t680 17.509
R8636 VSS.n541 VSS.t679 17.509
R8637 VSS.n584 VSS.t678 17.509
R8638 VSS.n587 VSS.t476 17.509
R8639 VSS.n559 VSS.t143 17.509
R8640 VSS.n547 VSS.t475 17.509
R8641 VSS.n625 VSS.t473 17.509
R8642 VSS.n640 VSS.t142 17.509
R8643 VSS.n669 VSS.t474 17.509
R8644 VSS.n680 VSS.t477 17.509
R8645 VSS.n700 VSS.t472 17.509
R8646 VSS.n574 VSS.t469 17.509
R8647 VSS.n618 VSS.t610 17.509
R8648 VSS.n603 VSS.t640 17.509
R8649 VSS.n529 VSS.t536 17.509
R8650 VSS.n551 VSS.t535 17.509
R8651 VSS.n663 VSS.t639 17.509
R8652 VSS.n690 VSS.t606 17.509
R8653 VSS.n707 VSS.t621 17.509
R8654 VSS.n609 VSS.t195 17.509
R8655 VSS.n554 VSS.t140 17.509
R8656 VSS.n612 VSS.t196 17.509
R8657 VSS.n582 VSS.t127 17.509
R8658 VSS.n523 VSS.t124 17.509
R8659 VSS.n657 VSS.t682 17.509
R8660 VSS.n505 VSS.t684 17.509
R8661 VSS.n716 VSS.t136 17.509
R8662 VSS.n622 VSS.t515 17.509
R8663 VSS.n557 VSS.t607 17.509
R8664 VSS.n579 VSS.t241 17.509
R8665 VSS.n686 VSS.t622 17.509
R8666 VSS.n713 VSS.t609 17.509
R8667 VSS.n660 VSS.t377 17.509
R8668 VSS.n526 VSS.t611 17.509
R8669 VSS.n606 VSS.t632 17.509
R8670 VSS.n537 VSS.t562 17.509
R8671 VSS.n567 VSS.t612 17.509
R8672 VSS.n590 VSS.t282 17.509
R8673 VSS.n632 VSS.t514 17.509
R8674 VSS.n514 VSS.t240 17.509
R8675 VSS.n507 VSS.t281 17.509
R8676 VSS.n499 VSS.t358 17.509
R8677 VSS.n491 VSS.t513 17.509
R8678 VSS.n250 VSS.t137 17.508
R8679 VSS.n199 VSS.t138 17.508
R8680 VSS.n206 VSS.t125 17.508
R8681 VSS.n229 VSS.t139 17.508
R8682 VSS.n235 VSS.t141 17.508
R8683 VSS.n242 VSS.t683 17.508
R8684 VSS.n222 VSS.t685 17.508
R8685 VSS.n215 VSS.t126 17.508
R8686 VSS.n615 VSS.t242 17.505
R8687 VSS.n645 VSS.t206 17.505
R8688 VSS.n565 VSS.t144 17.505
R8689 VSS.n704 VSS.t660 17.505
R8690 VSS.n676 VSS.t661 17.505
R8691 VSS.n654 VSS.t314 17.505
R8692 VSS.n542 VSS.t656 17.505
R8693 VSS.n585 VSS.t167 17.505
R8694 VSS.n588 VSS.t431 17.505
R8695 VSS.n560 VSS.t411 17.505
R8696 VSS.n548 VSS.t294 17.505
R8697 VSS.n626 VSS.t341 17.505
R8698 VSS.n641 VSS.t344 17.505
R8699 VSS.n670 VSS.t17 17.505
R8700 VSS.n681 VSS.t491 17.505
R8701 VSS.n701 VSS.t603 17.505
R8702 VSS.n573 VSS.t239 17.505
R8703 VSS.n617 VSS.t74 17.505
R8704 VSS.n602 VSS.t409 17.505
R8705 VSS.n528 VSS.t350 17.505
R8706 VSS.n550 VSS.t428 17.505
R8707 VSS.n662 VSS.t280 17.505
R8708 VSS.n689 VSS.t61 17.505
R8709 VSS.n706 VSS.t446 17.505
R8710 VSS.n608 VSS.t180 17.505
R8711 VSS.n553 VSS.t84 17.505
R8712 VSS.n611 VSS.t561 17.505
R8713 VSS.n581 VSS.t427 17.505
R8714 VSS.n522 VSS.t445 17.505
R8715 VSS.n656 VSS.t72 17.505
R8716 VSS.n504 VSS.t662 17.505
R8717 VSS.n715 VSS.t194 17.505
R8718 VSS.n621 VSS.t156 17.505
R8719 VSS.n556 VSS.t81 17.505
R8720 VSS.n578 VSS.t155 17.505
R8721 VSS.n685 VSS.t456 17.505
R8722 VSS.n712 VSS.t395 17.505
R8723 VSS.n659 VSS.t367 17.505
R8724 VSS.n525 VSS.t53 17.505
R8725 VSS.n605 VSS.t64 17.505
R8726 VSS.n538 VSS.t393 17.505
R8727 VSS.n568 VSS.t201 17.505
R8728 VSS.n591 VSS.t582 17.505
R8729 VSS.n633 VSS.t152 17.505
R8730 VSS.n515 VSS.t122 17.505
R8731 VSS.n508 VSS.t349 17.505
R8732 VSS.n498 VSS.t347 17.505
R8733 VSS.n490 VSS.t103 17.505
R8734 VSS.n251 VSS.t490 17.504
R8735 VSS.n200 VSS.t443 17.504
R8736 VSS.n207 VSS.t300 17.504
R8737 VSS.n230 VSS.t466 17.504
R8738 VSS.n236 VSS.t372 17.504
R8739 VSS.n243 VSS.t173 17.504
R8740 VSS.n223 VSS.t532 17.504
R8741 VSS.n216 VSS.t285 17.504
R8742 VSS.n426 VSS.t224 17.4
R8743 VSS.n426 VSS.t274 17.4
R8744 VSS.n364 VSS.t688 17.4
R8745 VSS.n364 VSS.t302 17.4
R8746 VSS.n312 VSS.t170 17.4
R8747 VSS.n312 VSS.t479 17.4
R8748 VSS.n263 VSS.t157 17.4
R8749 VSS.n263 VSS.t436 17.4
R8750 VSS.n169 VSS.t261 17.4
R8751 VSS.n169 VSS.t376 17.4
R8752 VSS.n117 VSS.t211 17.4
R8753 VSS.n117 VSS.t12 17.4
R8754 VSS.n434 VSS.t655 17.4
R8755 VSS.n434 VSS.t1 17.4
R8756 VSS.n63 VSS.t465 17.4
R8757 VSS.n63 VSS.t447 17.4
R8758 VSS.n338 VSS.t510 17.4
R8759 VSS.n338 VSS.t426 17.4
R8760 VSS.n291 VSS.t334 17.4
R8761 VSS.n291 VSS.t553 17.4
R8762 VSS.n114 VSS.t579 17.4
R8763 VSS.n114 VSS.t464 17.4
R8764 VSS.n450 VSS.t497 17.4
R8765 VSS.n450 VSS.t634 17.4
R8766 VSS.n386 VSS.t507 17.4
R8767 VSS.n386 VSS.t422 17.4
R8768 VSS.n275 VSS.t712 17.4
R8769 VSS.n275 VSS.t299 17.4
R8770 VSS.n382 VSS.t179 17.4
R8771 VSS.n382 VSS.t117 17.4
R8772 VSS.n374 VSS.t563 17.4
R8773 VSS.n374 VSS.t549 17.4
R8774 VSS.n446 VSS.t570 17.4
R8775 VSS.n446 VSS.t8 17.4
R8776 VSS.n439 VSS.t346 17.4
R8777 VSS.n439 VSS.t188 17.4
R8778 VSS.n334 VSS.t265 17.4
R8779 VSS.n334 VSS.t439 17.4
R8780 VSS.n322 VSS.t670 17.4
R8781 VSS.n322 VSS.t421 17.4
R8782 VSS.n286 VSS.t410 17.4
R8783 VSS.n286 VSS.t484 17.4
R8784 VSS.n268 VSS.t560 17.4
R8785 VSS.n268 VSS.t55 17.4
R8786 VSS.n598 VSS.t219 17.4
R8787 VSS.n598 VSS.t51 17.4
R8788 VSS.n595 VSS.t648 17.4
R8789 VSS.n595 VSS.t543 17.4
R8790 VSS.n576 VSS.t150 17.4
R8791 VSS.n576 VSS.t3 17.4
R8792 VSS.n600 VSS.t418 17.4
R8793 VSS.n600 VSS.t675 17.4
R8794 VSS.n562 VSS.t77 17.4
R8795 VSS.n562 VSS.t4 17.4
R8796 VSS.n535 VSS.t357 17.4
R8797 VSS.n535 VSS.t521 17.4
R8798 VSS.n531 VSS.t390 17.4
R8799 VSS.n531 VSS.t114 17.4
R8800 VSS.n649 VSS.t386 17.4
R8801 VSS.n649 VSS.t36 17.4
R8802 VSS.n61 VSS.t106 17.4
R8803 VSS.n61 VSS.t183 17.4
R8804 VSS.n329 VSS.t657 17.4
R8805 VSS.n329 VSS.t71 17.4
R8806 VSS.n314 VSS.t44 17.4
R8807 VSS.n314 VSS.t441 17.4
R8808 VSS.n162 VSS.t163 17.4
R8809 VSS.n162 VSS.t283 17.4
R8810 VSS.n27 VSS.t519 17.4
R8811 VSS.n27 VSS.t574 17.4
R8812 VSS.n431 VSS.t658 17.4
R8813 VSS.n431 VSS.t304 17.4
R8814 VSS.n366 VSS.t284 17.4
R8815 VSS.n366 VSS.t577 17.4
R8816 VSS.n280 VSS.t525 17.4
R8817 VSS.n280 VSS.t172 17.4
R8818 VSS.n359 VSS.t407 17.4
R8819 VSS.n359 VSS.t572 17.4
R8820 VSS.n421 VSS.t60 17.4
R8821 VSS.n421 VSS.t588 17.4
R8822 VSS.n464 VSS.t309 9.568
R8823 VSS.n396 VSS.t653 9.568
R8824 VSS.n95 VSS.t15 9.568
R8825 VSS.n153 VSS.t277 9.568
R8826 VSS.n17 VSS.t35 9.568
R8827 VSS.n50 VSS.t646 9.568
R8828 VSS.n90 VSS.t198 9.568
R8829 VSS.n132 VSS.t85 9.568
R8830 VSS.n407 VSS.t645 9.568
R8831 VSS.n108 VSS.t199 9.568
R8832 VSS.n131 VSS.t693 9.568
R8833 VSS.n471 VSS.t34 9.568
R8834 VSS.n11 VSS.t359 9.568
R8835 VSS.n44 VSS.t40 9.568
R8836 VSS.n84 VSS.t177 9.568
R8837 VSS.n142 VSS.t457 9.568
R8838 VSS.n460 VSS.t593 9.568
R8839 VSS.n78 VSS.t148 9.568
R8840 VSS.n148 VSS.t705 9.568
R8841 VSS.n38 VSS.t26 9.568
R8842 VSS.n102 VSS.t147 9.568
R8843 VSS.n469 VSS.t592 9.568
R8844 VSS.n136 VSS.t704 9.568
R8845 VSS.n402 VSS.t28 9.568
R8846 VSS.n284 VSS.t131 9.487
R8847 VSS.n332 VSS.t59 9.487
R8848 VSS.n379 VSS.t413 9.487
R8849 VSS.n423 VSS.t247 9.487
R8850 VSS.n361 VSS.t528 9.487
R8851 VSS.n120 VSS.t480 9.487
R8852 VSS.n179 VSS.t161 9.487
R8853 VSS.n358 VSS.t500 9.487
R8854 VSS.n121 VSS.t380 9.487
R8855 VSS.n180 VSS.t94 9.487
R8856 VSS.n420 VSS.t499 9.487
R8857 VSS.n357 VSS.t501 9.487
R8858 VSS.n299 VSS.t379 9.487
R8859 VSS.n178 VSS.t399 9.487
R8860 VSS.n25 VSS.t378 9.487
R8861 VSS.n60 VSS.t449 9.487
R8862 VSS.n328 VSS.t166 9.487
R8863 VSS.n283 VSS.t312 9.487
R8864 VSS.n327 VSS.t58 9.487
R8865 VSS.n282 VSS.t130 9.487
R8866 VSS.n59 VSS.t43 9.487
R8867 VSS.n26 VSS.t237 9.487
R8868 VSS.n444 VSS.t238 9.487
R8869 VSS.n36 VSS.t605 9.46
R8870 VSS.n546 VSS.t243 9.43
R8871 VSS.n652 VSS.t215 9.43
R8872 VSS.n262 VSS.t252 9.319
R8873 VSS.n193 VSS.t554 9.319
R8874 VSS.n260 VSS.t217 9.319
R8875 VSS.n478 VSS.t231 9.319
R8876 VSS.n477 VSS.t269 9.319
R8877 VSS.n194 VSS.t62 9.319
R8878 VSS.n261 VSS.t250 9.319
R8879 VSS.n257 VSS.t387 9.319
R8880 VSS.n195 VSS.t83 9.319
R8881 VSS.n9 VSS.t330 9.319
R8882 VSS.n258 VSS.t291 9.319
R8883 VSS.n8 VSS.t268 9.319
R8884 VSS.n196 VSS.t576 9.319
R8885 VSS.n424 VSS.t487 9.319
R8886 VSS.n362 VSS.t292 9.319
R8887 VSS.n259 VSS.t257 9.319
R8888 VSS.n300 VSS.t220 9.319
R8889 VSS.n665 VSS.t297 9.319
R8890 VSS.n674 VSS.t301 9.319
R8891 VSS.n503 VSS.t594 9.319
R8892 VSS.n668 VSS.t289 9.319
R8893 VSS.n696 VSS.t389 9.319
R8894 VSS.n709 VSS.t356 9.319
R8895 VSS.n119 VSS.t551 9.317
R8896 VSS.n363 VSS.t488 9.317
R8897 VSS.n425 VSS.t49 9.317
R8898 VSS.n615 VSS.t375 8.702
R8899 VSS.n614 VSS.t437 8.702
R8900 VSS.n645 VSS.t440 8.702
R8901 VSS.n644 VSS.t50 8.702
R8902 VSS.n565 VSS.t19 8.702
R8903 VSS.n564 VSS.t263 8.702
R8904 VSS.n704 VSS.t697 8.702
R8905 VSS.n703 VSS.t531 8.702
R8906 VSS.n676 VSS.t102 8.702
R8907 VSS.n675 VSS.t460 8.702
R8908 VSS.n654 VSS.t666 8.702
R8909 VSS.n653 VSS.t408 8.702
R8910 VSS.n542 VSS.t669 8.702
R8911 VSS.n541 VSS.t23 8.702
R8912 VSS.n585 VSS.t508 8.702
R8913 VSS.n584 VSS.t339 8.702
R8914 VSS.n588 VSS.t468 8.702
R8915 VSS.n587 VSS.t327 8.702
R8916 VSS.n560 VSS.t135 8.702
R8917 VSS.n559 VSS.t54 8.702
R8918 VSS.n548 VSS.t430 8.702
R8919 VSS.n547 VSS.t364 8.702
R8920 VSS.n626 VSS.t98 8.702
R8921 VSS.n625 VSS.t101 8.702
R8922 VSS.n641 VSS.t548 8.702
R8923 VSS.n640 VSS.t244 8.702
R8924 VSS.n670 VSS.t567 8.702
R8925 VSS.n669 VSS.t82 8.702
R8926 VSS.n681 VSS.t589 8.702
R8927 VSS.n680 VSS.t202 8.702
R8928 VSS.n701 VSS.t686 8.702
R8929 VSS.n700 VSS.t511 8.702
R8930 VSS.n574 VSS.t337 8.702
R8931 VSS.n573 VSS.t524 8.702
R8932 VSS.n618 VSS.t279 8.702
R8933 VSS.n617 VSS.t86 8.702
R8934 VSS.n603 VSS.t10 8.702
R8935 VSS.n602 VSS.t702 8.702
R8936 VSS.n529 VSS.t181 8.702
R8937 VSS.n528 VSS.t316 8.702
R8938 VSS.n551 VSS.t691 8.702
R8939 VSS.n550 VSS.t665 8.702
R8940 VSS.n663 VSS.t275 8.702
R8941 VSS.n662 VSS.t209 8.702
R8942 VSS.n690 VSS.t113 8.702
R8943 VSS.n689 VSS.t343 8.702
R8944 VSS.n707 VSS.t438 8.702
R8945 VSS.n706 VSS.t108 8.702
R8946 VSS.n609 VSS.t361 8.702
R8947 VSS.n608 VSS.t25 8.702
R8948 VSS.n554 VSS.t313 8.702
R8949 VSS.n553 VSS.t623 8.702
R8950 VSS.n612 VSS.t396 8.702
R8951 VSS.n611 VSS.t88 8.702
R8952 VSS.n582 VSS.t698 8.702
R8953 VSS.n581 VSS.t345 8.702
R8954 VSS.n523 VSS.t315 8.702
R8955 VSS.n522 VSS.t63 8.702
R8956 VSS.n657 VSS.t587 8.702
R8957 VSS.n656 VSS.t89 8.702
R8958 VSS.n505 VSS.t7 8.702
R8959 VSS.n504 VSS.t384 8.702
R8960 VSS.n716 VSS.t91 8.702
R8961 VSS.n715 VSS.t711 8.702
R8962 VSS.n622 VSS.t65 8.702
R8963 VSS.n621 VSS.t394 8.702
R8964 VSS.n557 VSS.t550 8.702
R8965 VSS.n556 VSS.t602 8.702
R8966 VSS.n579 VSS.t542 8.702
R8967 VSS.n578 VSS.t32 8.702
R8968 VSS.n686 VSS.t442 8.702
R8969 VSS.n685 VSS.t66 8.702
R8970 VSS.n713 VSS.t696 8.702
R8971 VSS.n712 VSS.t191 8.702
R8972 VSS.n660 VSS.t79 8.702
R8973 VSS.n659 VSS.t318 8.702
R8974 VSS.n526 VSS.t534 8.702
R8975 VSS.n525 VSS.t73 8.702
R8976 VSS.n606 VSS.t335 8.702
R8977 VSS.n605 VSS.t168 8.702
R8978 VSS.n537 VSS.t332 8.702
R8979 VSS.n538 VSS.t259 8.702
R8980 VSS.n567 VSS.t228 8.702
R8981 VSS.n568 VSS.t320 8.702
R8982 VSS.n590 VSS.t600 8.702
R8983 VSS.n591 VSS.t329 8.702
R8984 VSS.n632 VSS.t402 8.702
R8985 VSS.n633 VSS.t225 8.702
R8986 VSS.n514 VSS.t47 8.702
R8987 VSS.n515 VSS.t631 8.702
R8988 VSS.n507 VSS.t256 8.702
R8989 VSS.n508 VSS.t547 8.702
R8990 VSS.n499 VSS.t626 8.702
R8991 VSS.n498 VSS.t365 8.702
R8992 VSS.n491 VSS.t306 8.702
R8993 VSS.n490 VSS.t404 8.702
R8994 VSS.n251 VSS.t100 8.702
R8995 VSS.n200 VSS.t112 8.702
R8996 VSS.n207 VSS.t118 8.702
R8997 VSS.n230 VSS.t186 8.702
R8998 VSS.n236 VSS.t429 8.702
R8999 VSS.n243 VSS.t21 8.702
R9000 VSS.n223 VSS.t203 8.702
R9001 VSS.n216 VSS.t433 8.702
R9002 VSS.n250 VSS.t530 8.702
R9003 VSS.n199 VSS.t97 8.702
R9004 VSS.n206 VSS.t92 8.702
R9005 VSS.n229 VSS.t434 8.702
R9006 VSS.n235 VSS.t615 8.702
R9007 VSS.n242 VSS.t80 8.702
R9008 VSS.n222 VSS.t451 8.702
R9009 VSS.n215 VSS.t462 8.702
R9010 VSS.n184 VSS.t264 8.7
R9011 VSS.n184 VSS.t664 8.7
R9012 VSS.n452 VSS.t700 8.7
R9013 VSS.n452 VSS.t435 8.7
R9014 VSS.n30 VSS.t56 8.7
R9015 VSS.n30 VSS.t310 8.7
R9016 VSS.n388 VSS.t273 8.7
R9017 VSS.n388 VSS.t272 8.7
R9018 VSS.n66 VSS.t471 8.7
R9019 VSS.n66 VSS.t652 8.7
R9020 VSS.n343 VSS.t695 8.7
R9021 VSS.n343 VSS.t133 8.7
R9022 VSS.n304 VSS.t0 8.7
R9023 VSS.n304 VSS.t235 8.7
R9024 VSS.n174 VSS.t286 8.7
R9025 VSS.n174 VSS.t278 8.7
R9026 VSS.n159 VSS.t6 8.7
R9027 VSS.n159 VSS.t110 8.7
R9028 VSS.n191 VSS.t90 8.7
R9029 VSS.n191 VSS.t709 8.7
R9030 VSS.n666 VSS.t383 8.7
R9031 VSS.n666 VSS.t340 8.7
R9032 VSS.n533 VSS.t529 8.7
R9033 VSS.n533 VSS.t24 8.7
R9034 VSS.n544 VSS.t290 8.7
R9035 VSS.n544 VSS.t578 8.7
R9036 VSS.n520 VSS.t298 8.7
R9037 VSS.n520 VSS.t52 8.7
R9038 VSS.n710 VSS.t354 8.7
R9039 VSS.n710 VSS.t232 8.7
R9040 VSS.n693 VSS.t651 8.7
R9041 VSS.n693 VSS.t189 8.7
R9042 VSS.n678 VSS.t595 8.7
R9043 VSS.n678 VSS.t544 8.7
R9044 VSS.n571 VSS.t416 8.7
R9045 VSS.n571 VSS.t520 8.7
R9046 VSS.n346 VSS.t406 8.7
R9047 VSS.n346 VSS.t362 8.7
R9048 VSS.n301 VSS.t326 8.7
R9049 VSS.n301 VSS.t178 8.7
R9050 VSS.n56 VSS.t57 8.7
R9051 VSS.n56 VSS.t569 8.7
R9052 VSS.n74 VSS.t644 8.7
R9053 VSS.n74 VSS.t45 8.7
R9054 VSS.n33 VSS.t159 8.7
R9055 VSS.n33 VSS.t270 8.7
R9056 VSS.n22 VSS.t673 8.7
R9057 VSS.n22 VSS.t153 8.7
R9058 VSS.n189 VSS.t325 8.7
R9059 VSS.n189 VSS.t192 8.7
R9060 VSS.n171 VSS.t505 8.7
R9061 VSS.n171 VSS.t458 8.7
R9062 VSS.n295 VSS.t39 8.7
R9063 VSS.n295 VSS.t115 8.7
R9064 VSS.n187 VSS.t454 8.7
R9065 VSS.n187 VSS.t699 8.7
R9066 VSS.n316 VSS.t552 8.7
R9067 VSS.n316 VSS.t616 8.7
R9068 VSS.n340 VSS.t482 8.7
R9069 VSS.n340 VSS.t566 8.7
R9070 VSS.n455 VSS.t248 8.7
R9071 VSS.n455 VSS.t104 8.7
R9072 VSS.n428 VSS.t598 8.7
R9073 VSS.n428 VSS.t187 8.7
R9074 VSS.n391 VSS.t526 8.7
R9075 VSS.n391 VSS.t37 8.7
R9076 VSS.n368 VSS.t226 8.7
R9077 VSS.n368 VSS.t33 8.7
R9078 VSS.n128 VSS.t162 8.7
R9079 VSS.n128 VSS.t710 8.7
R9080 VSS.n270 VSS.t323 8.7
R9081 VSS.n270 VSS.t624 8.7
R9082 VSS.n417 VSS.t171 8.7
R9083 VSS.n417 VSS.t637 8.7
R9084 VSS.n414 VSS.t342 8.7
R9085 VSS.n414 VSS.t371 8.7
R9086 VSS.n351 VSS.t109 8.7
R9087 VSS.n351 VSS.t448 8.7
R9088 VSS.n354 VSS.t207 8.7
R9089 VSS.n354 VSS.t31 8.7
R9090 VSS.n125 VSS.t11 8.7
R9091 VSS.n125 VSS.t164 8.7
R9092 VSS.n122 VSS.t478 8.7
R9093 VSS.n122 VSS.t629 8.7
R9094 VSS.n181 VSS.t324 8.7
R9095 VSS.n181 VSS.t311 8.7
R9096 VSS.n265 VSS.t571 8.7
R9097 VSS.n265 VSS.t258 8.7
R9098 VSS.n4 VSS.t288 8.7
R9099 VSS.n4 VSS.t584 8.7
R9100 VSS.n2 VSS.t295 8.7
R9101 VSS.n2 VSS.t190 8.7
R9102 VSS.n480 VSS.t221 8.7
R9103 VSS.n480 VSS.t9 8.7
R9104 VSS.n0 VSS.t76 8.7
R9105 VSS.n0 VSS.t222 8.7
R9106 VSS.n487 VSS.t391 8.7
R9107 VSS.n487 VSS.t348 8.7
R9108 VSS.n483 VSS.t352 8.7
R9109 VSS.n483 VSS.t620 8.7
R9110 VSS.n720 VSS.t417 8.7
R9111 VSS.n720 VSS.t649 8.7
R9112 VSS.n6 VSS.t425 8.7
R9113 VSS.n6 VSS.t400 8.7
R9114 VSS.n539 VSS.n537 2.136
R9115 VSS.n569 VSS.n567 2.136
R9116 VSS.n592 VSS.n590 2.136
R9117 VSS.n634 VSS.n632 2.136
R9118 VSS.n516 VSS.n514 2.136
R9119 VSS.n509 VSS.n507 2.136
R9120 VSS.n638 VSS.n637 2.098
R9121 VSS.n539 VSS.n538 2.063
R9122 VSS.n569 VSS.n568 2.063
R9123 VSS.n592 VSS.n591 2.063
R9124 VSS.n634 VSS.n633 2.063
R9125 VSS.n516 VSS.n515 2.063
R9126 VSS.n509 VSS.n508 2.063
R9127 VSS.n616 VSS.n614 2.025
R9128 VSS.n646 VSS.n644 2.025
R9129 VSS.n566 VSS.n564 2.025
R9130 VSS.n705 VSS.n703 2.025
R9131 VSS.n677 VSS.n675 2.025
R9132 VSS.n655 VSS.n653 2.025
R9133 VSS.n543 VSS.n541 2.025
R9134 VSS.n586 VSS.n584 2.025
R9135 VSS.n589 VSS.n587 2.025
R9136 VSS.n561 VSS.n559 2.025
R9137 VSS.n549 VSS.n547 2.025
R9138 VSS.n627 VSS.n625 2.025
R9139 VSS.n642 VSS.n640 2.025
R9140 VSS.n671 VSS.n669 2.025
R9141 VSS.n682 VSS.n680 2.025
R9142 VSS.n702 VSS.n700 2.025
R9143 VSS.n575 VSS.n574 2.025
R9144 VSS.n619 VSS.n618 2.025
R9145 VSS.n604 VSS.n603 2.025
R9146 VSS.n530 VSS.n529 2.025
R9147 VSS.n552 VSS.n551 2.025
R9148 VSS.n664 VSS.n663 2.025
R9149 VSS.n691 VSS.n690 2.025
R9150 VSS.n708 VSS.n707 2.025
R9151 VSS.n610 VSS.n609 2.025
R9152 VSS.n555 VSS.n554 2.025
R9153 VSS.n613 VSS.n612 2.025
R9154 VSS.n583 VSS.n582 2.025
R9155 VSS.n524 VSS.n523 2.025
R9156 VSS.n658 VSS.n657 2.025
R9157 VSS.n506 VSS.n505 2.025
R9158 VSS.n717 VSS.n716 2.025
R9159 VSS.n623 VSS.n622 2.025
R9160 VSS.n558 VSS.n557 2.025
R9161 VSS.n580 VSS.n579 2.025
R9162 VSS.n687 VSS.n686 2.025
R9163 VSS.n714 VSS.n713 2.025
R9164 VSS.n661 VSS.n660 2.025
R9165 VSS.n527 VSS.n526 2.025
R9166 VSS.n607 VSS.n606 2.025
R9167 VSS.n500 VSS.n499 2.025
R9168 VSS.n492 VSS.n491 2.025
R9169 VSS.n252 VSS.n250 2.025
R9170 VSS.n201 VSS.n199 2.025
R9171 VSS.n208 VSS.n206 2.025
R9172 VSS.n231 VSS.n229 2.025
R9173 VSS.n237 VSS.n235 2.025
R9174 VSS.n244 VSS.n242 2.025
R9175 VSS.n224 VSS.n222 2.025
R9176 VSS.n217 VSS.n215 2.025
R9177 VSS.n616 VSS.n615 1.953
R9178 VSS.n646 VSS.n645 1.953
R9179 VSS.n566 VSS.n565 1.953
R9180 VSS.n705 VSS.n704 1.953
R9181 VSS.n677 VSS.n676 1.953
R9182 VSS.n655 VSS.n654 1.953
R9183 VSS.n543 VSS.n542 1.953
R9184 VSS.n586 VSS.n585 1.953
R9185 VSS.n589 VSS.n588 1.953
R9186 VSS.n561 VSS.n560 1.953
R9187 VSS.n549 VSS.n548 1.953
R9188 VSS.n627 VSS.n626 1.953
R9189 VSS.n642 VSS.n641 1.953
R9190 VSS.n671 VSS.n670 1.953
R9191 VSS.n682 VSS.n681 1.953
R9192 VSS.n702 VSS.n701 1.953
R9193 VSS.n575 VSS.n573 1.953
R9194 VSS.n619 VSS.n617 1.953
R9195 VSS.n604 VSS.n602 1.953
R9196 VSS.n530 VSS.n528 1.953
R9197 VSS.n552 VSS.n550 1.953
R9198 VSS.n664 VSS.n662 1.953
R9199 VSS.n691 VSS.n689 1.953
R9200 VSS.n708 VSS.n706 1.953
R9201 VSS.n610 VSS.n608 1.953
R9202 VSS.n555 VSS.n553 1.953
R9203 VSS.n613 VSS.n611 1.953
R9204 VSS.n583 VSS.n581 1.953
R9205 VSS.n524 VSS.n522 1.953
R9206 VSS.n658 VSS.n656 1.953
R9207 VSS.n506 VSS.n504 1.953
R9208 VSS.n717 VSS.n715 1.953
R9209 VSS.n623 VSS.n621 1.953
R9210 VSS.n558 VSS.n556 1.953
R9211 VSS.n580 VSS.n578 1.953
R9212 VSS.n687 VSS.n685 1.953
R9213 VSS.n714 VSS.n712 1.953
R9214 VSS.n661 VSS.n659 1.953
R9215 VSS.n527 VSS.n525 1.953
R9216 VSS.n607 VSS.n605 1.953
R9217 VSS.n500 VSS.n498 1.953
R9218 VSS.n492 VSS.n490 1.953
R9219 VSS.n252 VSS.n251 1.953
R9220 VSS.n201 VSS.n200 1.953
R9221 VSS.n208 VSS.n207 1.953
R9222 VSS.n231 VSS.n230 1.953
R9223 VSS.n237 VSS.n236 1.953
R9224 VSS.n244 VSS.n243 1.953
R9225 VSS.n224 VSS.n223 1.953
R9226 VSS.n217 VSS.n216 1.953
R9227 VSS.n453 VSS.n452 0.948
R9228 VSS.n31 VSS.n30 0.948
R9229 VSS.n389 VSS.n388 0.948
R9230 VSS.n67 VSS.n66 0.948
R9231 VSS.n344 VSS.n343 0.948
R9232 VSS.n305 VSS.n304 0.948
R9233 VSS.n175 VSS.n174 0.948
R9234 VSS.n160 VSS.n159 0.948
R9235 VSS.n667 VSS.n666 0.948
R9236 VSS.n534 VSS.n533 0.948
R9237 VSS.n545 VSS.n544 0.948
R9238 VSS.n521 VSS.n520 0.948
R9239 VSS.n711 VSS.n710 0.948
R9240 VSS.n694 VSS.n693 0.948
R9241 VSS.n679 VSS.n678 0.948
R9242 VSS.n572 VSS.n571 0.948
R9243 VSS.n347 VSS.n346 0.948
R9244 VSS.n302 VSS.n301 0.948
R9245 VSS.n57 VSS.n56 0.948
R9246 VSS.n75 VSS.n74 0.948
R9247 VSS.n34 VSS.n33 0.948
R9248 VSS.n23 VSS.n22 0.948
R9249 VSS.n172 VSS.n171 0.948
R9250 VSS.n296 VSS.n295 0.948
R9251 VSS.n317 VSS.n316 0.948
R9252 VSS.n341 VSS.n340 0.948
R9253 VSS.n456 VSS.n455 0.948
R9254 VSS.n429 VSS.n428 0.948
R9255 VSS.n392 VSS.n391 0.948
R9256 VSS.n369 VSS.n368 0.948
R9257 VSS.n129 VSS.n128 0.948
R9258 VSS.n271 VSS.n270 0.948
R9259 VSS.n418 VSS.n417 0.948
R9260 VSS.n415 VSS.n414 0.948
R9261 VSS.n352 VSS.n351 0.948
R9262 VSS.n355 VSS.n354 0.948
R9263 VSS.n126 VSS.n125 0.948
R9264 VSS.n123 VSS.n122 0.948
R9265 VSS.n182 VSS.n181 0.948
R9266 VSS.n266 VSS.n265 0.948
R9267 VSS.n5 VSS.n4 0.948
R9268 VSS.n3 VSS.n2 0.948
R9269 VSS.n481 VSS.n480 0.948
R9270 VSS.n1 VSS.n0 0.948
R9271 VSS.n488 VSS.n487 0.948
R9272 VSS.n484 VSS.n483 0.948
R9273 VSS.n721 VSS.n720 0.948
R9274 VSS.n7 VSS.n6 0.948
R9275 VSS.n185 VSS.n184 0.889
R9276 VSS.n192 VSS.n191 0.889
R9277 VSS.n190 VSS.n189 0.889
R9278 VSS.n188 VSS.n187 0.889
R9279 VSS.n315 VSS.n314 0.795
R9280 VSS.n367 VSS.n366 0.795
R9281 VSS.n281 VSS.n280 0.795
R9282 VSS.n62 VSS.n61 0.791
R9283 VSS.n330 VSS.n329 0.791
R9284 VSS.n163 VSS.n162 0.791
R9285 VSS.n427 VSS.n426 0.72
R9286 VSS.n365 VSS.n364 0.72
R9287 VSS.n313 VSS.n312 0.72
R9288 VSS.n264 VSS.n263 0.72
R9289 VSS.n170 VSS.n169 0.72
R9290 VSS.n118 VSS.n117 0.72
R9291 VSS.n435 VSS.n434 0.72
R9292 VSS.n64 VSS.n63 0.72
R9293 VSS.n339 VSS.n338 0.72
R9294 VSS.n292 VSS.n291 0.72
R9295 VSS.n115 VSS.n114 0.72
R9296 VSS.n451 VSS.n450 0.72
R9297 VSS.n387 VSS.n386 0.72
R9298 VSS.n276 VSS.n275 0.72
R9299 VSS.n383 VSS.n382 0.72
R9300 VSS.n375 VSS.n374 0.72
R9301 VSS.n447 VSS.n446 0.72
R9302 VSS.n440 VSS.n439 0.72
R9303 VSS.n335 VSS.n334 0.72
R9304 VSS.n323 VSS.n322 0.72
R9305 VSS.n287 VSS.n286 0.72
R9306 VSS.n269 VSS.n268 0.72
R9307 VSS.n28 VSS.n27 0.72
R9308 VSS.n432 VSS.n431 0.72
R9309 VSS.n360 VSS.n359 0.72
R9310 VSS.n422 VSS.n421 0.72
R9311 VSS.n599 VSS.n598 0.533
R9312 VSS.n601 VSS.n600 0.533
R9313 VSS.n563 VSS.n562 0.533
R9314 VSS.n532 VSS.n531 0.533
R9315 VSS.n650 VSS.n649 0.533
R9316 VSS.n596 VSS.n595 0.526
R9317 VSS.n577 VSS.n576 0.526
R9318 VSS.n536 VSS.n535 0.526
R9319 VSS.n672 VSS.n665 0.313
R9320 VSS.n639 VSS.n638 0.311
R9321 VSS.n697 VSS.n696 0.311
R9322 VSS.n319 VSS.n119 0.311
R9323 VSS.n371 VSS.n363 0.311
R9324 VSS.n433 VSS.n425 0.311
R9325 VSS.n683 VSS.n674 0.309
R9326 VSS.n695 VSS.n503 0.309
R9327 VSS.n672 VSS.n668 0.309
R9328 VSS.n718 VSS.n709 0.309
R9329 VSS.n274 VSS.n262 0.309
R9330 VSS.n255 VSS.n193 0.309
R9331 VSS.n274 VSS.n260 0.309
R9332 VSS.n479 VSS.n478 0.309
R9333 VSS.n479 VSS.n477 0.309
R9334 VSS.n255 VSS.n194 0.309
R9335 VSS.n274 VSS.n261 0.309
R9336 VSS.n274 VSS.n257 0.309
R9337 VSS.n255 VSS.n195 0.309
R9338 VSS.n479 VSS.n9 0.309
R9339 VSS.n479 VSS.n8 0.309
R9340 VSS.n255 VSS.n196 0.309
R9341 VSS.n433 VSS.n424 0.309
R9342 VSS.n371 VSS.n362 0.309
R9343 VSS.n274 VSS.n259 0.309
R9344 VSS.n319 VSS.n300 0.309
R9345 VSS.n274 VSS.n258 0.259
R9346 VSS.n433 VSS.n36 0.239
R9347 VSS.n651 VSS.n546 0.225
R9348 VSS.n672 VSS.n652 0.225
R9349 VSS VSS.n1 0.198
R9350 VSS VSS.n7 0.198
R9351 VSS VSS.n481 0.198
R9352 VSS VSS.n3 0.198
R9353 VSS VSS.n5 0.198
R9354 VSS.n672 VSS.n667 0.197
R9355 VSS.n651 VSS.n545 0.197
R9356 VSS.n672 VSS.n521 0.197
R9357 VSS.n718 VSS.n711 0.197
R9358 VSS.n695 VSS.n694 0.197
R9359 VSS.n683 VSS.n679 0.197
R9360 VSS.n651 VSS.n572 0.197
R9361 VSS.n651 VSS.n534 0.197
R9362 VSS.n489 VSS.n488 0.196
R9363 VSS.n485 VSS.n484 0.196
R9364 VSS.n722 VSS.n721 0.196
R9365 VSS.n651 VSS.n532 0.173
R9366 VSS.n648 VSS.n599 0.172
R9367 VSS.n648 VSS.n596 0.172
R9368 VSS.n648 VSS.n577 0.172
R9369 VSS.n648 VSS.n601 0.172
R9370 VSS.n651 VSS.n563 0.172
R9371 VSS.n651 VSS.n536 0.172
R9372 VSS.n651 VSS.n650 0.172
R9373 VSS.n319 VSS.n124 0.151
R9374 VSS.n433 VSS.n416 0.151
R9375 VSS.n371 VSS.n356 0.15
R9376 VSS.n177 VSS.n176 0.147
R9377 VSS.n433 VSS.n32 0.146
R9378 VSS.n69 VSS.n68 0.146
R9379 VSS.n307 VSS.n306 0.146
R9380 VSS.n319 VSS.n303 0.146
R9381 VSS.n371 VSS.n76 0.146
R9382 VSS.n433 VSS.n35 0.146
R9383 VSS.n274 VSS.n173 0.146
R9384 VSS.n319 VSS.n318 0.146
R9385 VSS.n350 VSS.n342 0.146
R9386 VSS.n476 VSS.n457 0.146
R9387 VSS.n433 VSS.n430 0.146
R9388 VSS.n413 VSS.n393 0.146
R9389 VSS.n371 VSS.n370 0.146
R9390 VSS.n298 VSS.n130 0.146
R9391 VSS.n274 VSS.n272 0.146
R9392 VSS.n433 VSS.n419 0.146
R9393 VSS.n371 VSS.n353 0.146
R9394 VSS.n319 VSS.n127 0.146
R9395 VSS.n274 VSS.n183 0.146
R9396 VSS.n274 VSS.n267 0.146
R9397 VSS.n274 VSS.n269 0.143
R9398 VSS.n274 VSS.n170 0.142
R9399 VSS.n319 VSS.n118 0.142
R9400 VSS.n476 VSS.n454 0.142
R9401 VSS.n413 VSS.n390 0.142
R9402 VSS.n350 VSS.n345 0.142
R9403 VSS.n413 VSS.n58 0.142
R9404 VSS.n298 VSS.n297 0.142
R9405 VSS.n445 VSS.n28 0.142
R9406 VSS.n371 VSS.n360 0.142
R9407 VSS.n433 VSS.n422 0.142
R9408 VSS.n65 VSS.n64 0.141
R9409 VSS.n350 VSS.n348 0.141
R9410 VSS.n298 VSS.n161 0.14
R9411 VSS.n476 VSS.n24 0.14
R9412 VSS.n433 VSS.n427 0.138
R9413 VSS.n371 VSS.n365 0.138
R9414 VSS.n319 VSS.n313 0.138
R9415 VSS.n274 VSS.n264 0.138
R9416 VSS.n436 VSS.n435 0.138
R9417 VSS.n433 VSS.n432 0.138
R9418 VSS.n277 VSS.n276 0.137
R9419 VSS.n376 VSS.n375 0.137
R9420 VSS.n413 VSS.n387 0.136
R9421 VSS.n441 VSS.n440 0.136
R9422 VSS.n476 VSS.n451 0.135
R9423 VSS.n288 VSS.n287 0.135
R9424 VSS.n350 VSS.n339 0.134
R9425 VSS.n116 VSS.n115 0.133
R9426 VSS.n448 VSS.n447 0.133
R9427 VSS.n324 VSS.n323 0.133
R9428 VSS.n336 VSS.n335 0.131
R9429 VSS.n293 VSS.n292 0.129
R9430 VSS.n384 VSS.n383 0.129
R9431 VSS.n350 VSS.n349 0.127
R9432 VSS.n454 VSS.n453 0.125
R9433 VSS.n32 VSS.n31 0.125
R9434 VSS.n390 VSS.n389 0.125
R9435 VSS.n68 VSS.n67 0.125
R9436 VSS.n345 VSS.n344 0.125
R9437 VSS.n306 VSS.n305 0.125
R9438 VSS.n176 VSS.n175 0.125
R9439 VSS.n161 VSS.n160 0.125
R9440 VSS.n348 VSS.n347 0.125
R9441 VSS.n303 VSS.n302 0.125
R9442 VSS.n58 VSS.n57 0.125
R9443 VSS.n76 VSS.n75 0.125
R9444 VSS.n35 VSS.n34 0.125
R9445 VSS.n24 VSS.n23 0.125
R9446 VSS.n173 VSS.n172 0.125
R9447 VSS.n297 VSS.n296 0.125
R9448 VSS.n318 VSS.n317 0.125
R9449 VSS.n342 VSS.n341 0.125
R9450 VSS.n457 VSS.n456 0.125
R9451 VSS.n430 VSS.n429 0.125
R9452 VSS.n393 VSS.n392 0.125
R9453 VSS.n370 VSS.n369 0.125
R9454 VSS.n130 VSS.n129 0.125
R9455 VSS.n272 VSS.n271 0.125
R9456 VSS.n419 VSS.n418 0.125
R9457 VSS.n416 VSS.n415 0.125
R9458 VSS.n353 VSS.n352 0.125
R9459 VSS.n356 VSS.n355 0.125
R9460 VSS.n127 VSS.n126 0.125
R9461 VSS.n124 VSS.n123 0.125
R9462 VSS.n183 VSS.n182 0.125
R9463 VSS.n267 VSS.n266 0.125
R9464 VSS.n298 VSS.n132 0.119
R9465 VSS.n476 VSS.n460 0.119
R9466 VSS.n96 VSS.n95 0.118
R9467 VSS.n476 VSS.n469 0.118
R9468 VSS.n298 VSS.n131 0.117
R9469 VSS.n109 VSS.n108 0.116
R9470 VSS.n12 VSS.n11 0.116
R9471 VSS.n45 VSS.n44 0.116
R9472 VSS.n85 VSS.n84 0.116
R9473 VSS.n143 VSS.n142 0.115
R9474 VSS.n39 VSS.n38 0.115
R9475 VSS.n51 VSS.n50 0.114
R9476 VSS.n91 VSS.n90 0.114
R9477 VSS.n137 VSS.n136 0.114
R9478 VSS.n465 VSS.n464 0.113
R9479 VSS.n154 VSS.n153 0.113
R9480 VSS.n408 VSS.n407 0.113
R9481 VSS.n472 VSS.n471 0.113
R9482 VSS.n403 VSS.n402 0.113
R9483 VSS.n79 VSS.n78 0.112
R9484 VSS.n397 VSS.n396 0.111
R9485 VSS.n103 VSS.n102 0.111
R9486 VSS.n18 VSS.n17 0.11
R9487 VSS.n149 VSS.n148 0.11
R9488 VSS.n718 VSS.n708 0.102
R9489 VSS.n683 VSS.n677 0.101
R9490 VSS.n648 VSS.n604 0.101
R9491 VSS.n648 VSS.n575 0.101
R9492 VSS.n672 VSS.n664 0.101
R9493 VSS.n651 VSS.n530 0.1
R9494 VSS.n651 VSS.n566 0.099
R9495 VSS.n651 VSS.n543 0.099
R9496 VSS.n651 VSS.n561 0.099
R9497 VSS.n651 VSS.n549 0.099
R9498 VSS.n648 VSS.n610 0.099
R9499 VSS.n651 VSS.n555 0.099
R9500 VSS.n648 VSS.n583 0.099
R9501 VSS.n651 VSS.n524 0.099
R9502 VSS.n672 VSS.n658 0.099
R9503 VSS.n718 VSS.n717 0.099
R9504 VSS.n651 VSS.n558 0.099
R9505 VSS.n718 VSS.n714 0.099
R9506 VSS.n672 VSS.n661 0.099
R9507 VSS.n651 VSS.n527 0.099
R9508 VSS.n684 VSS.n506 0.099
R9509 VSS.n651 VSS.n552 0.099
R9510 VSS.n718 VSS.n705 0.098
R9511 VSS.n672 VSS.n671 0.098
R9512 VSS.n628 VSS.n616 0.098
R9513 VSS.n672 VSS.n655 0.098
R9514 VSS.n718 VSS.n702 0.098
R9515 VSS.n648 VSS.n580 0.098
R9516 VSS.n648 VSS.n607 0.098
R9517 VSS.n628 VSS.n627 0.098
R9518 VSS.n648 VSS.n589 0.098
R9519 VSS.n648 VSS.n586 0.098
R9520 VSS.n683 VSS.n682 0.098
R9521 VSS.n688 VSS.n687 0.098
R9522 VSS.n643 VSS.n642 0.097
R9523 VSS.n629 VSS.n613 0.097
R9524 VSS.n620 VSS.n619 0.097
R9525 VSS.n624 VSS.n623 0.097
R9526 VSS.n647 VSS.n646 0.097
R9527 VSS.n692 VSS.n691 0.097
R9528 VSS.n253 VSS.n252 0.095
R9529 VSS.n202 VSS.n201 0.095
R9530 VSS.n209 VSS.n208 0.095
R9531 VSS.n232 VSS.n231 0.095
R9532 VSS.n238 VSS.n237 0.095
R9533 VSS.n245 VSS.n244 0.095
R9534 VSS.n225 VSS.n224 0.095
R9535 VSS.n501 VSS.n500 0.095
R9536 VSS.n493 VSS.n492 0.095
R9537 VSS.n218 VSS.n217 0.095
R9538 VSS.n635 VSS.n634 0.063
R9539 VSS.n570 VSS.n569 0.063
R9540 VSS.n540 VSS.n539 0.062
R9541 VSS.n256 VSS.n192 0.062
R9542 VSS.n256 VSS.n190 0.062
R9543 VSS.n256 VSS.n188 0.062
R9544 VSS.n186 VSS.n185 0.061
R9545 VSS.n593 VSS.n592 0.06
R9546 VSS.n517 VSS.n516 0.06
R9547 VSS.n510 VSS.n509 0.06
R9548 VSS.n381 VSS.n62 0.044
R9549 VSS.n333 VSS.n330 0.044
R9550 VSS.n319 VSS.n315 0.044
R9551 VSS.n298 VSS.n163 0.044
R9552 VSS.n371 VSS.n367 0.044
R9553 VSS.n285 VSS.n281 0.044
R9554 VSS.n465 VSS.n463 0.04
R9555 VSS.n137 VSS.n135 0.04
R9556 VSS.n699 VSS.n698 0.029
R9557 VSS.n512 VSS.n511 0.029
R9558 VSS.n476 VSS.n459 0.022
R9559 VSS.n274 VSS.n273 0.022
R9560 VSS.n319 VSS.n120 0.021
R9561 VSS.n433 VSS.n423 0.02
R9562 VSS.n371 VSS.n361 0.02
R9563 VSS.n399 VSS.n398 0.018
R9564 VSS.n99 VSS.n98 0.018
R9565 VSS.n411 VSS.n410 0.018
R9566 VSS.n111 VSS.n110 0.018
R9567 VSS.n474 VSS.n473 0.018
R9568 VSS.n87 VSS.n86 0.018
R9569 VSS.n145 VSS.n144 0.018
R9570 VSS.n151 VSS.n150 0.018
R9571 VSS.n433 VSS.n420 0.018
R9572 VSS.n371 VSS.n357 0.018
R9573 VSS.n319 VSS.n299 0.018
R9574 VSS.n274 VSS.n178 0.018
R9575 VSS.n274 VSS.n179 0.018
R9576 VSS.n371 VSS.n358 0.018
R9577 VSS.n319 VSS.n121 0.018
R9578 VSS.n274 VSS.n180 0.018
R9579 VSS.n445 VSS.n444 0.017
R9580 VSS.n166 VSS.n165 0.016
R9581 VSS.n285 VSS.n284 0.015
R9582 VSS.n333 VSS.n332 0.015
R9583 VSS.n381 VSS.n379 0.015
R9584 VSS.n445 VSS.n25 0.015
R9585 VSS.n381 VSS.n60 0.015
R9586 VSS.n333 VSS.n328 0.015
R9587 VSS.n285 VSS.n283 0.015
R9588 VSS.n333 VSS.n327 0.015
R9589 VSS.n285 VSS.n282 0.015
R9590 VSS.n381 VSS.n59 0.015
R9591 VSS.n445 VSS.n26 0.015
R9592 VSS.n350 VSS.n113 0.012
R9593 VSS.n412 VSS.n409 0.012
R9594 VSS.n72 VSS.n71 0.012
R9595 VSS.n310 VSS.n309 0.012
R9596 VSS.n413 VSS.n394 0.011
R9597 VSS.n476 VSS.n458 0.011
R9598 VSS.n445 VSS.n438 0.011
R9599 VSS.n381 VSS.n373 0.011
R9600 VSS.n333 VSS.n321 0.011
R9601 VSS.n285 VSS.n279 0.011
R9602 VSS.n381 VSS.n378 0.011
R9603 VSS.n333 VSS.n326 0.011
R9604 VSS.n158 VSS.n157 0.011
R9605 VSS.n156 VSS.n154 0.01
R9606 VSS.n145 VSS.n143 0.007
R9607 VSS.n278 VSS.n277 0.007
R9608 VSS.n320 VSS.n116 0.007
R9609 VSS.n100 VSS.n97 0.006
R9610 VSS.n20 VSS.n18 0.006
R9611 VSS.n474 VSS.n472 0.006
R9612 VSS.n151 VSS.n149 0.006
R9613 VSS.n372 VSS.n65 0.006
R9614 VSS.n445 VSS.n443 0.006
R9615 VSS.n437 VSS.n436 0.005
R9616 VSS.n53 VSS.n51 0.005
R9617 VSS.n87 VSS.n85 0.005
R9618 VSS.n290 VSS.n166 0.005
R9619 VSS.n81 VSS.n79 0.005
R9620 VSS.n41 VSS.n39 0.005
R9621 VSS.n405 VSS.n403 0.005
R9622 VSS VSS.n719 0.005
R9623 VSS.n294 VSS.n293 0.004
R9624 VSS.n73 VSS.n72 0.004
R9625 VSS.n311 VSS.n310 0.004
R9626 VSS.n93 VSS.n91 0.004
R9627 VSS.n14 VSS.n12 0.004
R9628 VSS.n105 VSS.n103 0.004
R9629 VSS.n255 VSS.n254 0.004
R9630 VSS.n298 VSS.n164 0.004
R9631 VSS.n325 VSS.n324 0.004
R9632 VSS.n449 VSS.n448 0.004
R9633 VSS.n442 VSS.n441 0.004
R9634 VSS.n377 VSS.n376 0.004
R9635 VSS.n385 VSS.n384 0.004
R9636 VSS.n337 VSS.n336 0.004
R9637 VSS.n289 VSS.n288 0.004
R9638 VSS.n594 VSS.n593 0.003
R9639 VSS.n496 VSS.n493 0.003
R9640 VSS.n512 VSS.n510 0.003
R9641 VSS.n502 VSS.n501 0.003
R9642 VSS.n274 VSS.n177 0.003
R9643 VSS.n695 VSS.n692 0.003
R9644 VSS.n630 VSS.n629 0.003
R9645 VSS.n643 VSS.n639 0.003
R9646 VSS.n111 VSS.n109 0.003
R9647 VSS.n47 VSS.n45 0.003
R9648 VSS.n20 VSS.n19 0.003
R9649 VSS.n53 VSS.n52 0.003
R9650 VSS.n93 VSS.n92 0.003
R9651 VSS.n14 VSS.n13 0.003
R9652 VSS.n47 VSS.n46 0.003
R9653 VSS.n81 VSS.n80 0.003
R9654 VSS.n41 VSS.n40 0.003
R9655 VSS.n466 VSS.n465 0.003
R9656 VSS.n518 VSS.n517 0.002
R9657 VSS.n684 VSS.n683 0.002
R9658 VSS.n213 VSS.n212 0.002
R9659 VSS.n635 VSS.n631 0.002
R9660 VSS.n156 VSS.n155 0.002
R9661 VSS.n105 VSS.n104 0.002
R9662 VSS.n405 VSS.n404 0.002
R9663 VSS.n399 VSS.n397 0.002
R9664 VSS.n479 VSS.n476 0.002
R9665 VSS VSS.n479 0.002
R9666 VSS.n138 VSS.n137 0.002
R9667 VSS.n350 VSS.n88 0.001
R9668 VSS.n88 VSS.n87 0.001
R9669 VSS.n146 VSS.n145 0.001
R9670 VSS.n298 VSS.n146 0.001
R9671 VSS.n152 VSS.n151 0.001
R9672 VSS.n298 VSS.n152 0.001
R9673 VSS.n413 VSS.n412 0.001
R9674 VSS.n412 VSS.n411 0.001
R9675 VSS.n350 VSS.n112 0.001
R9676 VSS.n112 VSS.n111 0.001
R9677 VSS.n476 VSS.n475 0.001
R9678 VSS.n475 VSS.n474 0.001
R9679 VSS.n140 VSS.n139 0.001
R9680 VSS.n298 VSS.n140 0.001
R9681 VSS.n413 VSS.n55 0.001
R9682 VSS.n256 VSS.n186 0.001
R9683 VSS.n256 VSS.n255 0.001
R9684 VSS.n274 VSS.n256 0.001
R9685 VSS.n319 VSS.n298 0.001
R9686 VSS.n371 VSS.n350 0.001
R9687 VSS.n433 VSS.n413 0.001
R9688 VSS.n719 VSS.n718 0.001
R9689 VSS.n683 VSS.n673 0.001
R9690 VSS.n673 VSS.n672 0.001
R9691 VSS.n672 VSS.n651 0.001
R9692 VSS.n651 VSS.n648 0.001
R9693 VSS.n631 VSS.n630 0.001
R9694 VSS.n468 VSS.n467 0.001
R9695 VSS.n476 VSS.n468 0.001
R9696 VSS.n320 VSS.n319 0.001
R9697 VSS.n372 VSS.n371 0.001
R9698 VSS.n333 VSS.n320 0.001
R9699 VSS.n381 VSS.n372 0.001
R9700 VSS.n413 VSS.n400 0.001
R9701 VSS.n400 VSS.n399 0.001
R9702 VSS.n350 VSS.n100 0.001
R9703 VSS.n100 VSS.n99 0.001
R9704 VSS.n285 VSS.n168 0.001
R9705 VSS.n290 VSS.n167 0.001
R9706 VSS.n445 VSS.n29 0.001
R9707 VSS.n333 VSS.n331 0.001
R9708 VSS.n648 VSS.n597 0.001
R9709 VSS.n719 VSS.n497 0.001
R9710 VSS.n673 VSS.n513 0.001
R9711 VSS.n672 VSS.n519 0.001
R9712 VSS.n294 VSS.n290 0.001
R9713 VSS.n298 VSS.n294 0.001
R9714 VSS.n254 VSS.n253 0.001
R9715 VSS.n254 VSS.n202 0.001
R9716 VSS.n254 VSS.n209 0.001
R9717 VSS.n254 VSS.n232 0.001
R9718 VSS.n254 VSS.n238 0.001
R9719 VSS.n254 VSS.n245 0.001
R9720 VSS.n254 VSS.n225 0.001
R9721 VSS.n254 VSS.n218 0.001
R9722 VSS.n648 VSS.n643 0.001
R9723 VSS.n628 VSS.n620 0.001
R9724 VSS.n628 VSS.n624 0.001
R9725 VSS.n629 VSS.n628 0.001
R9726 VSS.n651 VSS.n540 0.001
R9727 VSS.n648 VSS.n647 0.001
R9728 VSS.n253 VSS.n249 0.001
R9729 VSS.n202 VSS.n198 0.001
R9730 VSS.n209 VSS.n205 0.001
R9731 VSS.n232 VSS.n228 0.001
R9732 VSS.n238 VSS.n234 0.001
R9733 VSS.n245 VSS.n241 0.001
R9734 VSS.n225 VSS.n221 0.001
R9735 VSS.n218 VSS.n214 0.001
R9736 VSS.n139 VSS.n133 0.001
R9737 VSS.n695 VSS.n688 0.001
R9738 VSS.n651 VSS.n570 0.001
R9739 VSS.n639 VSS.n635 0.001
R9740 VSS.n467 VSS.n461 0.001
R9741 VSS.n18 VSS.n16 0.001
R9742 VSS.n149 VSS.n147 0.001
R9743 VSS.n254 VSS.n226 0.001
R9744 VSS.n397 VSS.n395 0.001
R9745 VSS.n103 VSS.n101 0.001
R9746 VSS.n254 VSS.n246 0.001
R9747 VSS.n79 VSS.n77 0.001
R9748 VSS.n254 VSS.n219 0.001
R9749 VSS.n254 VSS.n203 0.001
R9750 VSS.n472 VSS.n470 0.001
R9751 VSS.n403 VSS.n401 0.001
R9752 VSS.n409 VSS.n408 0.001
R9753 VSS.n91 VSS.n89 0.001
R9754 VSS.n51 VSS.n49 0.001
R9755 VSS.n39 VSS.n37 0.001
R9756 VSS.n143 VSS.n141 0.001
R9757 VSS.n254 VSS.n210 0.001
R9758 VSS.n254 VSS.n211 0.001
R9759 VSS.n109 VSS.n107 0.001
R9760 VSS.n45 VSS.n43 0.001
R9761 VSS.n254 VSS.n247 0.001
R9762 VSS.n12 VSS.n10 0.001
R9763 VSS.n85 VSS.n83 0.001
R9764 VSS.n254 VSS.n239 0.001
R9765 VSS.n97 VSS.n96 0.001
R9766 VSS.n254 VSS.n197 0.001
R9767 VSS.n254 VSS.n204 0.001
R9768 VSS.n254 VSS.n233 0.001
R9769 VSS.n254 VSS.n240 0.001
R9770 VSS.n254 VSS.n220 0.001
R9771 VSS.n254 VSS.n248 0.001
R9772 VSS.n254 VSS.n227 0.001
R9773 VSS.n254 VSS.n213 0.001
R9774 VSS.n371 VSS.n73 0.001
R9775 VSS.n319 VSS.n311 0.001
R9776 VSS VSS.n489 0.001
R9777 VSS VSS.n485 0.001
R9778 VSS.n722 VSS 0.001
R9779 VSS VSS.n486 0.001
R9780 VSS VSS.n482 0.001
R9781 VSS.n718 VSS.n502 0.001
R9782 VSS.n673 VSS.n512 0.001
R9783 VSS.n719 VSS.n496 0.001
R9784 VSS.n648 VSS.n594 0.001
R9785 VSS.n695 VSS.n684 0.001
R9786 VSS.n718 VSS.n699 0.001
R9787 VSS.n672 VSS.n518 0.001
R9788 VSS.n466 VSS.n462 0.001
R9789 VSS.n467 VSS.n466 0.001
R9790 VSS.n70 VSS.n69 0.001
R9791 VSS.n371 VSS.n70 0.001
R9792 VSS.n308 VSS.n307 0.001
R9793 VSS.n319 VSS.n308 0.001
R9794 VSS.n298 VSS.n158 0.001
R9795 VSS.n476 VSS.n21 0.001
R9796 VSS.n413 VSS.n54 0.001
R9797 VSS.n350 VSS.n94 0.001
R9798 VSS.n437 VSS.n433 0.001
R9799 VSS.n278 VSS.n274 0.001
R9800 VSS.n476 VSS.n15 0.001
R9801 VSS.n413 VSS.n48 0.001
R9802 VSS.n350 VSS.n82 0.001
R9803 VSS.n413 VSS.n42 0.001
R9804 VSS.n385 VSS.n381 0.001
R9805 VSS.n381 VSS.n380 0.001
R9806 VSS.n350 VSS.n106 0.001
R9807 VSS.n449 VSS.n445 0.001
R9808 VSS.n337 VSS.n333 0.001
R9809 VSS.n289 VSS.n285 0.001
R9810 VSS.n138 VSS.n134 0.001
R9811 VSS.n139 VSS.n138 0.001
R9812 VSS.n413 VSS.n406 0.001
R9813 VSS.n290 VSS.n289 0.001
R9814 VSS.n350 VSS.n337 0.001
R9815 VSS.n413 VSS.n385 0.001
R9816 VSS.n476 VSS.n449 0.001
R9817 VSS.n697 VSS.n695 0.001
R9818 VSS.n718 VSS.n697 0.001
R9819 VSS.n406 VSS.n405 0.001
R9820 VSS.n333 VSS.n325 0.001
R9821 VSS.n445 VSS.n442 0.001
R9822 VSS.n106 VSS.n105 0.001
R9823 VSS.n381 VSS.n377 0.001
R9824 VSS.n42 VSS.n41 0.001
R9825 VSS.n82 VSS.n81 0.001
R9826 VSS.n48 VSS.n47 0.001
R9827 VSS.n15 VSS.n14 0.001
R9828 VSS.n285 VSS.n278 0.001
R9829 VSS.n445 VSS.n437 0.001
R9830 VSS.n94 VSS.n93 0.001
R9831 VSS.n54 VSS.n53 0.001
R9832 VSS.n21 VSS.n20 0.001
R9833 VSS.n158 VSS.n156 0.001
R9834 a_59280_15743.n1 a_59280_15743.t6 318.922
R9835 a_59280_15743.n0 a_59280_15743.t5 273.935
R9836 a_59280_15743.n0 a_59280_15743.t7 273.935
R9837 a_59280_15743.n1 a_59280_15743.t4 269.116
R9838 a_59280_15743.n4 a_59280_15743.n3 193.227
R9839 a_59280_15743.t6 a_59280_15743.n0 179.142
R9840 a_59280_15743.n2 a_59280_15743.n1 106.999
R9841 a_59280_15743.n3 a_59280_15743.t0 28.568
R9842 a_59280_15743.n4 a_59280_15743.t1 28.565
R9843 a_59280_15743.t2 a_59280_15743.n4 28.565
R9844 a_59280_15743.n2 a_59280_15743.t3 18.149
R9845 a_59280_15743.n3 a_59280_15743.n2 3.726
R9846 a_42301_n1318.n7 a_42301_n1318.n6 861.987
R9847 a_42301_n1318.n6 a_42301_n1318.n5 560.726
R9848 a_42301_n1318.t4 a_42301_n1318.t12 415.315
R9849 a_42301_n1318.t5 a_42301_n1318.t6 415.315
R9850 a_42301_n1318.n2 a_42301_n1318.t14 394.151
R9851 a_42301_n1318.n5 a_42301_n1318.t19 294.653
R9852 a_42301_n1318.n1 a_42301_n1318.t18 269.523
R9853 a_42301_n1318.t14 a_42301_n1318.n1 269.523
R9854 a_42301_n1318.n9 a_42301_n1318.t4 217.716
R9855 a_42301_n1318.n8 a_42301_n1318.t16 214.335
R9856 a_42301_n1318.t12 a_42301_n1318.n8 214.335
R9857 a_42301_n1318.n0 a_42301_n1318.t7 214.335
R9858 a_42301_n1318.t6 a_42301_n1318.n0 214.335
R9859 a_42301_n1318.n7 a_42301_n1318.t5 198.921
R9860 a_42301_n1318.n3 a_42301_n1318.t17 198.043
R9861 a_42301_n1318.n12 a_42301_n1318.n11 192.754
R9862 a_42301_n1318.n1 a_42301_n1318.t10 160.666
R9863 a_42301_n1318.n5 a_42301_n1318.t8 111.663
R9864 a_42301_n1318.n4 a_42301_n1318.n2 97.816
R9865 a_42301_n1318.n3 a_42301_n1318.t13 93.989
R9866 a_42301_n1318.n8 a_42301_n1318.t9 80.333
R9867 a_42301_n1318.n2 a_42301_n1318.t11 80.333
R9868 a_42301_n1318.n0 a_42301_n1318.t15 80.333
R9869 a_42301_n1318.n6 a_42301_n1318.n4 65.07
R9870 a_42301_n1318.n11 a_42301_n1318.t2 28.568
R9871 a_42301_n1318.n12 a_42301_n1318.t1 28.565
R9872 a_42301_n1318.t0 a_42301_n1318.n12 28.565
R9873 a_42301_n1318.n10 a_42301_n1318.t3 18.827
R9874 a_42301_n1318.n9 a_42301_n1318.n7 16.411
R9875 a_42301_n1318.n4 a_42301_n1318.n3 6.615
R9876 a_42301_n1318.n10 a_42301_n1318.n9 4.997
R9877 a_42301_n1318.n11 a_42301_n1318.n10 1.105
R9878 a_44682_3363.t0 a_44682_3363.t1 17.4
R9879 a_63527_6198.n0 a_63527_6198.t9 214.335
R9880 a_63527_6198.t8 a_63527_6198.n0 214.335
R9881 a_63527_6198.n1 a_63527_6198.t8 143.851
R9882 a_63527_6198.n1 a_63527_6198.t10 135.658
R9883 a_63527_6198.n0 a_63527_6198.t7 80.333
R9884 a_63527_6198.n2 a_63527_6198.t6 28.565
R9885 a_63527_6198.n2 a_63527_6198.t5 28.565
R9886 a_63527_6198.n4 a_63527_6198.t4 28.565
R9887 a_63527_6198.n4 a_63527_6198.t2 28.565
R9888 a_63527_6198.t0 a_63527_6198.n7 28.565
R9889 a_63527_6198.n7 a_63527_6198.t1 28.565
R9890 a_63527_6198.n6 a_63527_6198.t3 9.714
R9891 a_63527_6198.n7 a_63527_6198.n6 1.003
R9892 a_63527_6198.n5 a_63527_6198.n3 0.833
R9893 a_63527_6198.n3 a_63527_6198.n2 0.653
R9894 a_63527_6198.n5 a_63527_6198.n4 0.653
R9895 a_63527_6198.n6 a_63527_6198.n5 0.341
R9896 a_63527_6198.n3 a_63527_6198.n1 0.032
R9897 a_64117_5761.n4 a_64117_5761.n3 563.136
R9898 a_64117_5761.t4 a_64117_5761.t14 437.233
R9899 a_64117_5761.t15 a_64117_5761.n1 313.873
R9900 a_64117_5761.n3 a_64117_5761.t6 294.986
R9901 a_64117_5761.n0 a_64117_5761.t8 272.288
R9902 a_64117_5761.n6 a_64117_5761.t4 217.824
R9903 a_64117_5761.n5 a_64117_5761.t12 214.686
R9904 a_64117_5761.t14 a_64117_5761.n5 214.686
R9905 a_64117_5761.n9 a_64117_5761.n8 192.754
R9906 a_64117_5761.n2 a_64117_5761.t15 190.152
R9907 a_64117_5761.n2 a_64117_5761.t5 190.152
R9908 a_64117_5761.n4 a_64117_5761.t11 178.973
R9909 a_64117_5761.n0 a_64117_5761.t13 160.666
R9910 a_64117_5761.n1 a_64117_5761.t10 160.666
R9911 a_64117_5761.n6 a_64117_5761.n4 133.838
R9912 a_64117_5761.n3 a_64117_5761.t7 110.859
R9913 a_64117_5761.n1 a_64117_5761.n0 96.129
R9914 a_64117_5761.t11 a_64117_5761.n2 80.333
R9915 a_64117_5761.n5 a_64117_5761.t9 80.333
R9916 a_64117_5761.n8 a_64117_5761.t0 28.568
R9917 a_64117_5761.t2 a_64117_5761.n9 28.565
R9918 a_64117_5761.n9 a_64117_5761.t1 28.565
R9919 a_64117_5761.n7 a_64117_5761.t3 18.824
R9920 a_64117_5761.n7 a_64117_5761.n6 5.567
R9921 a_64117_5761.n8 a_64117_5761.n7 1.105
R9922 a_70513_4160.n0 a_70513_4160.t2 14.282
R9923 a_70513_4160.t0 a_70513_4160.n0 14.282
R9924 a_70513_4160.n0 a_70513_4160.n1 258.161
R9925 a_70513_4160.n1 a_70513_4160.t1 14.283
R9926 a_70513_4160.n1 a_70513_4160.n5 0.852
R9927 a_70513_4160.n5 a_70513_4160.n6 4.366
R9928 a_70513_4160.n6 a_70513_4160.n7 258.161
R9929 a_70513_4160.n7 a_70513_4160.t7 14.282
R9930 a_70513_4160.n7 a_70513_4160.t5 14.282
R9931 a_70513_4160.n6 a_70513_4160.t6 14.283
R9932 a_70513_4160.n5 a_70513_4160.n4 73.514
R9933 a_70513_4160.n4 a_70513_4160.t8 1551.5
R9934 a_70513_4160.t8 a_70513_4160.n3 656.576
R9935 a_70513_4160.n3 a_70513_4160.t4 8.7
R9936 a_70513_4160.n3 a_70513_4160.t3 8.7
R9937 a_70513_4160.n4 a_70513_4160.t10 224.129
R9938 a_70513_4160.t10 a_70513_4160.n2 207.225
R9939 a_70513_4160.n2 a_70513_4160.t9 207.225
R9940 a_70513_4160.n2 a_70513_4160.t11 80.333
R9941 a_7957_1259.n3 a_7957_1259.t4 867.497
R9942 a_7957_1259.n3 a_7957_1259.t5 615.911
R9943 a_7957_1259.n2 a_7957_1259.t6 286.438
R9944 a_7957_1259.n2 a_7957_1259.t7 286.438
R9945 a_7957_1259.n10 a_7957_1259.n9 185.55
R9946 a_7957_1259.t4 a_7957_1259.n2 160.666
R9947 a_7957_1259.n8 a_7957_1259.n7 109.481
R9948 a_7957_1259.n9 a_7957_1259.t1 28.568
R9949 a_7957_1259.t2 a_7957_1259.n10 28.565
R9950 a_7957_1259.n10 a_7957_1259.t0 28.565
R9951 a_7957_1259.n8 a_7957_1259.t3 20.393
R9952 a_7957_1259.n4 a_7957_1259.n3 15.739
R9953 a_7957_1259.n9 a_7957_1259.n8 1.834
R9954 a_7957_1259.n7 a_7957_1259.n6 0.09
R9955 a_7957_1259.n6 a_7957_1259.n5 0.075
R9956 a_7957_1259.n1 a_7957_1259.n0 0.001
R9957 a_7957_1259.n5 a_7957_1259.n4 0.001
R9958 a_7957_1259.n4 a_7957_1259.n1 0.001
R9959 a_45279_16157.n6 a_45279_16157.n5 501.28
R9960 a_45279_16157.t7 a_45279_16157.t13 437.233
R9961 a_45279_16157.t15 a_45279_16157.t17 415.315
R9962 a_45279_16157.t8 a_45279_16157.n3 313.873
R9963 a_45279_16157.n5 a_45279_16157.t4 294.986
R9964 a_45279_16157.n2 a_45279_16157.t9 272.288
R9965 a_45279_16157.n6 a_45279_16157.t6 236.009
R9966 a_45279_16157.n9 a_45279_16157.t7 216.627
R9967 a_45279_16157.n7 a_45279_16157.t15 216.111
R9968 a_45279_16157.n8 a_45279_16157.t16 214.686
R9969 a_45279_16157.t13 a_45279_16157.n8 214.686
R9970 a_45279_16157.n1 a_45279_16157.t11 214.335
R9971 a_45279_16157.t17 a_45279_16157.n1 214.335
R9972 a_45279_16157.n4 a_45279_16157.t5 190.152
R9973 a_45279_16157.n4 a_45279_16157.t8 190.152
R9974 a_45279_16157.n2 a_45279_16157.t19 160.666
R9975 a_45279_16157.n3 a_45279_16157.t18 160.666
R9976 a_45279_16157.n7 a_45279_16157.n6 148.428
R9977 a_45279_16157.n5 a_45279_16157.t10 110.859
R9978 a_45279_16157.n3 a_45279_16157.n2 96.129
R9979 a_45279_16157.n8 a_45279_16157.t14 80.333
R9980 a_45279_16157.n1 a_45279_16157.t12 80.333
R9981 a_45279_16157.t6 a_45279_16157.n4 80.333
R9982 a_45279_16157.t0 a_45279_16157.n11 28.57
R9983 a_45279_16157.n0 a_45279_16157.t3 28.565
R9984 a_45279_16157.n0 a_45279_16157.t2 28.565
R9985 a_45279_16157.n11 a_45279_16157.t1 17.638
R9986 a_45279_16157.n10 a_45279_16157.n9 5.589
R9987 a_45279_16157.n9 a_45279_16157.n7 2.923
R9988 a_45279_16157.n10 a_45279_16157.n0 0.693
R9989 a_45279_16157.n11 a_45279_16157.n10 0.597
R9990 a_46175_15029.t0 a_46175_15029.t1 17.4
R9991 a_54665_15740.n1 a_54665_15740.t4 318.922
R9992 a_54665_15740.n0 a_54665_15740.t7 273.935
R9993 a_54665_15740.n0 a_54665_15740.t5 273.935
R9994 a_54665_15740.n1 a_54665_15740.t6 269.116
R9995 a_54665_15740.n4 a_54665_15740.n3 193.227
R9996 a_54665_15740.t4 a_54665_15740.n0 179.142
R9997 a_54665_15740.n2 a_54665_15740.n1 106.999
R9998 a_54665_15740.n3 a_54665_15740.t3 28.568
R9999 a_54665_15740.n4 a_54665_15740.t1 28.565
R10000 a_54665_15740.t0 a_54665_15740.n4 28.565
R10001 a_54665_15740.n2 a_54665_15740.t2 18.149
R10002 a_54665_15740.n3 a_54665_15740.n2 3.726
R10003 a_54253_15766.n0 a_54253_15766.t8 14.282
R10004 a_54253_15766.t0 a_54253_15766.n0 14.282
R10005 a_54253_15766.n0 a_54253_15766.n9 1.511
R10006 a_54253_15766.n9 a_54253_15766.n5 0.227
R10007 a_54253_15766.n9 a_54253_15766.n6 0.669
R10008 a_54253_15766.n6 a_54253_15766.n7 0.001
R10009 a_54253_15766.n6 a_54253_15766.n8 267.767
R10010 a_54253_15766.n8 a_54253_15766.t1 14.282
R10011 a_54253_15766.n8 a_54253_15766.t5 14.282
R10012 a_54253_15766.n7 a_54253_15766.t6 14.282
R10013 a_54253_15766.n7 a_54253_15766.t7 14.282
R10014 a_54253_15766.n5 a_54253_15766.n2 0.2
R10015 a_54253_15766.n5 a_54253_15766.n4 0.575
R10016 a_54253_15766.n4 a_54253_15766.t2 16.058
R10017 a_54253_15766.n4 a_54253_15766.n3 0.999
R10018 a_54253_15766.n3 a_54253_15766.t4 14.282
R10019 a_54253_15766.n3 a_54253_15766.t3 14.282
R10020 a_54253_15766.n2 a_54253_15766.n1 0.999
R10021 a_54253_15766.n1 a_54253_15766.t10 14.282
R10022 a_54253_15766.n1 a_54253_15766.t11 14.282
R10023 a_54253_15766.n2 a_54253_15766.t9 16.058
R10024 a_52710_16433.n0 a_52710_16433.n12 90.436
R10025 a_52710_16433.t5 a_52710_16433.n0 14.282
R10026 a_52710_16433.n0 a_52710_16433.t6 14.282
R10027 a_52710_16433.n12 a_52710_16433.n9 74.302
R10028 a_52710_16433.n9 a_52710_16433.n11 50.575
R10029 a_52710_16433.n11 a_52710_16433.n10 157.665
R10030 a_52710_16433.n10 a_52710_16433.t4 8.7
R10031 a_52710_16433.n10 a_52710_16433.t3 8.7
R10032 a_52710_16433.n9 a_52710_16433.n8 90.416
R10033 a_52710_16433.n8 a_52710_16433.t7 14.282
R10034 a_52710_16433.n8 a_52710_16433.t0 14.282
R10035 a_52710_16433.n11 a_52710_16433.n7 122.746
R10036 a_52710_16433.n7 a_52710_16433.t2 14.282
R10037 a_52710_16433.n7 a_52710_16433.t1 14.282
R10038 a_52710_16433.n12 a_52710_16433.n1 342.688
R10039 a_52710_16433.n1 a_52710_16433.n6 126.566
R10040 a_52710_16433.n6 a_52710_16433.t15 294.653
R10041 a_52710_16433.n6 a_52710_16433.t13 111.663
R10042 a_52710_16433.n1 a_52710_16433.n5 552.333
R10043 a_52710_16433.n5 a_52710_16433.n4 6.615
R10044 a_52710_16433.n4 a_52710_16433.t11 93.989
R10045 a_52710_16433.n4 a_52710_16433.t12 198.043
R10046 a_52710_16433.n5 a_52710_16433.n3 97.816
R10047 a_52710_16433.n3 a_52710_16433.t10 80.333
R10048 a_52710_16433.n3 a_52710_16433.t9 394.151
R10049 a_52710_16433.t9 a_52710_16433.n2 269.523
R10050 a_52710_16433.n2 a_52710_16433.t8 160.666
R10051 a_52710_16433.n2 a_52710_16433.t14 269.523
R10052 B[6].n6 B[6].t28 5229.8
R10053 B[6].t23 B[6].t27 800.875
R10054 B[6].n12 B[6].n6 692.057
R10055 B[6].n22 B[6].n21 648.993
R10056 B[6].n17 B[6].n16 618.566
R10057 B[6].n11 B[6].n7 592.056
R10058 B[6].t16 B[6].t0 437.233
R10059 B[6].t19 B[6].t29 437.233
R10060 B[6].t2 B[6].t9 415.315
R10061 B[6].t28 B[6].t10 415.315
R10062 B[6].t24 B[6].t1 415.315
R10063 B[6].t34 B[6].n14 313.873
R10064 B[6].t6 B[6].n9 313.069
R10065 B[6].n7 B[6].t30 294.986
R10066 B[6].n20 B[6].t21 284.688
R10067 B[6].n16 B[6].t35 273.077
R10068 B[6].n13 B[6].t33 272.288
R10069 B[6].n8 B[6].t13 271.484
R10070 B[6].n4 B[6].t24 220.313
R10071 B[6].n5 B[6].t16 219.163
R10072 B[6].n19 B[6].t2 217.532
R10073 B[6].n4 B[6].t19 217.194
R10074 B[6].n1 B[6].t3 214.686
R10075 B[6].t0 B[6].n1 214.686
R10076 B[6].n3 B[6].t14 214.686
R10077 B[6].t29 B[6].n3 214.686
R10078 B[6].n0 B[6].t38 214.335
R10079 B[6].t10 B[6].n0 214.335
R10080 B[6].n2 B[6].t18 214.335
R10081 B[6].t1 B[6].n2 214.335
R10082 B[6].n18 B[6].t39 214.335
R10083 B[6].t9 B[6].n18 214.335
R10084 B[6].n17 B[6].t5 204.679
R10085 B[6].n11 B[6].t25 204.672
R10086 B[6].n21 B[6].t23 192.799
R10087 B[6].n10 B[6].t6 190.955
R10088 B[6].n10 B[6].t31 190.955
R10089 B[6].n15 B[6].t17 190.152
R10090 B[6].n15 B[6].t34 190.152
R10091 B[6].n9 B[6].t37 160.666
R10092 B[6].n8 B[6].t20 160.666
R10093 B[6].n13 B[6].t32 160.666
R10094 B[6].n14 B[6].t11 160.666
R10095 B[6].n20 B[6].t22 160.666
R10096 B[6].n16 B[6].t7 137.369
R10097 B[6].n7 B[6].t26 110.859
R10098 B[6].n9 B[6].n8 96.129
R10099 B[6].n14 B[6].n13 96.129
R10100 B[6].n21 B[6].n20 91.889
R10101 B[6].n0 B[6].t12 80.333
R10102 B[6].n1 B[6].t4 80.333
R10103 B[6].n2 B[6].t36 80.333
R10104 B[6].n3 B[6].t15 80.333
R10105 B[6].t25 B[6].n10 80.333
R10106 B[6].n18 B[6].t8 80.333
R10107 B[6].t5 B[6].n15 80.333
R10108 B[6].n19 B[6].n17 51.824
R10109 B[6] B[6].n23 47.217
R10110 B[6].n12 B[6].n11 46.161
R10111 B[6].n23 B[6].n12 34.775
R10112 B[6].n23 B[6].n22 24.272
R10113 B[6].n6 B[6].n5 23.931
R10114 B[6].n5 B[6].n4 11.749
R10115 B[6].n22 B[6].n19 6.378
R10116 a_54914_n1762.n2 a_54914_n1762.t10 214.335
R10117 a_54914_n1762.t8 a_54914_n1762.n2 214.335
R10118 a_54914_n1762.n3 a_54914_n1762.t8 143.85
R10119 a_54914_n1762.n3 a_54914_n1762.t7 135.66
R10120 a_54914_n1762.n2 a_54914_n1762.t9 80.333
R10121 a_54914_n1762.n4 a_54914_n1762.t6 28.565
R10122 a_54914_n1762.n4 a_54914_n1762.t5 28.565
R10123 a_54914_n1762.n0 a_54914_n1762.t0 28.565
R10124 a_54914_n1762.n0 a_54914_n1762.t1 28.565
R10125 a_54914_n1762.t4 a_54914_n1762.n7 28.565
R10126 a_54914_n1762.n7 a_54914_n1762.t2 28.565
R10127 a_54914_n1762.n1 a_54914_n1762.t3 9.714
R10128 a_54914_n1762.n1 a_54914_n1762.n0 1.003
R10129 a_54914_n1762.n6 a_54914_n1762.n5 0.836
R10130 a_54914_n1762.n7 a_54914_n1762.n6 0.653
R10131 a_54914_n1762.n5 a_54914_n1762.n4 0.65
R10132 a_54914_n1762.n6 a_54914_n1762.n1 0.341
R10133 a_54914_n1762.n5 a_54914_n1762.n3 0.032
R10134 a_44405_8194.n6 a_44405_8194.n5 501.28
R10135 a_44405_8194.t10 a_44405_8194.t7 437.233
R10136 a_44405_8194.t8 a_44405_8194.t5 415.315
R10137 a_44405_8194.t13 a_44405_8194.n3 313.873
R10138 a_44405_8194.n5 a_44405_8194.t19 294.986
R10139 a_44405_8194.n2 a_44405_8194.t11 272.288
R10140 a_44405_8194.n6 a_44405_8194.t4 236.01
R10141 a_44405_8194.n9 a_44405_8194.t10 216.627
R10142 a_44405_8194.n7 a_44405_8194.t8 216.111
R10143 a_44405_8194.n8 a_44405_8194.t18 214.686
R10144 a_44405_8194.t7 a_44405_8194.n8 214.686
R10145 a_44405_8194.n1 a_44405_8194.t9 214.335
R10146 a_44405_8194.t5 a_44405_8194.n1 214.335
R10147 a_44405_8194.n4 a_44405_8194.t13 190.152
R10148 a_44405_8194.n4 a_44405_8194.t14 190.152
R10149 a_44405_8194.n2 a_44405_8194.t6 160.666
R10150 a_44405_8194.n3 a_44405_8194.t16 160.666
R10151 a_44405_8194.n7 a_44405_8194.n6 148.428
R10152 a_44405_8194.n5 a_44405_8194.t17 110.859
R10153 a_44405_8194.n3 a_44405_8194.n2 96.129
R10154 a_44405_8194.n8 a_44405_8194.t12 80.333
R10155 a_44405_8194.n1 a_44405_8194.t15 80.333
R10156 a_44405_8194.t4 a_44405_8194.n4 80.333
R10157 a_44405_8194.n0 a_44405_8194.t3 28.57
R10158 a_44405_8194.n11 a_44405_8194.t2 28.565
R10159 a_44405_8194.t0 a_44405_8194.n11 28.565
R10160 a_44405_8194.n0 a_44405_8194.t1 17.638
R10161 a_44405_8194.n10 a_44405_8194.n9 12.318
R10162 a_44405_8194.n9 a_44405_8194.n7 2.923
R10163 a_44405_8194.n11 a_44405_8194.n10 0.69
R10164 a_44405_8194.n10 a_44405_8194.n0 0.6
R10165 a_48548_6884.n1 a_48548_6884.t4 318.922
R10166 a_48548_6884.n0 a_48548_6884.t5 274.739
R10167 a_48548_6884.n0 a_48548_6884.t7 274.739
R10168 a_48548_6884.n1 a_48548_6884.t6 269.116
R10169 a_48548_6884.t4 a_48548_6884.n0 179.946
R10170 a_48548_6884.n2 a_48548_6884.n1 105.178
R10171 a_48548_6884.n3 a_48548_6884.t0 29.444
R10172 a_48548_6884.t2 a_48548_6884.n4 28.565
R10173 a_48548_6884.n4 a_48548_6884.t1 28.565
R10174 a_48548_6884.n2 a_48548_6884.t3 18.145
R10175 a_48548_6884.n3 a_48548_6884.n2 2.878
R10176 a_48548_6884.n4 a_48548_6884.n3 0.764
R10177 a_3591_21596.n0 a_3591_21596.n9 167.433
R10178 a_3591_21596.n0 a_3591_21596.t6 14.282
R10179 a_3591_21596.t0 a_3591_21596.n0 14.282
R10180 a_3591_21596.n9 a_3591_21596.n8 77.784
R10181 a_3591_21596.n8 a_3591_21596.n6 77.456
R10182 a_3591_21596.n6 a_3591_21596.n4 77.456
R10183 a_3591_21596.n4 a_3591_21596.n2 75.815
R10184 a_3591_21596.n9 a_3591_21596.t1 104.259
R10185 a_3591_21596.n8 a_3591_21596.n7 89.977
R10186 a_3591_21596.n7 a_3591_21596.t2 14.282
R10187 a_3591_21596.n7 a_3591_21596.t8 14.282
R10188 a_3591_21596.n6 a_3591_21596.n5 89.977
R10189 a_3591_21596.n5 a_3591_21596.t7 14.282
R10190 a_3591_21596.n5 a_3591_21596.t9 14.282
R10191 a_3591_21596.n4 a_3591_21596.n3 89.977
R10192 a_3591_21596.n3 a_3591_21596.t10 14.282
R10193 a_3591_21596.n3 a_3591_21596.t11 14.282
R10194 a_3591_21596.n2 a_3591_21596.t5 104.259
R10195 a_3591_21596.n2 a_3591_21596.n1 167.433
R10196 a_3591_21596.n1 a_3591_21596.t4 14.282
R10197 a_3591_21596.n1 a_3591_21596.t3 14.282
R10198 A[6].n35 A[6].n25 2865.54
R10199 A[6].n21 A[6].t36 2858.78
R10200 A[6].n25 A[6].n21 2573.2
R10201 A[6].n8 A[6].n7 2321.13
R10202 A[6].n17 A[6].n16 1027.63
R10203 A[6].n17 A[6].t10 990.34
R10204 A[6].n16 A[6].t31 867.497
R10205 A[6].n16 A[6].t37 591.811
R10206 A[6].t2 A[6].t57 575.234
R10207 A[6].n30 A[6].n29 535.449
R10208 A[6].t19 A[6].t32 437.233
R10209 A[6].t36 A[6].t14 437.233
R10210 A[6].t17 A[6].t26 437.233
R10211 A[6].t3 A[6].t7 437.233
R10212 A[6].n36 A[6].n18 435.722
R10213 A[6].t9 A[6].t58 415.315
R10214 A[6].t59 A[6].t5 415.315
R10215 A[6].t18 A[6].t52 415.315
R10216 A[6].n5 A[6].n4 412.11
R10217 A[6].n17 A[6].t45 408.211
R10218 A[6].n2 A[6].t28 394.151
R10219 A[6].t47 A[6].n27 313.873
R10220 A[6].n29 A[6].t40 294.986
R10221 A[6].n4 A[6].t25 294.653
R10222 A[6].n14 A[6].t0 286.438
R10223 A[6].n14 A[6].t15 286.438
R10224 A[6].n15 A[6].t6 286.438
R10225 A[6].n15 A[6].t33 286.438
R10226 A[6].n10 A[6].t43 284.688
R10227 A[6].n26 A[6].t53 272.288
R10228 A[6].n1 A[6].t23 269.523
R10229 A[6].t28 A[6].n1 269.523
R10230 A[6].n30 A[6].t46 245.184
R10231 A[6].n24 A[6].t18 238.523
R10232 A[6].n5 A[6].n3 224.13
R10233 A[6].n12 A[6].t19 222.529
R10234 A[6].n32 A[6].t3 218.627
R10235 A[6].n24 A[6].t59 217.897
R10236 A[6].n21 A[6].t9 217.528
R10237 A[6].n34 A[6].t17 217.023
R10238 A[6].n9 A[6].t35 214.686
R10239 A[6].t32 A[6].n9 214.686
R10240 A[6].n20 A[6].t20 214.686
R10241 A[6].t14 A[6].n20 214.686
R10242 A[6].n33 A[6].t30 214.686
R10243 A[6].t26 A[6].n33 214.686
R10244 A[6].n31 A[6].t16 214.686
R10245 A[6].t7 A[6].n31 214.686
R10246 A[6].n19 A[6].t29 214.335
R10247 A[6].t58 A[6].n19 214.335
R10248 A[6].n22 A[6].t13 214.335
R10249 A[6].t5 A[6].n22 214.335
R10250 A[6].n23 A[6].t56 214.335
R10251 A[6].t52 A[6].n23 214.335
R10252 A[6].n0 A[6].t50 198.043
R10253 A[6].n28 A[6].t44 190.152
R10254 A[6].n28 A[6].t47 190.152
R10255 A[6].n6 A[6].t42 185.301
R10256 A[6].n6 A[6].t8 185.301
R10257 A[6].n12 A[6].n11 181.968
R10258 A[6].t10 A[6].n14 160.666
R10259 A[6].t31 A[6].n15 160.666
R10260 A[6].n1 A[6].t49 160.666
R10261 A[6].n10 A[6].t1 160.666
R10262 A[6].n11 A[6].t2 160.666
R10263 A[6].n26 A[6].t51 160.666
R10264 A[6].n27 A[6].t38 160.666
R10265 A[6].n8 A[6].n5 142.366
R10266 A[6].n7 A[6].t21 137.369
R10267 A[6].n11 A[6].n10 115.593
R10268 A[6].n4 A[6].t41 111.663
R10269 A[6].n29 A[6].t55 110.859
R10270 A[6].n6 A[6].t11 107.646
R10271 A[6].n3 A[6].n2 97.816
R10272 A[6].n27 A[6].n26 96.129
R10273 A[6].n0 A[6].t24 93.989
R10274 A[6].n2 A[6].t48 80.333
R10275 A[6].n9 A[6].t34 80.333
R10276 A[6].n19 A[6].t4 80.333
R10277 A[6].n20 A[6].t22 80.333
R10278 A[6].n22 A[6].t39 80.333
R10279 A[6].n23 A[6].t54 80.333
R10280 A[6].n33 A[6].t27 80.333
R10281 A[6].t46 A[6].n28 80.333
R10282 A[6].n31 A[6].t12 80.333
R10283 A[6].n7 A[6].n6 61.856
R10284 A[6] A[6].n36 48.497
R10285 A[6].n13 A[6].n12 38.951
R10286 A[6].n35 A[6].n34 37.965
R10287 A[6].n18 A[6].n17 34.1
R10288 A[6].n13 A[6].n8 31.43
R10289 A[6].n32 A[6].n30 14.9
R10290 A[6].n18 A[6].n13 10.125
R10291 A[6].n3 A[6].n0 6.615
R10292 A[6].n36 A[6].n35 3.16
R10293 A[6].n34 A[6].n32 2.599
R10294 A[6].n25 A[6].n24 0.274
R10295 a_9867_21592.n0 a_9867_21592.t4 14.282
R10296 a_9867_21592.t3 a_9867_21592.n0 14.282
R10297 a_9867_21592.n0 a_9867_21592.n9 89.977
R10298 a_9867_21592.n9 a_9867_21592.n7 77.784
R10299 a_9867_21592.n9 a_9867_21592.n6 77.456
R10300 a_9867_21592.n6 a_9867_21592.n4 77.456
R10301 a_9867_21592.n4 a_9867_21592.n2 75.815
R10302 a_9867_21592.n7 a_9867_21592.n8 167.433
R10303 a_9867_21592.n8 a_9867_21592.t5 14.282
R10304 a_9867_21592.n8 a_9867_21592.t6 14.282
R10305 a_9867_21592.n7 a_9867_21592.t7 104.259
R10306 a_9867_21592.n6 a_9867_21592.n5 89.977
R10307 a_9867_21592.n5 a_9867_21592.t11 14.282
R10308 a_9867_21592.n5 a_9867_21592.t10 14.282
R10309 a_9867_21592.n4 a_9867_21592.n3 89.977
R10310 a_9867_21592.n3 a_9867_21592.t8 14.282
R10311 a_9867_21592.n3 a_9867_21592.t9 14.282
R10312 a_9867_21592.n2 a_9867_21592.t2 104.259
R10313 a_9867_21592.n2 a_9867_21592.n1 167.433
R10314 a_9867_21592.n1 a_9867_21592.t1 14.282
R10315 a_9867_21592.n1 a_9867_21592.t0 14.282
R10316 a_48124_21370.n0 a_48124_21370.t3 14.282
R10317 a_48124_21370.t0 a_48124_21370.n0 14.282
R10318 a_48124_21370.n0 a_48124_21370.n12 90.416
R10319 a_48124_21370.n12 a_48124_21370.n11 50.575
R10320 a_48124_21370.n12 a_48124_21370.n8 74.302
R10321 a_48124_21370.n11 a_48124_21370.n10 157.665
R10322 a_48124_21370.n10 a_48124_21370.t7 8.7
R10323 a_48124_21370.n10 a_48124_21370.t6 8.7
R10324 a_48124_21370.n11 a_48124_21370.n9 122.999
R10325 a_48124_21370.n9 a_48124_21370.t4 14.282
R10326 a_48124_21370.n9 a_48124_21370.t5 14.282
R10327 a_48124_21370.n8 a_48124_21370.n7 90.436
R10328 a_48124_21370.n7 a_48124_21370.t1 14.282
R10329 a_48124_21370.n7 a_48124_21370.t2 14.282
R10330 a_48124_21370.n8 a_48124_21370.n1 342.688
R10331 a_48124_21370.n1 a_48124_21370.n6 126.566
R10332 a_48124_21370.n6 a_48124_21370.t12 294.653
R10333 a_48124_21370.n6 a_48124_21370.t8 111.663
R10334 a_48124_21370.n1 a_48124_21370.n5 552.333
R10335 a_48124_21370.n5 a_48124_21370.n4 6.615
R10336 a_48124_21370.n4 a_48124_21370.t14 93.989
R10337 a_48124_21370.n5 a_48124_21370.n3 97.816
R10338 a_48124_21370.n3 a_48124_21370.t15 80.333
R10339 a_48124_21370.n3 a_48124_21370.t9 394.151
R10340 a_48124_21370.t9 a_48124_21370.n2 269.523
R10341 a_48124_21370.n2 a_48124_21370.t10 160.666
R10342 a_48124_21370.n2 a_48124_21370.t11 269.523
R10343 a_48124_21370.n4 a_48124_21370.t13 198.043
R10344 a_49477_22063.n2 a_49477_22063.t7 318.922
R10345 a_49477_22063.n1 a_49477_22063.t6 273.935
R10346 a_49477_22063.n1 a_49477_22063.t5 273.935
R10347 a_49477_22063.n2 a_49477_22063.t4 269.116
R10348 a_49477_22063.n4 a_49477_22063.n0 193.227
R10349 a_49477_22063.t7 a_49477_22063.n1 179.142
R10350 a_49477_22063.n3 a_49477_22063.n2 106.999
R10351 a_49477_22063.t2 a_49477_22063.n4 28.568
R10352 a_49477_22063.n0 a_49477_22063.t0 28.565
R10353 a_49477_22063.n0 a_49477_22063.t1 28.565
R10354 a_49477_22063.n3 a_49477_22063.t3 18.149
R10355 a_49477_22063.n4 a_49477_22063.n3 3.726
R10356 A[2].n12 A[2].n11 3389.21
R10357 A[2].n17 A[2].n16 1131.17
R10358 A[2].n17 A[2].t21 990.34
R10359 A[2].n16 A[2].t17 867.497
R10360 A[2].n16 A[2].t43 591.811
R10361 A[2].t42 A[2].t15 573.627
R10362 A[2].n23 A[2].n22 535.449
R10363 A[2].n28 A[2].n18 500.512
R10364 A[2].t12 A[2].t22 437.233
R10365 A[2].t38 A[2].t41 437.233
R10366 A[2].t0 A[2].t3 437.233
R10367 A[2].n9 A[2].n8 412.11
R10368 A[2].n17 A[2].t7 408.211
R10369 A[2].n6 A[2].t13 394.151
R10370 A[2].t33 A[2].n20 313.873
R10371 A[2].n22 A[2].t26 294.986
R10372 A[2].n8 A[2].t36 294.653
R10373 A[2].n14 A[2].t20 286.438
R10374 A[2].n14 A[2].t40 286.438
R10375 A[2].n15 A[2].t16 286.438
R10376 A[2].n15 A[2].t32 286.438
R10377 A[2].n1 A[2].t24 285.543
R10378 A[2].n19 A[2].t8 272.288
R10379 A[2].n5 A[2].t1 269.523
R10380 A[2].t13 A[2].n5 269.523
R10381 A[2].n23 A[2].t6 245.184
R10382 A[2].n9 A[2].n7 224.13
R10383 A[2].n3 A[2].t12 220.881
R10384 A[2].n25 A[2].t0 218.628
R10385 A[2].n27 A[2].t38 217.024
R10386 A[2].n0 A[2].t19 214.686
R10387 A[2].t22 A[2].n0 214.686
R10388 A[2].n26 A[2].t10 214.686
R10389 A[2].t41 A[2].n26 214.686
R10390 A[2].n24 A[2].t35 214.686
R10391 A[2].t3 A[2].n24 214.686
R10392 A[2].n4 A[2].t4 198.043
R10393 A[2].n21 A[2].t33 190.152
R10394 A[2].n21 A[2].t14 190.152
R10395 A[2].n10 A[2].t39 186.908
R10396 A[2].n10 A[2].t28 186.908
R10397 A[2].n3 A[2].n2 182.197
R10398 A[2].n1 A[2].t27 160.666
R10399 A[2].n2 A[2].t42 160.666
R10400 A[2].n5 A[2].t31 160.666
R10401 A[2].t21 A[2].n14 160.666
R10402 A[2].t17 A[2].n15 160.666
R10403 A[2].n19 A[2].t9 160.666
R10404 A[2].n20 A[2].t11 160.666
R10405 A[2].n12 A[2].n9 141.534
R10406 A[2].n11 A[2].t5 140.583
R10407 A[2].n18 A[2].n17 129.415
R10408 A[2].n2 A[2].n1 114.089
R10409 A[2].n8 A[2].t25 111.663
R10410 A[2].n22 A[2].t34 110.859
R10411 A[2].n10 A[2].t2 109.253
R10412 A[2].n7 A[2].n6 97.816
R10413 A[2].n20 A[2].n19 96.129
R10414 A[2].n4 A[2].t30 93.989
R10415 A[2].n0 A[2].t18 80.333
R10416 A[2].n6 A[2].t29 80.333
R10417 A[2].n26 A[2].t23 80.333
R10418 A[2].t6 A[2].n21 80.333
R10419 A[2].n24 A[2].t37 80.333
R10420 A[2].n11 A[2].n10 61.856
R10421 A[2] A[2].n28 45.457
R10422 A[2].n13 A[2].n3 31.383
R10423 A[2].n28 A[2].n27 29.008
R10424 A[2].n25 A[2].n23 14.9
R10425 A[2].n18 A[2].n13 12.997
R10426 A[2].n13 A[2].n12 11.766
R10427 A[2].n7 A[2].n4 6.615
R10428 A[2].n27 A[2].n25 2.599
R10429 a_52762_21071.n4 a_52762_21071.t10 214.335
R10430 a_52762_21071.t7 a_52762_21071.n4 214.335
R10431 a_52762_21071.n5 a_52762_21071.t7 143.851
R10432 a_52762_21071.n5 a_52762_21071.t8 135.658
R10433 a_52762_21071.n4 a_52762_21071.t9 80.333
R10434 a_52762_21071.n0 a_52762_21071.t3 28.565
R10435 a_52762_21071.n0 a_52762_21071.t4 28.565
R10436 a_52762_21071.n2 a_52762_21071.t1 28.565
R10437 a_52762_21071.n2 a_52762_21071.t5 28.565
R10438 a_52762_21071.t0 a_52762_21071.n7 28.565
R10439 a_52762_21071.n7 a_52762_21071.t2 28.565
R10440 a_52762_21071.n1 a_52762_21071.t6 9.714
R10441 a_52762_21071.n1 a_52762_21071.n0 1.003
R10442 a_52762_21071.n6 a_52762_21071.n3 0.833
R10443 a_52762_21071.n3 a_52762_21071.n2 0.653
R10444 a_52762_21071.n7 a_52762_21071.n6 0.653
R10445 a_52762_21071.n3 a_52762_21071.n1 0.341
R10446 a_52762_21071.n6 a_52762_21071.n5 0.032
R10447 a_52999_20434.t0 a_52999_20434.t1 17.4
R10448 a_30152_10818.n1 a_30152_10818.t7 318.119
R10449 a_30152_10818.n1 a_30152_10818.t4 269.919
R10450 a_30152_10818.n0 a_30152_10818.t5 267.256
R10451 a_30152_10818.n0 a_30152_10818.t6 267.256
R10452 a_30152_10818.n4 a_30152_10818.n3 193.227
R10453 a_30152_10818.t7 a_30152_10818.n0 160.666
R10454 a_30152_10818.n2 a_30152_10818.n1 106.999
R10455 a_30152_10818.n3 a_30152_10818.t1 28.568
R10456 a_30152_10818.t0 a_30152_10818.n4 28.565
R10457 a_30152_10818.n4 a_30152_10818.t3 28.565
R10458 a_30152_10818.n2 a_30152_10818.t2 18.149
R10459 a_30152_10818.n3 a_30152_10818.n2 3.726
R10460 a_30645_10037.t0 a_30645_10037.n0 14.282
R10461 a_30645_10037.n0 a_30645_10037.t1 14.282
R10462 a_30645_10037.n0 a_30645_10037.n16 90.436
R10463 a_30645_10037.n16 a_30645_10037.n2 74.302
R10464 a_30645_10037.n2 a_30645_10037.n4 50.575
R10465 a_30645_10037.n4 a_30645_10037.n5 110.084
R10466 a_30645_10037.n16 a_30645_10037.n6 206.242
R10467 a_30645_10037.n6 a_30645_10037.n8 16.411
R10468 a_30645_10037.n8 a_30645_10037.t10 198.921
R10469 a_30645_10037.t10 a_30645_10037.t11 415.315
R10470 a_30645_10037.t11 a_30645_10037.n15 214.335
R10471 a_30645_10037.n15 a_30645_10037.t13 80.333
R10472 a_30645_10037.n15 a_30645_10037.t14 214.335
R10473 a_30645_10037.n8 a_30645_10037.n14 861.987
R10474 a_30645_10037.n14 a_30645_10037.n9 560.726
R10475 a_30645_10037.n14 a_30645_10037.n13 65.07
R10476 a_30645_10037.n13 a_30645_10037.n12 6.615
R10477 a_30645_10037.n12 a_30645_10037.t17 93.989
R10478 a_30645_10037.n13 a_30645_10037.n11 97.816
R10479 a_30645_10037.n11 a_30645_10037.t18 80.333
R10480 a_30645_10037.n11 a_30645_10037.t21 394.151
R10481 a_30645_10037.t21 a_30645_10037.n10 269.523
R10482 a_30645_10037.n10 a_30645_10037.t8 160.666
R10483 a_30645_10037.n10 a_30645_10037.t9 269.523
R10484 a_30645_10037.n12 a_30645_10037.t16 198.043
R10485 a_30645_10037.n9 a_30645_10037.t20 294.653
R10486 a_30645_10037.n9 a_30645_10037.t19 111.663
R10487 a_30645_10037.n6 a_30645_10037.t12 217.716
R10488 a_30645_10037.t12 a_30645_10037.t22 415.315
R10489 a_30645_10037.t22 a_30645_10037.n7 214.335
R10490 a_30645_10037.n7 a_30645_10037.t23 80.333
R10491 a_30645_10037.n7 a_30645_10037.t15 214.335
R10492 a_30645_10037.n5 a_30645_10037.t5 14.282
R10493 a_30645_10037.n5 a_30645_10037.t3 14.282
R10494 a_30645_10037.n4 a_30645_10037.n3 157.665
R10495 a_30645_10037.n3 a_30645_10037.t7 8.7
R10496 a_30645_10037.n3 a_30645_10037.t4 8.7
R10497 a_30645_10037.n2 a_30645_10037.n1 90.416
R10498 a_30645_10037.n1 a_30645_10037.t2 14.282
R10499 a_30645_10037.n1 a_30645_10037.t6 14.282
R10500 a_31377_10037.t0 a_31377_10037.t1 379.845
R10501 A[4].n29 A[4].n28 2886.86
R10502 A[4].n16 A[4].n6 1956.22
R10503 A[4].n6 A[4].n4 1494.07
R10504 A[4].n20 A[4].n19 1074.41
R10505 A[4].n20 A[4].t19 990.34
R10506 A[4].n19 A[4].t33 867.497
R10507 A[4].n36 A[4].n35 660.71
R10508 A[4].n19 A[4].t24 591.811
R10509 A[4].t59 A[4].t17 576.841
R10510 A[4].n11 A[4].n10 535.449
R10511 A[4].t46 A[4].t57 437.233
R10512 A[4].t45 A[4].t42 437.233
R10513 A[4].t48 A[4].t40 437.233
R10514 A[4].t39 A[4].t41 437.233
R10515 A[4].t9 A[4].t1 437.233
R10516 A[4].t43 A[4].t3 437.233
R10517 A[4].t21 A[4].t49 415.315
R10518 A[4].n26 A[4].n25 412.11
R10519 A[4].n20 A[4].t4 408.211
R10520 A[4].n23 A[4].t18 394.151
R10521 A[4].t28 A[4].n8 313.873
R10522 A[4].n10 A[4].t51 294.986
R10523 A[4].n25 A[4].t15 294.653
R10524 A[4].n17 A[4].t16 286.438
R10525 A[4].n17 A[4].t20 286.438
R10526 A[4].n18 A[4].t32 286.438
R10527 A[4].n18 A[4].t38 286.438
R10528 A[4].n31 A[4].t54 284.688
R10529 A[4].n7 A[4].t29 272.288
R10530 A[4].n22 A[4].t7 269.523
R10531 A[4].t18 A[4].n22 269.523
R10532 A[4].n11 A[4].t26 245.184
R10533 A[4].n3 A[4].t48 224.833
R10534 A[4].n26 A[4].n24 224.13
R10535 A[4].n33 A[4].t46 221.772
R10536 A[4].n4 A[4].t21 219.944
R10537 A[4].n13 A[4].t43 218.627
R10538 A[4].n6 A[4].t39 217.054
R10539 A[4].n15 A[4].t9 217.023
R10540 A[4].n3 A[4].t45 216.198
R10541 A[4].n30 A[4].t13 214.686
R10542 A[4].t57 A[4].n30 214.686
R10543 A[4].n2 A[4].t22 214.686
R10544 A[4].t42 A[4].n2 214.686
R10545 A[4].n1 A[4].t36 214.686
R10546 A[4].t40 A[4].n1 214.686
R10547 A[4].n5 A[4].t31 214.686
R10548 A[4].t41 A[4].n5 214.686
R10549 A[4].n14 A[4].t44 214.686
R10550 A[4].t1 A[4].n14 214.686
R10551 A[4].n12 A[4].t34 214.686
R10552 A[4].t3 A[4].n12 214.686
R10553 A[4].n0 A[4].t53 214.335
R10554 A[4].t49 A[4].n0 214.335
R10555 A[4].n21 A[4].t14 198.043
R10556 A[4].n9 A[4].t58 190.152
R10557 A[4].n9 A[4].t28 190.152
R10558 A[4].n27 A[4].t0 185.301
R10559 A[4].n27 A[4].t52 185.301
R10560 A[4].n33 A[4].n32 182.459
R10561 A[4].t19 A[4].n17 160.666
R10562 A[4].t33 A[4].n18 160.666
R10563 A[4].n31 A[4].t56 160.666
R10564 A[4].n32 A[4].t59 160.666
R10565 A[4].n22 A[4].t37 160.666
R10566 A[4].n7 A[4].t10 160.666
R10567 A[4].n8 A[4].t6 160.666
R10568 A[4].n29 A[4].n26 141.986
R10569 A[4].n28 A[4].t2 140.583
R10570 A[4].n32 A[4].n31 115.593
R10571 A[4].n25 A[4].t30 111.663
R10572 A[4].n10 A[4].t47 110.859
R10573 A[4].n27 A[4].t25 107.646
R10574 A[4].n24 A[4].n23 97.816
R10575 A[4].n8 A[4].n7 96.129
R10576 A[4].n21 A[4].t11 93.989
R10577 A[4].n30 A[4].t8 80.333
R10578 A[4].n23 A[4].t35 80.333
R10579 A[4].n0 A[4].t50 80.333
R10580 A[4].n2 A[4].t55 80.333
R10581 A[4].n1 A[4].t12 80.333
R10582 A[4].n5 A[4].t23 80.333
R10583 A[4].n14 A[4].t27 80.333
R10584 A[4].t26 A[4].n9 80.333
R10585 A[4].n12 A[4].t5 80.333
R10586 A[4].n28 A[4].n27 61.856
R10587 A[4].n16 A[4].n15 53.076
R10588 A[4] A[4].n36 53.033
R10589 A[4].n4 A[4].n3 34.046
R10590 A[4].n34 A[4].n33 33.949
R10591 A[4].n35 A[4].n20 21.17
R10592 A[4].n34 A[4].n29 19.007
R10593 A[4].n13 A[4].n11 14.9
R10594 A[4].n35 A[4].n34 11.896
R10595 A[4].n24 A[4].n21 6.615
R10596 A[4].n36 A[4].n16 4.819
R10597 A[4].n15 A[4].n13 2.599
R10598 a_5331_6357.n1 a_5331_6357.t7 990.34
R10599 a_5331_6357.n1 a_5331_6357.t5 408.211
R10600 a_5331_6357.n0 a_5331_6357.t4 286.438
R10601 a_5331_6357.n0 a_5331_6357.t6 286.438
R10602 a_5331_6357.n4 a_5331_6357.n3 197.272
R10603 a_5331_6357.t7 a_5331_6357.n0 160.666
R10604 a_5331_6357.n3 a_5331_6357.t0 28.568
R10605 a_5331_6357.t2 a_5331_6357.n4 28.565
R10606 a_5331_6357.n4 a_5331_6357.t1 28.565
R10607 a_5331_6357.n2 a_5331_6357.n1 25.661
R10608 a_5331_6357.n2 a_5331_6357.t3 18.103
R10609 a_5331_6357.n3 a_5331_6357.n2 0.459
R10610 a_53343_23888.t6 a_53343_23888.t5 800.071
R10611 a_53343_23888.n2 a_53343_23888.n1 659.097
R10612 a_53343_23888.n0 a_53343_23888.t4 285.109
R10613 a_53343_23888.n1 a_53343_23888.t6 193.602
R10614 a_53343_23888.n4 a_53343_23888.n3 192.754
R10615 a_53343_23888.n0 a_53343_23888.t7 160.666
R10616 a_53343_23888.n1 a_53343_23888.n0 91.507
R10617 a_53343_23888.n3 a_53343_23888.t3 28.568
R10618 a_53343_23888.n4 a_53343_23888.t2 28.565
R10619 a_53343_23888.t1 a_53343_23888.n4 28.565
R10620 a_53343_23888.n2 a_53343_23888.t0 19.061
R10621 a_53343_23888.n3 a_53343_23888.n2 1.005
R10622 a_55078_24197.n0 a_55078_24197.t1 14.282
R10623 a_55078_24197.n0 a_55078_24197.t5 14.282
R10624 a_55078_24197.n1 a_55078_24197.t2 14.282
R10625 a_55078_24197.n1 a_55078_24197.t0 14.282
R10626 a_55078_24197.n3 a_55078_24197.t4 14.282
R10627 a_55078_24197.t3 a_55078_24197.n3 14.282
R10628 a_55078_24197.n3 a_55078_24197.n2 2.546
R10629 a_55078_24197.n2 a_55078_24197.n1 2.367
R10630 a_55078_24197.n2 a_55078_24197.n0 0.001
R10631 a_51813_16162.n6 a_51813_16162.n5 501.28
R10632 a_51813_16162.t5 a_51813_16162.t15 437.233
R10633 a_51813_16162.t4 a_51813_16162.t12 415.315
R10634 a_51813_16162.t19 a_51813_16162.n3 313.873
R10635 a_51813_16162.n5 a_51813_16162.t18 294.986
R10636 a_51813_16162.n2 a_51813_16162.t14 272.288
R10637 a_51813_16162.n6 a_51813_16162.t11 236.009
R10638 a_51813_16162.n9 a_51813_16162.t5 216.627
R10639 a_51813_16162.n7 a_51813_16162.t4 216.111
R10640 a_51813_16162.n8 a_51813_16162.t17 214.686
R10641 a_51813_16162.t15 a_51813_16162.n8 214.686
R10642 a_51813_16162.n1 a_51813_16162.t7 214.335
R10643 a_51813_16162.t12 a_51813_16162.n1 214.335
R10644 a_51813_16162.n4 a_51813_16162.t8 190.152
R10645 a_51813_16162.n4 a_51813_16162.t19 190.152
R10646 a_51813_16162.n2 a_51813_16162.t13 160.666
R10647 a_51813_16162.n3 a_51813_16162.t10 160.666
R10648 a_51813_16162.n7 a_51813_16162.n6 148.428
R10649 a_51813_16162.n5 a_51813_16162.t6 110.859
R10650 a_51813_16162.n3 a_51813_16162.n2 96.129
R10651 a_51813_16162.n8 a_51813_16162.t16 80.333
R10652 a_51813_16162.n1 a_51813_16162.t9 80.333
R10653 a_51813_16162.t11 a_51813_16162.n4 80.333
R10654 a_51813_16162.n0 a_51813_16162.t3 28.57
R10655 a_51813_16162.n11 a_51813_16162.t2 28.565
R10656 a_51813_16162.t1 a_51813_16162.n11 28.565
R10657 a_51813_16162.n0 a_51813_16162.t0 17.638
R10658 a_51813_16162.n10 a_51813_16162.n9 5.55
R10659 a_51813_16162.n9 a_51813_16162.n7 2.923
R10660 a_51813_16162.n11 a_51813_16162.n10 0.693
R10661 a_51813_16162.n10 a_51813_16162.n0 0.597
R10662 a_56502_14835.t0 a_56502_14835.t1 17.4
R10663 a_61518_24201.t8 a_61518_24201.n2 404.877
R10664 a_61518_24201.n1 a_61518_24201.t7 210.902
R10665 a_61518_24201.n3 a_61518_24201.t8 136.943
R10666 a_61518_24201.n2 a_61518_24201.n1 107.801
R10667 a_61518_24201.n1 a_61518_24201.t6 80.333
R10668 a_61518_24201.n2 a_61518_24201.t5 80.333
R10669 a_61518_24201.n0 a_61518_24201.t4 17.4
R10670 a_61518_24201.n0 a_61518_24201.t1 17.4
R10671 a_61518_24201.n4 a_61518_24201.t2 15.032
R10672 a_61518_24201.t0 a_61518_24201.n5 14.282
R10673 a_61518_24201.n5 a_61518_24201.t3 14.282
R10674 a_61518_24201.n5 a_61518_24201.n4 1.65
R10675 a_61518_24201.n3 a_61518_24201.n0 0.672
R10676 a_61518_24201.n4 a_61518_24201.n3 0.665
R10677 a_61782_23618.t5 a_61782_23618.t7 800.071
R10678 a_61782_23618.n3 a_61782_23618.n2 672.951
R10679 a_61782_23618.n1 a_61782_23618.t4 285.109
R10680 a_61782_23618.n2 a_61782_23618.t5 193.602
R10681 a_61782_23618.n1 a_61782_23618.t6 160.666
R10682 a_61782_23618.n2 a_61782_23618.n1 91.507
R10683 a_61782_23618.t2 a_61782_23618.n4 28.57
R10684 a_61782_23618.n0 a_61782_23618.t0 28.565
R10685 a_61782_23618.n0 a_61782_23618.t1 28.565
R10686 a_61782_23618.n4 a_61782_23618.t3 17.638
R10687 a_61782_23618.n3 a_61782_23618.n0 0.69
R10688 a_61782_23618.n4 a_61782_23618.n3 0.6
R10689 A[7].n10 A[7].n9 2069.93
R10690 A[7].n1 A[7].t22 990.34
R10691 A[7].t38 A[7].t32 573.627
R10692 A[7].n21 A[7].n20 535.449
R10693 A[7].t3 A[7].t10 437.233
R10694 A[7].t16 A[7].t23 437.233
R10695 A[7].t8 A[7].t29 437.233
R10696 A[7].n26 A[7].n16 433.641
R10697 A[7].n7 A[7].n6 412.11
R10698 A[7].n1 A[7].t26 408.211
R10699 A[7].n4 A[7].t7 394.151
R10700 A[7].t28 A[7].n18 313.873
R10701 A[7].n20 A[7].t19 294.986
R10702 A[7].n6 A[7].t6 294.653
R10703 A[7].n0 A[7].t27 286.438
R10704 A[7].n0 A[7].t36 286.438
R10705 A[7].n12 A[7].t31 285.543
R10706 A[7].n17 A[7].t14 272.288
R10707 A[7].n3 A[7].t33 269.523
R10708 A[7].t7 A[7].n3 269.523
R10709 A[7].n21 A[7].t11 245.184
R10710 A[7].n7 A[7].n5 224.13
R10711 A[7].n14 A[7].t3 223.33
R10712 A[7].n23 A[7].t8 218.627
R10713 A[7].n25 A[7].t16 217.023
R10714 A[7].n11 A[7].t13 214.686
R10715 A[7].t10 A[7].n11 214.686
R10716 A[7].n24 A[7].t0 214.686
R10717 A[7].t23 A[7].n24 214.686
R10718 A[7].n22 A[7].t2 214.686
R10719 A[7].t29 A[7].n22 214.686
R10720 A[7].n2 A[7].t20 198.043
R10721 A[7].n19 A[7].t9 190.152
R10722 A[7].n19 A[7].t28 190.152
R10723 A[7].n8 A[7].t39 185.301
R10724 A[7].n8 A[7].t35 185.301
R10725 A[7].n14 A[7].n13 181.056
R10726 A[7].t22 A[7].n0 160.666
R10727 A[7].n3 A[7].t18 160.666
R10728 A[7].n12 A[7].t37 160.666
R10729 A[7].n13 A[7].t38 160.666
R10730 A[7].n17 A[7].t4 160.666
R10731 A[7].n18 A[7].t1 160.666
R10732 A[7].n10 A[7].n7 142.556
R10733 A[7].n9 A[7].t25 137.369
R10734 A[7].n13 A[7].n12 114.089
R10735 A[7].n6 A[7].t15 111.663
R10736 A[7].n20 A[7].t5 110.859
R10737 A[7].n8 A[7].t21 107.646
R10738 A[7].n5 A[7].n4 97.816
R10739 A[7].n18 A[7].n17 96.129
R10740 A[7].n2 A[7].t34 93.989
R10741 A[7].n4 A[7].t17 80.333
R10742 A[7].n11 A[7].t12 80.333
R10743 A[7].n24 A[7].t24 80.333
R10744 A[7].t11 A[7].n19 80.333
R10745 A[7].n22 A[7].t30 80.333
R10746 A[7].n9 A[7].n8 61.856
R10747 A[7] A[7].n26 49.563
R10748 A[7].n16 A[7].n1 48.482
R10749 A[7].n15 A[7].n14 42.073
R10750 A[7].n26 A[7].n25 32.836
R10751 A[7].n15 A[7].n10 32.163
R10752 A[7].n23 A[7].n21 14.9
R10753 A[7].n16 A[7].n15 9.006
R10754 A[7].n5 A[7].n2 6.615
R10755 A[7].n25 A[7].n23 2.599
R10756 a_42770_18699.n0 a_42770_18699.t10 214.335
R10757 a_42770_18699.t9 a_42770_18699.n0 214.335
R10758 a_42770_18699.n1 a_42770_18699.t9 143.851
R10759 a_42770_18699.n1 a_42770_18699.t8 135.658
R10760 a_42770_18699.n0 a_42770_18699.t7 80.333
R10761 a_42770_18699.n4 a_42770_18699.t3 28.565
R10762 a_42770_18699.n4 a_42770_18699.t1 28.565
R10763 a_42770_18699.n2 a_42770_18699.t6 28.565
R10764 a_42770_18699.n2 a_42770_18699.t5 28.565
R10765 a_42770_18699.n7 a_42770_18699.t2 28.565
R10766 a_42770_18699.t0 a_42770_18699.n7 28.565
R10767 a_42770_18699.n5 a_42770_18699.t4 9.714
R10768 a_42770_18699.n5 a_42770_18699.n4 1.003
R10769 a_42770_18699.n6 a_42770_18699.n3 0.833
R10770 a_42770_18699.n3 a_42770_18699.n2 0.653
R10771 a_42770_18699.n7 a_42770_18699.n6 0.653
R10772 a_42770_18699.n6 a_42770_18699.n5 0.341
R10773 a_42770_18699.n3 a_42770_18699.n1 0.032
R10774 a_62375_18703.n0 a_62375_18703.t8 214.335
R10775 a_62375_18703.t10 a_62375_18703.n0 214.335
R10776 a_62375_18703.n1 a_62375_18703.t10 143.851
R10777 a_62375_18703.n1 a_62375_18703.t7 135.658
R10778 a_62375_18703.n0 a_62375_18703.t9 80.333
R10779 a_62375_18703.n2 a_62375_18703.t3 28.565
R10780 a_62375_18703.n2 a_62375_18703.t4 28.565
R10781 a_62375_18703.n4 a_62375_18703.t5 28.565
R10782 a_62375_18703.n4 a_62375_18703.t2 28.565
R10783 a_62375_18703.n7 a_62375_18703.t1 28.565
R10784 a_62375_18703.t0 a_62375_18703.n7 28.565
R10785 a_62375_18703.n3 a_62375_18703.t6 9.714
R10786 a_62375_18703.n3 a_62375_18703.n2 1.003
R10787 a_62375_18703.n6 a_62375_18703.n5 0.833
R10788 a_62375_18703.n5 a_62375_18703.n4 0.653
R10789 a_62375_18703.n7 a_62375_18703.n6 0.653
R10790 a_62375_18703.n5 a_62375_18703.n3 0.341
R10791 a_62375_18703.n6 a_62375_18703.n1 0.032
R10792 a_47794_3876.t6 a_47794_3876.n3 404.877
R10793 a_47794_3876.n2 a_47794_3876.t7 210.902
R10794 a_47794_3876.n4 a_47794_3876.t6 136.943
R10795 a_47794_3876.n3 a_47794_3876.n2 107.801
R10796 a_47794_3876.n2 a_47794_3876.t5 80.333
R10797 a_47794_3876.n3 a_47794_3876.t8 80.333
R10798 a_47794_3876.n1 a_47794_3876.t1 17.4
R10799 a_47794_3876.n1 a_47794_3876.t2 17.4
R10800 a_47794_3876.t0 a_47794_3876.n5 15.032
R10801 a_47794_3876.n0 a_47794_3876.t3 14.282
R10802 a_47794_3876.n0 a_47794_3876.t4 14.282
R10803 a_47794_3876.n5 a_47794_3876.n0 1.65
R10804 a_47794_3876.n4 a_47794_3876.n1 0.672
R10805 a_47794_3876.n5 a_47794_3876.n4 0.665
R10806 a_59635_6910.n0 a_59635_6910.t1 14.282
R10807 a_59635_6910.t0 a_59635_6910.n0 14.282
R10808 a_59635_6910.n0 a_59635_6910.n12 90.436
R10809 a_59635_6910.n8 a_59635_6910.n11 50.575
R10810 a_59635_6910.n12 a_59635_6910.n8 74.302
R10811 a_59635_6910.n11 a_59635_6910.n10 157.665
R10812 a_59635_6910.n10 a_59635_6910.t4 8.7
R10813 a_59635_6910.n10 a_59635_6910.t7 8.7
R10814 a_59635_6910.n11 a_59635_6910.n9 122.999
R10815 a_59635_6910.n9 a_59635_6910.t6 14.282
R10816 a_59635_6910.n9 a_59635_6910.t5 14.282
R10817 a_59635_6910.n8 a_59635_6910.n7 90.416
R10818 a_59635_6910.n7 a_59635_6910.t3 14.282
R10819 a_59635_6910.n7 a_59635_6910.t2 14.282
R10820 a_59635_6910.n12 a_59635_6910.n1 342.688
R10821 a_59635_6910.n1 a_59635_6910.n6 126.566
R10822 a_59635_6910.n6 a_59635_6910.t9 294.653
R10823 a_59635_6910.n6 a_59635_6910.t14 111.663
R10824 a_59635_6910.n1 a_59635_6910.n5 552.333
R10825 a_59635_6910.n5 a_59635_6910.n4 6.615
R10826 a_59635_6910.n4 a_59635_6910.t12 93.989
R10827 a_59635_6910.n5 a_59635_6910.n3 97.816
R10828 a_59635_6910.n3 a_59635_6910.t10 80.333
R10829 a_59635_6910.n3 a_59635_6910.t11 394.151
R10830 a_59635_6910.t11 a_59635_6910.n2 269.523
R10831 a_59635_6910.n2 a_59635_6910.t8 160.666
R10832 a_59635_6910.n2 a_59635_6910.t13 269.523
R10833 a_59635_6910.n4 a_59635_6910.t15 198.043
R10834 a_61415_6910.t3 a_61415_6910.n0 14.282
R10835 a_61415_6910.n0 a_61415_6910.t4 14.282
R10836 a_61415_6910.n0 a_61415_6910.n9 0.999
R10837 a_61415_6910.n9 a_61415_6910.n6 0.575
R10838 a_61415_6910.n6 a_61415_6910.n8 0.2
R10839 a_61415_6910.n8 a_61415_6910.t8 16.058
R10840 a_61415_6910.n8 a_61415_6910.n7 0.999
R10841 a_61415_6910.n7 a_61415_6910.t9 14.282
R10842 a_61415_6910.n7 a_61415_6910.t10 14.282
R10843 a_61415_6910.n9 a_61415_6910.t5 16.058
R10844 a_61415_6910.n6 a_61415_6910.n4 0.227
R10845 a_61415_6910.n4 a_61415_6910.n5 1.511
R10846 a_61415_6910.n5 a_61415_6910.t1 14.282
R10847 a_61415_6910.n5 a_61415_6910.t2 14.282
R10848 a_61415_6910.n4 a_61415_6910.n1 0.669
R10849 a_61415_6910.n1 a_61415_6910.n2 0.001
R10850 a_61415_6910.n1 a_61415_6910.n3 267.767
R10851 a_61415_6910.n3 a_61415_6910.t11 14.282
R10852 a_61415_6910.n3 a_61415_6910.t7 14.282
R10853 a_61415_6910.n2 a_61415_6910.t0 14.282
R10854 a_61415_6910.n2 a_61415_6910.t6 14.282
R10855 a_44460_6616.n0 a_44460_6616.t7 214.335
R10856 a_44460_6616.t10 a_44460_6616.n0 214.335
R10857 a_44460_6616.n1 a_44460_6616.t10 143.851
R10858 a_44460_6616.n1 a_44460_6616.t8 135.658
R10859 a_44460_6616.n0 a_44460_6616.t9 80.333
R10860 a_44460_6616.n2 a_44460_6616.t5 28.565
R10861 a_44460_6616.n2 a_44460_6616.t4 28.565
R10862 a_44460_6616.n4 a_44460_6616.t6 28.565
R10863 a_44460_6616.n4 a_44460_6616.t2 28.565
R10864 a_44460_6616.t0 a_44460_6616.n7 28.565
R10865 a_44460_6616.n7 a_44460_6616.t1 28.565
R10866 a_44460_6616.n6 a_44460_6616.t3 9.714
R10867 a_44460_6616.n7 a_44460_6616.n6 1.003
R10868 a_44460_6616.n5 a_44460_6616.n3 0.833
R10869 a_44460_6616.n3 a_44460_6616.n2 0.653
R10870 a_44460_6616.n5 a_44460_6616.n4 0.653
R10871 a_44460_6616.n6 a_44460_6616.n5 0.341
R10872 a_44460_6616.n3 a_44460_6616.n1 0.032
R10873 a_53816_17942.t6 a_53816_17942.n2 404.877
R10874 a_53816_17942.n1 a_53816_17942.t8 210.902
R10875 a_53816_17942.n3 a_53816_17942.t6 136.949
R10876 a_53816_17942.n2 a_53816_17942.n1 107.801
R10877 a_53816_17942.n1 a_53816_17942.t5 80.333
R10878 a_53816_17942.n2 a_53816_17942.t7 80.333
R10879 a_53816_17942.n0 a_53816_17942.t4 17.4
R10880 a_53816_17942.n0 a_53816_17942.t0 17.4
R10881 a_53816_17942.n4 a_53816_17942.t3 15.032
R10882 a_53816_17942.n5 a_53816_17942.t2 14.282
R10883 a_53816_17942.t1 a_53816_17942.n5 14.282
R10884 a_53816_17942.n5 a_53816_17942.n4 1.65
R10885 a_53816_17942.n3 a_53816_17942.n0 0.657
R10886 a_53816_17942.n4 a_53816_17942.n3 0.614
R10887 a_52749_18576.t7 a_52749_18576.t4 800.071
R10888 a_52749_18576.n3 a_52749_18576.n2 672.95
R10889 a_52749_18576.n1 a_52749_18576.t5 285.109
R10890 a_52749_18576.n2 a_52749_18576.t7 193.602
R10891 a_52749_18576.n1 a_52749_18576.t6 160.666
R10892 a_52749_18576.n2 a_52749_18576.n1 91.507
R10893 a_52749_18576.n0 a_52749_18576.t1 28.57
R10894 a_52749_18576.t2 a_52749_18576.n4 28.565
R10895 a_52749_18576.n4 a_52749_18576.t0 28.565
R10896 a_52749_18576.n0 a_52749_18576.t3 17.638
R10897 a_52749_18576.n4 a_52749_18576.n3 0.693
R10898 a_52749_18576.n3 a_52749_18576.n0 0.597
R10899 B[0].t7 B[0].t23 802.481
R10900 B[0].n3 B[0].n1 653.736
R10901 B[0].n8 B[0].n7 618.566
R10902 B[0].n14 B[0].n10 592.056
R10903 B[0].t16 B[0].t21 415.315
R10904 B[0].t12 B[0].n5 313.873
R10905 B[0].t18 B[0].n12 313.069
R10906 B[0].n10 B[0].t0 294.986
R10907 B[0].n0 B[0].t5 284.688
R10908 B[0].n7 B[0].t3 273.077
R10909 B[0].n4 B[0].t10 272.288
R10910 B[0].n11 B[0].t19 271.484
R10911 B[0].n3 B[0].t16 218.405
R10912 B[0].n2 B[0].t14 214.335
R10913 B[0].t21 B[0].n2 214.335
R10914 B[0].n8 B[0].t17 204.679
R10915 B[0].n14 B[0].t9 204.672
R10916 B[0].n1 B[0].t7 192.799
R10917 B[0].n13 B[0].t18 190.955
R10918 B[0].n13 B[0].t22 190.955
R10919 B[0].n6 B[0].t1 190.152
R10920 B[0].n6 B[0].t12 190.152
R10921 B[0].n0 B[0].t6 160.666
R10922 B[0].n4 B[0].t15 160.666
R10923 B[0].n5 B[0].t8 160.666
R10924 B[0].n12 B[0].t4 160.666
R10925 B[0].n11 B[0].t11 160.666
R10926 B[0].n7 B[0].t13 137.369
R10927 B[0].n10 B[0].t2 110.859
R10928 B[0].n5 B[0].n4 96.129
R10929 B[0].n12 B[0].n11 96.129
R10930 B[0].n1 B[0].n0 91.889
R10931 B[0].n2 B[0].t20 80.333
R10932 B[0].t17 B[0].n6 80.333
R10933 B[0].t9 B[0].n13 80.333
R10934 B[0] B[0].n15 49.826
R10935 B[0].n9 B[0].n8 49.449
R10936 B[0].n15 B[0].n14 48.886
R10937 B[0].n15 B[0].n9 2.694
R10938 B[0].n9 B[0].n3 0.639
R10939 a_31379_12341.t0 a_31379_12341.t1 17.4
R10940 a_4857_n2637.n1 a_4857_n2637.t5 867.497
R10941 a_4857_n2637.n1 a_4857_n2637.t7 615.911
R10942 a_4857_n2637.n0 a_4857_n2637.t4 286.438
R10943 a_4857_n2637.n0 a_4857_n2637.t6 286.438
R10944 a_4857_n2637.n4 a_4857_n2637.n3 185.55
R10945 a_4857_n2637.t5 a_4857_n2637.n0 160.666
R10946 a_4857_n2637.n3 a_4857_n2637.t2 28.568
R10947 a_4857_n2637.n4 a_4857_n2637.t3 28.565
R10948 a_4857_n2637.t1 a_4857_n2637.n4 28.565
R10949 a_4857_n2637.n2 a_4857_n2637.n1 22.356
R10950 a_4857_n2637.n2 a_4857_n2637.t0 20.393
R10951 a_4857_n2637.n3 a_4857_n2637.n2 2.038
R10952 a_3983_n2152.n0 a_3983_n2152.n9 167.433
R10953 a_3983_n2152.n0 a_3983_n2152.t1 14.282
R10954 a_3983_n2152.t0 a_3983_n2152.n0 14.282
R10955 a_3983_n2152.n9 a_3983_n2152.n8 75.815
R10956 a_3983_n2152.n8 a_3983_n2152.n6 77.456
R10957 a_3983_n2152.n6 a_3983_n2152.n4 77.456
R10958 a_3983_n2152.n4 a_3983_n2152.n2 77.784
R10959 a_3983_n2152.n9 a_3983_n2152.t2 104.259
R10960 a_3983_n2152.n8 a_3983_n2152.n7 89.977
R10961 a_3983_n2152.n7 a_3983_n2152.t3 14.282
R10962 a_3983_n2152.n7 a_3983_n2152.t10 14.282
R10963 a_3983_n2152.n6 a_3983_n2152.n5 89.977
R10964 a_3983_n2152.n5 a_3983_n2152.t11 14.282
R10965 a_3983_n2152.n5 a_3983_n2152.t7 14.282
R10966 a_3983_n2152.n4 a_3983_n2152.n3 89.977
R10967 a_3983_n2152.n3 a_3983_n2152.t8 14.282
R10968 a_3983_n2152.n3 a_3983_n2152.t9 14.282
R10969 a_3983_n2152.n2 a_3983_n2152.t6 104.259
R10970 a_3983_n2152.n2 a_3983_n2152.n1 167.433
R10971 a_3983_n2152.n1 a_3983_n2152.t5 14.282
R10972 a_3983_n2152.n1 a_3983_n2152.t4 14.282
R10973 a_4332_n2152.t1 a_4332_n2152.n0 14.283
R10974 a_4332_n2152.n0 a_4332_n2152.n7 4.366
R10975 a_4332_n2152.n7 a_4332_n2152.n5 0.852
R10976 a_4332_n2152.n5 a_4332_n2152.n6 258.161
R10977 a_4332_n2152.n6 a_4332_n2152.t4 14.282
R10978 a_4332_n2152.n6 a_4332_n2152.t3 14.282
R10979 a_4332_n2152.n5 a_4332_n2152.t2 14.283
R10980 a_4332_n2152.n7 a_4332_n2152.n4 97.614
R10981 a_4332_n2152.n4 a_4332_n2152.t9 200.029
R10982 a_4332_n2152.t9 a_4332_n2152.n3 206.421
R10983 a_4332_n2152.n3 a_4332_n2152.t8 80.333
R10984 a_4332_n2152.n3 a_4332_n2152.t10 206.421
R10985 a_4332_n2152.n4 a_4332_n2152.t11 1527.4
R10986 a_4332_n2152.t11 a_4332_n2152.n2 657.379
R10987 a_4332_n2152.n2 a_4332_n2152.t5 8.7
R10988 a_4332_n2152.n2 a_4332_n2152.t0 8.7
R10989 a_4332_n2152.n0 a_4332_n2152.n1 258.161
R10990 a_4332_n2152.n1 a_4332_n2152.t6 14.282
R10991 a_4332_n2152.n1 a_4332_n2152.t7 14.282
R10992 a_45049_1913.t7 a_45049_1913.t4 574.43
R10993 a_45049_1913.n0 a_45049_1913.t5 285.109
R10994 a_45049_1913.n2 a_45049_1913.n1 211.136
R10995 a_45049_1913.n4 a_45049_1913.n3 192.754
R10996 a_45049_1913.n0 a_45049_1913.t6 160.666
R10997 a_45049_1913.n1 a_45049_1913.t7 160.666
R10998 a_45049_1913.n1 a_45049_1913.n0 114.829
R10999 a_45049_1913.n3 a_45049_1913.t2 28.568
R11000 a_45049_1913.n4 a_45049_1913.t3 28.565
R11001 a_45049_1913.t1 a_45049_1913.n4 28.565
R11002 a_45049_1913.n2 a_45049_1913.t0 19.084
R11003 a_45049_1913.n3 a_45049_1913.n2 1.051
R11004 a_1735_13585.n3 a_1735_13585.t7 448.381
R11005 a_1735_13585.n2 a_1735_13585.t6 286.438
R11006 a_1735_13585.n2 a_1735_13585.t5 286.438
R11007 a_1735_13585.n1 a_1735_13585.t4 247.69
R11008 a_1735_13585.n4 a_1735_13585.n0 182.117
R11009 a_1735_13585.t7 a_1735_13585.n2 160.666
R11010 a_1735_13585.t0 a_1735_13585.n4 28.568
R11011 a_1735_13585.n0 a_1735_13585.t3 28.565
R11012 a_1735_13585.n0 a_1735_13585.t2 28.565
R11013 a_1735_13585.n1 a_1735_13585.t1 18.127
R11014 a_1735_13585.n3 a_1735_13585.n1 4.036
R11015 a_1735_13585.n4 a_1735_13585.n3 0.937
R11016 a_1680_13125.t0 a_1680_13125.t1 17.4
R11017 a_556_13728.t0 a_556_13728.n0 14.283
R11018 a_556_13728.n0 a_556_13728.n5 0.852
R11019 a_556_13728.n5 a_556_13728.n6 4.366
R11020 a_556_13728.n6 a_556_13728.n7 258.161
R11021 a_556_13728.n7 a_556_13728.t5 14.282
R11022 a_556_13728.n7 a_556_13728.t4 14.282
R11023 a_556_13728.n6 a_556_13728.t6 14.283
R11024 a_556_13728.n5 a_556_13728.n4 97.614
R11025 a_556_13728.n4 a_556_13728.t9 200.029
R11026 a_556_13728.t9 a_556_13728.n3 206.421
R11027 a_556_13728.n3 a_556_13728.t10 80.333
R11028 a_556_13728.n3 a_556_13728.t11 206.421
R11029 a_556_13728.n4 a_556_13728.t8 1527.4
R11030 a_556_13728.t8 a_556_13728.n2 657.379
R11031 a_556_13728.n2 a_556_13728.t3 8.7
R11032 a_556_13728.n2 a_556_13728.t7 8.7
R11033 a_556_13728.n0 a_556_13728.n1 258.161
R11034 a_556_13728.n1 a_556_13728.t1 14.282
R11035 a_556_13728.n1 a_556_13728.t2 14.282
R11036 opcode[2].n1 opcode[2].t10 1374.12
R11037 opcode[2].n8 opcode[2].t53 1374.12
R11038 opcode[2].n13 opcode[2].t24 1374.12
R11039 opcode[2].n18 opcode[2].t59 1374.12
R11040 opcode[2].n23 opcode[2].t21 1374.12
R11041 opcode[2].n28 opcode[2].t12 1374.12
R11042 opcode[2].n33 opcode[2].t36 1374.12
R11043 opcode[2].n38 opcode[2].t7 1374.12
R11044 opcode[2].n3 opcode[2].t9 623.291
R11045 opcode[2].n6 opcode[2].t33 623.291
R11046 opcode[2].n11 opcode[2].t56 623.291
R11047 opcode[2].n16 opcode[2].t2 623.291
R11048 opcode[2].n21 opcode[2].t30 623.291
R11049 opcode[2].n26 opcode[2].t61 623.291
R11050 opcode[2].n31 opcode[2].t17 623.291
R11051 opcode[2].n36 opcode[2].t19 623.291
R11052 opcode[2].n3 opcode[2].t44 610.283
R11053 opcode[2].n6 opcode[2].t22 610.283
R11054 opcode[2].n11 opcode[2].t52 610.283
R11055 opcode[2].n16 opcode[2].t27 610.283
R11056 opcode[2].n21 opcode[2].t35 610.283
R11057 opcode[2].n26 opcode[2].t32 610.283
R11058 opcode[2].n31 opcode[2].t63 610.283
R11059 opcode[2].n36 opcode[2].t42 610.283
R11060 opcode[2].n40 opcode[2].n39 490.666
R11061 opcode[2].n43 opcode[2].n42 333.008
R11062 opcode[2].n42 opcode[2].n41 327.284
R11063 opcode[2].n44 opcode[2].n43 327.284
R11064 opcode[2].n46 opcode[2].n45 326.243
R11065 opcode[2].n45 opcode[2].n44 326.139
R11066 opcode[2].n1 opcode[2].t49 326.034
R11067 opcode[2].n8 opcode[2].t58 326.034
R11068 opcode[2].n13 opcode[2].t25 326.034
R11069 opcode[2].n18 opcode[2].t26 326.034
R11070 opcode[2].n23 opcode[2].t37 326.034
R11071 opcode[2].n28 opcode[2].t28 326.034
R11072 opcode[2].n33 opcode[2].t39 326.034
R11073 opcode[2].n38 opcode[2].t48 326.034
R11074 opcode[2].n41 opcode[2].n40 325.931
R11075 opcode[2].n2 opcode[2].t34 286.438
R11076 opcode[2].n2 opcode[2].t41 286.438
R11077 opcode[2].n5 opcode[2].t51 286.438
R11078 opcode[2].n5 opcode[2].t54 286.438
R11079 opcode[2].n10 opcode[2].t11 286.438
R11080 opcode[2].n10 opcode[2].t57 286.438
R11081 opcode[2].n15 opcode[2].t20 286.438
R11082 opcode[2].n15 opcode[2].t47 286.438
R11083 opcode[2].n20 opcode[2].t15 286.438
R11084 opcode[2].n20 opcode[2].t5 286.438
R11085 opcode[2].n25 opcode[2].t18 286.438
R11086 opcode[2].n25 opcode[2].t43 286.438
R11087 opcode[2].n30 opcode[2].t40 286.438
R11088 opcode[2].n30 opcode[2].t45 286.438
R11089 opcode[2].n35 opcode[2].t55 286.438
R11090 opcode[2].n35 opcode[2].t62 286.438
R11091 opcode[2] opcode[2].n46 221.469
R11092 opcode[2].n0 opcode[2].t6 206.421
R11093 opcode[2].t49 opcode[2].n0 206.421
R11094 opcode[2].n7 opcode[2].t0 206.421
R11095 opcode[2].t58 opcode[2].n7 206.421
R11096 opcode[2].n12 opcode[2].t8 206.421
R11097 opcode[2].t25 opcode[2].n12 206.421
R11098 opcode[2].n17 opcode[2].t46 206.421
R11099 opcode[2].t26 opcode[2].n17 206.421
R11100 opcode[2].n22 opcode[2].t13 206.421
R11101 opcode[2].t37 opcode[2].n22 206.421
R11102 opcode[2].n27 opcode[2].t14 206.421
R11103 opcode[2].t28 opcode[2].n27 206.421
R11104 opcode[2].n32 opcode[2].t60 206.421
R11105 opcode[2].t39 opcode[2].n32 206.421
R11106 opcode[2].n37 opcode[2].t4 206.421
R11107 opcode[2].t48 opcode[2].n37 206.421
R11108 opcode[2].n45 opcode[2].n9 171.411
R11109 opcode[2].n41 opcode[2].n29 164.146
R11110 opcode[2].n44 opcode[2].n14 164.04
R11111 opcode[2].n40 opcode[2].n34 162.638
R11112 opcode[2].n42 opcode[2].n24 161.961
R11113 opcode[2].t9 opcode[2].n2 160.666
R11114 opcode[2].t33 opcode[2].n5 160.666
R11115 opcode[2].t56 opcode[2].n10 160.666
R11116 opcode[2].t2 opcode[2].n15 160.666
R11117 opcode[2].t30 opcode[2].n20 160.666
R11118 opcode[2].t61 opcode[2].n25 160.666
R11119 opcode[2].t17 opcode[2].n30 160.666
R11120 opcode[2].t19 opcode[2].n35 160.666
R11121 opcode[2].n43 opcode[2].n19 157.479
R11122 opcode[2].n46 opcode[2].n4 155.498
R11123 opcode[2].n0 opcode[2].t31 80.333
R11124 opcode[2].n7 opcode[2].t23 80.333
R11125 opcode[2].n12 opcode[2].t50 80.333
R11126 opcode[2].n17 opcode[2].t1 80.333
R11127 opcode[2].n22 opcode[2].t38 80.333
R11128 opcode[2].n27 opcode[2].t3 80.333
R11129 opcode[2].n32 opcode[2].t16 80.333
R11130 opcode[2].n37 opcode[2].t29 80.333
R11131 opcode[2] opcode[2].n47 17.018
R11132 opcode[2].n47 opcode[2] 16.924
R11133 opcode[2].n9 opcode[2].n6 1.617
R11134 opcode[2].n14 opcode[2].n11 1.617
R11135 opcode[2].n19 opcode[2].n16 1.617
R11136 opcode[2].n24 opcode[2].n21 1.617
R11137 opcode[2].n29 opcode[2].n26 1.617
R11138 opcode[2].n34 opcode[2].n31 1.617
R11139 opcode[2].n39 opcode[2].n36 1.617
R11140 opcode[2].n4 opcode[2].n3 1.616
R11141 opcode[2].n47 opcode[2] 1.144
R11142 opcode[2].n47 opcode[2] 1.137
R11143 opcode[2].n4 opcode[2].n1 0.003
R11144 opcode[2].n9 opcode[2].n8 0.003
R11145 opcode[2].n14 opcode[2].n13 0.003
R11146 opcode[2].n19 opcode[2].n18 0.003
R11147 opcode[2].n24 opcode[2].n23 0.003
R11148 opcode[2].n29 opcode[2].n28 0.003
R11149 opcode[2].n34 opcode[2].n33 0.003
R11150 opcode[2].n39 opcode[2].n38 0.003
R11151 a_3392_1740.n2 a_3392_1740.t7 448.382
R11152 a_3392_1740.n1 a_3392_1740.t4 286.438
R11153 a_3392_1740.n1 a_3392_1740.t5 286.438
R11154 a_3392_1740.n0 a_3392_1740.t6 247.69
R11155 a_3392_1740.n4 a_3392_1740.n3 182.117
R11156 a_3392_1740.t7 a_3392_1740.n1 160.666
R11157 a_3392_1740.n3 a_3392_1740.t0 28.568
R11158 a_3392_1740.t2 a_3392_1740.n4 28.565
R11159 a_3392_1740.n4 a_3392_1740.t1 28.565
R11160 a_3392_1740.n0 a_3392_1740.t3 18.127
R11161 a_3392_1740.n2 a_3392_1740.n0 4.039
R11162 a_3392_1740.n3 a_3392_1740.n2 0.937
R11163 a_4183_8966.t0 a_4183_8966.n0 14.282
R11164 a_4183_8966.n0 a_4183_8966.t6 14.282
R11165 a_4183_8966.n0 a_4183_8966.n8 90.416
R11166 a_4183_8966.n8 a_4183_8966.n5 74.302
R11167 a_4183_8966.n8 a_4183_8966.n7 50.575
R11168 a_4183_8966.n7 a_4183_8966.n6 157.665
R11169 a_4183_8966.n6 a_4183_8966.t3 8.7
R11170 a_4183_8966.n6 a_4183_8966.t5 8.7
R11171 a_4183_8966.n5 a_4183_8966.n4 90.436
R11172 a_4183_8966.n4 a_4183_8966.t2 14.282
R11173 a_4183_8966.n4 a_4183_8966.t1 14.282
R11174 a_4183_8966.n7 a_4183_8966.n3 122.746
R11175 a_4183_8966.n3 a_4183_8966.t4 14.282
R11176 a_4183_8966.n3 a_4183_8966.t7 14.282
R11177 a_4183_8966.n5 a_4183_8966.n1 1832.15
R11178 a_4183_8966.n1 a_4183_8966.t10 591.811
R11179 a_4183_8966.n1 a_4183_8966.t11 867.497
R11180 a_4183_8966.t11 a_4183_8966.n2 160.666
R11181 a_4183_8966.n2 a_4183_8966.t8 286.438
R11182 a_4183_8966.n2 a_4183_8966.t9 286.438
R11183 a_3710_8262.t0 a_3710_8262.n0 14.282
R11184 a_3710_8262.n0 a_3710_8262.t2 14.282
R11185 a_3710_8262.n0 a_3710_8262.n1 258.161
R11186 a_3710_8262.n1 a_3710_8262.n5 0.852
R11187 a_3710_8262.n5 a_3710_8262.n6 4.366
R11188 a_3710_8262.n6 a_3710_8262.n7 258.161
R11189 a_3710_8262.n7 a_3710_8262.t4 14.282
R11190 a_3710_8262.n7 a_3710_8262.t7 14.282
R11191 a_3710_8262.n6 a_3710_8262.t6 14.283
R11192 a_3710_8262.n5 a_3710_8262.n4 97.614
R11193 a_3710_8262.n4 a_3710_8262.t10 200.029
R11194 a_3710_8262.t10 a_3710_8262.n3 206.421
R11195 a_3710_8262.n3 a_3710_8262.t8 80.333
R11196 a_3710_8262.n3 a_3710_8262.t11 206.421
R11197 a_3710_8262.n4 a_3710_8262.t9 1527.4
R11198 a_3710_8262.t9 a_3710_8262.n2 657.379
R11199 a_3710_8262.n2 a_3710_8262.t5 8.7
R11200 a_3710_8262.n2 a_3710_8262.t3 8.7
R11201 a_3710_8262.n1 a_3710_8262.t1 14.283
R11202 a_4243_8992.t0 a_4243_8992.n0 14.282
R11203 a_4243_8992.n0 a_4243_8992.t2 14.282
R11204 a_4243_8992.n7 a_4243_8992.n8 77.784
R11205 a_4243_8992.n5 a_4243_8992.n7 77.456
R11206 a_4243_8992.n3 a_4243_8992.n5 77.456
R11207 a_4243_8992.n1 a_4243_8992.n3 75.815
R11208 a_4243_8992.n0 a_4243_8992.n1 167.433
R11209 a_4243_8992.n8 a_4243_8992.n9 167.433
R11210 a_4243_8992.n9 a_4243_8992.t5 14.282
R11211 a_4243_8992.n9 a_4243_8992.t4 14.282
R11212 a_4243_8992.n8 a_4243_8992.t6 104.259
R11213 a_4243_8992.n7 a_4243_8992.n6 89.977
R11214 a_4243_8992.n6 a_4243_8992.t3 14.282
R11215 a_4243_8992.n6 a_4243_8992.t7 14.282
R11216 a_4243_8992.n5 a_4243_8992.n4 89.977
R11217 a_4243_8992.n4 a_4243_8992.t11 14.282
R11218 a_4243_8992.n4 a_4243_8992.t8 14.282
R11219 a_4243_8992.n3 a_4243_8992.n2 89.977
R11220 a_4243_8992.n2 a_4243_8992.t10 14.282
R11221 a_4243_8992.n2 a_4243_8992.t9 14.282
R11222 a_4243_8992.n1 a_4243_8992.t1 104.259
R11223 a_70513_7304.t1 a_70513_7304.n0 14.283
R11224 a_70513_7304.n0 a_70513_7304.n7 258.161
R11225 a_70513_7304.n7 a_70513_7304.t2 14.282
R11226 a_70513_7304.n7 a_70513_7304.t3 14.282
R11227 a_70513_7304.n0 a_70513_7304.n4 0.852
R11228 a_70513_7304.n4 a_70513_7304.n5 4.366
R11229 a_70513_7304.n5 a_70513_7304.n6 258.161
R11230 a_70513_7304.n6 a_70513_7304.t6 14.282
R11231 a_70513_7304.n6 a_70513_7304.t7 14.282
R11232 a_70513_7304.n5 a_70513_7304.t4 14.283
R11233 a_70513_7304.n4 a_70513_7304.n3 73.514
R11234 a_70513_7304.n3 a_70513_7304.t11 1551.5
R11235 a_70513_7304.t11 a_70513_7304.n2 656.576
R11236 a_70513_7304.n2 a_70513_7304.t5 8.7
R11237 a_70513_7304.n2 a_70513_7304.t0 8.7
R11238 a_70513_7304.n3 a_70513_7304.t8 224.129
R11239 a_70513_7304.t8 a_70513_7304.n1 207.225
R11240 a_70513_7304.n1 a_70513_7304.t10 207.225
R11241 a_70513_7304.n1 a_70513_7304.t9 80.333
R11242 a_11101_1259.n3 a_11101_1259.t5 867.497
R11243 a_11101_1259.n3 a_11101_1259.t4 615.911
R11244 a_11101_1259.n2 a_11101_1259.t6 286.438
R11245 a_11101_1259.n2 a_11101_1259.t7 286.438
R11246 a_11101_1259.n10 a_11101_1259.n9 185.55
R11247 a_11101_1259.t5 a_11101_1259.n2 160.666
R11248 a_11101_1259.n8 a_11101_1259.n7 109.11
R11249 a_11101_1259.t2 a_11101_1259.n10 28.568
R11250 a_11101_1259.n9 a_11101_1259.t0 28.565
R11251 a_11101_1259.n9 a_11101_1259.t1 28.565
R11252 a_11101_1259.n8 a_11101_1259.t3 20.393
R11253 a_11101_1259.n4 a_11101_1259.n3 15.739
R11254 a_11101_1259.n10 a_11101_1259.n8 1.835
R11255 a_11101_1259.n7 a_11101_1259.n6 0.069
R11256 a_11101_1259.n6 a_11101_1259.n5 0.058
R11257 a_11101_1259.n1 a_11101_1259.n0 0.001
R11258 a_11101_1259.n5 a_11101_1259.n4 0.001
R11259 a_11101_1259.n4 a_11101_1259.n1 0.001
R11260 a_1745_8119.n2 a_1745_8119.t5 448.381
R11261 a_1745_8119.n1 a_1745_8119.t6 286.438
R11262 a_1745_8119.n1 a_1745_8119.t4 286.438
R11263 a_1745_8119.n0 a_1745_8119.t7 247.69
R11264 a_1745_8119.n4 a_1745_8119.n3 182.117
R11265 a_1745_8119.t5 a_1745_8119.n1 160.666
R11266 a_1745_8119.n3 a_1745_8119.t2 28.568
R11267 a_1745_8119.n4 a_1745_8119.t3 28.565
R11268 a_1745_8119.t0 a_1745_8119.n4 28.565
R11269 a_1745_8119.n0 a_1745_8119.t1 18.127
R11270 a_1745_8119.n2 a_1745_8119.n0 4.036
R11271 a_1745_8119.n3 a_1745_8119.n2 0.937
R11272 a_1099_8992.n0 a_1099_8992.n9 167.433
R11273 a_1099_8992.n0 a_1099_8992.t1 14.282
R11274 a_1099_8992.t0 a_1099_8992.n0 14.282
R11275 a_1099_8992.n9 a_1099_8992.n8 77.784
R11276 a_1099_8992.n8 a_1099_8992.n6 77.456
R11277 a_1099_8992.n6 a_1099_8992.n4 77.456
R11278 a_1099_8992.n4 a_1099_8992.n2 75.815
R11279 a_1099_8992.n9 a_1099_8992.t2 104.259
R11280 a_1099_8992.n8 a_1099_8992.n7 89.977
R11281 a_1099_8992.n7 a_1099_8992.t10 14.282
R11282 a_1099_8992.n7 a_1099_8992.t9 14.282
R11283 a_1099_8992.n6 a_1099_8992.n5 89.977
R11284 a_1099_8992.n5 a_1099_8992.t11 14.282
R11285 a_1099_8992.n5 a_1099_8992.t6 14.282
R11286 a_1099_8992.n4 a_1099_8992.n3 89.977
R11287 a_1099_8992.n3 a_1099_8992.t7 14.282
R11288 a_1099_8992.n3 a_1099_8992.t8 14.282
R11289 a_1099_8992.n2 a_1099_8992.t4 104.259
R11290 a_1099_8992.n2 a_1099_8992.n1 167.433
R11291 a_1099_8992.n1 a_1099_8992.t3 14.282
R11292 a_1099_8992.n1 a_1099_8992.t5 14.282
R11293 a_566_8262.t0 a_566_8262.n0 14.282
R11294 a_566_8262.n0 a_566_8262.t2 14.282
R11295 a_566_8262.n0 a_566_8262.n1 258.161
R11296 a_566_8262.n1 a_566_8262.n5 0.852
R11297 a_566_8262.n5 a_566_8262.n6 4.366
R11298 a_566_8262.n6 a_566_8262.n7 258.161
R11299 a_566_8262.n7 a_566_8262.t4 14.282
R11300 a_566_8262.n7 a_566_8262.t5 14.282
R11301 a_566_8262.n6 a_566_8262.t6 14.283
R11302 a_566_8262.n5 a_566_8262.n4 97.614
R11303 a_566_8262.n4 a_566_8262.t10 200.029
R11304 a_566_8262.t10 a_566_8262.n3 206.421
R11305 a_566_8262.n3 a_566_8262.t9 80.333
R11306 a_566_8262.n3 a_566_8262.t11 206.421
R11307 a_566_8262.n4 a_566_8262.t8 1527.4
R11308 a_566_8262.t8 a_566_8262.n2 657.379
R11309 a_566_8262.n2 a_566_8262.t3 8.7
R11310 a_566_8262.n2 a_566_8262.t7 8.7
R11311 a_566_8262.n1 a_566_8262.t1 14.283
R11312 a_54879_11969.n2 a_54879_11969.t7 214.335
R11313 a_54879_11969.t9 a_54879_11969.n2 214.335
R11314 a_54879_11969.n3 a_54879_11969.t9 143.851
R11315 a_54879_11969.n3 a_54879_11969.t8 135.658
R11316 a_54879_11969.n2 a_54879_11969.t10 80.333
R11317 a_54879_11969.n4 a_54879_11969.t0 28.565
R11318 a_54879_11969.n4 a_54879_11969.t1 28.565
R11319 a_54879_11969.n0 a_54879_11969.t4 28.565
R11320 a_54879_11969.n0 a_54879_11969.t5 28.565
R11321 a_54879_11969.t2 a_54879_11969.n7 28.565
R11322 a_54879_11969.n7 a_54879_11969.t6 28.565
R11323 a_54879_11969.n1 a_54879_11969.t3 9.714
R11324 a_54879_11969.n1 a_54879_11969.n0 1.003
R11325 a_54879_11969.n6 a_54879_11969.n5 0.833
R11326 a_54879_11969.n5 a_54879_11969.n4 0.653
R11327 a_54879_11969.n7 a_54879_11969.n6 0.653
R11328 a_54879_11969.n6 a_54879_11969.n1 0.341
R11329 a_54879_11969.n5 a_54879_11969.n3 0.032
R11330 a_55469_11532.n5 a_55469_11532.n4 535.449
R11331 a_55469_11532.t13 a_55469_11532.t12 437.233
R11332 a_55469_11532.t9 a_55469_11532.t5 437.233
R11333 a_55469_11532.t14 a_55469_11532.n2 313.873
R11334 a_55469_11532.n4 a_55469_11532.t8 294.986
R11335 a_55469_11532.n1 a_55469_11532.t18 272.288
R11336 a_55469_11532.n5 a_55469_11532.t10 245.184
R11337 a_55469_11532.n7 a_55469_11532.t9 218.628
R11338 a_55469_11532.n9 a_55469_11532.t13 217.024
R11339 a_55469_11532.n8 a_55469_11532.t16 214.686
R11340 a_55469_11532.t12 a_55469_11532.n8 214.686
R11341 a_55469_11532.n6 a_55469_11532.t4 214.686
R11342 a_55469_11532.t5 a_55469_11532.n6 214.686
R11343 a_55469_11532.n11 a_55469_11532.n0 192.754
R11344 a_55469_11532.n3 a_55469_11532.t14 190.152
R11345 a_55469_11532.n3 a_55469_11532.t17 190.152
R11346 a_55469_11532.n1 a_55469_11532.t11 160.666
R11347 a_55469_11532.n2 a_55469_11532.t7 160.666
R11348 a_55469_11532.n4 a_55469_11532.t19 110.859
R11349 a_55469_11532.n2 a_55469_11532.n1 96.129
R11350 a_55469_11532.n8 a_55469_11532.t6 80.333
R11351 a_55469_11532.t10 a_55469_11532.n3 80.333
R11352 a_55469_11532.n6 a_55469_11532.t15 80.333
R11353 a_55469_11532.t2 a_55469_11532.n11 28.568
R11354 a_55469_11532.n0 a_55469_11532.t0 28.565
R11355 a_55469_11532.n0 a_55469_11532.t1 28.565
R11356 a_55469_11532.n10 a_55469_11532.t3 18.823
R11357 a_55469_11532.n7 a_55469_11532.n5 14.9
R11358 a_55469_11532.n10 a_55469_11532.n9 3.074
R11359 a_55469_11532.n9 a_55469_11532.n7 2.599
R11360 a_55469_11532.n11 a_55469_11532.n10 1.105
R11361 opcode[1].n51 opcode[1].t56 1374.48
R11362 opcode[1].n46 opcode[1].t127 1374.48
R11363 opcode[1].n41 opcode[1].t117 1374.48
R11364 opcode[1].n63 opcode[1].t25 1374.48
R11365 opcode[1].n68 opcode[1].t8 1374.48
R11366 opcode[1].n73 opcode[1].t55 1374.48
R11367 opcode[1].n82 opcode[1].t4 1374.48
R11368 opcode[1].n88 opcode[1].t3 1374.48
R11369 opcode[1].n1 opcode[1].t0 1374.12
R11370 opcode[1].n4 opcode[1].t126 1374.12
R11371 opcode[1].n7 opcode[1].t116 1374.12
R11372 opcode[1].n10 opcode[1].t10 1374.12
R11373 opcode[1].n13 opcode[1].t48 1374.12
R11374 opcode[1].n16 opcode[1].t61 1374.12
R11375 opcode[1].n19 opcode[1].t77 1374.12
R11376 opcode[1].n22 opcode[1].t112 1374.12
R11377 opcode[1].n38 opcode[1].t93 623.291
R11378 opcode[1].n36 opcode[1].t39 623.291
R11379 opcode[1].n34 opcode[1].t50 623.291
R11380 opcode[1].n32 opcode[1].t88 623.291
R11381 opcode[1].n30 opcode[1].t21 623.291
R11382 opcode[1].n28 opcode[1].t47 623.291
R11383 opcode[1].n26 opcode[1].t20 623.291
R11384 opcode[1].n24 opcode[1].t69 623.291
R11385 opcode[1].n54 opcode[1].t111 622.488
R11386 opcode[1].n48 opcode[1].t70 622.488
R11387 opcode[1].n43 opcode[1].t75 622.488
R11388 opcode[1].n65 opcode[1].t114 622.488
R11389 opcode[1].n70 opcode[1].t5 622.488
R11390 opcode[1].n75 opcode[1].t2 622.488
R11391 opcode[1].n78 opcode[1].t103 622.488
R11392 opcode[1].n90 opcode[1].t34 622.488
R11393 opcode[1].n38 opcode[1].t119 610.283
R11394 opcode[1].n36 opcode[1].t46 610.283
R11395 opcode[1].n34 opcode[1].t124 610.283
R11396 opcode[1].n32 opcode[1].t38 610.283
R11397 opcode[1].n30 opcode[1].t62 610.283
R11398 opcode[1].n28 opcode[1].t76 610.283
R11399 opcode[1].n26 opcode[1].t98 610.283
R11400 opcode[1].n24 opcode[1].t1 610.283
R11401 opcode[1].n54 opcode[1].t78 610.283
R11402 opcode[1].n48 opcode[1].t44 610.283
R11403 opcode[1].n43 opcode[1].t19 610.283
R11404 opcode[1].n65 opcode[1].t89 610.283
R11405 opcode[1].n70 opcode[1].t52 610.283
R11406 opcode[1].n75 opcode[1].t83 610.283
R11407 opcode[1].n78 opcode[1].t40 610.283
R11408 opcode[1].n90 opcode[1].t110 610.283
R11409 opcode[1].n1 opcode[1].t90 326.034
R11410 opcode[1].n4 opcode[1].t125 326.034
R11411 opcode[1].n7 opcode[1].t59 326.034
R11412 opcode[1].n10 opcode[1].t109 326.034
R11413 opcode[1].n13 opcode[1].t37 326.034
R11414 opcode[1].n16 opcode[1].t45 326.034
R11415 opcode[1].n19 opcode[1].t17 326.034
R11416 opcode[1].n22 opcode[1].t67 326.034
R11417 opcode[1].n51 opcode[1].t118 325.68
R11418 opcode[1].n46 opcode[1].t92 325.68
R11419 opcode[1].n41 opcode[1].t101 325.68
R11420 opcode[1].n63 opcode[1].t123 325.68
R11421 opcode[1].n68 opcode[1].t121 325.68
R11422 opcode[1].n73 opcode[1].t31 325.68
R11423 opcode[1].n82 opcode[1].t86 325.68
R11424 opcode[1].n88 opcode[1].t12 325.68
R11425 opcode[1].n53 opcode[1].t23 287.241
R11426 opcode[1].n53 opcode[1].t53 287.241
R11427 opcode[1].n47 opcode[1].t81 287.241
R11428 opcode[1].n47 opcode[1].t9 287.241
R11429 opcode[1].n42 opcode[1].t99 287.241
R11430 opcode[1].n42 opcode[1].t66 287.241
R11431 opcode[1].n64 opcode[1].t36 287.241
R11432 opcode[1].n64 opcode[1].t63 287.241
R11433 opcode[1].n69 opcode[1].t73 287.241
R11434 opcode[1].n69 opcode[1].t95 287.241
R11435 opcode[1].n74 opcode[1].t68 287.241
R11436 opcode[1].n74 opcode[1].t29 287.241
R11437 opcode[1].n77 opcode[1].t16 287.241
R11438 opcode[1].n77 opcode[1].t51 287.241
R11439 opcode[1].n89 opcode[1].t113 287.241
R11440 opcode[1].n89 opcode[1].t84 287.241
R11441 opcode[1].n2 opcode[1].t87 286.438
R11442 opcode[1].n2 opcode[1].t97 286.438
R11443 opcode[1].n5 opcode[1].t120 286.438
R11444 opcode[1].n5 opcode[1].t42 286.438
R11445 opcode[1].n8 opcode[1].t49 286.438
R11446 opcode[1].n8 opcode[1].t96 286.438
R11447 opcode[1].n11 opcode[1].t85 286.438
R11448 opcode[1].n11 opcode[1].t94 286.438
R11449 opcode[1].n14 opcode[1].t35 286.438
R11450 opcode[1].n14 opcode[1].t58 286.438
R11451 opcode[1].n17 opcode[1].t43 286.438
R11452 opcode[1].n17 opcode[1].t74 286.438
R11453 opcode[1].n20 opcode[1].t14 286.438
R11454 opcode[1].n20 opcode[1].t24 286.438
R11455 opcode[1].n23 opcode[1].t65 286.438
R11456 opcode[1].n23 opcode[1].t106 286.438
R11457 opcode[1].n50 opcode[1].t15 207.225
R11458 opcode[1].t118 opcode[1].n50 207.225
R11459 opcode[1].n45 opcode[1].t11 207.225
R11460 opcode[1].t92 opcode[1].n45 207.225
R11461 opcode[1].n40 opcode[1].t32 207.225
R11462 opcode[1].t101 opcode[1].n40 207.225
R11463 opcode[1].n62 opcode[1].t64 207.225
R11464 opcode[1].t123 opcode[1].n62 207.225
R11465 opcode[1].n67 opcode[1].t60 207.225
R11466 opcode[1].t121 opcode[1].n67 207.225
R11467 opcode[1].n72 opcode[1].t91 207.225
R11468 opcode[1].t31 opcode[1].n72 207.225
R11469 opcode[1].n81 opcode[1].t6 207.225
R11470 opcode[1].t86 opcode[1].n81 207.225
R11471 opcode[1].n87 opcode[1].t22 207.225
R11472 opcode[1].t12 opcode[1].n87 207.225
R11473 opcode[1].n0 opcode[1].t102 206.421
R11474 opcode[1].t90 opcode[1].n0 206.421
R11475 opcode[1].n3 opcode[1].t100 206.421
R11476 opcode[1].t125 opcode[1].n3 206.421
R11477 opcode[1].n6 opcode[1].t18 206.421
R11478 opcode[1].t59 opcode[1].n6 206.421
R11479 opcode[1].n9 opcode[1].t54 206.421
R11480 opcode[1].t109 opcode[1].n9 206.421
R11481 opcode[1].n12 opcode[1].t115 206.421
R11482 opcode[1].t37 opcode[1].n12 206.421
R11483 opcode[1].n15 opcode[1].t122 206.421
R11484 opcode[1].t45 opcode[1].n15 206.421
R11485 opcode[1].n18 opcode[1].t28 206.421
R11486 opcode[1].t17 opcode[1].n18 206.421
R11487 opcode[1].n21 opcode[1].t26 206.421
R11488 opcode[1].t67 opcode[1].n21 206.421
R11489 opcode[1].t93 opcode[1].n2 160.666
R11490 opcode[1].t39 opcode[1].n5 160.666
R11491 opcode[1].t50 opcode[1].n8 160.666
R11492 opcode[1].t88 opcode[1].n11 160.666
R11493 opcode[1].t21 opcode[1].n14 160.666
R11494 opcode[1].t47 opcode[1].n17 160.666
R11495 opcode[1].t20 opcode[1].n20 160.666
R11496 opcode[1].t69 opcode[1].n23 160.666
R11497 opcode[1].t111 opcode[1].n53 160.666
R11498 opcode[1].t70 opcode[1].n47 160.666
R11499 opcode[1].t75 opcode[1].n42 160.666
R11500 opcode[1].t114 opcode[1].n64 160.666
R11501 opcode[1].t5 opcode[1].n69 160.666
R11502 opcode[1].t2 opcode[1].n74 160.666
R11503 opcode[1].t103 opcode[1].n77 160.666
R11504 opcode[1].t34 opcode[1].n89 160.666
R11505 opcode[1].n0 opcode[1].t107 80.333
R11506 opcode[1].n3 opcode[1].t105 80.333
R11507 opcode[1].n6 opcode[1].t57 80.333
R11508 opcode[1].n9 opcode[1].t104 80.333
R11509 opcode[1].n12 opcode[1].t33 80.333
R11510 opcode[1].n15 opcode[1].t41 80.333
R11511 opcode[1].n18 opcode[1].t7 80.333
R11512 opcode[1].n21 opcode[1].t30 80.333
R11513 opcode[1].n50 opcode[1].t72 80.333
R11514 opcode[1].n45 opcode[1].t71 80.333
R11515 opcode[1].n40 opcode[1].t82 80.333
R11516 opcode[1].n62 opcode[1].t80 80.333
R11517 opcode[1].n67 opcode[1].t79 80.333
R11518 opcode[1].n72 opcode[1].t13 80.333
R11519 opcode[1].n81 opcode[1].t27 80.333
R11520 opcode[1].n87 opcode[1].t108 80.333
R11521 opcode[1].n97 opcode[1].n96 57.595
R11522 opcode[1] opcode[1].n97 49.044
R11523 opcode[1].n97 opcode[1].n39 18.595
R11524 opcode[1].n92 opcode[1].n91 7.802
R11525 opcode[1].n60 opcode[1].n59 7.174
R11526 opcode[1].n94 opcode[1].n71 4.102
R11527 opcode[1].n93 opcode[1].n76 4.1
R11528 opcode[1].n60 opcode[1].n49 4.052
R11529 opcode[1].n61 opcode[1].n44 4.046
R11530 opcode[1].n95 opcode[1].n66 3.999
R11531 opcode[1].n92 opcode[1].n86 3.828
R11532 opcode[1].n95 opcode[1].n94 3.777
R11533 opcode[1].n94 opcode[1].n93 3.707
R11534 opcode[1].n61 opcode[1].n60 3.693
R11535 opcode[1].n93 opcode[1].n92 3.693
R11536 opcode[1].n96 opcode[1].n61 3.625
R11537 opcode[1].n32 opcode[1].n31 3.312
R11538 opcode[1].n30 opcode[1].n29 3.12
R11539 opcode[1].n26 opcode[1].n25 3.089
R11540 opcode[1].n34 opcode[1].n33 3.059
R11541 opcode[1].n38 opcode[1].n37 3.059
R11542 opcode[1].n36 opcode[1].n35 3.037
R11543 opcode[1].n28 opcode[1].n27 2.994
R11544 opcode[1].n55 opcode[1].n54 2.07
R11545 opcode[1].n79 opcode[1].n78 1.715
R11546 opcode[1].n35 opcode[1].n34 1.616
R11547 opcode[1].n29 opcode[1].n28 1.616
R11548 opcode[1].n49 opcode[1].n48 1.614
R11549 opcode[1].n44 opcode[1].n43 1.614
R11550 opcode[1].n66 opcode[1].n65 1.614
R11551 opcode[1].n71 opcode[1].n70 1.614
R11552 opcode[1].n76 opcode[1].n75 1.614
R11553 opcode[1].n91 opcode[1].n90 1.614
R11554 opcode[1].n39 opcode[1].n38 1.614
R11555 opcode[1].n37 opcode[1].n36 1.614
R11556 opcode[1].n33 opcode[1].n32 1.614
R11557 opcode[1].n31 opcode[1].n30 1.614
R11558 opcode[1].n27 opcode[1].n26 1.614
R11559 opcode[1].n25 opcode[1].n24 1.614
R11560 opcode[1].n86 opcode[1].n85 0.243
R11561 opcode[1].n59 opcode[1].n58 0.236
R11562 opcode[1].n58 opcode[1].n57 0.086
R11563 opcode[1].n96 opcode[1].n95 0.08
R11564 opcode[1].n85 opcode[1].n84 0.056
R11565 opcode[1].n49 opcode[1].n46 0.003
R11566 opcode[1].n44 opcode[1].n41 0.003
R11567 opcode[1].n66 opcode[1].n63 0.003
R11568 opcode[1].n71 opcode[1].n68 0.003
R11569 opcode[1].n76 opcode[1].n73 0.003
R11570 opcode[1].n91 opcode[1].n88 0.003
R11571 opcode[1].n39 opcode[1].n1 0.003
R11572 opcode[1].n37 opcode[1].n4 0.003
R11573 opcode[1].n33 opcode[1].n10 0.003
R11574 opcode[1].n31 opcode[1].n13 0.003
R11575 opcode[1].n27 opcode[1].n19 0.003
R11576 opcode[1].n25 opcode[1].n22 0.003
R11577 opcode[1].n35 opcode[1].n7 0.003
R11578 opcode[1].n29 opcode[1].n16 0.003
R11579 opcode[1].n57 opcode[1].n56 0.002
R11580 opcode[1].n84 opcode[1].n80 0.002
R11581 opcode[1].n52 opcode[1].n51 0.001
R11582 opcode[1].n83 opcode[1].n82 0.001
R11583 opcode[1].n80 opcode[1].n79 0.001
R11584 opcode[1].n56 opcode[1].n55 0.001
R11585 opcode[1].n57 opcode[1].n52 0.001
R11586 opcode[1].n84 opcode[1].n83 0.001
R11587 a_23777_10847.n3 a_23777_10847.t4 448.381
R11588 a_23777_10847.n2 a_23777_10847.t7 286.438
R11589 a_23777_10847.n2 a_23777_10847.t5 286.438
R11590 a_23777_10847.n1 a_23777_10847.t6 247.69
R11591 a_23777_10847.n4 a_23777_10847.n0 182.117
R11592 a_23777_10847.t4 a_23777_10847.n2 160.666
R11593 a_23777_10847.t2 a_23777_10847.n4 28.568
R11594 a_23777_10847.n0 a_23777_10847.t0 28.565
R11595 a_23777_10847.n0 a_23777_10847.t1 28.565
R11596 a_23777_10847.n1 a_23777_10847.t3 18.127
R11597 a_23777_10847.n3 a_23777_10847.n1 4.036
R11598 a_23777_10847.n4 a_23777_10847.n3 0.937
R11599 a_35594_7027.n7 a_35594_7027.n6 861.987
R11600 a_35594_7027.n6 a_35594_7027.n5 560.726
R11601 a_35594_7027.t11 a_35594_7027.t10 415.315
R11602 a_35594_7027.t17 a_35594_7027.t13 415.315
R11603 a_35594_7027.n2 a_35594_7027.t15 394.151
R11604 a_35594_7027.n5 a_35594_7027.t19 294.653
R11605 a_35594_7027.n1 a_35594_7027.t6 269.523
R11606 a_35594_7027.t15 a_35594_7027.n1 269.523
R11607 a_35594_7027.n9 a_35594_7027.t11 217.716
R11608 a_35594_7027.n8 a_35594_7027.t12 214.335
R11609 a_35594_7027.t10 a_35594_7027.n8 214.335
R11610 a_35594_7027.n0 a_35594_7027.t14 214.335
R11611 a_35594_7027.t13 a_35594_7027.n0 214.335
R11612 a_35594_7027.n7 a_35594_7027.t17 198.921
R11613 a_35594_7027.n3 a_35594_7027.t7 198.043
R11614 a_35594_7027.n12 a_35594_7027.n11 192.754
R11615 a_35594_7027.n1 a_35594_7027.t8 160.666
R11616 a_35594_7027.n5 a_35594_7027.t5 111.663
R11617 a_35594_7027.n4 a_35594_7027.n2 97.816
R11618 a_35594_7027.n3 a_35594_7027.t16 93.989
R11619 a_35594_7027.n8 a_35594_7027.t18 80.333
R11620 a_35594_7027.n2 a_35594_7027.t9 80.333
R11621 a_35594_7027.n0 a_35594_7027.t4 80.333
R11622 a_35594_7027.n6 a_35594_7027.n4 65.07
R11623 a_35594_7027.n11 a_35594_7027.t2 28.568
R11624 a_35594_7027.n12 a_35594_7027.t3 28.565
R11625 a_35594_7027.t0 a_35594_7027.n12 28.565
R11626 a_35594_7027.n10 a_35594_7027.t1 18.825
R11627 a_35594_7027.n9 a_35594_7027.n7 16.411
R11628 a_35594_7027.n4 a_35594_7027.n3 6.615
R11629 a_35594_7027.n10 a_35594_7027.n9 2.757
R11630 a_35594_7027.n11 a_35594_7027.n10 1.105
R11631 a_37916_8132.n0 a_37916_8132.t9 214.335
R11632 a_37916_8132.t8 a_37916_8132.n0 214.335
R11633 a_37916_8132.n1 a_37916_8132.t8 143.851
R11634 a_37916_8132.n1 a_37916_8132.t10 135.658
R11635 a_37916_8132.n0 a_37916_8132.t7 80.333
R11636 a_37916_8132.n2 a_37916_8132.t4 28.565
R11637 a_37916_8132.n2 a_37916_8132.t6 28.565
R11638 a_37916_8132.n4 a_37916_8132.t5 28.565
R11639 a_37916_8132.n4 a_37916_8132.t1 28.565
R11640 a_37916_8132.t0 a_37916_8132.n7 28.565
R11641 a_37916_8132.n7 a_37916_8132.t2 28.565
R11642 a_37916_8132.n6 a_37916_8132.t3 9.714
R11643 a_37916_8132.n7 a_37916_8132.n6 1.003
R11644 a_37916_8132.n5 a_37916_8132.n3 0.833
R11645 a_37916_8132.n3 a_37916_8132.n2 0.653
R11646 a_37916_8132.n5 a_37916_8132.n4 0.653
R11647 a_37916_8132.n6 a_37916_8132.n5 0.341
R11648 a_37916_8132.n3 a_37916_8132.n1 0.032
R11649 a_48542_1014.n1 a_48542_1014.t7 318.922
R11650 a_48542_1014.n0 a_48542_1014.t4 274.739
R11651 a_48542_1014.n0 a_48542_1014.t6 274.739
R11652 a_48542_1014.n1 a_48542_1014.t5 269.116
R11653 a_48542_1014.t7 a_48542_1014.n0 179.946
R11654 a_48542_1014.n2 a_48542_1014.n1 105.178
R11655 a_48542_1014.n3 a_48542_1014.t3 29.444
R11656 a_48542_1014.n4 a_48542_1014.t1 28.565
R11657 a_48542_1014.t0 a_48542_1014.n4 28.565
R11658 a_48542_1014.n2 a_48542_1014.t2 18.145
R11659 a_48542_1014.n3 a_48542_1014.n2 2.878
R11660 a_48542_1014.n4 a_48542_1014.n3 0.764
R11661 a_48248_1040.n0 a_48248_1040.n13 122.999
R11662 a_48248_1040.t0 a_48248_1040.n0 14.282
R11663 a_48248_1040.n0 a_48248_1040.t3 14.282
R11664 a_48248_1040.n13 a_48248_1040.n11 50.575
R11665 a_48248_1040.n11 a_48248_1040.n9 74.302
R11666 a_48248_1040.n13 a_48248_1040.n12 157.665
R11667 a_48248_1040.n12 a_48248_1040.t2 8.7
R11668 a_48248_1040.n12 a_48248_1040.t4 8.7
R11669 a_48248_1040.n11 a_48248_1040.n10 90.416
R11670 a_48248_1040.n10 a_48248_1040.t1 14.282
R11671 a_48248_1040.n10 a_48248_1040.t7 14.282
R11672 a_48248_1040.n9 a_48248_1040.n8 90.436
R11673 a_48248_1040.n8 a_48248_1040.t5 14.282
R11674 a_48248_1040.n8 a_48248_1040.t6 14.282
R11675 a_48248_1040.n9 a_48248_1040.n1 1712.43
R11676 a_48248_1040.n1 a_48248_1040.t17 217.826
R11677 a_48248_1040.n1 a_48248_1040.n6 133.839
R11678 a_48248_1040.t17 a_48248_1040.t16 437.233
R11679 a_48248_1040.t16 a_48248_1040.n7 214.686
R11680 a_48248_1040.n7 a_48248_1040.t9 80.333
R11681 a_48248_1040.n7 a_48248_1040.t13 214.686
R11682 a_48248_1040.n6 a_48248_1040.n2 563.136
R11683 a_48248_1040.n6 a_48248_1040.t12 178.973
R11684 a_48248_1040.t12 a_48248_1040.n5 80.333
R11685 a_48248_1040.n5 a_48248_1040.t19 190.152
R11686 a_48248_1040.n5 a_48248_1040.t18 190.152
R11687 a_48248_1040.t18 a_48248_1040.n4 313.873
R11688 a_48248_1040.n4 a_48248_1040.t10 160.666
R11689 a_48248_1040.n4 a_48248_1040.n3 96.129
R11690 a_48248_1040.n3 a_48248_1040.t14 160.666
R11691 a_48248_1040.n3 a_48248_1040.t8 272.288
R11692 a_48248_1040.n2 a_48248_1040.t15 294.986
R11693 a_48248_1040.n2 a_48248_1040.t11 110.859
R11694 a_48130_1040.t0 a_48130_1040.n7 16.058
R11695 a_48130_1040.n7 a_48130_1040.n5 0.575
R11696 a_48130_1040.n5 a_48130_1040.n9 0.2
R11697 a_48130_1040.n9 a_48130_1040.t10 16.058
R11698 a_48130_1040.n9 a_48130_1040.n8 0.999
R11699 a_48130_1040.n8 a_48130_1040.t11 14.282
R11700 a_48130_1040.n8 a_48130_1040.t9 14.282
R11701 a_48130_1040.n7 a_48130_1040.n6 0.999
R11702 a_48130_1040.n6 a_48130_1040.t2 14.282
R11703 a_48130_1040.n6 a_48130_1040.t1 14.282
R11704 a_48130_1040.n5 a_48130_1040.n3 0.227
R11705 a_48130_1040.n3 a_48130_1040.n4 1.511
R11706 a_48130_1040.n4 a_48130_1040.t6 14.282
R11707 a_48130_1040.n4 a_48130_1040.t8 14.282
R11708 a_48130_1040.n3 a_48130_1040.n0 0.669
R11709 a_48130_1040.n0 a_48130_1040.n1 0.001
R11710 a_48130_1040.n0 a_48130_1040.n2 267.767
R11711 a_48130_1040.n2 a_48130_1040.t3 14.282
R11712 a_48130_1040.n2 a_48130_1040.t5 14.282
R11713 a_48130_1040.n1 a_48130_1040.t7 14.282
R11714 a_48130_1040.n1 a_48130_1040.t4 14.282
R11715 a_54908_6842.n0 a_54908_6842.n13 122.999
R11716 a_54908_6842.t0 a_54908_6842.n0 14.282
R11717 a_54908_6842.n0 a_54908_6842.t2 14.282
R11718 a_54908_6842.n13 a_54908_6842.n11 50.575
R11719 a_54908_6842.n11 a_54908_6842.n9 74.302
R11720 a_54908_6842.n13 a_54908_6842.n12 157.665
R11721 a_54908_6842.n12 a_54908_6842.t1 8.7
R11722 a_54908_6842.n12 a_54908_6842.t6 8.7
R11723 a_54908_6842.n11 a_54908_6842.n10 90.416
R11724 a_54908_6842.n10 a_54908_6842.t3 14.282
R11725 a_54908_6842.n10 a_54908_6842.t4 14.282
R11726 a_54908_6842.n9 a_54908_6842.n8 90.436
R11727 a_54908_6842.n8 a_54908_6842.t7 14.282
R11728 a_54908_6842.n8 a_54908_6842.t5 14.282
R11729 a_54908_6842.n1 a_54908_6842.t17 217.826
R11730 a_54908_6842.n9 a_54908_6842.n1 277.579
R11731 a_54908_6842.n1 a_54908_6842.n6 133.839
R11732 a_54908_6842.t17 a_54908_6842.t10 437.233
R11733 a_54908_6842.t10 a_54908_6842.n7 214.686
R11734 a_54908_6842.n7 a_54908_6842.t18 80.333
R11735 a_54908_6842.n7 a_54908_6842.t8 214.686
R11736 a_54908_6842.n6 a_54908_6842.n2 563.136
R11737 a_54908_6842.n6 a_54908_6842.t11 178.973
R11738 a_54908_6842.t11 a_54908_6842.n5 80.333
R11739 a_54908_6842.n5 a_54908_6842.t16 190.152
R11740 a_54908_6842.n5 a_54908_6842.t15 190.152
R11741 a_54908_6842.t15 a_54908_6842.n4 313.873
R11742 a_54908_6842.n4 a_54908_6842.t9 160.666
R11743 a_54908_6842.n4 a_54908_6842.n3 96.129
R11744 a_54908_6842.n3 a_54908_6842.t12 160.666
R11745 a_54908_6842.n3 a_54908_6842.t19 272.288
R11746 a_54908_6842.n2 a_54908_6842.t14 294.986
R11747 a_54908_6842.n2 a_54908_6842.t13 110.859
R11748 a_67135_3808.n4 a_67135_3808.t9 214.335
R11749 a_67135_3808.t8 a_67135_3808.n4 214.335
R11750 a_67135_3808.n5 a_67135_3808.t8 143.851
R11751 a_67135_3808.n5 a_67135_3808.t7 135.658
R11752 a_67135_3808.n4 a_67135_3808.t10 80.333
R11753 a_67135_3808.n0 a_67135_3808.t2 28.565
R11754 a_67135_3808.n0 a_67135_3808.t4 28.565
R11755 a_67135_3808.n2 a_67135_3808.t1 28.565
R11756 a_67135_3808.n2 a_67135_3808.t3 28.565
R11757 a_67135_3808.n7 a_67135_3808.t6 28.565
R11758 a_67135_3808.t0 a_67135_3808.n7 28.565
R11759 a_67135_3808.n1 a_67135_3808.t5 9.714
R11760 a_67135_3808.n1 a_67135_3808.n0 1.003
R11761 a_67135_3808.n6 a_67135_3808.n3 0.833
R11762 a_67135_3808.n3 a_67135_3808.n2 0.653
R11763 a_67135_3808.n7 a_67135_3808.n6 0.653
R11764 a_67135_3808.n3 a_67135_3808.n1 0.341
R11765 a_67135_3808.n6 a_67135_3808.n5 0.032
R11766 a_48006_21370.n0 a_48006_21370.n1 0.001
R11767 a_48006_21370.n0 a_48006_21370.t9 14.282
R11768 a_48006_21370.t0 a_48006_21370.n0 14.282
R11769 a_48006_21370.n1 a_48006_21370.n9 267.767
R11770 a_48006_21370.n9 a_48006_21370.t1 14.282
R11771 a_48006_21370.n9 a_48006_21370.t11 14.282
R11772 a_48006_21370.n1 a_48006_21370.n7 0.669
R11773 a_48006_21370.n7 a_48006_21370.n8 1.511
R11774 a_48006_21370.n8 a_48006_21370.t8 14.282
R11775 a_48006_21370.n8 a_48006_21370.t10 14.282
R11776 a_48006_21370.n7 a_48006_21370.n6 0.227
R11777 a_48006_21370.n6 a_48006_21370.n3 0.575
R11778 a_48006_21370.n6 a_48006_21370.n5 0.2
R11779 a_48006_21370.n5 a_48006_21370.t4 16.058
R11780 a_48006_21370.n5 a_48006_21370.n4 0.999
R11781 a_48006_21370.n4 a_48006_21370.t2 14.282
R11782 a_48006_21370.n4 a_48006_21370.t3 14.282
R11783 a_48006_21370.n3 a_48006_21370.n2 0.999
R11784 a_48006_21370.n2 a_48006_21370.t7 14.282
R11785 a_48006_21370.n2 a_48006_21370.t5 14.282
R11786 a_48006_21370.n3 a_48006_21370.t6 16.058
R11787 a_1974_8339.n1 a_1974_8339.t5 990.34
R11788 a_1974_8339.n1 a_1974_8339.t4 408.211
R11789 a_1974_8339.n0 a_1974_8339.t6 286.438
R11790 a_1974_8339.n0 a_1974_8339.t7 286.438
R11791 a_1974_8339.n4 a_1974_8339.n3 197.272
R11792 a_1974_8339.t5 a_1974_8339.n0 160.666
R11793 a_1974_8339.n3 a_1974_8339.t1 28.568
R11794 a_1974_8339.n4 a_1974_8339.t0 28.565
R11795 a_1974_8339.t2 a_1974_8339.n4 28.565
R11796 a_1974_8339.n2 a_1974_8339.t3 18.092
R11797 a_1974_8339.n2 a_1974_8339.n1 6.447
R11798 a_1974_8339.n3 a_1974_8339.n2 0.459
R11799 a_1926_7659.t0 a_1926_7659.t1 17.4
R11800 B[5].n12 B[5].n6 973.987
R11801 B[5].t37 B[5].t2 800.874
R11802 B[5].n22 B[5].n21 649.333
R11803 B[5].n18 B[5].n17 618.566
R11804 B[5].n11 B[5].n7 592.056
R11805 B[5].t0 B[5].t27 437.233
R11806 B[5].t7 B[5].t25 437.233
R11807 B[5].t11 B[5].t23 415.315
R11808 B[5].t30 B[5].t26 415.315
R11809 B[5].t15 B[5].t8 415.315
R11810 B[5].t5 B[5].n15 313.873
R11811 B[5].t17 B[5].n9 313.069
R11812 B[5].n7 B[5].t6 294.986
R11813 B[5].n20 B[5].t29 285.543
R11814 B[5].n17 B[5].t13 273.077
R11815 B[5].n14 B[5].t3 272.288
R11816 B[5].n8 B[5].t4 271.484
R11817 B[5].n2 B[5].t15 240.379
R11818 B[5].n5 B[5].t7 227.856
R11819 B[5].n2 B[5].t30 218.339
R11820 B[5].n5 B[5].t0 218.225
R11821 B[5].n19 B[5].t11 217.527
R11822 B[5].n3 B[5].t9 214.686
R11823 B[5].t27 B[5].n3 214.686
R11824 B[5].n4 B[5].t20 214.686
R11825 B[5].t25 B[5].n4 214.686
R11826 B[5].n1 B[5].t32 214.335
R11827 B[5].t26 B[5].n1 214.335
R11828 B[5].n0 B[5].t34 214.335
R11829 B[5].t8 B[5].n0 214.335
R11830 B[5].n13 B[5].t19 214.335
R11831 B[5].t23 B[5].n13 214.335
R11832 B[5].n18 B[5].t16 204.679
R11833 B[5].n11 B[5].t12 204.672
R11834 B[5].n21 B[5].t37 194.406
R11835 B[5].n10 B[5].t17 190.955
R11836 B[5].n10 B[5].t1 190.955
R11837 B[5].n16 B[5].t38 190.152
R11838 B[5].n16 B[5].t5 190.152
R11839 B[5].n9 B[5].t10 160.666
R11840 B[5].n8 B[5].t36 160.666
R11841 B[5].n14 B[5].t14 160.666
R11842 B[5].n15 B[5].t35 160.666
R11843 B[5].n20 B[5].t18 160.666
R11844 B[5].n17 B[5].t31 137.369
R11845 B[5].n7 B[5].t39 110.859
R11846 B[5].n9 B[5].n8 96.129
R11847 B[5].n15 B[5].n14 96.129
R11848 B[5].n21 B[5].n20 91.137
R11849 B[5].n1 B[5].t28 80.333
R11850 B[5].n0 B[5].t33 80.333
R11851 B[5].n3 B[5].t24 80.333
R11852 B[5].n4 B[5].t22 80.333
R11853 B[5].t12 B[5].n10 80.333
R11854 B[5].n13 B[5].t21 80.333
R11855 B[5].t16 B[5].n16 80.333
R11856 B[5].n19 B[5].n18 51.128
R11857 B[5] B[5].n23 48.831
R11858 B[5].n12 B[5].n11 46.001
R11859 B[5].n23 B[5].n12 29.459
R11860 B[5].n6 B[5].n2 28.897
R11861 B[5].n23 B[5].n22 19.593
R11862 B[5].n6 B[5].n5 7.414
R11863 B[5].n22 B[5].n19 5.864
R11864 a_41711_n1755.n0 a_41711_n1755.t9 214.335
R11865 a_41711_n1755.t7 a_41711_n1755.n0 214.335
R11866 a_41711_n1755.n1 a_41711_n1755.t7 143.85
R11867 a_41711_n1755.n1 a_41711_n1755.t10 135.66
R11868 a_41711_n1755.n0 a_41711_n1755.t8 80.333
R11869 a_41711_n1755.n2 a_41711_n1755.t4 28.565
R11870 a_41711_n1755.n2 a_41711_n1755.t5 28.565
R11871 a_41711_n1755.n4 a_41711_n1755.t6 28.565
R11872 a_41711_n1755.n4 a_41711_n1755.t1 28.565
R11873 a_41711_n1755.n7 a_41711_n1755.t2 28.565
R11874 a_41711_n1755.t3 a_41711_n1755.n7 28.565
R11875 a_41711_n1755.n6 a_41711_n1755.t0 9.714
R11876 a_41711_n1755.n7 a_41711_n1755.n6 1.003
R11877 a_41711_n1755.n5 a_41711_n1755.n3 0.836
R11878 a_41711_n1755.n5 a_41711_n1755.n4 0.653
R11879 a_41711_n1755.n3 a_41711_n1755.n2 0.65
R11880 a_41711_n1755.n6 a_41711_n1755.n5 0.341
R11881 a_41711_n1755.n3 a_41711_n1755.n1 0.032
R11882 a_41948_n1318.t0 a_41948_n1318.t1 17.4
R11883 a_30647_12105.t0 a_30647_12105.n0 14.282
R11884 a_30647_12105.n0 a_30647_12105.t2 14.282
R11885 a_30647_12105.n4 a_30647_12105.n2 74.302
R11886 a_30647_12105.n6 a_30647_12105.n4 50.575
R11887 a_30647_12105.n0 a_30647_12105.n6 110.084
R11888 a_30647_12105.n2 a_30647_12105.n7 201.691
R11889 a_30647_12105.n7 a_30647_12105.n9 16.411
R11890 a_30647_12105.n9 a_30647_12105.t17 198.921
R11891 a_30647_12105.t17 a_30647_12105.t18 415.315
R11892 a_30647_12105.t18 a_30647_12105.n16 214.335
R11893 a_30647_12105.n16 a_30647_12105.t21 80.333
R11894 a_30647_12105.n16 a_30647_12105.t22 214.335
R11895 a_30647_12105.n9 a_30647_12105.n15 861.987
R11896 a_30647_12105.n15 a_30647_12105.n10 560.726
R11897 a_30647_12105.n15 a_30647_12105.n14 65.07
R11898 a_30647_12105.n14 a_30647_12105.n13 6.615
R11899 a_30647_12105.n13 a_30647_12105.t10 93.989
R11900 a_30647_12105.n14 a_30647_12105.n12 97.816
R11901 a_30647_12105.n12 a_30647_12105.t11 80.333
R11902 a_30647_12105.n12 a_30647_12105.t15 394.151
R11903 a_30647_12105.t15 a_30647_12105.n11 269.523
R11904 a_30647_12105.n11 a_30647_12105.t16 160.666
R11905 a_30647_12105.n11 a_30647_12105.t19 269.523
R11906 a_30647_12105.n13 a_30647_12105.t9 198.043
R11907 a_30647_12105.n10 a_30647_12105.t12 294.653
R11908 a_30647_12105.n10 a_30647_12105.t13 111.663
R11909 a_30647_12105.n7 a_30647_12105.t20 217.716
R11910 a_30647_12105.t20 a_30647_12105.t14 415.315
R11911 a_30647_12105.t14 a_30647_12105.n8 214.335
R11912 a_30647_12105.n8 a_30647_12105.t23 80.333
R11913 a_30647_12105.n8 a_30647_12105.t8 214.335
R11914 a_30647_12105.n6 a_30647_12105.n5 157.665
R11915 a_30647_12105.n5 a_30647_12105.t7 8.7
R11916 a_30647_12105.n5 a_30647_12105.t1 8.7
R11917 a_30647_12105.n4 a_30647_12105.n3 90.416
R11918 a_30647_12105.n3 a_30647_12105.t6 14.282
R11919 a_30647_12105.n3 a_30647_12105.t3 14.282
R11920 a_30647_12105.n2 a_30647_12105.n1 90.436
R11921 a_30647_12105.n1 a_30647_12105.t4 14.282
R11922 a_30647_12105.n1 a_30647_12105.t5 14.282
R11923 a_39706_24333.n0 a_39706_24333.t9 214.335
R11924 a_39706_24333.t7 a_39706_24333.n0 214.335
R11925 a_39706_24333.n1 a_39706_24333.t7 143.851
R11926 a_39706_24333.n1 a_39706_24333.t10 135.658
R11927 a_39706_24333.n0 a_39706_24333.t8 80.333
R11928 a_39706_24333.n2 a_39706_24333.t6 28.565
R11929 a_39706_24333.n2 a_39706_24333.t4 28.565
R11930 a_39706_24333.n4 a_39706_24333.t5 28.565
R11931 a_39706_24333.n4 a_39706_24333.t1 28.565
R11932 a_39706_24333.t0 a_39706_24333.n7 28.565
R11933 a_39706_24333.n7 a_39706_24333.t2 28.565
R11934 a_39706_24333.n6 a_39706_24333.t3 9.714
R11935 a_39706_24333.n7 a_39706_24333.n6 1.003
R11936 a_39706_24333.n5 a_39706_24333.n3 0.833
R11937 a_39706_24333.n3 a_39706_24333.n2 0.653
R11938 a_39706_24333.n5 a_39706_24333.n4 0.653
R11939 a_39706_24333.n6 a_39706_24333.n5 0.341
R11940 a_39706_24333.n3 a_39706_24333.n1 0.032
R11941 a_70513_19926.t0 a_70513_19926.n0 14.282
R11942 a_70513_19926.n0 a_70513_19926.t1 14.282
R11943 a_70513_19926.n0 a_70513_19926.n1 258.161
R11944 a_70513_19926.n1 a_70513_19926.n7 4.366
R11945 a_70513_19926.n7 a_70513_19926.n5 0.852
R11946 a_70513_19926.n5 a_70513_19926.n6 258.161
R11947 a_70513_19926.n6 a_70513_19926.t4 14.282
R11948 a_70513_19926.n6 a_70513_19926.t6 14.282
R11949 a_70513_19926.n5 a_70513_19926.t5 14.283
R11950 a_70513_19926.n7 a_70513_19926.n4 73.514
R11951 a_70513_19926.n4 a_70513_19926.t11 1551.5
R11952 a_70513_19926.t11 a_70513_19926.n3 656.576
R11953 a_70513_19926.n3 a_70513_19926.t2 8.7
R11954 a_70513_19926.n3 a_70513_19926.t7 8.7
R11955 a_70513_19926.n4 a_70513_19926.t9 224.129
R11956 a_70513_19926.t9 a_70513_19926.n2 207.225
R11957 a_70513_19926.n2 a_70513_19926.t8 207.225
R11958 a_70513_19926.n2 a_70513_19926.t10 80.333
R11959 a_70513_19926.n1 a_70513_19926.t3 14.283
R11960 a_23723_1259.n1 a_23723_1259.t7 867.497
R11961 a_23723_1259.n1 a_23723_1259.t6 615.911
R11962 a_23723_1259.n0 a_23723_1259.t5 286.438
R11963 a_23723_1259.n0 a_23723_1259.t4 286.438
R11964 a_23723_1259.n4 a_23723_1259.n3 185.55
R11965 a_23723_1259.t7 a_23723_1259.n0 160.666
R11966 a_23723_1259.n2 a_23723_1259.n1 135.283
R11967 a_23723_1259.n3 a_23723_1259.t1 28.568
R11968 a_23723_1259.t2 a_23723_1259.n4 28.565
R11969 a_23723_1259.n4 a_23723_1259.t0 28.565
R11970 a_23723_1259.n2 a_23723_1259.t3 20.393
R11971 a_23723_1259.n3 a_23723_1259.n2 1.831
R11972 a_49832_23623.n6 a_49832_23623.n5 501.28
R11973 a_49832_23623.t11 a_49832_23623.t12 437.233
R11974 a_49832_23623.t15 a_49832_23623.t17 415.315
R11975 a_49832_23623.t7 a_49832_23623.n3 313.873
R11976 a_49832_23623.n5 a_49832_23623.t6 294.986
R11977 a_49832_23623.n2 a_49832_23623.t16 272.288
R11978 a_49832_23623.n6 a_49832_23623.t19 236.01
R11979 a_49832_23623.n9 a_49832_23623.t11 216.627
R11980 a_49832_23623.n7 a_49832_23623.t15 216.111
R11981 a_49832_23623.n8 a_49832_23623.t9 214.686
R11982 a_49832_23623.t12 a_49832_23623.n8 214.686
R11983 a_49832_23623.n1 a_49832_23623.t4 214.335
R11984 a_49832_23623.t17 a_49832_23623.n1 214.335
R11985 a_49832_23623.n4 a_49832_23623.t7 190.152
R11986 a_49832_23623.n4 a_49832_23623.t5 190.152
R11987 a_49832_23623.n2 a_49832_23623.t13 160.666
R11988 a_49832_23623.n3 a_49832_23623.t14 160.666
R11989 a_49832_23623.n7 a_49832_23623.n6 148.428
R11990 a_49832_23623.n5 a_49832_23623.t8 110.859
R11991 a_49832_23623.n3 a_49832_23623.n2 96.129
R11992 a_49832_23623.n8 a_49832_23623.t10 80.333
R11993 a_49832_23623.n1 a_49832_23623.t18 80.333
R11994 a_49832_23623.t19 a_49832_23623.n4 80.333
R11995 a_49832_23623.t1 a_49832_23623.n11 28.57
R11996 a_49832_23623.n0 a_49832_23623.t3 28.565
R11997 a_49832_23623.n0 a_49832_23623.t2 28.565
R11998 a_49832_23623.n11 a_49832_23623.t0 17.638
R11999 a_49832_23623.n10 a_49832_23623.n9 5.6
R12000 a_49832_23623.n9 a_49832_23623.n7 2.923
R12001 a_49832_23623.n10 a_49832_23623.n0 0.69
R12002 a_49832_23623.n11 a_49832_23623.n10 0.6
R12003 a_47579_22063.n2 a_47579_22063.t7 318.922
R12004 a_47579_22063.n1 a_47579_22063.t6 273.935
R12005 a_47579_22063.n1 a_47579_22063.t5 273.935
R12006 a_47579_22063.n2 a_47579_22063.t4 269.116
R12007 a_47579_22063.n4 a_47579_22063.n0 193.227
R12008 a_47579_22063.t7 a_47579_22063.n1 179.142
R12009 a_47579_22063.n3 a_47579_22063.n2 106.999
R12010 a_47579_22063.t2 a_47579_22063.n4 28.568
R12011 a_47579_22063.n0 a_47579_22063.t0 28.565
R12012 a_47579_22063.n0 a_47579_22063.t1 28.565
R12013 a_47579_22063.n3 a_47579_22063.t3 18.149
R12014 a_47579_22063.n4 a_47579_22063.n3 3.726
R12015 a_48124_20638.t0 a_48124_20638.t1 380.209
R12016 a_16274_8992.n1 a_16274_8992.t7 990.34
R12017 a_16274_8992.n1 a_16274_8992.t6 408.211
R12018 a_16274_8992.n0 a_16274_8992.t5 286.438
R12019 a_16274_8992.n0 a_16274_8992.t4 286.438
R12020 a_16274_8992.n4 a_16274_8992.n3 185.55
R12021 a_16274_8992.t7 a_16274_8992.n0 160.666
R12022 a_16274_8992.n3 a_16274_8992.t3 28.568
R12023 a_16274_8992.t0 a_16274_8992.n4 28.565
R12024 a_16274_8992.n4 a_16274_8992.t1 28.565
R12025 a_16274_8992.n2 a_16274_8992.t2 21.5
R12026 a_16274_8992.n2 a_16274_8992.n1 12.946
R12027 a_16274_8992.n3 a_16274_8992.n2 1.537
R12028 a_16855_11724.n0 a_16855_11724.t5 14.282
R12029 a_16855_11724.t0 a_16855_11724.n0 14.282
R12030 a_16855_11724.n0 a_16855_11724.n9 89.977
R12031 a_16855_11724.n6 a_16855_11724.n7 77.784
R12032 a_16855_11724.n4 a_16855_11724.n6 77.456
R12033 a_16855_11724.n9 a_16855_11724.n4 77.456
R12034 a_16855_11724.n9 a_16855_11724.n2 75.815
R12035 a_16855_11724.n7 a_16855_11724.n8 167.433
R12036 a_16855_11724.n8 a_16855_11724.t3 14.282
R12037 a_16855_11724.n8 a_16855_11724.t2 14.282
R12038 a_16855_11724.n7 a_16855_11724.t1 104.259
R12039 a_16855_11724.n6 a_16855_11724.n5 89.977
R12040 a_16855_11724.n5 a_16855_11724.t8 14.282
R12041 a_16855_11724.n5 a_16855_11724.t7 14.282
R12042 a_16855_11724.n4 a_16855_11724.n3 89.977
R12043 a_16855_11724.n3 a_16855_11724.t6 14.282
R12044 a_16855_11724.n3 a_16855_11724.t4 14.282
R12045 a_16855_11724.n2 a_16855_11724.t10 104.259
R12046 a_16855_11724.n2 a_16855_11724.n1 167.433
R12047 a_16855_11724.n1 a_16855_11724.t9 14.282
R12048 a_16855_11724.n1 a_16855_11724.t11 14.282
R12049 a_556_10994.t0 a_556_10994.n0 14.283
R12050 a_556_10994.n0 a_556_10994.n5 0.852
R12051 a_556_10994.n5 a_556_10994.n6 4.366
R12052 a_556_10994.n6 a_556_10994.n7 258.161
R12053 a_556_10994.n7 a_556_10994.t7 14.282
R12054 a_556_10994.n7 a_556_10994.t4 14.282
R12055 a_556_10994.n6 a_556_10994.t5 14.283
R12056 a_556_10994.n5 a_556_10994.n4 97.614
R12057 a_556_10994.n4 a_556_10994.t8 200.029
R12058 a_556_10994.t8 a_556_10994.n3 206.421
R12059 a_556_10994.n3 a_556_10994.t10 80.333
R12060 a_556_10994.n3 a_556_10994.t11 206.421
R12061 a_556_10994.n4 a_556_10994.t9 1527.4
R12062 a_556_10994.t9 a_556_10994.n2 657.379
R12063 a_556_10994.n2 a_556_10994.t2 8.7
R12064 a_556_10994.n2 a_556_10994.t6 8.7
R12065 a_556_10994.n0 a_556_10994.n1 258.161
R12066 a_556_10994.n1 a_556_10994.t1 14.282
R12067 a_556_10994.n1 a_556_10994.t3 14.282
R12068 a_1916_10391.t0 a_1916_10391.t1 17.4
R12069 a_16805_8966.t0 a_16805_8966.n0 14.282
R12070 a_16805_8966.n0 a_16805_8966.t3 14.282
R12071 a_16805_8966.n0 a_16805_8966.n8 122.747
R12072 a_16805_8966.n4 a_16805_8966.n6 74.302
R12073 a_16805_8966.n8 a_16805_8966.n4 50.575
R12074 a_16805_8966.n8 a_16805_8966.n7 157.665
R12075 a_16805_8966.n7 a_16805_8966.t4 8.7
R12076 a_16805_8966.n7 a_16805_8966.t1 8.7
R12077 a_16805_8966.n6 a_16805_8966.n5 90.436
R12078 a_16805_8966.n5 a_16805_8966.t5 14.282
R12079 a_16805_8966.n5 a_16805_8966.t7 14.282
R12080 a_16805_8966.n4 a_16805_8966.n3 90.416
R12081 a_16805_8966.n3 a_16805_8966.t6 14.282
R12082 a_16805_8966.n3 a_16805_8966.t2 14.282
R12083 a_16805_8966.n6 a_16805_8966.n1 953.188
R12084 a_16805_8966.n1 a_16805_8966.t8 591.811
R12085 a_16805_8966.n1 a_16805_8966.t10 867.497
R12086 a_16805_8966.t10 a_16805_8966.n2 160.666
R12087 a_16805_8966.n2 a_16805_8966.t11 286.438
R12088 a_16805_8966.n2 a_16805_8966.t9 286.438
R12089 a_17456_7659.t0 a_17456_7659.t1 17.4
R12090 a_7464_n2148.t0 a_7464_n2148.n0 14.282
R12091 a_7464_n2148.n0 a_7464_n2148.t1 14.282
R12092 a_7464_n2148.n0 a_7464_n2148.n1 258.161
R12093 a_7464_n2148.n1 a_7464_n2148.t2 14.283
R12094 a_7464_n2148.n1 a_7464_n2148.n5 0.852
R12095 a_7464_n2148.n5 a_7464_n2148.n6 4.366
R12096 a_7464_n2148.n6 a_7464_n2148.n7 258.161
R12097 a_7464_n2148.n7 a_7464_n2148.t6 14.282
R12098 a_7464_n2148.n7 a_7464_n2148.t7 14.282
R12099 a_7464_n2148.n6 a_7464_n2148.t5 14.283
R12100 a_7464_n2148.n5 a_7464_n2148.n4 97.614
R12101 a_7464_n2148.n4 a_7464_n2148.t9 200.029
R12102 a_7464_n2148.t9 a_7464_n2148.n3 206.421
R12103 a_7464_n2148.n3 a_7464_n2148.t8 80.333
R12104 a_7464_n2148.n3 a_7464_n2148.t11 206.421
R12105 a_7464_n2148.n4 a_7464_n2148.t10 1527.4
R12106 a_7464_n2148.t10 a_7464_n2148.n2 657.379
R12107 a_7464_n2148.n2 a_7464_n2148.t3 8.7
R12108 a_7464_n2148.n2 a_7464_n2148.t4 8.7
R12109 Y[5].n1 Y[5].n0 185.55
R12110 Y[5].n1 Y[5].t1 28.568
R12111 Y[5].n0 Y[5].t2 28.565
R12112 Y[5].n0 Y[5].t0 28.565
R12113 Y[5].n2 Y[5].t3 20.393
R12114 Y[5].n2 Y[5].n1 1.827
R12115 Y[5] Y[5].n2 1.789
R12116 a_17511_8119.n2 a_17511_8119.t4 448.381
R12117 a_17511_8119.n1 a_17511_8119.t5 286.438
R12118 a_17511_8119.n1 a_17511_8119.t6 286.438
R12119 a_17511_8119.n0 a_17511_8119.t7 247.69
R12120 a_17511_8119.n4 a_17511_8119.n3 182.117
R12121 a_17511_8119.t4 a_17511_8119.n1 160.666
R12122 a_17511_8119.n3 a_17511_8119.t1 28.568
R12123 a_17511_8119.n4 a_17511_8119.t2 28.565
R12124 a_17511_8119.t0 a_17511_8119.n4 28.565
R12125 a_17511_8119.n0 a_17511_8119.t3 18.127
R12126 a_17511_8119.n2 a_17511_8119.n0 4.036
R12127 a_17511_8119.n3 a_17511_8119.n2 0.937
R12128 a_16332_8262.n0 a_16332_8262.t2 14.282
R12129 a_16332_8262.t0 a_16332_8262.n0 14.282
R12130 a_16332_8262.n0 a_16332_8262.n1 258.161
R12131 a_16332_8262.n1 a_16332_8262.n5 0.852
R12132 a_16332_8262.n5 a_16332_8262.n6 4.366
R12133 a_16332_8262.n6 a_16332_8262.n7 258.161
R12134 a_16332_8262.n7 a_16332_8262.t4 14.282
R12135 a_16332_8262.n7 a_16332_8262.t5 14.282
R12136 a_16332_8262.n6 a_16332_8262.t6 14.283
R12137 a_16332_8262.n5 a_16332_8262.n4 97.614
R12138 a_16332_8262.n4 a_16332_8262.t8 200.029
R12139 a_16332_8262.t8 a_16332_8262.n3 206.421
R12140 a_16332_8262.n3 a_16332_8262.t10 80.333
R12141 a_16332_8262.n3 a_16332_8262.t9 206.421
R12142 a_16332_8262.n4 a_16332_8262.t11 1527.4
R12143 a_16332_8262.t11 a_16332_8262.n2 657.379
R12144 a_16332_8262.n2 a_16332_8262.t3 8.7
R12145 a_16332_8262.n2 a_16332_8262.t7 8.7
R12146 a_16332_8262.n1 a_16332_8262.t1 14.283
R12147 a_16865_8992.t3 a_16865_8992.n0 14.282
R12148 a_16865_8992.n0 a_16865_8992.t9 14.282
R12149 a_16865_8992.n0 a_16865_8992.n9 89.977
R12150 a_16865_8992.n6 a_16865_8992.n7 77.784
R12151 a_16865_8992.n9 a_16865_8992.n6 77.456
R12152 a_16865_8992.n9 a_16865_8992.n4 77.456
R12153 a_16865_8992.n4 a_16865_8992.n2 75.815
R12154 a_16865_8992.n7 a_16865_8992.n8 167.433
R12155 a_16865_8992.n8 a_16865_8992.t2 14.282
R12156 a_16865_8992.n8 a_16865_8992.t1 14.282
R12157 a_16865_8992.n7 a_16865_8992.t0 104.259
R12158 a_16865_8992.n6 a_16865_8992.n5 89.977
R12159 a_16865_8992.n5 a_16865_8992.t11 14.282
R12160 a_16865_8992.n5 a_16865_8992.t7 14.282
R12161 a_16865_8992.n4 a_16865_8992.n3 89.977
R12162 a_16865_8992.n3 a_16865_8992.t10 14.282
R12163 a_16865_8992.n3 a_16865_8992.t8 14.282
R12164 a_16865_8992.n2 a_16865_8992.t4 104.259
R12165 a_16865_8992.n2 a_16865_8992.n1 167.433
R12166 a_16865_8992.n1 a_16865_8992.t6 14.282
R12167 a_16865_8992.n1 a_16865_8992.t5 14.282
R12168 a_30150_n1593.n1 a_30150_n1593.t6 318.119
R12169 a_30150_n1593.n1 a_30150_n1593.t7 269.919
R12170 a_30150_n1593.n0 a_30150_n1593.t5 267.256
R12171 a_30150_n1593.n0 a_30150_n1593.t4 267.256
R12172 a_30150_n1593.n4 a_30150_n1593.n3 193.227
R12173 a_30150_n1593.t6 a_30150_n1593.n0 160.666
R12174 a_30150_n1593.n2 a_30150_n1593.n1 106.999
R12175 a_30150_n1593.n3 a_30150_n1593.t1 28.568
R12176 a_30150_n1593.t0 a_30150_n1593.n4 28.565
R12177 a_30150_n1593.n4 a_30150_n1593.t3 28.565
R12178 a_30150_n1593.n2 a_30150_n1593.t2 18.149
R12179 a_30150_n1593.n3 a_30150_n1593.n2 3.726
R12180 a_30643_n2374.t1 a_30643_n2374.n0 14.282
R12181 a_30643_n2374.n0 a_30643_n2374.t4 14.282
R12182 a_30643_n2374.n0 a_30643_n2374.n16 90.416
R12183 a_30643_n2374.n16 a_30643_n2374.n2 74.302
R12184 a_30643_n2374.n16 a_30643_n2374.n4 50.575
R12185 a_30643_n2374.n4 a_30643_n2374.n5 110.084
R12186 a_30643_n2374.n2 a_30643_n2374.n6 664.97
R12187 a_30643_n2374.n6 a_30643_n2374.n8 16.411
R12188 a_30643_n2374.n8 a_30643_n2374.t9 198.921
R12189 a_30643_n2374.t9 a_30643_n2374.t20 415.315
R12190 a_30643_n2374.t20 a_30643_n2374.n15 214.335
R12191 a_30643_n2374.n15 a_30643_n2374.t19 80.333
R12192 a_30643_n2374.n15 a_30643_n2374.t14 214.335
R12193 a_30643_n2374.n8 a_30643_n2374.n14 861.987
R12194 a_30643_n2374.n14 a_30643_n2374.n9 560.726
R12195 a_30643_n2374.n14 a_30643_n2374.n13 65.07
R12196 a_30643_n2374.n13 a_30643_n2374.n12 6.615
R12197 a_30643_n2374.n12 a_30643_n2374.t16 93.989
R12198 a_30643_n2374.n12 a_30643_n2374.t17 198.043
R12199 a_30643_n2374.n13 a_30643_n2374.n11 97.816
R12200 a_30643_n2374.n11 a_30643_n2374.t8 80.333
R12201 a_30643_n2374.n11 a_30643_n2374.t23 394.151
R12202 a_30643_n2374.t23 a_30643_n2374.n10 269.523
R12203 a_30643_n2374.n10 a_30643_n2374.t22 160.666
R12204 a_30643_n2374.n10 a_30643_n2374.t21 269.523
R12205 a_30643_n2374.n9 a_30643_n2374.t18 294.653
R12206 a_30643_n2374.n9 a_30643_n2374.t11 111.663
R12207 a_30643_n2374.n6 a_30643_n2374.t15 217.716
R12208 a_30643_n2374.t15 a_30643_n2374.t13 415.315
R12209 a_30643_n2374.t13 a_30643_n2374.n7 214.335
R12210 a_30643_n2374.n7 a_30643_n2374.t12 80.333
R12211 a_30643_n2374.n7 a_30643_n2374.t10 214.335
R12212 a_30643_n2374.n5 a_30643_n2374.t5 14.282
R12213 a_30643_n2374.n5 a_30643_n2374.t7 14.282
R12214 a_30643_n2374.n4 a_30643_n2374.n3 157.665
R12215 a_30643_n2374.n3 a_30643_n2374.t0 8.7
R12216 a_30643_n2374.n3 a_30643_n2374.t6 8.7
R12217 a_30643_n2374.n2 a_30643_n2374.n1 90.436
R12218 a_30643_n2374.n1 a_30643_n2374.t3 14.282
R12219 a_30643_n2374.n1 a_30643_n2374.t2 14.282
R12220 a_29950_n2431.t0 a_29950_n2431.n0 14.282
R12221 a_29950_n2431.n0 a_29950_n2431.t3 14.282
R12222 a_29950_n2431.n1 a_29950_n2431.n9 0.001
R12223 a_29950_n2431.n0 a_29950_n2431.n1 267.767
R12224 a_29950_n2431.n9 a_29950_n2431.t2 14.282
R12225 a_29950_n2431.n9 a_29950_n2431.t4 14.282
R12226 a_29950_n2431.n1 a_29950_n2431.n7 0.669
R12227 a_29950_n2431.n7 a_29950_n2431.n8 1.511
R12228 a_29950_n2431.n8 a_29950_n2431.t5 14.282
R12229 a_29950_n2431.n8 a_29950_n2431.t1 14.282
R12230 a_29950_n2431.n7 a_29950_n2431.n6 0.227
R12231 a_29950_n2431.n6 a_29950_n2431.n5 0.2
R12232 a_29950_n2431.n6 a_29950_n2431.n3 0.575
R12233 a_29950_n2431.n5 a_29950_n2431.t8 16.058
R12234 a_29950_n2431.n5 a_29950_n2431.n4 0.999
R12235 a_29950_n2431.n4 a_29950_n2431.t7 14.282
R12236 a_29950_n2431.n4 a_29950_n2431.t6 14.282
R12237 a_29950_n2431.n3 a_29950_n2431.n2 0.999
R12238 a_29950_n2431.n2 a_29950_n2431.t11 14.282
R12239 a_29950_n2431.n2 a_29950_n2431.t9 14.282
R12240 a_29950_n2431.n3 a_29950_n2431.t10 16.058
R12241 a_53005_1041.n0 a_53005_1041.n12 122.999
R12242 a_53005_1041.t1 a_53005_1041.n0 14.282
R12243 a_53005_1041.n0 a_53005_1041.t2 14.282
R12244 a_53005_1041.n12 a_53005_1041.n10 50.575
R12245 a_53005_1041.n10 a_53005_1041.n8 74.302
R12246 a_53005_1041.n12 a_53005_1041.n11 157.665
R12247 a_53005_1041.n11 a_53005_1041.t4 8.7
R12248 a_53005_1041.n11 a_53005_1041.t0 8.7
R12249 a_53005_1041.n10 a_53005_1041.n9 90.416
R12250 a_53005_1041.n9 a_53005_1041.t3 14.282
R12251 a_53005_1041.n9 a_53005_1041.t5 14.282
R12252 a_53005_1041.n8 a_53005_1041.n7 90.436
R12253 a_53005_1041.n7 a_53005_1041.t7 14.282
R12254 a_53005_1041.n7 a_53005_1041.t6 14.282
R12255 a_53005_1041.n8 a_53005_1041.n1 342.688
R12256 a_53005_1041.n1 a_53005_1041.n6 126.566
R12257 a_53005_1041.n6 a_53005_1041.t9 294.653
R12258 a_53005_1041.n6 a_53005_1041.t13 111.663
R12259 a_53005_1041.n1 a_53005_1041.n5 552.333
R12260 a_53005_1041.n5 a_53005_1041.n4 6.615
R12261 a_53005_1041.n4 a_53005_1041.t14 93.989
R12262 a_53005_1041.n5 a_53005_1041.n3 97.816
R12263 a_53005_1041.n3 a_53005_1041.t10 80.333
R12264 a_53005_1041.n3 a_53005_1041.t12 394.151
R12265 a_53005_1041.t12 a_53005_1041.n2 269.523
R12266 a_53005_1041.n2 a_53005_1041.t11 160.666
R12267 a_53005_1041.n2 a_53005_1041.t8 269.523
R12268 a_53005_1041.n4 a_53005_1041.t15 198.043
R12269 a_54785_1041.n0 a_54785_1041.t4 14.282
R12270 a_54785_1041.t0 a_54785_1041.n0 14.282
R12271 a_54785_1041.n0 a_54785_1041.n9 0.999
R12272 a_54785_1041.n6 a_54785_1041.n8 0.575
R12273 a_54785_1041.n9 a_54785_1041.n6 0.2
R12274 a_54785_1041.n9 a_54785_1041.t5 16.058
R12275 a_54785_1041.n8 a_54785_1041.n7 0.999
R12276 a_54785_1041.n7 a_54785_1041.t8 14.282
R12277 a_54785_1041.n7 a_54785_1041.t7 14.282
R12278 a_54785_1041.n8 a_54785_1041.t6 16.058
R12279 a_54785_1041.n6 a_54785_1041.n4 0.227
R12280 a_54785_1041.n4 a_54785_1041.n5 1.511
R12281 a_54785_1041.n5 a_54785_1041.t9 14.282
R12282 a_54785_1041.n5 a_54785_1041.t10 14.282
R12283 a_54785_1041.n4 a_54785_1041.n1 0.669
R12284 a_54785_1041.n1 a_54785_1041.n2 0.001
R12285 a_54785_1041.n1 a_54785_1041.n3 267.767
R12286 a_54785_1041.n3 a_54785_1041.t2 14.282
R12287 a_54785_1041.n3 a_54785_1041.t1 14.282
R12288 a_54785_1041.n2 a_54785_1041.t11 14.282
R12289 a_54785_1041.n2 a_54785_1041.t3 14.282
R12290 opcode[0].n1 opcode[0].t95 1374.12
R12291 opcode[0].n4 opcode[0].t92 1374.12
R12292 opcode[0].n7 opcode[0].t107 1374.12
R12293 opcode[0].n10 opcode[0].t38 1374.12
R12294 opcode[0].n13 opcode[0].t18 1374.12
R12295 opcode[0].n16 opcode[0].t3 1374.12
R12296 opcode[0].n19 opcode[0].t64 1374.12
R12297 opcode[0].n22 opcode[0].t6 1374.12
R12298 opcode[0].n41 opcode[0].t71 1374.12
R12299 opcode[0].n44 opcode[0].t67 1374.12
R12300 opcode[0].n47 opcode[0].t220 1374.12
R12301 opcode[0].n50 opcode[0].t14 1374.12
R12302 opcode[0].n53 opcode[0].t141 1374.12
R12303 opcode[0].n56 opcode[0].t178 1374.12
R12304 opcode[0].n59 opcode[0].t133 1374.12
R12305 opcode[0].n62 opcode[0].t197 1374.12
R12306 opcode[0].n148 opcode[0].t192 1374.12
R12307 opcode[0].n152 opcode[0].t270 1374.12
R12308 opcode[0].n155 opcode[0].t24 1374.12
R12309 opcode[0].n158 opcode[0].t175 1374.12
R12310 opcode[0].n161 opcode[0].t26 1374.12
R12311 opcode[0].n164 opcode[0].t142 1374.12
R12312 opcode[0].n167 opcode[0].t126 1374.12
R12313 opcode[0].n170 opcode[0].t194 1374.12
R12314 opcode[0].n38 opcode[0].t215 623.291
R12315 opcode[0].n36 opcode[0].t65 623.291
R12316 opcode[0].n34 opcode[0].t54 623.291
R12317 opcode[0].n32 opcode[0].t271 623.291
R12318 opcode[0].n30 opcode[0].t149 623.291
R12319 opcode[0].n28 opcode[0].t253 623.291
R12320 opcode[0].n26 opcode[0].t196 623.291
R12321 opcode[0].n24 opcode[0].t117 623.291
R12322 opcode[0].n78 opcode[0].t233 623.291
R12323 opcode[0].n76 opcode[0].t108 623.291
R12324 opcode[0].n74 opcode[0].t130 623.291
R12325 opcode[0].n72 opcode[0].t229 623.291
R12326 opcode[0].n70 opcode[0].t81 623.291
R12327 opcode[0].n68 opcode[0].t121 623.291
R12328 opcode[0].n66 opcode[0].t80 623.291
R12329 opcode[0].n64 opcode[0].t171 623.291
R12330 opcode[0].n150 opcode[0].t187 623.291
R12331 opcode[0].n184 opcode[0].t11 623.291
R12332 opcode[0].n182 opcode[0].t120 623.291
R12333 opcode[0].n180 opcode[0].t217 623.291
R12334 opcode[0].n178 opcode[0].t70 623.291
R12335 opcode[0].n176 opcode[0].t139 623.291
R12336 opcode[0].n174 opcode[0].t44 623.291
R12337 opcode[0].n172 opcode[0].t131 623.291
R12338 opcode[0].n38 opcode[0].t186 610.283
R12339 opcode[0].n36 opcode[0].t182 610.283
R12340 opcode[0].n34 opcode[0].t19 610.283
R12341 opcode[0].n32 opcode[0].t213 610.283
R12342 opcode[0].n30 opcode[0].t189 610.283
R12343 opcode[0].n28 opcode[0].t168 610.283
R12344 opcode[0].n26 opcode[0].t261 610.283
R12345 opcode[0].n24 opcode[0].t75 610.283
R12346 opcode[0].n78 opcode[0].t49 610.283
R12347 opcode[0].n76 opcode[0].t136 610.283
R12348 opcode[0].n74 opcode[0].t267 610.283
R12349 opcode[0].n72 opcode[0].t45 610.283
R12350 opcode[0].n70 opcode[0].t179 610.283
R12351 opcode[0].n68 opcode[0].t216 610.283
R12352 opcode[0].n66 opcode[0].t170 610.283
R12353 opcode[0].n64 opcode[0].t5 610.283
R12354 opcode[0].n150 opcode[0].t235 610.283
R12355 opcode[0].n184 opcode[0].t22 610.283
R12356 opcode[0].n182 opcode[0].t57 610.283
R12357 opcode[0].n180 opcode[0].t254 610.283
R12358 opcode[0].n178 opcode[0].t87 610.283
R12359 opcode[0].n176 opcode[0].t180 610.283
R12360 opcode[0].n174 opcode[0].t162 610.283
R12361 opcode[0].n172 opcode[0].t237 610.283
R12362 opcode[0].n86 opcode[0].n85 501.28
R12363 opcode[0].t42 opcode[0].t46 437.233
R12364 opcode[0].n137 opcode[0].n132 436.21
R12365 opcode[0].n131 opcode[0].n126 436.21
R12366 opcode[0].n125 opcode[0].n120 436.21
R12367 opcode[0].n119 opcode[0].n114 436.21
R12368 opcode[0].n113 opcode[0].n108 436.21
R12369 opcode[0].n107 opcode[0].n102 436.21
R12370 opcode[0].n101 opcode[0].n96 436.21
R12371 opcode[0].n95 opcode[0].n90 436.21
R12372 opcode[0].t224 opcode[0].t230 415.315
R12373 opcode[0].n135 opcode[0].t76 393.348
R12374 opcode[0].n129 opcode[0].t252 393.348
R12375 opcode[0].n123 opcode[0].t242 393.348
R12376 opcode[0].n117 opcode[0].t53 393.348
R12377 opcode[0].n111 opcode[0].t174 393.348
R12378 opcode[0].n105 opcode[0].t7 393.348
R12379 opcode[0].n99 opcode[0].t98 393.348
R12380 opcode[0].n93 opcode[0].t154 393.348
R12381 opcode[0].n1 opcode[0].t181 326.034
R12382 opcode[0].n4 opcode[0].t221 326.034
R12383 opcode[0].n7 opcode[0].t199 326.034
R12384 opcode[0].n10 opcode[0].t128 326.034
R12385 opcode[0].n13 opcode[0].t27 326.034
R12386 opcode[0].n16 opcode[0].t10 326.034
R12387 opcode[0].n19 opcode[0].t158 326.034
R12388 opcode[0].n22 opcode[0].t86 326.034
R12389 opcode[0].n41 opcode[0].t231 326.034
R12390 opcode[0].n44 opcode[0].t47 326.034
R12391 opcode[0].n47 opcode[0].t156 326.034
R12392 opcode[0].n50 opcode[0].t264 326.034
R12393 opcode[0].n53 opcode[0].t106 326.034
R12394 opcode[0].n56 opcode[0].t115 326.034
R12395 opcode[0].n59 opcode[0].t73 326.034
R12396 opcode[0].n62 opcode[0].t167 326.034
R12397 opcode[0].n148 opcode[0].t218 326.034
R12398 opcode[0].n152 opcode[0].t34 326.034
R12399 opcode[0].n155 opcode[0].t249 326.034
R12400 opcode[0].n158 opcode[0].t209 326.034
R12401 opcode[0].n161 opcode[0].t99 326.034
R12402 opcode[0].n164 opcode[0].t166 326.034
R12403 opcode[0].n167 opcode[0].t66 326.034
R12404 opcode[0].n170 opcode[0].t157 326.034
R12405 opcode[0].t144 opcode[0].n83 313.873
R12406 opcode[0].n85 opcode[0].t105 294.986
R12407 opcode[0].n132 opcode[0].t25 294.653
R12408 opcode[0].n126 opcode[0].t234 294.653
R12409 opcode[0].n120 opcode[0].t185 294.653
R12410 opcode[0].n114 opcode[0].t12 294.653
R12411 opcode[0].n108 opcode[0].t122 294.653
R12412 opcode[0].n102 opcode[0].t227 294.653
R12413 opcode[0].n96 opcode[0].t245 294.653
R12414 opcode[0].n90 opcode[0].t20 294.653
R12415 opcode[0].n2 opcode[0].t33 286.438
R12416 opcode[0].n2 opcode[0].t119 286.438
R12417 opcode[0].n5 opcode[0].t243 286.438
R12418 opcode[0].n5 opcode[0].t269 286.438
R12419 opcode[0].n8 opcode[0].t145 286.438
R12420 opcode[0].n8 opcode[0].t169 286.438
R12421 opcode[0].n11 opcode[0].t69 286.438
R12422 opcode[0].n11 opcode[0].t165 286.438
R12423 opcode[0].n14 opcode[0].t146 286.438
R12424 opcode[0].n14 opcode[0].t1 286.438
R12425 opcode[0].n17 opcode[0].t123 286.438
R12426 opcode[0].n17 opcode[0].t257 286.438
R12427 opcode[0].n20 opcode[0].t17 286.438
R12428 opcode[0].n20 opcode[0].t102 286.438
R12429 opcode[0].n23 opcode[0].t212 286.438
R12430 opcode[0].n23 opcode[0].t247 286.438
R12431 opcode[0].n42 opcode[0].t226 286.438
R12432 opcode[0].n42 opcode[0].t244 286.438
R12433 opcode[0].n45 opcode[0].t37 286.438
R12434 opcode[0].n45 opcode[0].t112 286.438
R12435 opcode[0].n48 opcode[0].t124 286.438
R12436 opcode[0].n48 opcode[0].t241 286.438
R12437 opcode[0].n51 opcode[0].t219 286.438
R12438 opcode[0].n51 opcode[0].t236 286.438
R12439 opcode[0].n54 opcode[0].t104 286.438
R12440 opcode[0].n54 opcode[0].t153 286.438
R12441 opcode[0].n57 opcode[0].t113 286.438
R12442 opcode[0].n57 opcode[0].t193 286.438
R12443 opcode[0].n60 opcode[0].t72 286.438
R12444 opcode[0].n60 opcode[0].t85 286.438
R12445 opcode[0].n63 opcode[0].t164 286.438
R12446 opcode[0].n63 opcode[0].t260 286.438
R12447 opcode[0].n149 opcode[0].t184 286.438
R12448 opcode[0].n149 opcode[0].t195 286.438
R12449 opcode[0].n153 opcode[0].t32 286.438
R12450 opcode[0].n153 opcode[0].t74 286.438
R12451 opcode[0].n156 opcode[0].t51 286.438
R12452 opcode[0].n156 opcode[0].t36 286.438
R12453 opcode[0].n159 opcode[0].t206 286.438
R12454 opcode[0].n159 opcode[0].t223 286.438
R12455 opcode[0].n162 opcode[0].t63 286.438
R12456 opcode[0].n162 opcode[0].t78 286.438
R12457 opcode[0].n165 opcode[0].t62 286.438
R12458 opcode[0].n165 opcode[0].t250 286.438
R12459 opcode[0].n168 opcode[0].t39 286.438
R12460 opcode[0].n168 opcode[0].t50 286.438
R12461 opcode[0].n171 opcode[0].t125 286.438
R12462 opcode[0].n171 opcode[0].t137 286.438
R12463 opcode[0].n82 opcode[0].t138 272.288
R12464 opcode[0].n134 opcode[0].t239 270.326
R12465 opcode[0].t76 opcode[0].n134 270.326
R12466 opcode[0].n128 opcode[0].t118 270.326
R12467 opcode[0].t252 opcode[0].n128 270.326
R12468 opcode[0].n122 opcode[0].t91 270.326
R12469 opcode[0].t242 opcode[0].n122 270.326
R12470 opcode[0].n116 opcode[0].t176 270.326
R12471 opcode[0].t53 opcode[0].n116 270.326
R12472 opcode[0].n110 opcode[0].t240 270.326
R12473 opcode[0].t174 opcode[0].n110 270.326
R12474 opcode[0].n104 opcode[0].t52 270.326
R12475 opcode[0].t7 opcode[0].n104 270.326
R12476 opcode[0].n98 opcode[0].t228 270.326
R12477 opcode[0].t98 opcode[0].n98 270.326
R12478 opcode[0].n92 opcode[0].t23 270.326
R12479 opcode[0].t154 opcode[0].n92 270.326
R12480 opcode[0].n137 opcode[0].n136 248.23
R12481 opcode[0].n131 opcode[0].n130 248.23
R12482 opcode[0].n125 opcode[0].n124 248.23
R12483 opcode[0].n119 opcode[0].n118 248.23
R12484 opcode[0].n113 opcode[0].n112 248.23
R12485 opcode[0].n107 opcode[0].n106 248.23
R12486 opcode[0].n101 opcode[0].n100 248.23
R12487 opcode[0].n95 opcode[0].n94 248.23
R12488 opcode[0].n86 opcode[0].t147 236.01
R12489 opcode[0].n89 opcode[0].t42 216.627
R12490 opcode[0].n87 opcode[0].t224 216.111
R12491 opcode[0].n88 opcode[0].t248 214.686
R12492 opcode[0].t46 opcode[0].n88 214.686
R12493 opcode[0].n81 opcode[0].t246 214.335
R12494 opcode[0].t230 opcode[0].n81 214.335
R12495 opcode[0].n0 opcode[0].t4 206.421
R12496 opcode[0].t181 opcode[0].n0 206.421
R12497 opcode[0].n3 opcode[0].t0 206.421
R12498 opcode[0].t221 opcode[0].n3 206.421
R12499 opcode[0].n6 opcode[0].t183 206.421
R12500 opcode[0].t199 opcode[0].n6 206.421
R12501 opcode[0].n9 opcode[0].t103 206.421
R12502 opcode[0].t128 opcode[0].n9 206.421
R12503 opcode[0].n12 opcode[0].t9 206.421
R12504 opcode[0].t27 opcode[0].n12 206.421
R12505 opcode[0].n15 opcode[0].t268 206.421
R12506 opcode[0].t10 opcode[0].n15 206.421
R12507 opcode[0].n18 opcode[0].t263 206.421
R12508 opcode[0].t158 opcode[0].n18 206.421
R12509 opcode[0].n21 opcode[0].t258 206.421
R12510 opcode[0].t86 opcode[0].n21 206.421
R12511 opcode[0].n40 opcode[0].t255 206.421
R12512 opcode[0].t231 opcode[0].n40 206.421
R12513 opcode[0].n43 opcode[0].t251 206.421
R12514 opcode[0].t47 opcode[0].n43 206.421
R12515 opcode[0].n46 opcode[0].t77 206.421
R12516 opcode[0].t156 opcode[0].n46 206.421
R12517 opcode[0].n49 opcode[0].t143 206.421
R12518 opcode[0].t264 opcode[0].n49 206.421
R12519 opcode[0].n52 opcode[0].t13 206.421
R12520 opcode[0].t106 opcode[0].n52 206.421
R12521 opcode[0].n55 opcode[0].t41 206.421
R12522 opcode[0].t115 opcode[0].n55 206.421
R12523 opcode[0].n58 opcode[0].t94 206.421
R12524 opcode[0].t73 opcode[0].n58 206.421
R12525 opcode[0].n61 opcode[0].t90 206.421
R12526 opcode[0].t167 opcode[0].n61 206.421
R12527 opcode[0].n147 opcode[0].t200 206.421
R12528 opcode[0].t218 opcode[0].n147 206.421
R12529 opcode[0].n151 opcode[0].t198 206.421
R12530 opcode[0].t34 opcode[0].n151 206.421
R12531 opcode[0].n154 opcode[0].t155 206.421
R12532 opcode[0].t249 opcode[0].n154 206.421
R12533 opcode[0].n157 opcode[0].t134 206.421
R12534 opcode[0].t209 opcode[0].n157 206.421
R12535 opcode[0].n160 opcode[0].t8 206.421
R12536 opcode[0].t99 opcode[0].n160 206.421
R12537 opcode[0].n163 opcode[0].t84 206.421
R12538 opcode[0].t166 opcode[0].n163 206.421
R12539 opcode[0].n166 opcode[0].t2 206.421
R12540 opcode[0].t66 opcode[0].n166 206.421
R12541 opcode[0].n169 opcode[0].t55 206.421
R12542 opcode[0].t157 opcode[0].n169 206.421
R12543 opcode[0].n133 opcode[0].t191 197.241
R12544 opcode[0].n127 opcode[0].t28 197.241
R12545 opcode[0].n121 opcode[0].t83 197.241
R12546 opcode[0].n115 opcode[0].t163 197.241
R12547 opcode[0].n109 opcode[0].t225 197.241
R12548 opcode[0].n103 opcode[0].t43 197.241
R12549 opcode[0].n97 opcode[0].t48 197.241
R12550 opcode[0].n91 opcode[0].t129 197.241
R12551 opcode[0].n84 opcode[0].t144 190.152
R12552 opcode[0].n84 opcode[0].t232 190.152
R12553 opcode[0].t215 opcode[0].n2 160.666
R12554 opcode[0].t65 opcode[0].n5 160.666
R12555 opcode[0].t54 opcode[0].n8 160.666
R12556 opcode[0].t271 opcode[0].n11 160.666
R12557 opcode[0].t149 opcode[0].n14 160.666
R12558 opcode[0].t253 opcode[0].n17 160.666
R12559 opcode[0].t196 opcode[0].n20 160.666
R12560 opcode[0].t117 opcode[0].n23 160.666
R12561 opcode[0].t233 opcode[0].n42 160.666
R12562 opcode[0].t108 opcode[0].n45 160.666
R12563 opcode[0].t130 opcode[0].n48 160.666
R12564 opcode[0].t229 opcode[0].n51 160.666
R12565 opcode[0].t81 opcode[0].n54 160.666
R12566 opcode[0].t121 opcode[0].n57 160.666
R12567 opcode[0].t80 opcode[0].n60 160.666
R12568 opcode[0].t171 opcode[0].n63 160.666
R12569 opcode[0].n82 opcode[0].t214 160.666
R12570 opcode[0].n83 opcode[0].t188 160.666
R12571 opcode[0].n134 opcode[0].t114 160.666
R12572 opcode[0].n128 opcode[0].t140 160.666
R12573 opcode[0].n122 opcode[0].t116 160.666
R12574 opcode[0].n116 opcode[0].t16 160.666
R12575 opcode[0].n110 opcode[0].t61 160.666
R12576 opcode[0].n104 opcode[0].t159 160.666
R12577 opcode[0].n98 opcode[0].t56 160.666
R12578 opcode[0].n92 opcode[0].t127 160.666
R12579 opcode[0].t187 opcode[0].n149 160.666
R12580 opcode[0].t11 opcode[0].n153 160.666
R12581 opcode[0].t120 opcode[0].n156 160.666
R12582 opcode[0].t217 opcode[0].n159 160.666
R12583 opcode[0].t70 opcode[0].n162 160.666
R12584 opcode[0].t139 opcode[0].n165 160.666
R12585 opcode[0].t44 opcode[0].n168 160.666
R12586 opcode[0].t131 opcode[0].n171 160.666
R12587 opcode[0].n87 opcode[0].n86 148.428
R12588 opcode[0].n138 opcode[0].n137 121.522
R12589 opcode[0].n144 opcode[0].n95 119.477
R12590 opcode[0].n143 opcode[0].n101 118.483
R12591 opcode[0].n140 opcode[0].n119 118.277
R12592 opcode[0].n141 opcode[0].n113 118.275
R12593 opcode[0].n142 opcode[0].n107 118.132
R12594 opcode[0].n138 opcode[0].n131 118.08
R12595 opcode[0].n139 opcode[0].n125 118.08
R12596 opcode[0].n132 opcode[0].t211 111.663
R12597 opcode[0].n126 opcode[0].t202 111.663
R12598 opcode[0].n120 opcode[0].t58 111.663
R12599 opcode[0].n114 opcode[0].t152 111.663
R12600 opcode[0].n108 opcode[0].t208 111.663
R12601 opcode[0].n102 opcode[0].t35 111.663
R12602 opcode[0].n96 opcode[0].t30 111.663
R12603 opcode[0].n90 opcode[0].t97 111.663
R12604 opcode[0].n85 opcode[0].t148 110.859
R12605 opcode[0].n136 opcode[0].n135 97.816
R12606 opcode[0].n130 opcode[0].n129 97.816
R12607 opcode[0].n124 opcode[0].n123 97.816
R12608 opcode[0].n118 opcode[0].n117 97.816
R12609 opcode[0].n112 opcode[0].n111 97.816
R12610 opcode[0].n106 opcode[0].n105 97.816
R12611 opcode[0].n100 opcode[0].n99 97.816
R12612 opcode[0].n94 opcode[0].n93 97.816
R12613 opcode[0].n83 opcode[0].n82 96.129
R12614 opcode[0].n133 opcode[0].t29 93.989
R12615 opcode[0].n127 opcode[0].t190 93.989
R12616 opcode[0].n121 opcode[0].t265 93.989
R12617 opcode[0].n115 opcode[0].t135 93.989
R12618 opcode[0].n109 opcode[0].t109 93.989
R12619 opcode[0].n103 opcode[0].t205 93.989
R12620 opcode[0].n97 opcode[0].t210 93.989
R12621 opcode[0].n91 opcode[0].t15 93.989
R12622 opcode[0].n0 opcode[0].t177 80.333
R12623 opcode[0].n3 opcode[0].t172 80.333
R12624 opcode[0].n6 opcode[0].t21 80.333
R12625 opcode[0].n9 opcode[0].t222 80.333
R12626 opcode[0].n12 opcode[0].t110 80.333
R12627 opcode[0].n15 opcode[0].t88 80.333
R12628 opcode[0].n18 opcode[0].t266 80.333
R12629 opcode[0].n21 opcode[0].t151 80.333
R12630 opcode[0].n40 opcode[0].t262 80.333
R12631 opcode[0].n43 opcode[0].t259 80.333
R12632 opcode[0].n46 opcode[0].t150 80.333
R12633 opcode[0].n49 opcode[0].t256 80.333
R12634 opcode[0].n52 opcode[0].t101 80.333
R12635 opcode[0].n55 opcode[0].t111 80.333
R12636 opcode[0].n58 opcode[0].t68 80.333
R12637 opcode[0].n61 opcode[0].t96 80.333
R12638 opcode[0].n88 opcode[0].t40 80.333
R12639 opcode[0].n81 opcode[0].t238 80.333
R12640 opcode[0].t147 opcode[0].n84 80.333
R12641 opcode[0].n135 opcode[0].t132 80.333
R12642 opcode[0].n129 opcode[0].t79 80.333
R12643 opcode[0].n123 opcode[0].t204 80.333
R12644 opcode[0].n117 opcode[0].t31 80.333
R12645 opcode[0].n111 opcode[0].t82 80.333
R12646 opcode[0].n105 opcode[0].t161 80.333
R12647 opcode[0].n99 opcode[0].t100 80.333
R12648 opcode[0].n93 opcode[0].t173 80.333
R12649 opcode[0].n147 opcode[0].t207 80.333
R12650 opcode[0].n151 opcode[0].t203 80.333
R12651 opcode[0].n154 opcode[0].t160 80.333
R12652 opcode[0].n157 opcode[0].t201 80.333
R12653 opcode[0].n160 opcode[0].t93 80.333
R12654 opcode[0].n163 opcode[0].t89 80.333
R12655 opcode[0].n166 opcode[0].t60 80.333
R12656 opcode[0].n169 opcode[0].t59 80.333
R12657 opcode[0] opcode[0].n188 46.46
R12658 opcode[0].n146 opcode[0].n80 17.359
R12659 opcode[0].n145 opcode[0].n144 11.636
R12660 opcode[0].n136 opcode[0].n133 6.615
R12661 opcode[0].n130 opcode[0].n127 6.615
R12662 opcode[0].n124 opcode[0].n121 6.615
R12663 opcode[0].n118 opcode[0].n115 6.615
R12664 opcode[0].n112 opcode[0].n109 6.615
R12665 opcode[0].n106 opcode[0].n103 6.615
R12666 opcode[0].n100 opcode[0].n97 6.615
R12667 opcode[0].n94 opcode[0].n91 6.615
R12668 opcode[0].n80 opcode[0].n79 4.765
R12669 opcode[0].n80 opcode[0].n39 3.91
R12670 opcode[0].n144 opcode[0].n143 3.481
R12671 opcode[0].n141 opcode[0].n140 3.446
R12672 opcode[0].n139 opcode[0].n138 3.446
R12673 opcode[0].n140 opcode[0].n139 3.445
R12674 opcode[0].n142 opcode[0].n141 3.44
R12675 opcode[0].n143 opcode[0].n142 3.433
R12676 opcode[0].n145 opcode[0].n89 3.293
R12677 opcode[0].n180 opcode[0].n179 3.277
R12678 opcode[0].n72 opcode[0].n71 3.143
R12679 opcode[0].n32 opcode[0].n31 3.102
R12680 opcode[0].n70 opcode[0].n69 3.059
R12681 opcode[0].n78 opcode[0].n77 3.059
R12682 opcode[0].n174 opcode[0].n173 3.059
R12683 opcode[0].n182 opcode[0].n181 3.059
R12684 opcode[0].n186 opcode[0].n185 3.058
R12685 opcode[0].n66 opcode[0].n65 3.037
R12686 opcode[0].n74 opcode[0].n73 3.037
R12687 opcode[0].n178 opcode[0].n177 3.028
R12688 opcode[0].n68 opcode[0].n67 3.022
R12689 opcode[0].n76 opcode[0].n75 3.022
R12690 opcode[0].n30 opcode[0].n29 3.021
R12691 opcode[0].n38 opcode[0].n37 3.021
R12692 opcode[0].n146 opcode[0].n145 3.016
R12693 opcode[0].n26 opcode[0].n25 2.998
R12694 opcode[0].n34 opcode[0].n33 2.998
R12695 opcode[0].n28 opcode[0].n27 2.985
R12696 opcode[0].n36 opcode[0].n35 2.984
R12697 opcode[0].n89 opcode[0].n87 2.923
R12698 opcode[0].n184 opcode[0].n183 2.922
R12699 opcode[0].n176 opcode[0].n175 2.917
R12700 opcode[0].n188 opcode[0].n146 2.581
R12701 opcode[0].n187 opcode[0].n186 1.616
R12702 opcode[0].n173 opcode[0].n172 1.614
R12703 opcode[0].n79 opcode[0].n78 1.614
R12704 opcode[0].n77 opcode[0].n76 1.614
R12705 opcode[0].n71 opcode[0].n70 1.614
R12706 opcode[0].n69 opcode[0].n68 1.614
R12707 opcode[0].n183 opcode[0].n182 1.614
R12708 opcode[0].n181 opcode[0].n180 1.614
R12709 opcode[0].n175 opcode[0].n174 1.614
R12710 opcode[0].n179 opcode[0].n178 1.613
R12711 opcode[0].n177 opcode[0].n176 1.61
R12712 opcode[0].n185 opcode[0].n184 1.608
R12713 opcode[0].n39 opcode[0].n38 1.595
R12714 opcode[0].n37 opcode[0].n36 1.595
R12715 opcode[0].n31 opcode[0].n30 1.595
R12716 opcode[0].n29 opcode[0].n28 1.595
R12717 opcode[0].n75 opcode[0].n74 1.541
R12718 opcode[0].n73 opcode[0].n72 1.541
R12719 opcode[0].n67 opcode[0].n66 1.541
R12720 opcode[0].n65 opcode[0].n64 1.541
R12721 opcode[0].n35 opcode[0].n34 1.523
R12722 opcode[0].n33 opcode[0].n32 1.523
R12723 opcode[0].n27 opcode[0].n26 1.523
R12724 opcode[0].n25 opcode[0].n24 1.523
R12725 opcode[0].n188 opcode[0].n187 1.017
R12726 opcode[0].n35 opcode[0].n7 0.003
R12727 opcode[0].n33 opcode[0].n10 0.003
R12728 opcode[0].n27 opcode[0].n19 0.003
R12729 opcode[0].n25 opcode[0].n22 0.003
R12730 opcode[0].n75 opcode[0].n47 0.003
R12731 opcode[0].n73 opcode[0].n50 0.003
R12732 opcode[0].n67 opcode[0].n59 0.003
R12733 opcode[0].n65 opcode[0].n62 0.003
R12734 opcode[0].n39 opcode[0].n1 0.003
R12735 opcode[0].n37 opcode[0].n4 0.003
R12736 opcode[0].n31 opcode[0].n13 0.003
R12737 opcode[0].n29 opcode[0].n16 0.003
R12738 opcode[0].n79 opcode[0].n41 0.003
R12739 opcode[0].n77 opcode[0].n44 0.003
R12740 opcode[0].n71 opcode[0].n53 0.003
R12741 opcode[0].n69 opcode[0].n56 0.003
R12742 opcode[0].n187 opcode[0].n148 0.003
R12743 opcode[0].n185 opcode[0].n152 0.003
R12744 opcode[0].n183 opcode[0].n155 0.003
R12745 opcode[0].n181 opcode[0].n158 0.003
R12746 opcode[0].n179 opcode[0].n161 0.003
R12747 opcode[0].n177 opcode[0].n164 0.003
R12748 opcode[0].n175 opcode[0].n167 0.003
R12749 opcode[0].n173 opcode[0].n170 0.003
R12750 opcode[0].n186 opcode[0].n150 0.001
R12751 a_20643_8115.n2 a_20643_8115.t6 448.381
R12752 a_20643_8115.n1 a_20643_8115.t7 286.438
R12753 a_20643_8115.n1 a_20643_8115.t5 286.438
R12754 a_20643_8115.n0 a_20643_8115.t4 247.69
R12755 a_20643_8115.n4 a_20643_8115.n3 182.117
R12756 a_20643_8115.t6 a_20643_8115.n1 160.666
R12757 a_20643_8115.n3 a_20643_8115.t0 28.568
R12758 a_20643_8115.n4 a_20643_8115.t1 28.565
R12759 a_20643_8115.t2 a_20643_8115.n4 28.565
R12760 a_20643_8115.n0 a_20643_8115.t3 18.127
R12761 a_20643_8115.n2 a_20643_8115.n0 4.036
R12762 a_20643_8115.n3 a_20643_8115.n2 0.937
R12763 B[7].t16 B[7].t17 799.268
R12764 B[7].n9 B[7].n1 648.503
R12765 B[7].n7 B[7].n6 618.566
R12766 B[7].n14 B[7].n10 592.056
R12767 B[7].t1 B[7].t5 415.315
R12768 B[7].t10 B[7].n4 313.873
R12769 B[7].t13 B[7].n12 313.069
R12770 B[7].n10 B[7].t14 294.986
R12771 B[7].n0 B[7].t9 285.543
R12772 B[7].n6 B[7].t12 273.077
R12773 B[7].n3 B[7].t4 272.288
R12774 B[7].n11 B[7].t6 271.484
R12775 B[7].n8 B[7].t1 217.471
R12776 B[7].n2 B[7].t22 214.335
R12777 B[7].t5 B[7].n2 214.335
R12778 B[7].n7 B[7].t23 204.679
R12779 B[7].n14 B[7].t21 204.672
R12780 B[7].n1 B[7].t16 194.406
R12781 B[7].n13 B[7].t13 190.955
R12782 B[7].n13 B[7].t7 190.955
R12783 B[7].n5 B[7].t8 190.152
R12784 B[7].n5 B[7].t10 190.152
R12785 B[7].n12 B[7].t2 160.666
R12786 B[7].n11 B[7].t15 160.666
R12787 B[7].n0 B[7].t11 160.666
R12788 B[7].n3 B[7].t18 160.666
R12789 B[7].n4 B[7].t3 160.666
R12790 B[7].n6 B[7].t19 137.369
R12791 B[7].n10 B[7].t20 110.859
R12792 B[7].n12 B[7].n11 96.129
R12793 B[7].n4 B[7].n3 96.129
R12794 B[7].n1 B[7].n0 91.137
R12795 B[7].n15 B[7].n14 85.657
R12796 B[7].t21 B[7].n13 80.333
R12797 B[7].n2 B[7].t0 80.333
R12798 B[7].t23 B[7].n5 80.333
R12799 B[7].n8 B[7].n7 61.582
R12800 B[7] B[7].n15 47.62
R12801 B[7].n15 B[7].n9 36.576
R12802 B[7].n9 B[7].n8 6.998
R12803 a_13849_16387.n0 a_13849_16387.t8 214.335
R12804 a_13849_16387.t7 a_13849_16387.n0 214.335
R12805 a_13849_16387.n1 a_13849_16387.t7 143.851
R12806 a_13849_16387.n1 a_13849_16387.t10 135.658
R12807 a_13849_16387.n0 a_13849_16387.t9 80.333
R12808 a_13849_16387.n2 a_13849_16387.t3 28.565
R12809 a_13849_16387.n2 a_13849_16387.t4 28.565
R12810 a_13849_16387.n4 a_13849_16387.t5 28.565
R12811 a_13849_16387.n4 a_13849_16387.t1 28.565
R12812 a_13849_16387.t2 a_13849_16387.n7 28.565
R12813 a_13849_16387.n7 a_13849_16387.t0 28.565
R12814 a_13849_16387.n3 a_13849_16387.t6 9.714
R12815 a_13849_16387.n3 a_13849_16387.n2 1.003
R12816 a_13849_16387.n6 a_13849_16387.n5 0.833
R12817 a_13849_16387.n5 a_13849_16387.n4 0.653
R12818 a_13849_16387.n7 a_13849_16387.n6 0.653
R12819 a_13849_16387.n5 a_13849_16387.n3 0.341
R12820 a_13849_16387.n6 a_13849_16387.n1 0.032
R12821 a_63532_11802.n0 a_63532_11802.t8 214.335
R12822 a_63532_11802.t10 a_63532_11802.n0 214.335
R12823 a_63532_11802.n1 a_63532_11802.t10 143.851
R12824 a_63532_11802.n1 a_63532_11802.t9 135.658
R12825 a_63532_11802.n0 a_63532_11802.t7 80.333
R12826 a_63532_11802.n2 a_63532_11802.t0 28.565
R12827 a_63532_11802.n2 a_63532_11802.t1 28.565
R12828 a_63532_11802.n4 a_63532_11802.t2 28.565
R12829 a_63532_11802.n4 a_63532_11802.t6 28.565
R12830 a_63532_11802.n7 a_63532_11802.t5 28.565
R12831 a_63532_11802.t4 a_63532_11802.n7 28.565
R12832 a_63532_11802.n6 a_63532_11802.t3 9.714
R12833 a_63532_11802.n7 a_63532_11802.n6 1.003
R12834 a_63532_11802.n5 a_63532_11802.n3 0.833
R12835 a_63532_11802.n3 a_63532_11802.n2 0.653
R12836 a_63532_11802.n5 a_63532_11802.n4 0.653
R12837 a_63532_11802.n6 a_63532_11802.n5 0.341
R12838 a_63532_11802.n3 a_63532_11802.n1 0.032
R12839 a_51695_9365.t5 a_51695_9365.t6 800.071
R12840 a_51695_9365.n2 a_51695_9365.n1 659.097
R12841 a_51695_9365.n0 a_51695_9365.t7 285.109
R12842 a_51695_9365.n1 a_51695_9365.t5 193.602
R12843 a_51695_9365.n4 a_51695_9365.n3 192.754
R12844 a_51695_9365.n0 a_51695_9365.t4 160.666
R12845 a_51695_9365.n1 a_51695_9365.n0 91.507
R12846 a_51695_9365.n3 a_51695_9365.t2 28.568
R12847 a_51695_9365.t0 a_51695_9365.n4 28.565
R12848 a_51695_9365.n4 a_51695_9365.t1 28.565
R12849 a_51695_9365.n2 a_51695_9365.t3 19.061
R12850 a_51695_9365.n3 a_51695_9365.n2 1.005
R12851 a_53430_9674.n0 a_53430_9674.t4 14.282
R12852 a_53430_9674.n0 a_53430_9674.t2 14.282
R12853 a_53430_9674.n1 a_53430_9674.t3 14.282
R12854 a_53430_9674.n1 a_53430_9674.t5 14.282
R12855 a_53430_9674.n3 a_53430_9674.t1 14.282
R12856 a_53430_9674.t0 a_53430_9674.n3 14.282
R12857 a_53430_9674.n3 a_53430_9674.n2 2.546
R12858 a_53430_9674.n2 a_53430_9674.n1 2.367
R12859 a_53430_9674.n2 a_53430_9674.n0 0.001
R12860 a_498_11724.n2 a_498_11724.t4 990.34
R12861 a_498_11724.n2 a_498_11724.t7 408.211
R12862 a_498_11724.n1 a_498_11724.t5 286.438
R12863 a_498_11724.n1 a_498_11724.t6 286.438
R12864 a_498_11724.n4 a_498_11724.n0 185.55
R12865 a_498_11724.t4 a_498_11724.n1 160.666
R12866 a_498_11724.t2 a_498_11724.n4 28.568
R12867 a_498_11724.n0 a_498_11724.t0 28.565
R12868 a_498_11724.n0 a_498_11724.t1 28.565
R12869 a_498_11724.n3 a_498_11724.t3 21.376
R12870 a_498_11724.n3 a_498_11724.n2 10.434
R12871 a_498_11724.n4 a_498_11724.n3 1.537
R12872 a_807_1740.t0 a_807_1740.n0 14.282
R12873 a_807_1740.n0 a_807_1740.t7 14.282
R12874 a_807_1740.n0 a_807_1740.n9 89.977
R12875 a_807_1740.n6 a_807_1740.n7 75.815
R12876 a_807_1740.n9 a_807_1740.n6 77.456
R12877 a_807_1740.n9 a_807_1740.n4 77.456
R12878 a_807_1740.n4 a_807_1740.n2 77.784
R12879 a_807_1740.n7 a_807_1740.n8 167.433
R12880 a_807_1740.n8 a_807_1740.t10 14.282
R12881 a_807_1740.n8 a_807_1740.t11 14.282
R12882 a_807_1740.n7 a_807_1740.t9 104.259
R12883 a_807_1740.n6 a_807_1740.n5 89.977
R12884 a_807_1740.n5 a_807_1740.t2 14.282
R12885 a_807_1740.n5 a_807_1740.t1 14.282
R12886 a_807_1740.n4 a_807_1740.n3 89.977
R12887 a_807_1740.n3 a_807_1740.t8 14.282
R12888 a_807_1740.n3 a_807_1740.t6 14.282
R12889 a_807_1740.n2 a_807_1740.t3 104.259
R12890 a_807_1740.n2 a_807_1740.n1 167.433
R12891 a_807_1740.n1 a_807_1740.t5 14.282
R12892 a_807_1740.n1 a_807_1740.t4 14.282
R12893 a_10519_8988.n0 a_10519_8988.n9 167.433
R12894 a_10519_8988.n0 a_10519_8988.t4 14.282
R12895 a_10519_8988.t3 a_10519_8988.n0 14.282
R12896 a_10519_8988.n9 a_10519_8988.n8 77.784
R12897 a_10519_8988.n8 a_10519_8988.n6 77.456
R12898 a_10519_8988.n6 a_10519_8988.n4 77.456
R12899 a_10519_8988.n4 a_10519_8988.n2 75.815
R12900 a_10519_8988.n9 a_10519_8988.t5 104.259
R12901 a_10519_8988.n8 a_10519_8988.n7 89.977
R12902 a_10519_8988.n7 a_10519_8988.t1 14.282
R12903 a_10519_8988.n7 a_10519_8988.t0 14.282
R12904 a_10519_8988.n6 a_10519_8988.n5 89.977
R12905 a_10519_8988.n5 a_10519_8988.t2 14.282
R12906 a_10519_8988.n5 a_10519_8988.t11 14.282
R12907 a_10519_8988.n4 a_10519_8988.n3 89.977
R12908 a_10519_8988.n3 a_10519_8988.t10 14.282
R12909 a_10519_8988.n3 a_10519_8988.t6 14.282
R12910 a_10519_8988.n2 a_10519_8988.t9 104.259
R12911 a_10519_8988.n2 a_10519_8988.n1 167.433
R12912 a_10519_8988.n1 a_10519_8988.t7 14.282
R12913 a_10519_8988.n1 a_10519_8988.t8 14.282
R12914 a_57739_6616.n4 a_57739_6616.t7 214.335
R12915 a_57739_6616.t10 a_57739_6616.n4 214.335
R12916 a_57739_6616.n5 a_57739_6616.t10 143.851
R12917 a_57739_6616.n5 a_57739_6616.t8 135.658
R12918 a_57739_6616.n4 a_57739_6616.t9 80.333
R12919 a_57739_6616.n0 a_57739_6616.t0 28.565
R12920 a_57739_6616.n0 a_57739_6616.t2 28.565
R12921 a_57739_6616.n2 a_57739_6616.t5 28.565
R12922 a_57739_6616.n2 a_57739_6616.t1 28.565
R12923 a_57739_6616.n7 a_57739_6616.t6 28.565
R12924 a_57739_6616.t4 a_57739_6616.n7 28.565
R12925 a_57739_6616.n1 a_57739_6616.t3 9.714
R12926 a_57739_6616.n1 a_57739_6616.n0 1.003
R12927 a_57739_6616.n6 a_57739_6616.n3 0.833
R12928 a_57739_6616.n3 a_57739_6616.n2 0.653
R12929 a_57739_6616.n7 a_57739_6616.n6 0.653
R12930 a_57739_6616.n3 a_57739_6616.n1 0.341
R12931 a_57739_6616.n6 a_57739_6616.n5 0.032
R12932 a_58329_6179.t7 a_58329_6179.t6 574.43
R12933 a_58329_6179.n1 a_58329_6179.t4 285.109
R12934 a_58329_6179.n3 a_58329_6179.n2 197.217
R12935 a_58329_6179.n4 a_58329_6179.n0 192.754
R12936 a_58329_6179.n1 a_58329_6179.t5 160.666
R12937 a_58329_6179.n2 a_58329_6179.t7 160.666
R12938 a_58329_6179.n2 a_58329_6179.n1 114.829
R12939 a_58329_6179.t2 a_58329_6179.n4 28.568
R12940 a_58329_6179.n0 a_58329_6179.t1 28.565
R12941 a_58329_6179.n0 a_58329_6179.t0 28.565
R12942 a_58329_6179.n3 a_58329_6179.t3 18.838
R12943 a_58329_6179.n4 a_58329_6179.n3 1.129
R12944 a_41507_3295.n8 a_41507_3295.n7 861.987
R12945 a_41507_3295.n7 a_41507_3295.n6 560.726
R12946 a_41507_3295.t13 a_41507_3295.t12 415.315
R12947 a_41507_3295.t5 a_41507_3295.t14 415.315
R12948 a_41507_3295.n3 a_41507_3295.t9 394.151
R12949 a_41507_3295.n6 a_41507_3295.t19 294.653
R12950 a_41507_3295.n2 a_41507_3295.t11 269.523
R12951 a_41507_3295.t9 a_41507_3295.n2 269.523
R12952 a_41507_3295.n10 a_41507_3295.t13 217.716
R12953 a_41507_3295.n9 a_41507_3295.t16 214.335
R12954 a_41507_3295.t12 a_41507_3295.n9 214.335
R12955 a_41507_3295.n1 a_41507_3295.t17 214.335
R12956 a_41507_3295.t14 a_41507_3295.n1 214.335
R12957 a_41507_3295.n8 a_41507_3295.t5 198.921
R12958 a_41507_3295.n4 a_41507_3295.t10 198.043
R12959 a_41507_3295.n2 a_41507_3295.t18 160.666
R12960 a_41507_3295.n6 a_41507_3295.t7 111.663
R12961 a_41507_3295.n5 a_41507_3295.n3 97.816
R12962 a_41507_3295.n4 a_41507_3295.t4 93.989
R12963 a_41507_3295.n9 a_41507_3295.t6 80.333
R12964 a_41507_3295.n3 a_41507_3295.t15 80.333
R12965 a_41507_3295.n1 a_41507_3295.t8 80.333
R12966 a_41507_3295.n7 a_41507_3295.n5 65.07
R12967 a_41507_3295.n0 a_41507_3295.t2 28.57
R12968 a_41507_3295.n12 a_41507_3295.t3 28.565
R12969 a_41507_3295.t0 a_41507_3295.n12 28.565
R12970 a_41507_3295.n0 a_41507_3295.t1 17.638
R12971 a_41507_3295.n10 a_41507_3295.n8 16.411
R12972 a_41507_3295.n11 a_41507_3295.n10 8.712
R12973 a_41507_3295.n5 a_41507_3295.n4 6.615
R12974 a_41507_3295.n12 a_41507_3295.n11 0.69
R12975 a_41507_3295.n11 a_41507_3295.n0 0.6
R12976 a_45811_7603.n1 a_45811_7603.t7 318.922
R12977 a_45811_7603.n0 a_45811_7603.t5 273.935
R12978 a_45811_7603.n0 a_45811_7603.t6 273.935
R12979 a_45811_7603.n1 a_45811_7603.t4 269.116
R12980 a_45811_7603.n4 a_45811_7603.n3 193.227
R12981 a_45811_7603.t7 a_45811_7603.n0 179.142
R12982 a_45811_7603.n2 a_45811_7603.n1 106.999
R12983 a_45811_7603.n3 a_45811_7603.t1 28.568
R12984 a_45811_7603.n4 a_45811_7603.t0 28.565
R12985 a_45811_7603.t2 a_45811_7603.n4 28.565
R12986 a_45811_7603.n2 a_45811_7603.t3 18.149
R12987 a_45811_7603.n3 a_45811_7603.n2 3.726
R12988 a_18447_5326.n1 a_18447_5326.t4 318.922
R12989 a_18447_5326.n0 a_18447_5326.t5 273.935
R12990 a_18447_5326.n0 a_18447_5326.t7 273.935
R12991 a_18447_5326.n1 a_18447_5326.t6 269.116
R12992 a_18447_5326.n4 a_18447_5326.n3 193.227
R12993 a_18447_5326.t4 a_18447_5326.n0 179.142
R12994 a_18447_5326.n2 a_18447_5326.n1 106.999
R12995 a_18447_5326.n3 a_18447_5326.t0 28.568
R12996 a_18447_5326.t2 a_18447_5326.n4 28.565
R12997 a_18447_5326.n4 a_18447_5326.t1 28.565
R12998 a_18447_5326.n2 a_18447_5326.t3 18.149
R12999 a_18447_5326.n3 a_18447_5326.n2 3.726
R13000 a_18035_5352.t0 a_18035_5352.n0 14.282
R13001 a_18035_5352.n0 a_18035_5352.t7 14.282
R13002 a_18035_5352.n0 a_18035_5352.n9 0.999
R13003 a_18035_5352.n9 a_18035_5352.n6 0.2
R13004 a_18035_5352.n6 a_18035_5352.n8 0.575
R13005 a_18035_5352.n8 a_18035_5352.t1 16.058
R13006 a_18035_5352.n8 a_18035_5352.n7 0.999
R13007 a_18035_5352.n7 a_18035_5352.t2 14.282
R13008 a_18035_5352.n7 a_18035_5352.t3 14.282
R13009 a_18035_5352.n9 a_18035_5352.t8 16.058
R13010 a_18035_5352.n6 a_18035_5352.n4 0.227
R13011 a_18035_5352.n4 a_18035_5352.n5 1.511
R13012 a_18035_5352.n5 a_18035_5352.t5 14.282
R13013 a_18035_5352.n5 a_18035_5352.t4 14.282
R13014 a_18035_5352.n4 a_18035_5352.n1 0.669
R13015 a_18035_5352.n1 a_18035_5352.n2 0.001
R13016 a_18035_5352.n1 a_18035_5352.n3 267.767
R13017 a_18035_5352.n3 a_18035_5352.t10 14.282
R13018 a_18035_5352.n3 a_18035_5352.t11 14.282
R13019 a_18035_5352.n2 a_18035_5352.t9 14.282
R13020 a_18035_5352.n2 a_18035_5352.t6 14.282
R13021 a_13661_8966.n0 a_13661_8966.t7 14.282
R13022 a_13661_8966.t0 a_13661_8966.n0 14.282
R13023 a_13661_8966.n0 a_13661_8966.n8 90.436
R13024 a_13661_8966.n8 a_13661_8966.n5 74.302
R13025 a_13661_8966.n5 a_13661_8966.n7 50.575
R13026 a_13661_8966.n7 a_13661_8966.n6 157.665
R13027 a_13661_8966.n6 a_13661_8966.t5 8.7
R13028 a_13661_8966.n6 a_13661_8966.t1 8.7
R13029 a_13661_8966.n5 a_13661_8966.n4 90.416
R13030 a_13661_8966.n4 a_13661_8966.t6 14.282
R13031 a_13661_8966.n4 a_13661_8966.t3 14.282
R13032 a_13661_8966.n7 a_13661_8966.n3 122.746
R13033 a_13661_8966.n3 a_13661_8966.t4 14.282
R13034 a_13661_8966.n3 a_13661_8966.t2 14.282
R13035 a_13661_8966.n8 a_13661_8966.n1 1161.26
R13036 a_13661_8966.n1 a_13661_8966.t11 591.811
R13037 a_13661_8966.n1 a_13661_8966.t10 867.497
R13038 a_13661_8966.t10 a_13661_8966.n2 160.666
R13039 a_13661_8966.n2 a_13661_8966.t9 286.438
R13040 a_13661_8966.n2 a_13661_8966.t8 286.438
R13041 a_7381_20723.n2 a_7381_20723.t6 448.381
R13042 a_7381_20723.n1 a_7381_20723.t5 286.438
R13043 a_7381_20723.n1 a_7381_20723.t7 286.438
R13044 a_7381_20723.n0 a_7381_20723.t4 247.69
R13045 a_7381_20723.n4 a_7381_20723.n3 182.117
R13046 a_7381_20723.t6 a_7381_20723.n1 160.666
R13047 a_7381_20723.n3 a_7381_20723.t0 28.568
R13048 a_7381_20723.n4 a_7381_20723.t1 28.565
R13049 a_7381_20723.t2 a_7381_20723.n4 28.565
R13050 a_7381_20723.n0 a_7381_20723.t3 18.127
R13051 a_7381_20723.n2 a_7381_20723.n0 4.036
R13052 a_7381_20723.n3 a_7381_20723.n2 0.937
R13053 a_41066_22066.n2 a_41066_22066.t6 318.922
R13054 a_41066_22066.n1 a_41066_22066.t5 273.935
R13055 a_41066_22066.n1 a_41066_22066.t7 273.935
R13056 a_41066_22066.n2 a_41066_22066.t4 269.116
R13057 a_41066_22066.n4 a_41066_22066.n0 193.227
R13058 a_41066_22066.t6 a_41066_22066.n1 179.142
R13059 a_41066_22066.n3 a_41066_22066.n2 106.999
R13060 a_41066_22066.t2 a_41066_22066.n4 28.568
R13061 a_41066_22066.n0 a_41066_22066.t0 28.565
R13062 a_41066_22066.n0 a_41066_22066.t1 28.565
R13063 a_41066_22066.n3 a_41066_22066.t3 18.149
R13064 a_41066_22066.n4 a_41066_22066.n3 3.726
R13065 a_7315_8962.t0 a_7315_8962.n0 14.282
R13066 a_7315_8962.n0 a_7315_8962.t1 14.282
R13067 a_7315_8962.n0 a_7315_8962.n8 90.416
R13068 a_7315_8962.n8 a_7315_8962.n5 74.302
R13069 a_7315_8962.n8 a_7315_8962.n7 50.575
R13070 a_7315_8962.n7 a_7315_8962.n6 157.665
R13071 a_7315_8962.n6 a_7315_8962.t4 8.7
R13072 a_7315_8962.n6 a_7315_8962.t7 8.7
R13073 a_7315_8962.n5 a_7315_8962.n4 90.436
R13074 a_7315_8962.n4 a_7315_8962.t5 14.282
R13075 a_7315_8962.n4 a_7315_8962.t6 14.282
R13076 a_7315_8962.n7 a_7315_8962.n3 122.746
R13077 a_7315_8962.n3 a_7315_8962.t3 14.282
R13078 a_7315_8962.n3 a_7315_8962.t2 14.282
R13079 a_7315_8962.n5 a_7315_8962.n1 1617.45
R13080 a_7315_8962.n1 a_7315_8962.t11 591.811
R13081 a_7315_8962.n1 a_7315_8962.t8 867.497
R13082 a_7315_8962.t8 a_7315_8962.n2 160.666
R13083 a_7315_8962.n2 a_7315_8962.t10 286.438
R13084 a_7315_8962.n2 a_7315_8962.t9 286.438
R13085 a_7375_8988.t3 a_7375_8988.n0 14.282
R13086 a_7375_8988.n0 a_7375_8988.t5 14.282
R13087 a_7375_8988.n7 a_7375_8988.n8 77.784
R13088 a_7375_8988.n5 a_7375_8988.n7 77.456
R13089 a_7375_8988.n3 a_7375_8988.n5 77.456
R13090 a_7375_8988.n1 a_7375_8988.n3 75.815
R13091 a_7375_8988.n0 a_7375_8988.n1 167.433
R13092 a_7375_8988.n8 a_7375_8988.n9 167.433
R13093 a_7375_8988.n9 a_7375_8988.t10 14.282
R13094 a_7375_8988.n9 a_7375_8988.t8 14.282
R13095 a_7375_8988.n8 a_7375_8988.t9 104.259
R13096 a_7375_8988.n7 a_7375_8988.n6 89.977
R13097 a_7375_8988.n6 a_7375_8988.t2 14.282
R13098 a_7375_8988.n6 a_7375_8988.t1 14.282
R13099 a_7375_8988.n5 a_7375_8988.n4 89.977
R13100 a_7375_8988.n4 a_7375_8988.t0 14.282
R13101 a_7375_8988.n4 a_7375_8988.t6 14.282
R13102 a_7375_8988.n3 a_7375_8988.n2 89.977
R13103 a_7375_8988.n2 a_7375_8988.t11 14.282
R13104 a_7375_8988.n2 a_7375_8988.t7 14.282
R13105 a_7375_8988.n1 a_7375_8988.t4 104.259
R13106 a_6842_8258.t2 a_6842_8258.n0 14.282
R13107 a_6842_8258.n0 a_6842_8258.t7 14.282
R13108 a_6842_8258.n0 a_6842_8258.n1 258.161
R13109 a_6842_8258.n1 a_6842_8258.t3 14.283
R13110 a_6842_8258.n1 a_6842_8258.n7 4.366
R13111 a_6842_8258.n7 a_6842_8258.n5 0.852
R13112 a_6842_8258.n5 a_6842_8258.n6 258.161
R13113 a_6842_8258.n6 a_6842_8258.t6 14.282
R13114 a_6842_8258.n6 a_6842_8258.t4 14.282
R13115 a_6842_8258.n5 a_6842_8258.t5 14.283
R13116 a_6842_8258.n7 a_6842_8258.n4 97.614
R13117 a_6842_8258.n4 a_6842_8258.t8 200.029
R13118 a_6842_8258.t8 a_6842_8258.n3 206.421
R13119 a_6842_8258.n3 a_6842_8258.t11 80.333
R13120 a_6842_8258.n3 a_6842_8258.t10 206.421
R13121 a_6842_8258.n4 a_6842_8258.t9 1527.4
R13122 a_6842_8258.t9 a_6842_8258.n2 657.379
R13123 a_6842_8258.n2 a_6842_8258.t0 8.7
R13124 a_6842_8258.n2 a_6842_8258.t1 8.7
R13125 a_41697_1042.n0 a_41697_1042.t1 14.282
R13126 a_41697_1042.t0 a_41697_1042.n0 14.282
R13127 a_41697_1042.n0 a_41697_1042.n15 90.436
R13128 a_41697_1042.n11 a_41697_1042.n14 50.575
R13129 a_41697_1042.n15 a_41697_1042.n11 74.302
R13130 a_41697_1042.n14 a_41697_1042.n13 157.665
R13131 a_41697_1042.n13 a_41697_1042.t3 8.7
R13132 a_41697_1042.n13 a_41697_1042.t7 8.7
R13133 a_41697_1042.n14 a_41697_1042.n12 122.999
R13134 a_41697_1042.n12 a_41697_1042.t5 14.282
R13135 a_41697_1042.n12 a_41697_1042.t4 14.282
R13136 a_41697_1042.n11 a_41697_1042.n10 90.416
R13137 a_41697_1042.n10 a_41697_1042.t2 14.282
R13138 a_41697_1042.n10 a_41697_1042.t6 14.282
R13139 a_41697_1042.n15 a_41697_1042.n9 220.358
R13140 a_41697_1042.n9 a_41697_1042.n2 2.596
R13141 a_41697_1042.n2 a_41697_1042.t22 218.628
R13142 a_41697_1042.t22 a_41697_1042.t14 437.233
R13143 a_41697_1042.t14 a_41697_1042.n8 214.686
R13144 a_41697_1042.n8 a_41697_1042.t18 80.333
R13145 a_41697_1042.n8 a_41697_1042.t16 214.686
R13146 a_41697_1042.n2 a_41697_1042.n3 14.9
R13147 a_41697_1042.n3 a_41697_1042.n7 535.449
R13148 a_41697_1042.n7 a_41697_1042.t21 294.986
R13149 a_41697_1042.n7 a_41697_1042.t13 110.859
R13150 a_41697_1042.n3 a_41697_1042.t23 245.184
R13151 a_41697_1042.t23 a_41697_1042.n6 80.333
R13152 a_41697_1042.n6 a_41697_1042.t19 190.152
R13153 a_41697_1042.n6 a_41697_1042.t17 190.152
R13154 a_41697_1042.t17 a_41697_1042.n5 313.873
R13155 a_41697_1042.n5 a_41697_1042.t12 160.666
R13156 a_41697_1042.n5 a_41697_1042.n4 96.129
R13157 a_41697_1042.n4 a_41697_1042.t20 160.666
R13158 a_41697_1042.n4 a_41697_1042.t10 272.288
R13159 a_41697_1042.n9 a_41697_1042.t11 217.023
R13160 a_41697_1042.t11 a_41697_1042.t9 437.233
R13161 a_41697_1042.t9 a_41697_1042.n1 214.686
R13162 a_41697_1042.n1 a_41697_1042.t15 80.333
R13163 a_41697_1042.n1 a_41697_1042.t8 214.686
R13164 a_44445_4000.n4 a_44445_4000.t8 214.335
R13165 a_44445_4000.t10 a_44445_4000.n4 214.335
R13166 a_44445_4000.n5 a_44445_4000.t10 143.851
R13167 a_44445_4000.n5 a_44445_4000.t9 135.658
R13168 a_44445_4000.n4 a_44445_4000.t7 80.333
R13169 a_44445_4000.n0 a_44445_4000.t4 28.565
R13170 a_44445_4000.n0 a_44445_4000.t6 28.565
R13171 a_44445_4000.n2 a_44445_4000.t1 28.565
R13172 a_44445_4000.n2 a_44445_4000.t5 28.565
R13173 a_44445_4000.n7 a_44445_4000.t0 28.565
R13174 a_44445_4000.t2 a_44445_4000.n7 28.565
R13175 a_44445_4000.n1 a_44445_4000.t3 9.714
R13176 a_44445_4000.n1 a_44445_4000.n0 1.003
R13177 a_44445_4000.n6 a_44445_4000.n3 0.833
R13178 a_44445_4000.n3 a_44445_4000.n2 0.653
R13179 a_44445_4000.n7 a_44445_4000.n6 0.653
R13180 a_44445_4000.n3 a_44445_4000.n1 0.341
R13181 a_44445_4000.n6 a_44445_4000.n5 0.032
R13182 a_64122_11365.n2 a_64122_11365.n1 2062.97
R13183 a_64122_11365.n1 a_64122_11365.t4 989.744
R13184 a_64122_11365.n1 a_64122_11365.t7 408.806
R13185 a_64122_11365.n0 a_64122_11365.t5 287.241
R13186 a_64122_11365.n0 a_64122_11365.t6 287.241
R13187 a_64122_11365.n4 a_64122_11365.n3 192.754
R13188 a_64122_11365.t4 a_64122_11365.n0 160.666
R13189 a_64122_11365.n3 a_64122_11365.t1 28.568
R13190 a_64122_11365.t2 a_64122_11365.n4 28.565
R13191 a_64122_11365.n4 a_64122_11365.t0 28.565
R13192 a_64122_11365.n2 a_64122_11365.t3 19.164
R13193 a_64122_11365.n3 a_64122_11365.n2 1.101
R13194 a_70513_20044.n0 a_70513_20044.t8 14.282
R13195 a_70513_20044.t0 a_70513_20044.n0 14.282
R13196 a_70513_20044.n0 a_70513_20044.n9 89.977
R13197 a_70513_20044.n4 a_70513_20044.n2 77.784
R13198 a_70513_20044.n9 a_70513_20044.n4 77.456
R13199 a_70513_20044.n9 a_70513_20044.n6 77.456
R13200 a_70513_20044.n6 a_70513_20044.n7 75.815
R13201 a_70513_20044.n7 a_70513_20044.n8 167.433
R13202 a_70513_20044.n8 a_70513_20044.t11 14.282
R13203 a_70513_20044.n8 a_70513_20044.t10 14.282
R13204 a_70513_20044.n7 a_70513_20044.t9 104.259
R13205 a_70513_20044.n6 a_70513_20044.n5 89.977
R13206 a_70513_20044.n5 a_70513_20044.t1 14.282
R13207 a_70513_20044.n5 a_70513_20044.t2 14.282
R13208 a_70513_20044.n4 a_70513_20044.n3 89.977
R13209 a_70513_20044.n3 a_70513_20044.t7 14.282
R13210 a_70513_20044.n3 a_70513_20044.t6 14.282
R13211 a_70513_20044.n2 a_70513_20044.t5 104.259
R13212 a_70513_20044.n2 a_70513_20044.n1 167.433
R13213 a_70513_20044.n1 a_70513_20044.t4 14.282
R13214 a_70513_20044.n1 a_70513_20044.t3 14.282
R13215 a_1713_n2637.n1 a_1713_n2637.t4 867.497
R13216 a_1713_n2637.n1 a_1713_n2637.t6 615.911
R13217 a_1713_n2637.n0 a_1713_n2637.t7 286.438
R13218 a_1713_n2637.n0 a_1713_n2637.t5 286.438
R13219 a_1713_n2637.n4 a_1713_n2637.n3 185.55
R13220 a_1713_n2637.t4 a_1713_n2637.n0 160.666
R13221 a_1713_n2637.n3 a_1713_n2637.t2 28.568
R13222 a_1713_n2637.t0 a_1713_n2637.n4 28.565
R13223 a_1713_n2637.n4 a_1713_n2637.t1 28.565
R13224 a_1713_n2637.n2 a_1713_n2637.n1 22.215
R13225 a_1713_n2637.n2 a_1713_n2637.t3 20.397
R13226 a_1713_n2637.n3 a_1713_n2637.n2 1.838
R13227 a_1188_n2152.t0 a_1188_n2152.n0 14.283
R13228 a_1188_n2152.n0 a_1188_n2152.n7 4.366
R13229 a_1188_n2152.n7 a_1188_n2152.n5 0.852
R13230 a_1188_n2152.n5 a_1188_n2152.n6 258.161
R13231 a_1188_n2152.n6 a_1188_n2152.t3 14.282
R13232 a_1188_n2152.n6 a_1188_n2152.t5 14.282
R13233 a_1188_n2152.n5 a_1188_n2152.t4 14.283
R13234 a_1188_n2152.n7 a_1188_n2152.n4 97.614
R13235 a_1188_n2152.n4 a_1188_n2152.t11 200.029
R13236 a_1188_n2152.t11 a_1188_n2152.n3 206.421
R13237 a_1188_n2152.n3 a_1188_n2152.t10 80.333
R13238 a_1188_n2152.n3 a_1188_n2152.t9 206.421
R13239 a_1188_n2152.n4 a_1188_n2152.t8 1527.4
R13240 a_1188_n2152.t8 a_1188_n2152.n2 657.379
R13241 a_1188_n2152.n2 a_1188_n2152.t7 8.7
R13242 a_1188_n2152.n2 a_1188_n2152.t6 8.7
R13243 a_1188_n2152.n0 a_1188_n2152.n1 258.161
R13244 a_1188_n2152.n1 a_1188_n2152.t1 14.282
R13245 a_1188_n2152.n1 a_1188_n2152.t2 14.282
R13246 a_839_n2152.t0 a_839_n2152.n0 14.282
R13247 a_839_n2152.n0 a_839_n2152.t1 14.282
R13248 a_839_n2152.n0 a_839_n2152.n9 89.977
R13249 a_839_n2152.n9 a_839_n2152.n7 75.815
R13250 a_839_n2152.n9 a_839_n2152.n6 77.456
R13251 a_839_n2152.n6 a_839_n2152.n4 77.456
R13252 a_839_n2152.n4 a_839_n2152.n2 77.784
R13253 a_839_n2152.n7 a_839_n2152.n8 167.433
R13254 a_839_n2152.n8 a_839_n2152.t3 14.282
R13255 a_839_n2152.n8 a_839_n2152.t4 14.282
R13256 a_839_n2152.n7 a_839_n2152.t5 104.259
R13257 a_839_n2152.n6 a_839_n2152.n5 89.977
R13258 a_839_n2152.n5 a_839_n2152.t2 14.282
R13259 a_839_n2152.n5 a_839_n2152.t9 14.282
R13260 a_839_n2152.n4 a_839_n2152.n3 89.977
R13261 a_839_n2152.n3 a_839_n2152.t10 14.282
R13262 a_839_n2152.n3 a_839_n2152.t11 14.282
R13263 a_839_n2152.n2 a_839_n2152.t6 104.259
R13264 a_839_n2152.n2 a_839_n2152.n1 167.433
R13265 a_839_n2152.n1 a_839_n2152.t8 14.282
R13266 a_839_n2152.n1 a_839_n2152.t7 14.282
R13267 a_51054_2325.n6 a_51054_2325.n5 501.28
R13268 a_51054_2325.t13 a_51054_2325.t14 437.233
R13269 a_51054_2325.t6 a_51054_2325.t11 415.315
R13270 a_51054_2325.t10 a_51054_2325.n3 313.873
R13271 a_51054_2325.n5 a_51054_2325.t19 294.986
R13272 a_51054_2325.n2 a_51054_2325.t16 272.288
R13273 a_51054_2325.n6 a_51054_2325.t18 236.01
R13274 a_51054_2325.n9 a_51054_2325.t13 216.627
R13275 a_51054_2325.n7 a_51054_2325.t6 216.111
R13276 a_51054_2325.n8 a_51054_2325.t7 214.686
R13277 a_51054_2325.t14 a_51054_2325.n8 214.686
R13278 a_51054_2325.n1 a_51054_2325.t4 214.335
R13279 a_51054_2325.t11 a_51054_2325.n1 214.335
R13280 a_51054_2325.n4 a_51054_2325.t10 190.152
R13281 a_51054_2325.n4 a_51054_2325.t15 190.152
R13282 a_51054_2325.n2 a_51054_2325.t12 160.666
R13283 a_51054_2325.n3 a_51054_2325.t5 160.666
R13284 a_51054_2325.n7 a_51054_2325.n6 148.428
R13285 a_51054_2325.n5 a_51054_2325.t9 110.859
R13286 a_51054_2325.n3 a_51054_2325.n2 96.129
R13287 a_51054_2325.n8 a_51054_2325.t17 80.333
R13288 a_51054_2325.n1 a_51054_2325.t8 80.333
R13289 a_51054_2325.t18 a_51054_2325.n4 80.333
R13290 a_51054_2325.n0 a_51054_2325.t2 28.57
R13291 a_51054_2325.n11 a_51054_2325.t3 28.565
R13292 a_51054_2325.t0 a_51054_2325.n11 28.565
R13293 a_51054_2325.n0 a_51054_2325.t1 17.638
R13294 a_51054_2325.n10 a_51054_2325.n9 6.64
R13295 a_51054_2325.n9 a_51054_2325.n7 2.923
R13296 a_51054_2325.n11 a_51054_2325.n10 0.69
R13297 a_51054_2325.n10 a_51054_2325.n0 0.6
R13298 a_51109_747.n0 a_51109_747.t7 214.335
R13299 a_51109_747.t9 a_51109_747.n0 214.335
R13300 a_51109_747.n1 a_51109_747.t9 143.851
R13301 a_51109_747.n1 a_51109_747.t10 135.658
R13302 a_51109_747.n0 a_51109_747.t8 80.333
R13303 a_51109_747.n2 a_51109_747.t5 28.565
R13304 a_51109_747.n2 a_51109_747.t4 28.565
R13305 a_51109_747.n4 a_51109_747.t3 28.565
R13306 a_51109_747.n4 a_51109_747.t6 28.565
R13307 a_51109_747.t1 a_51109_747.n7 28.565
R13308 a_51109_747.n7 a_51109_747.t2 28.565
R13309 a_51109_747.n6 a_51109_747.t0 9.714
R13310 a_51109_747.n7 a_51109_747.n6 1.003
R13311 a_51109_747.n5 a_51109_747.n3 0.833
R13312 a_51109_747.n3 a_51109_747.n2 0.653
R13313 a_51109_747.n5 a_51109_747.n4 0.653
R13314 a_51109_747.n6 a_51109_747.n5 0.341
R13315 a_51109_747.n3 a_51109_747.n1 0.032
R13316 a_56850_21339.n1 a_56850_21339.t7 318.922
R13317 a_56850_21339.n0 a_56850_21339.t5 274.739
R13318 a_56850_21339.n0 a_56850_21339.t6 274.739
R13319 a_56850_21339.n1 a_56850_21339.t4 269.116
R13320 a_56850_21339.t7 a_56850_21339.n0 179.946
R13321 a_56850_21339.n2 a_56850_21339.n1 105.178
R13322 a_56850_21339.t2 a_56850_21339.n4 29.444
R13323 a_56850_21339.n3 a_56850_21339.t0 28.565
R13324 a_56850_21339.n3 a_56850_21339.t1 28.565
R13325 a_56850_21339.n2 a_56850_21339.t3 18.145
R13326 a_56850_21339.n4 a_56850_21339.n2 2.878
R13327 a_56850_21339.n4 a_56850_21339.n3 0.764
R13328 a_35012_10049.n2 a_35012_10049.t9 214.335
R13329 a_35012_10049.t7 a_35012_10049.n2 214.335
R13330 a_35012_10049.n3 a_35012_10049.t7 143.851
R13331 a_35012_10049.n3 a_35012_10049.t10 135.658
R13332 a_35012_10049.n2 a_35012_10049.t8 80.333
R13333 a_35012_10049.n4 a_35012_10049.t2 28.565
R13334 a_35012_10049.n4 a_35012_10049.t1 28.565
R13335 a_35012_10049.n0 a_35012_10049.t5 28.565
R13336 a_35012_10049.n0 a_35012_10049.t4 28.565
R13337 a_35012_10049.t0 a_35012_10049.n7 28.565
R13338 a_35012_10049.n7 a_35012_10049.t3 28.565
R13339 a_35012_10049.n1 a_35012_10049.t6 9.714
R13340 a_35012_10049.n1 a_35012_10049.n0 1.003
R13341 a_35012_10049.n6 a_35012_10049.n5 0.833
R13342 a_35012_10049.n5 a_35012_10049.n4 0.653
R13343 a_35012_10049.n7 a_35012_10049.n6 0.653
R13344 a_35012_10049.n6 a_35012_10049.n1 0.341
R13345 a_35012_10049.n5 a_35012_10049.n3 0.032
R13346 a_35602_9612.n4 a_35602_9612.n3 535.449
R13347 a_35602_9612.t16 a_35602_9612.t15 437.233
R13348 a_35602_9612.t18 a_35602_9612.t8 437.233
R13349 a_35602_9612.t11 a_35602_9612.n1 313.873
R13350 a_35602_9612.n3 a_35602_9612.t12 294.986
R13351 a_35602_9612.n0 a_35602_9612.t14 272.288
R13352 a_35602_9612.n4 a_35602_9612.t4 245.184
R13353 a_35602_9612.n6 a_35602_9612.t18 218.628
R13354 a_35602_9612.n8 a_35602_9612.t16 217.024
R13355 a_35602_9612.n7 a_35602_9612.t9 214.686
R13356 a_35602_9612.t15 a_35602_9612.n7 214.686
R13357 a_35602_9612.n5 a_35602_9612.t19 214.686
R13358 a_35602_9612.t8 a_35602_9612.n5 214.686
R13359 a_35602_9612.n11 a_35602_9612.n10 192.754
R13360 a_35602_9612.n2 a_35602_9612.t11 190.152
R13361 a_35602_9612.n2 a_35602_9612.t13 190.152
R13362 a_35602_9612.n0 a_35602_9612.t10 160.666
R13363 a_35602_9612.n1 a_35602_9612.t6 160.666
R13364 a_35602_9612.n3 a_35602_9612.t17 110.859
R13365 a_35602_9612.n1 a_35602_9612.n0 96.129
R13366 a_35602_9612.n7 a_35602_9612.t5 80.333
R13367 a_35602_9612.t4 a_35602_9612.n2 80.333
R13368 a_35602_9612.n5 a_35602_9612.t7 80.333
R13369 a_35602_9612.n10 a_35602_9612.t0 28.568
R13370 a_35602_9612.n11 a_35602_9612.t1 28.565
R13371 a_35602_9612.t2 a_35602_9612.n11 28.565
R13372 a_35602_9612.n9 a_35602_9612.t3 18.726
R13373 a_35602_9612.n6 a_35602_9612.n4 14.9
R13374 a_35602_9612.n8 a_35602_9612.n6 2.599
R13375 a_35602_9612.n9 a_35602_9612.n8 2.514
R13376 a_35602_9612.n10 a_35602_9612.n9 1.123
R13377 B[1].t9 B[1].t12 800.875
R13378 B[1].n9 B[1].n1 654.791
R13379 B[1].n7 B[1].n6 618.566
R13380 B[1].n14 B[1].n10 592.056
R13381 B[1].t8 B[1].t14 415.315
R13382 B[1].t20 B[1].n4 313.873
R13383 B[1].t10 B[1].n12 313.069
R13384 B[1].n10 B[1].t13 294.986
R13385 B[1].n0 B[1].t17 284.688
R13386 B[1].n6 B[1].t2 273.077
R13387 B[1].n3 B[1].t19 272.288
R13388 B[1].n11 B[1].t11 271.484
R13389 B[1].n8 B[1].t8 217.528
R13390 B[1].n2 B[1].t5 214.335
R13391 B[1].t14 B[1].n2 214.335
R13392 B[1].n7 B[1].t3 204.679
R13393 B[1].n14 B[1].t23 204.672
R13394 B[1].n1 B[1].t9 192.799
R13395 B[1].n13 B[1].t10 190.955
R13396 B[1].n13 B[1].t15 190.955
R13397 B[1].n5 B[1].t22 190.152
R13398 B[1].n5 B[1].t20 190.152
R13399 B[1].n3 B[1].t16 160.666
R13400 B[1].n4 B[1].t21 160.666
R13401 B[1].n0 B[1].t0 160.666
R13402 B[1].n12 B[1].t4 160.666
R13403 B[1].n11 B[1].t1 160.666
R13404 B[1].n6 B[1].t6 137.369
R13405 B[1].n10 B[1].t18 110.859
R13406 B[1].n4 B[1].n3 96.129
R13407 B[1].n12 B[1].n11 96.129
R13408 B[1].n1 B[1].n0 91.889
R13409 B[1].n2 B[1].t7 80.333
R13410 B[1].t3 B[1].n5 80.333
R13411 B[1].t23 B[1].n13 80.333
R13412 B[1].n15 B[1].n14 57.39
R13413 B[1].n8 B[1].n7 49.906
R13414 B[1] B[1].n15 49.362
R13415 B[1].n15 B[1].n9 11.093
R13416 B[1].n9 B[1].n8 0.414
R13417 a_11640_16408.n0 a_11640_16408.t5 14.282
R13418 a_11640_16408.n0 a_11640_16408.t1 14.282
R13419 a_11640_16408.n1 a_11640_16408.t2 14.282
R13420 a_11640_16408.n1 a_11640_16408.t0 14.282
R13421 a_11640_16408.n3 a_11640_16408.t4 14.282
R13422 a_11640_16408.t3 a_11640_16408.n3 14.282
R13423 a_11640_16408.n3 a_11640_16408.n2 2.538
R13424 a_11640_16408.n2 a_11640_16408.n1 2.375
R13425 a_11640_16408.n2 a_11640_16408.n0 0.001
R13426 a_46176_16428.n0 a_46176_16428.n12 90.436
R13427 a_46176_16428.t0 a_46176_16428.n0 14.282
R13428 a_46176_16428.n0 a_46176_16428.t1 14.282
R13429 a_46176_16428.n12 a_46176_16428.n9 74.302
R13430 a_46176_16428.n9 a_46176_16428.n11 50.575
R13431 a_46176_16428.n11 a_46176_16428.n10 157.665
R13432 a_46176_16428.n10 a_46176_16428.t7 8.7
R13433 a_46176_16428.n10 a_46176_16428.t6 8.7
R13434 a_46176_16428.n9 a_46176_16428.n8 90.416
R13435 a_46176_16428.n8 a_46176_16428.t2 14.282
R13436 a_46176_16428.n8 a_46176_16428.t3 14.282
R13437 a_46176_16428.n11 a_46176_16428.n7 122.746
R13438 a_46176_16428.n7 a_46176_16428.t4 14.282
R13439 a_46176_16428.n7 a_46176_16428.t5 14.282
R13440 a_46176_16428.n12 a_46176_16428.n1 342.688
R13441 a_46176_16428.n1 a_46176_16428.n6 126.566
R13442 a_46176_16428.n6 a_46176_16428.t9 294.653
R13443 a_46176_16428.n6 a_46176_16428.t14 111.663
R13444 a_46176_16428.n1 a_46176_16428.n5 552.333
R13445 a_46176_16428.n5 a_46176_16428.n4 6.615
R13446 a_46176_16428.n4 a_46176_16428.t8 93.989
R13447 a_46176_16428.n4 a_46176_16428.t10 198.043
R13448 a_46176_16428.n5 a_46176_16428.n3 97.816
R13449 a_46176_16428.n3 a_46176_16428.t15 80.333
R13450 a_46176_16428.n3 a_46176_16428.t13 394.151
R13451 a_46176_16428.t13 a_46176_16428.n2 269.523
R13452 a_46176_16428.n2 a_46176_16428.t12 160.666
R13453 a_46176_16428.n2 a_46176_16428.t11 269.523
R13454 a_46233_15735.n1 a_46233_15735.t7 318.922
R13455 a_46233_15735.n0 a_46233_15735.t6 273.935
R13456 a_46233_15735.n0 a_46233_15735.t4 273.935
R13457 a_46233_15735.n1 a_46233_15735.t5 269.116
R13458 a_46233_15735.n4 a_46233_15735.n3 193.227
R13459 a_46233_15735.t7 a_46233_15735.n0 179.142
R13460 a_46233_15735.n2 a_46233_15735.n1 106.999
R13461 a_46233_15735.n3 a_46233_15735.t1 28.568
R13462 a_46233_15735.t2 a_46233_15735.n4 28.565
R13463 a_46233_15735.n4 a_46233_15735.t0 28.565
R13464 a_46233_15735.n2 a_46233_15735.t3 18.149
R13465 a_46233_15735.n3 a_46233_15735.n2 3.726
R13466 a_59929_3874.t5 a_59929_3874.n2 404.877
R13467 a_59929_3874.n1 a_59929_3874.t6 210.902
R13468 a_59929_3874.n3 a_59929_3874.t5 136.943
R13469 a_59929_3874.n2 a_59929_3874.n1 107.801
R13470 a_59929_3874.n1 a_59929_3874.t7 80.333
R13471 a_59929_3874.n2 a_59929_3874.t8 80.333
R13472 a_59929_3874.n0 a_59929_3874.t2 17.4
R13473 a_59929_3874.n0 a_59929_3874.t0 17.4
R13474 a_59929_3874.n4 a_59929_3874.t3 15.032
R13475 a_59929_3874.n5 a_59929_3874.t4 14.282
R13476 a_59929_3874.t1 a_59929_3874.n5 14.282
R13477 a_59929_3874.n5 a_59929_3874.n4 1.65
R13478 a_59929_3874.n3 a_59929_3874.n0 0.672
R13479 a_59929_3874.n4 a_59929_3874.n3 0.665
R13480 a_60193_3291.t6 a_60193_3291.t7 800.071
R13481 a_60193_3291.n3 a_60193_3291.n2 672.951
R13482 a_60193_3291.n1 a_60193_3291.t5 285.109
R13483 a_60193_3291.n2 a_60193_3291.t6 193.602
R13484 a_60193_3291.n1 a_60193_3291.t4 160.666
R13485 a_60193_3291.n2 a_60193_3291.n1 91.507
R13486 a_60193_3291.n0 a_60193_3291.t0 28.57
R13487 a_60193_3291.t2 a_60193_3291.n4 28.565
R13488 a_60193_3291.n4 a_60193_3291.t1 28.565
R13489 a_60193_3291.n0 a_60193_3291.t3 17.638
R13490 a_60193_3291.n4 a_60193_3291.n3 0.69
R13491 a_60193_3291.n3 a_60193_3291.n0 0.6
R13492 a_62660_24205.t6 a_62660_24205.n3 404.877
R13493 a_62660_24205.n2 a_62660_24205.t5 210.902
R13494 a_62660_24205.n4 a_62660_24205.t6 136.943
R13495 a_62660_24205.n3 a_62660_24205.n2 107.801
R13496 a_62660_24205.n2 a_62660_24205.t8 80.333
R13497 a_62660_24205.n3 a_62660_24205.t7 80.333
R13498 a_62660_24205.n1 a_62660_24205.t0 17.4
R13499 a_62660_24205.n1 a_62660_24205.t4 17.4
R13500 a_62660_24205.t1 a_62660_24205.n5 15.032
R13501 a_62660_24205.n0 a_62660_24205.t3 14.282
R13502 a_62660_24205.n0 a_62660_24205.t2 14.282
R13503 a_62660_24205.n5 a_62660_24205.n0 1.65
R13504 a_62660_24205.n4 a_62660_24205.n1 0.672
R13505 a_62660_24205.n5 a_62660_24205.n4 0.665
R13506 a_58326_16165.n6 a_58326_16165.n5 501.28
R13507 a_58326_16165.t8 a_58326_16165.t12 437.233
R13508 a_58326_16165.t15 a_58326_16165.t7 415.315
R13509 a_58326_16165.t10 a_58326_16165.n3 313.873
R13510 a_58326_16165.n5 a_58326_16165.t17 294.986
R13511 a_58326_16165.n2 a_58326_16165.t11 272.288
R13512 a_58326_16165.n6 a_58326_16165.t9 236.009
R13513 a_58326_16165.n9 a_58326_16165.t8 216.627
R13514 a_58326_16165.n7 a_58326_16165.t15 216.111
R13515 a_58326_16165.n8 a_58326_16165.t16 214.686
R13516 a_58326_16165.t12 a_58326_16165.n8 214.686
R13517 a_58326_16165.n1 a_58326_16165.t18 214.335
R13518 a_58326_16165.t7 a_58326_16165.n1 214.335
R13519 a_58326_16165.n4 a_58326_16165.t19 190.152
R13520 a_58326_16165.n4 a_58326_16165.t10 190.152
R13521 a_58326_16165.n2 a_58326_16165.t5 160.666
R13522 a_58326_16165.n3 a_58326_16165.t4 160.666
R13523 a_58326_16165.n7 a_58326_16165.n6 148.428
R13524 a_58326_16165.n5 a_58326_16165.t14 110.859
R13525 a_58326_16165.n3 a_58326_16165.n2 96.129
R13526 a_58326_16165.n8 a_58326_16165.t13 80.333
R13527 a_58326_16165.n1 a_58326_16165.t6 80.333
R13528 a_58326_16165.t9 a_58326_16165.n4 80.333
R13529 a_58326_16165.n0 a_58326_16165.t1 28.57
R13530 a_58326_16165.t2 a_58326_16165.n11 28.565
R13531 a_58326_16165.n11 a_58326_16165.t0 28.565
R13532 a_58326_16165.n0 a_58326_16165.t3 17.638
R13533 a_58326_16165.n10 a_58326_16165.n9 10.943
R13534 a_58326_16165.n9 a_58326_16165.n7 2.923
R13535 a_58326_16165.n11 a_58326_16165.n10 0.69
R13536 a_58326_16165.n10 a_58326_16165.n0 0.6
R13537 a_779_n2178.n2 a_779_n2178.t6 990.34
R13538 a_779_n2178.n2 a_779_n2178.t4 408.211
R13539 a_779_n2178.n1 a_779_n2178.t5 286.438
R13540 a_779_n2178.n1 a_779_n2178.t7 286.438
R13541 a_779_n2178.n4 a_779_n2178.n0 185.55
R13542 a_779_n2178.t6 a_779_n2178.n1 160.666
R13543 a_779_n2178.t1 a_779_n2178.n4 28.568
R13544 a_779_n2178.n0 a_779_n2178.t3 28.565
R13545 a_779_n2178.n0 a_779_n2178.t2 28.565
R13546 a_779_n2178.n3 a_779_n2178.t0 21.583
R13547 a_779_n2178.n3 a_779_n2178.n2 18.186
R13548 a_779_n2178.n4 a_779_n2178.n3 1.537
R13549 a_1424_n3485.t0 a_1424_n3485.t1 17.4
R13550 a_45939_15761.n0 a_45939_15761.n8 90.436
R13551 a_45939_15761.t0 a_45939_15761.n0 14.282
R13552 a_45939_15761.n0 a_45939_15761.t1 14.282
R13553 a_45939_15761.n8 a_45939_15761.n5 74.302
R13554 a_45939_15761.n5 a_45939_15761.n7 50.575
R13555 a_45939_15761.n7 a_45939_15761.n6 157.665
R13556 a_45939_15761.n6 a_45939_15761.t3 8.7
R13557 a_45939_15761.n6 a_45939_15761.t7 8.7
R13558 a_45939_15761.n5 a_45939_15761.n4 90.416
R13559 a_45939_15761.n4 a_45939_15761.t2 14.282
R13560 a_45939_15761.n4 a_45939_15761.t5 14.282
R13561 a_45939_15761.n7 a_45939_15761.n3 122.746
R13562 a_45939_15761.n3 a_45939_15761.t4 14.282
R13563 a_45939_15761.n3 a_45939_15761.t6 14.282
R13564 a_45939_15761.n8 a_45939_15761.n1 294.955
R13565 a_45939_15761.t8 a_45939_15761.n2 160.666
R13566 a_45939_15761.n1 a_45939_15761.t8 867.393
R13567 a_45939_15761.n2 a_45939_15761.t11 287.241
R13568 a_45939_15761.n2 a_45939_15761.t9 287.241
R13569 a_45939_15761.n1 a_45939_15761.t10 545.094
R13570 a_45821_15761.t0 a_45821_15761.n7 16.058
R13571 a_45821_15761.n7 a_45821_15761.n5 0.2
R13572 a_45821_15761.n5 a_45821_15761.n9 0.575
R13573 a_45821_15761.n9 a_45821_15761.t11 16.058
R13574 a_45821_15761.n9 a_45821_15761.n8 0.999
R13575 a_45821_15761.n8 a_45821_15761.t10 14.282
R13576 a_45821_15761.n8 a_45821_15761.t9 14.282
R13577 a_45821_15761.n7 a_45821_15761.n6 0.999
R13578 a_45821_15761.n6 a_45821_15761.t1 14.282
R13579 a_45821_15761.n6 a_45821_15761.t2 14.282
R13580 a_45821_15761.n5 a_45821_15761.n3 0.227
R13581 a_45821_15761.n3 a_45821_15761.n4 1.511
R13582 a_45821_15761.n4 a_45821_15761.t7 14.282
R13583 a_45821_15761.n4 a_45821_15761.t6 14.282
R13584 a_45821_15761.n3 a_45821_15761.n0 0.669
R13585 a_45821_15761.n0 a_45821_15761.n1 0.001
R13586 a_45821_15761.n0 a_45821_15761.n2 267.767
R13587 a_45821_15761.n2 a_45821_15761.t4 14.282
R13588 a_45821_15761.n2 a_45821_15761.t3 14.282
R13589 a_45821_15761.n1 a_45821_15761.t5 14.282
R13590 a_45821_15761.n1 a_45821_15761.t8 14.282
R13591 a_6832_13724.t0 a_6832_13724.n0 14.283
R13592 a_6832_13724.n0 a_6832_13724.n5 0.852
R13593 a_6832_13724.n5 a_6832_13724.n6 4.366
R13594 a_6832_13724.n6 a_6832_13724.n7 258.161
R13595 a_6832_13724.n7 a_6832_13724.t5 14.282
R13596 a_6832_13724.n7 a_6832_13724.t6 14.282
R13597 a_6832_13724.n6 a_6832_13724.t4 14.283
R13598 a_6832_13724.n5 a_6832_13724.n4 97.614
R13599 a_6832_13724.n4 a_6832_13724.t9 200.029
R13600 a_6832_13724.t9 a_6832_13724.n3 206.421
R13601 a_6832_13724.n3 a_6832_13724.t10 80.333
R13602 a_6832_13724.n3 a_6832_13724.t11 206.421
R13603 a_6832_13724.n4 a_6832_13724.t8 1527.4
R13604 a_6832_13724.t8 a_6832_13724.n2 657.379
R13605 a_6832_13724.n2 a_6832_13724.t7 8.7
R13606 a_6832_13724.n2 a_6832_13724.t3 8.7
R13607 a_6832_13724.n0 a_6832_13724.n1 258.161
R13608 a_6832_13724.n1 a_6832_13724.t1 14.282
R13609 a_6832_13724.n1 a_6832_13724.t2 14.282
R13610 a_6774_14454.n2 a_6774_14454.t5 867.497
R13611 a_6774_14454.n2 a_6774_14454.t7 591.811
R13612 a_6774_14454.n1 a_6774_14454.t4 286.438
R13613 a_6774_14454.n1 a_6774_14454.t6 286.438
R13614 a_6774_14454.n4 a_6774_14454.n0 185.55
R13615 a_6774_14454.t5 a_6774_14454.n1 160.666
R13616 a_6774_14454.t2 a_6774_14454.n4 28.568
R13617 a_6774_14454.n0 a_6774_14454.t0 28.565
R13618 a_6774_14454.n0 a_6774_14454.t1 28.565
R13619 a_6774_14454.n3 a_6774_14454.n2 25.434
R13620 a_6774_14454.n3 a_6774_14454.t3 22.077
R13621 a_6774_14454.n4 a_6774_14454.n3 1.628
R13622 B[4].n15 B[4].t26 1361.95
R13623 B[4].n14 B[4].t38 1211.76
R13624 B[4].t29 B[4].t3 802.481
R13625 B[4].n9 B[4].n8 650.496
R13626 B[4].n4 B[4].n3 618.566
R13627 B[4].n20 B[4].n16 592.056
R13628 B[4].n15 B[4].t4 561.041
R13629 B[4].t26 B[4].t17 437.233
R13630 B[4].t4 B[4].t35 437.233
R13631 B[4].t20 B[4].t33 415.315
R13632 B[4].t38 B[4].t22 415.315
R13633 B[4].t37 B[4].t34 415.315
R13634 B[4].t13 B[4].n1 313.873
R13635 B[4].t27 B[4].n18 313.069
R13636 B[4].n16 B[4].t18 294.986
R13637 B[4].n7 B[4].t7 284.688
R13638 B[4].n3 B[4].t23 273.077
R13639 B[4].n0 B[4].t11 272.288
R13640 B[4].n17 B[4].t14 271.484
R13641 B[4].n14 B[4].t37 219.359
R13642 B[4].n6 B[4].t20 217.534
R13643 B[4].n10 B[4].t5 214.686
R13644 B[4].t17 B[4].n10 214.686
R13645 B[4].n11 B[4].t28 214.686
R13646 B[4].t35 B[4].n11 214.686
R13647 B[4].n5 B[4].t16 214.335
R13648 B[4].t33 B[4].n5 214.335
R13649 B[4].n12 B[4].t25 214.335
R13650 B[4].t22 B[4].n12 214.335
R13651 B[4].n13 B[4].t39 214.335
R13652 B[4].t34 B[4].n13 214.335
R13653 B[4].n4 B[4].t24 204.679
R13654 B[4].n20 B[4].t12 204.672
R13655 B[4].n8 B[4].t29 192.799
R13656 B[4].n19 B[4].t27 190.955
R13657 B[4].n19 B[4].t8 190.955
R13658 B[4].n2 B[4].t9 190.152
R13659 B[4].n2 B[4].t13 190.152
R13660 B[4].n0 B[4].t1 160.666
R13661 B[4].n1 B[4].t0 160.666
R13662 B[4].n7 B[4].t15 160.666
R13663 B[4].n18 B[4].t21 160.666
R13664 B[4].n17 B[4].t2 160.666
R13665 B[4].n3 B[4].t19 137.369
R13666 B[4].n16 B[4].t6 110.859
R13667 B[4].n1 B[4].n0 96.129
R13668 B[4].n18 B[4].n17 96.129
R13669 B[4].n8 B[4].n7 91.889
R13670 B[4].n5 B[4].t31 80.333
R13671 B[4].t24 B[4].n2 80.333
R13672 B[4].n10 B[4].t30 80.333
R13673 B[4].n11 B[4].t32 80.333
R13674 B[4].n12 B[4].t10 80.333
R13675 B[4].n13 B[4].t36 80.333
R13676 B[4].t12 B[4].n19 80.333
R13677 B[4].n21 B[4].n20 52.607
R13678 B[4].n6 B[4].n4 50.196
R13679 B[4] B[4].n22 48.804
R13680 B[4].n22 B[4].n21 18.66
R13681 B[4].n22 B[4].n9 15.841
R13682 B[4].n9 B[4].n6 5.535
R13683 B[4].n21 B[4].n15 1.607
R13684 B[4].n15 B[4].n14 1.018
R13685 a_15966_5352.n0 a_15966_5352.t4 14.282
R13686 a_15966_5352.t3 a_15966_5352.n0 14.282
R13687 a_15966_5352.n0 a_15966_5352.n9 0.999
R13688 a_15966_5352.n9 a_15966_5352.n6 0.2
R13689 a_15966_5352.n6 a_15966_5352.n8 0.575
R13690 a_15966_5352.n8 a_15966_5352.t11 16.058
R13691 a_15966_5352.n8 a_15966_5352.n7 0.999
R13692 a_15966_5352.n7 a_15966_5352.t9 14.282
R13693 a_15966_5352.n7 a_15966_5352.t8 14.282
R13694 a_15966_5352.n9 a_15966_5352.t10 16.058
R13695 a_15966_5352.n6 a_15966_5352.n4 0.227
R13696 a_15966_5352.n4 a_15966_5352.n5 1.511
R13697 a_15966_5352.n5 a_15966_5352.t5 14.282
R13698 a_15966_5352.n5 a_15966_5352.t6 14.282
R13699 a_15966_5352.n4 a_15966_5352.n1 0.669
R13700 a_15966_5352.n1 a_15966_5352.n2 0.001
R13701 a_15966_5352.n1 a_15966_5352.n3 267.767
R13702 a_15966_5352.n3 a_15966_5352.t2 14.282
R13703 a_15966_5352.n3 a_15966_5352.t1 14.282
R13704 a_15966_5352.n2 a_15966_5352.t0 14.282
R13705 a_15966_5352.n2 a_15966_5352.t7 14.282
R13706 a_70513_4278.t0 a_70513_4278.n9 104.259
R13707 a_70513_4278.n9 a_70513_4278.n2 77.784
R13708 a_70513_4278.n2 a_70513_4278.n4 77.456
R13709 a_70513_4278.n4 a_70513_4278.n6 77.456
R13710 a_70513_4278.n6 a_70513_4278.n7 75.815
R13711 a_70513_4278.n7 a_70513_4278.n8 167.433
R13712 a_70513_4278.n8 a_70513_4278.t4 14.282
R13713 a_70513_4278.n8 a_70513_4278.t5 14.282
R13714 a_70513_4278.n7 a_70513_4278.t3 104.259
R13715 a_70513_4278.n6 a_70513_4278.n5 89.977
R13716 a_70513_4278.n5 a_70513_4278.t6 14.282
R13717 a_70513_4278.n5 a_70513_4278.t7 14.282
R13718 a_70513_4278.n4 a_70513_4278.n3 89.977
R13719 a_70513_4278.n3 a_70513_4278.t9 14.282
R13720 a_70513_4278.n3 a_70513_4278.t8 14.282
R13721 a_70513_4278.n2 a_70513_4278.n1 89.977
R13722 a_70513_4278.n1 a_70513_4278.t10 14.282
R13723 a_70513_4278.n1 a_70513_4278.t11 14.282
R13724 a_70513_4278.n9 a_70513_4278.n0 167.433
R13725 a_70513_4278.n0 a_70513_4278.t1 14.282
R13726 a_70513_4278.n0 a_70513_4278.t2 14.282
R13727 A[0].n15 A[0].n3 4143.01
R13728 A[0].n1 A[0].t4 867.497
R13729 A[0].n1 A[0].t27 591.811
R13730 A[0].t22 A[0].t10 576.841
R13731 A[0].n21 A[0].n20 535.449
R13732 A[0].n26 A[0].n16 497.047
R13733 A[0].t20 A[0].t30 437.233
R13734 A[0].t11 A[0].t3 437.233
R13735 A[0].t8 A[0].t34 437.233
R13736 A[0].n13 A[0].n12 412.11
R13737 A[0].n10 A[0].t6 394.151
R13738 A[0].t32 A[0].n18 313.873
R13739 A[0].n20 A[0].t25 294.986
R13740 A[0].n12 A[0].t23 294.653
R13741 A[0].n0 A[0].t2 286.438
R13742 A[0].n0 A[0].t5 286.438
R13743 A[0].n4 A[0].t14 284.688
R13744 A[0].n17 A[0].t29 272.288
R13745 A[0].n9 A[0].t38 269.523
R13746 A[0].t6 A[0].n9 269.523
R13747 A[0].n21 A[0].t35 245.184
R13748 A[0].n13 A[0].n11 224.13
R13749 A[0].n23 A[0].t8 218.628
R13750 A[0].n7 A[0].t20 217.073
R13751 A[0].n25 A[0].t11 217.024
R13752 A[0].n6 A[0].t9 214.686
R13753 A[0].t30 A[0].n6 214.686
R13754 A[0].n24 A[0].t39 214.686
R13755 A[0].t3 A[0].n24 214.686
R13756 A[0].n22 A[0].t28 214.686
R13757 A[0].t34 A[0].n22 214.686
R13758 A[0].n8 A[0].t24 198.043
R13759 A[0].n19 A[0].t32 190.152
R13760 A[0].n19 A[0].t37 190.152
R13761 A[0].n7 A[0].n5 185.868
R13762 A[0].n2 A[0].t13 185.301
R13763 A[0].n2 A[0].t1 185.301
R13764 A[0].t4 A[0].n0 160.666
R13765 A[0].n9 A[0].t15 160.666
R13766 A[0].n4 A[0].t17 160.666
R13767 A[0].n5 A[0].t22 160.666
R13768 A[0].n17 A[0].t26 160.666
R13769 A[0].n18 A[0].t7 160.666
R13770 A[0].n3 A[0].t16 140.583
R13771 A[0].n14 A[0].n13 138.41
R13772 A[0].n5 A[0].n4 115.593
R13773 A[0].n12 A[0].t18 111.663
R13774 A[0].n20 A[0].t36 110.859
R13775 A[0].n2 A[0].t21 107.646
R13776 A[0].n11 A[0].n10 97.816
R13777 A[0].n18 A[0].n17 96.129
R13778 A[0].n8 A[0].t12 93.989
R13779 A[0].n10 A[0].t19 80.333
R13780 A[0].n6 A[0].t33 80.333
R13781 A[0].n24 A[0].t0 80.333
R13782 A[0].t35 A[0].n19 80.333
R13783 A[0].n22 A[0].t31 80.333
R13784 A[0].n3 A[0].n2 61.856
R13785 A[0] A[0].n26 45.108
R13786 A[0].n16 A[0].n1 22.594
R13787 A[0].n16 A[0].n15 16.366
R13788 A[0].n23 A[0].n21 14.9
R13789 A[0].n26 A[0].n25 9.838
R13790 A[0].n14 A[0].n7 6.82
R13791 A[0].n11 A[0].n8 6.615
R13792 A[0].n25 A[0].n23 2.599
R13793 A[0].n15 A[0].n14 0.001
R13794 a_38506_7695.t7 a_38506_7695.t5 574.43
R13795 a_38506_7695.n0 a_38506_7695.t4 285.109
R13796 a_38506_7695.n2 a_38506_7695.n1 211.136
R13797 a_38506_7695.n4 a_38506_7695.n3 192.754
R13798 a_38506_7695.n0 a_38506_7695.t6 160.666
R13799 a_38506_7695.n1 a_38506_7695.t7 160.666
R13800 a_38506_7695.n1 a_38506_7695.n0 114.829
R13801 a_38506_7695.n3 a_38506_7695.t0 28.568
R13802 a_38506_7695.t2 a_38506_7695.n4 28.565
R13803 a_38506_7695.n4 a_38506_7695.t1 28.565
R13804 a_38506_7695.n2 a_38506_7695.t3 19.084
R13805 a_38506_7695.n3 a_38506_7695.n2 1.051
R13806 a_30645_5900.t0 a_30645_5900.n0 14.282
R13807 a_30645_5900.n0 a_30645_5900.t2 14.282
R13808 a_30645_5900.n0 a_30645_5900.n16 90.436
R13809 a_30645_5900.n16 a_30645_5900.n2 74.302
R13810 a_30645_5900.n2 a_30645_5900.n4 50.575
R13811 a_30645_5900.n4 a_30645_5900.n5 110.084
R13812 a_30645_5900.n16 a_30645_5900.n6 214.569
R13813 a_30645_5900.n6 a_30645_5900.n8 16.411
R13814 a_30645_5900.n8 a_30645_5900.t17 198.921
R13815 a_30645_5900.t17 a_30645_5900.t15 415.315
R13816 a_30645_5900.t15 a_30645_5900.n15 214.335
R13817 a_30645_5900.n15 a_30645_5900.t16 80.333
R13818 a_30645_5900.n15 a_30645_5900.t18 214.335
R13819 a_30645_5900.n8 a_30645_5900.n14 861.987
R13820 a_30645_5900.n14 a_30645_5900.n9 560.726
R13821 a_30645_5900.n14 a_30645_5900.n13 65.07
R13822 a_30645_5900.n13 a_30645_5900.n12 6.615
R13823 a_30645_5900.n12 a_30645_5900.t12 93.989
R13824 a_30645_5900.n13 a_30645_5900.n11 97.816
R13825 a_30645_5900.n11 a_30645_5900.t13 80.333
R13826 a_30645_5900.n11 a_30645_5900.t20 394.151
R13827 a_30645_5900.t20 a_30645_5900.n10 269.523
R13828 a_30645_5900.n10 a_30645_5900.t21 160.666
R13829 a_30645_5900.n10 a_30645_5900.t22 269.523
R13830 a_30645_5900.n12 a_30645_5900.t10 198.043
R13831 a_30645_5900.n9 a_30645_5900.t23 294.653
R13832 a_30645_5900.n9 a_30645_5900.t14 111.663
R13833 a_30645_5900.n6 a_30645_5900.t19 217.716
R13834 a_30645_5900.t19 a_30645_5900.t8 415.315
R13835 a_30645_5900.t8 a_30645_5900.n7 214.335
R13836 a_30645_5900.n7 a_30645_5900.t9 80.333
R13837 a_30645_5900.n7 a_30645_5900.t11 214.335
R13838 a_30645_5900.n5 a_30645_5900.t7 14.282
R13839 a_30645_5900.n5 a_30645_5900.t4 14.282
R13840 a_30645_5900.n4 a_30645_5900.n3 157.665
R13841 a_30645_5900.n3 a_30645_5900.t1 8.7
R13842 a_30645_5900.n3 a_30645_5900.t5 8.7
R13843 a_30645_5900.n2 a_30645_5900.n1 90.416
R13844 a_30645_5900.n1 a_30645_5900.t3 14.282
R13845 a_30645_5900.n1 a_30645_5900.t6 14.282
R13846 a_59311_24329.n2 a_59311_24329.t10 214.335
R13847 a_59311_24329.t8 a_59311_24329.n2 214.335
R13848 a_59311_24329.n3 a_59311_24329.t8 143.851
R13849 a_59311_24329.n3 a_59311_24329.t7 135.658
R13850 a_59311_24329.n2 a_59311_24329.t9 80.333
R13851 a_59311_24329.n4 a_59311_24329.t0 28.565
R13852 a_59311_24329.n4 a_59311_24329.t1 28.565
R13853 a_59311_24329.n0 a_59311_24329.t5 28.565
R13854 a_59311_24329.n0 a_59311_24329.t6 28.565
R13855 a_59311_24329.t2 a_59311_24329.n7 28.565
R13856 a_59311_24329.n7 a_59311_24329.t4 28.565
R13857 a_59311_24329.n1 a_59311_24329.t3 9.714
R13858 a_59311_24329.n1 a_59311_24329.n0 1.003
R13859 a_59311_24329.n6 a_59311_24329.n5 0.833
R13860 a_59311_24329.n5 a_59311_24329.n4 0.653
R13861 a_59311_24329.n7 a_59311_24329.n6 0.653
R13862 a_59311_24329.n6 a_59311_24329.n1 0.341
R13863 a_59311_24329.n5 a_59311_24329.n3 0.032
R13864 a_51815_16459.n1 a_51815_16459.t5 318.922
R13865 a_51815_16459.n0 a_51815_16459.t4 274.739
R13866 a_51815_16459.n0 a_51815_16459.t6 274.739
R13867 a_51815_16459.n1 a_51815_16459.t7 269.116
R13868 a_51815_16459.t5 a_51815_16459.n0 179.946
R13869 a_51815_16459.n2 a_51815_16459.n1 105.178
R13870 a_51815_16459.t2 a_51815_16459.n4 29.444
R13871 a_51815_16459.n3 a_51815_16459.t0 28.565
R13872 a_51815_16459.n3 a_51815_16459.t1 28.565
R13873 a_51815_16459.n2 a_51815_16459.t3 18.145
R13874 a_51815_16459.n4 a_51815_16459.n2 2.878
R13875 a_51815_16459.n4 a_51815_16459.n3 0.764
R13876 a_52355_15766.n0 a_52355_15766.t4 14.282
R13877 a_52355_15766.t3 a_52355_15766.n0 14.282
R13878 a_52355_15766.n0 a_52355_15766.n9 0.999
R13879 a_52355_15766.n9 a_52355_15766.n6 0.2
R13880 a_52355_15766.n6 a_52355_15766.n8 0.575
R13881 a_52355_15766.n8 a_52355_15766.t11 16.058
R13882 a_52355_15766.n8 a_52355_15766.n7 0.999
R13883 a_52355_15766.n7 a_52355_15766.t9 14.282
R13884 a_52355_15766.n7 a_52355_15766.t10 14.282
R13885 a_52355_15766.n9 a_52355_15766.t5 16.058
R13886 a_52355_15766.n6 a_52355_15766.n4 0.227
R13887 a_52355_15766.n4 a_52355_15766.n5 1.511
R13888 a_52355_15766.n5 a_52355_15766.t2 14.282
R13889 a_52355_15766.n5 a_52355_15766.t1 14.282
R13890 a_52355_15766.n4 a_52355_15766.n1 0.669
R13891 a_52355_15766.n1 a_52355_15766.n2 0.001
R13892 a_52355_15766.n1 a_52355_15766.n3 267.767
R13893 a_52355_15766.n3 a_52355_15766.t8 14.282
R13894 a_52355_15766.n3 a_52355_15766.t7 14.282
R13895 a_52355_15766.n2 a_52355_15766.t6 14.282
R13896 a_52355_15766.n2 a_52355_15766.t0 14.282
R13897 a_52473_15766.n0 a_52473_15766.t2 14.282
R13898 a_52473_15766.t5 a_52473_15766.n0 14.282
R13899 a_52473_15766.n0 a_52473_15766.n8 90.416
R13900 a_52473_15766.n8 a_52473_15766.n5 74.302
R13901 a_52473_15766.n8 a_52473_15766.n7 50.575
R13902 a_52473_15766.n7 a_52473_15766.n6 157.665
R13903 a_52473_15766.n6 a_52473_15766.t1 8.7
R13904 a_52473_15766.n6 a_52473_15766.t0 8.7
R13905 a_52473_15766.n5 a_52473_15766.n4 90.436
R13906 a_52473_15766.n4 a_52473_15766.t4 14.282
R13907 a_52473_15766.n4 a_52473_15766.t3 14.282
R13908 a_52473_15766.n7 a_52473_15766.n3 122.746
R13909 a_52473_15766.n3 a_52473_15766.t6 14.282
R13910 a_52473_15766.n3 a_52473_15766.t7 14.282
R13911 a_52473_15766.n5 a_52473_15766.n1 275.913
R13912 a_52473_15766.t10 a_52473_15766.n2 160.666
R13913 a_52473_15766.n1 a_52473_15766.t10 867.393
R13914 a_52473_15766.n2 a_52473_15766.t9 287.241
R13915 a_52473_15766.n2 a_52473_15766.t8 287.241
R13916 a_52473_15766.n1 a_52473_15766.t11 545.094
R13917 a_42177_23622.t7 a_42177_23622.t6 800.071
R13918 a_42177_23622.n3 a_42177_23622.n2 672.951
R13919 a_42177_23622.n1 a_42177_23622.t5 285.109
R13920 a_42177_23622.n2 a_42177_23622.t7 193.602
R13921 a_42177_23622.n1 a_42177_23622.t4 160.666
R13922 a_42177_23622.n2 a_42177_23622.n1 91.507
R13923 a_42177_23622.t0 a_42177_23622.n4 28.57
R13924 a_42177_23622.n0 a_42177_23622.t3 28.565
R13925 a_42177_23622.n0 a_42177_23622.t2 28.565
R13926 a_42177_23622.n4 a_42177_23622.t1 17.638
R13927 a_42177_23622.n3 a_42177_23622.n0 0.69
R13928 a_42177_23622.n4 a_42177_23622.n3 0.6
R13929 a_43173_24209.n0 a_43173_24209.t3 14.282
R13930 a_43173_24209.n0 a_43173_24209.t2 14.282
R13931 a_43173_24209.n1 a_43173_24209.t4 14.282
R13932 a_43173_24209.n1 a_43173_24209.t5 14.282
R13933 a_43173_24209.n3 a_43173_24209.t1 14.282
R13934 a_43173_24209.t0 a_43173_24209.n3 14.282
R13935 a_43173_24209.n3 a_43173_24209.n2 2.546
R13936 a_43173_24209.n2 a_43173_24209.n1 2.367
R13937 a_43173_24209.n2 a_43173_24209.n0 0.001
R13938 a_54113_22058.n2 a_54113_22058.t4 318.922
R13939 a_54113_22058.n1 a_54113_22058.t7 273.935
R13940 a_54113_22058.n1 a_54113_22058.t5 273.935
R13941 a_54113_22058.n2 a_54113_22058.t6 269.116
R13942 a_54113_22058.n4 a_54113_22058.n0 193.227
R13943 a_54113_22058.t4 a_54113_22058.n1 179.142
R13944 a_54113_22058.n3 a_54113_22058.n2 106.999
R13945 a_54113_22058.t0 a_54113_22058.n4 28.568
R13946 a_54113_22058.n0 a_54113_22058.t2 28.565
R13947 a_54113_22058.n0 a_54113_22058.t1 28.565
R13948 a_54113_22058.n3 a_54113_22058.t3 18.149
R13949 a_54113_22058.n4 a_54113_22058.n3 3.726
R13950 a_54658_21365.n0 a_54658_21365.n12 122.999
R13951 a_54658_21365.t2 a_54658_21365.n0 14.282
R13952 a_54658_21365.n0 a_54658_21365.t4 14.282
R13953 a_54658_21365.n12 a_54658_21365.n10 50.575
R13954 a_54658_21365.n10 a_54658_21365.n8 74.302
R13955 a_54658_21365.n12 a_54658_21365.n11 157.665
R13956 a_54658_21365.n11 a_54658_21365.t1 8.7
R13957 a_54658_21365.n11 a_54658_21365.t0 8.7
R13958 a_54658_21365.n10 a_54658_21365.n9 90.416
R13959 a_54658_21365.n9 a_54658_21365.t3 14.282
R13960 a_54658_21365.n9 a_54658_21365.t5 14.282
R13961 a_54658_21365.n8 a_54658_21365.n7 90.436
R13962 a_54658_21365.n7 a_54658_21365.t7 14.282
R13963 a_54658_21365.n7 a_54658_21365.t6 14.282
R13964 a_54658_21365.n8 a_54658_21365.n1 342.688
R13965 a_54658_21365.n1 a_54658_21365.n6 126.566
R13966 a_54658_21365.n6 a_54658_21365.t10 294.653
R13967 a_54658_21365.n6 a_54658_21365.t9 111.663
R13968 a_54658_21365.n1 a_54658_21365.n5 552.333
R13969 a_54658_21365.n5 a_54658_21365.n4 6.615
R13970 a_54658_21365.n4 a_54658_21365.t15 93.989
R13971 a_54658_21365.n5 a_54658_21365.n3 97.816
R13972 a_54658_21365.n3 a_54658_21365.t8 80.333
R13973 a_54658_21365.n3 a_54658_21365.t11 394.151
R13974 a_54658_21365.t11 a_54658_21365.n2 269.523
R13975 a_54658_21365.n2 a_54658_21365.t12 160.666
R13976 a_54658_21365.n2 a_54658_21365.t13 269.523
R13977 a_54658_21365.n4 a_54658_21365.t14 198.043
R13978 a_54540_21365.n0 a_54540_21365.n9 1.511
R13979 a_54540_21365.t0 a_54540_21365.n0 14.282
R13980 a_54540_21365.n0 a_54540_21365.t1 14.282
R13981 a_54540_21365.n9 a_54540_21365.n5 0.227
R13982 a_54540_21365.n9 a_54540_21365.n6 0.669
R13983 a_54540_21365.n6 a_54540_21365.n7 0.001
R13984 a_54540_21365.n6 a_54540_21365.n8 267.767
R13985 a_54540_21365.n8 a_54540_21365.t7 14.282
R13986 a_54540_21365.n8 a_54540_21365.t6 14.282
R13987 a_54540_21365.n7 a_54540_21365.t2 14.282
R13988 a_54540_21365.n7 a_54540_21365.t8 14.282
R13989 a_54540_21365.n5 a_54540_21365.n2 0.575
R13990 a_54540_21365.n5 a_54540_21365.n4 0.2
R13991 a_54540_21365.n4 a_54540_21365.t10 16.058
R13992 a_54540_21365.n4 a_54540_21365.n3 0.999
R13993 a_54540_21365.n3 a_54540_21365.t9 14.282
R13994 a_54540_21365.n3 a_54540_21365.t11 14.282
R13995 a_54540_21365.n2 a_54540_21365.n1 0.999
R13996 a_54540_21365.n1 a_54540_21365.t5 14.282
R13997 a_54540_21365.n1 a_54540_21365.t4 14.282
R13998 a_54540_21365.n2 a_54540_21365.t3 16.058
R13999 a_6827_15753.t5 a_6827_15753.n2 405.372
R14000 a_6827_15753.n1 a_6827_15753.t7 207.38
R14001 a_6827_15753.n3 a_6827_15753.t5 138.556
R14002 a_6827_15753.n2 a_6827_15753.n1 112.003
R14003 a_6827_15753.n1 a_6827_15753.t8 80.333
R14004 a_6827_15753.n2 a_6827_15753.t6 80.333
R14005 a_6827_15753.n0 a_6827_15753.t1 17.4
R14006 a_6827_15753.n0 a_6827_15753.t0 17.4
R14007 a_6827_15753.n4 a_6827_15753.t4 15.029
R14008 a_6827_15753.n5 a_6827_15753.t3 14.282
R14009 a_6827_15753.t2 a_6827_15753.n5 14.282
R14010 a_6827_15753.n5 a_6827_15753.n4 1.647
R14011 a_6827_15753.n3 a_6827_15753.n0 0.664
R14012 a_6827_15753.n4 a_6827_15753.n3 0.614
R14013 a_6887_15819.n2 a_6887_15819.t4 990.34
R14014 a_6887_15819.n3 a_6887_15819.n2 903.227
R14015 a_6887_15819.n2 a_6887_15819.t6 408.211
R14016 a_6887_15819.n1 a_6887_15819.t7 286.438
R14017 a_6887_15819.n1 a_6887_15819.t5 286.438
R14018 a_6887_15819.t4 a_6887_15819.n1 160.666
R14019 a_6887_15819.n4 a_6887_15819.n3 97.311
R14020 a_6887_15819.n3 a_6887_15819.n0 94.754
R14021 a_6887_15819.t2 a_6887_15819.n4 28.568
R14022 a_6887_15819.n0 a_6887_15819.t0 28.565
R14023 a_6887_15819.n0 a_6887_15819.t1 28.565
R14024 a_6887_15819.n4 a_6887_15819.t3 17.64
R14025 a_8021_8115.n3 a_8021_8115.t4 448.381
R14026 a_8021_8115.n2 a_8021_8115.t5 286.438
R14027 a_8021_8115.n2 a_8021_8115.t6 286.438
R14028 a_8021_8115.n1 a_8021_8115.t7 247.69
R14029 a_8021_8115.n4 a_8021_8115.n0 182.117
R14030 a_8021_8115.t4 a_8021_8115.n2 160.666
R14031 a_8021_8115.t2 a_8021_8115.n4 28.568
R14032 a_8021_8115.n0 a_8021_8115.t1 28.565
R14033 a_8021_8115.n0 a_8021_8115.t0 28.565
R14034 a_8021_8115.n1 a_8021_8115.t3 18.127
R14035 a_8021_8115.n3 a_8021_8115.n1 4.036
R14036 a_8021_8115.n4 a_8021_8115.n3 0.937
R14037 a_6774_11720.n2 a_6774_11720.t6 990.34
R14038 a_6774_11720.n2 a_6774_11720.t7 408.211
R14039 a_6774_11720.n1 a_6774_11720.t4 286.438
R14040 a_6774_11720.n1 a_6774_11720.t5 286.438
R14041 a_6774_11720.n4 a_6774_11720.n0 185.55
R14042 a_6774_11720.t6 a_6774_11720.n1 160.666
R14043 a_6774_11720.n3 a_6774_11720.n2 31.762
R14044 a_6774_11720.t1 a_6774_11720.n4 28.568
R14045 a_6774_11720.n0 a_6774_11720.t3 28.565
R14046 a_6774_11720.n0 a_6774_11720.t2 28.565
R14047 a_6774_11720.n3 a_6774_11720.t0 21.376
R14048 a_6774_11720.n4 a_6774_11720.n3 1.637
R14049 a_7083_1744.n0 a_7083_1744.t8 14.282
R14050 a_7083_1744.t6 a_7083_1744.n0 14.282
R14051 a_7083_1744.n7 a_7083_1744.n8 75.815
R14052 a_7083_1744.n5 a_7083_1744.n7 77.456
R14053 a_7083_1744.n3 a_7083_1744.n5 77.456
R14054 a_7083_1744.n1 a_7083_1744.n3 77.784
R14055 a_7083_1744.n0 a_7083_1744.n1 167.433
R14056 a_7083_1744.n8 a_7083_1744.n9 167.433
R14057 a_7083_1744.n9 a_7083_1744.t2 14.282
R14058 a_7083_1744.n9 a_7083_1744.t0 14.282
R14059 a_7083_1744.n8 a_7083_1744.t1 104.259
R14060 a_7083_1744.n7 a_7083_1744.n6 89.977
R14061 a_7083_1744.n6 a_7083_1744.t10 14.282
R14062 a_7083_1744.n6 a_7083_1744.t11 14.282
R14063 a_7083_1744.n5 a_7083_1744.n4 89.977
R14064 a_7083_1744.n4 a_7083_1744.t9 14.282
R14065 a_7083_1744.n4 a_7083_1744.t5 14.282
R14066 a_7083_1744.n3 a_7083_1744.n2 89.977
R14067 a_7083_1744.n2 a_7083_1744.t4 14.282
R14068 a_7083_1744.n2 a_7083_1744.t3 14.282
R14069 a_7083_1744.n1 a_7083_1744.t7 104.259
R14070 a_51059_8126.n17 a_51059_8126.n16 538.835
R14071 a_51059_8126.n9 a_51059_8126.n8 501.28
R14072 a_51059_8126.t18 a_51059_8126.t19 437.233
R14073 a_51059_8126.t14 a_51059_8126.t11 415.315
R14074 a_51059_8126.t4 a_51059_8126.n6 313.873
R14075 a_51059_8126.n8 a_51059_8126.t15 294.986
R14076 a_51059_8126.n5 a_51059_8126.t7 272.288
R14077 a_51059_8126.n9 a_51059_8126.t13 236.01
R14078 a_51059_8126.n12 a_51059_8126.t18 216.627
R14079 a_51059_8126.n10 a_51059_8126.t14 216.111
R14080 a_51059_8126.n11 a_51059_8126.t12 214.686
R14081 a_51059_8126.t19 a_51059_8126.n11 214.686
R14082 a_51059_8126.n4 a_51059_8126.t17 214.335
R14083 a_51059_8126.t11 a_51059_8126.n4 214.335
R14084 a_51059_8126.n19 a_51059_8126.n18 192.754
R14085 a_51059_8126.n7 a_51059_8126.t4 190.152
R14086 a_51059_8126.n7 a_51059_8126.t6 190.152
R14087 a_51059_8126.n5 a_51059_8126.t16 160.666
R14088 a_51059_8126.n6 a_51059_8126.t10 160.666
R14089 a_51059_8126.n10 a_51059_8126.n9 148.428
R14090 a_51059_8126.n8 a_51059_8126.t5 110.859
R14091 a_51059_8126.n6 a_51059_8126.n5 96.129
R14092 a_51059_8126.n11 a_51059_8126.t9 80.333
R14093 a_51059_8126.n4 a_51059_8126.t8 80.333
R14094 a_51059_8126.t13 a_51059_8126.n7 80.333
R14095 a_51059_8126.n18 a_51059_8126.t2 28.568
R14096 a_51059_8126.n19 a_51059_8126.t3 28.565
R14097 a_51059_8126.t0 a_51059_8126.n19 28.565
R14098 a_51059_8126.n17 a_51059_8126.t1 18.514
R14099 a_51059_8126.n16 a_51059_8126.n15 4.161
R14100 a_51059_8126.n12 a_51059_8126.n10 2.923
R14101 a_51059_8126.n18 a_51059_8126.n17 1.177
R14102 a_51059_8126.n13 a_51059_8126.n12 0.707
R14103 a_51059_8126.n15 a_51059_8126.n14 0.078
R14104 a_51059_8126.n1 a_51059_8126.n0 0.045
R14105 a_51059_8126.n3 a_51059_8126.n2 0.006
R14106 a_51059_8126.n15 a_51059_8126.n1 0.003
R14107 a_51059_8126.n13 a_51059_8126.n3 0.002
R14108 a_51059_8126.n15 a_51059_8126.n13 0.001
R14109 a_55202_6816.n1 a_55202_6816.t7 318.922
R14110 a_55202_6816.n0 a_55202_6816.t4 274.739
R14111 a_55202_6816.n0 a_55202_6816.t5 274.739
R14112 a_55202_6816.n1 a_55202_6816.t6 269.116
R14113 a_55202_6816.t7 a_55202_6816.n0 179.946
R14114 a_55202_6816.n2 a_55202_6816.n1 105.178
R14115 a_55202_6816.n3 a_55202_6816.t1 29.444
R14116 a_55202_6816.n4 a_55202_6816.t0 28.565
R14117 a_55202_6816.t2 a_55202_6816.n4 28.565
R14118 a_55202_6816.n2 a_55202_6816.t3 18.145
R14119 a_55202_6816.n3 a_55202_6816.n2 2.878
R14120 a_55202_6816.n4 a_55202_6816.n3 0.764
R14121 a_11505_15751.t8 a_11505_15751.n2 404.877
R14122 a_11505_15751.n1 a_11505_15751.t5 210.902
R14123 a_11505_15751.n3 a_11505_15751.t8 136.949
R14124 a_11505_15751.n2 a_11505_15751.n1 107.801
R14125 a_11505_15751.n1 a_11505_15751.t6 80.333
R14126 a_11505_15751.n2 a_11505_15751.t7 80.333
R14127 a_11505_15751.n0 a_11505_15751.t4 17.4
R14128 a_11505_15751.n0 a_11505_15751.t0 17.4
R14129 a_11505_15751.n4 a_11505_15751.t2 15.036
R14130 a_11505_15751.t1 a_11505_15751.n5 14.282
R14131 a_11505_15751.n5 a_11505_15751.t3 14.282
R14132 a_11505_15751.n5 a_11505_15751.n4 1.654
R14133 a_11505_15751.n3 a_11505_15751.n0 0.657
R14134 a_11505_15751.n4 a_11505_15751.n3 0.614
R14135 a_11565_15824.n3 a_11565_15824.n1 2881.06
R14136 a_11565_15824.n1 a_11565_15824.t6 990.34
R14137 a_11565_15824.n1 a_11565_15824.t5 408.211
R14138 a_11565_15824.n0 a_11565_15824.t4 286.438
R14139 a_11565_15824.n0 a_11565_15824.t7 286.438
R14140 a_11565_15824.t6 a_11565_15824.n0 160.666
R14141 a_11565_15824.n4 a_11565_15824.n3 112.943
R14142 a_11565_15824.n3 a_11565_15824.n2 112.94
R14143 a_11565_15824.n2 a_11565_15824.t0 28.568
R14144 a_11565_15824.n4 a_11565_15824.t1 28.565
R14145 a_11565_15824.t2 a_11565_15824.n4 28.565
R14146 a_11565_15824.n2 a_11565_15824.t3 17.64
R14147 a_40101_6796.n1 a_40101_6796.t5 318.922
R14148 a_40101_6796.n0 a_40101_6796.t6 274.739
R14149 a_40101_6796.n0 a_40101_6796.t7 274.739
R14150 a_40101_6796.n1 a_40101_6796.t4 269.116
R14151 a_40101_6796.t5 a_40101_6796.n0 179.946
R14152 a_40101_6796.n2 a_40101_6796.n1 107.263
R14153 a_40101_6796.n3 a_40101_6796.t0 29.444
R14154 a_40101_6796.t2 a_40101_6796.n4 28.565
R14155 a_40101_6796.n4 a_40101_6796.t1 28.565
R14156 a_40101_6796.n2 a_40101_6796.t3 18.145
R14157 a_40101_6796.n3 a_40101_6796.n2 2.878
R14158 a_40101_6796.n4 a_40101_6796.n3 0.764
R14159 a_70455_n1231.n3 a_70455_n1231.t5 448.381
R14160 a_70455_n1231.n2 a_70455_n1231.t4 287.241
R14161 a_70455_n1231.n2 a_70455_n1231.t6 287.241
R14162 a_70455_n1231.n1 a_70455_n1231.t7 247.733
R14163 a_70455_n1231.n4 a_70455_n1231.n0 182.117
R14164 a_70455_n1231.t5 a_70455_n1231.n2 160.666
R14165 a_70455_n1231.t2 a_70455_n1231.n4 28.568
R14166 a_70455_n1231.n0 a_70455_n1231.t0 28.565
R14167 a_70455_n1231.n0 a_70455_n1231.t1 28.565
R14168 a_70455_n1231.n1 a_70455_n1231.t3 18.127
R14169 a_70455_n1231.n3 a_70455_n1231.n1 4.036
R14170 a_70455_n1231.n4 a_70455_n1231.n3 0.937
R14171 a_70455_1913.n2 a_70455_1913.t6 448.381
R14172 a_70455_1913.n1 a_70455_1913.t7 287.241
R14173 a_70455_1913.n1 a_70455_1913.t5 287.241
R14174 a_70455_1913.n0 a_70455_1913.t4 247.733
R14175 a_70455_1913.n4 a_70455_1913.n3 182.117
R14176 a_70455_1913.t6 a_70455_1913.n1 160.666
R14177 a_70455_1913.n3 a_70455_1913.t0 28.568
R14178 a_70455_1913.n4 a_70455_1913.t1 28.565
R14179 a_70455_1913.t2 a_70455_1913.n4 28.565
R14180 a_70455_1913.n0 a_70455_1913.t3 18.127
R14181 a_70455_1913.n2 a_70455_1913.n0 4.036
R14182 a_70455_1913.n3 a_70455_1913.n2 0.937
R14183 a_48815_11511.n5 a_48815_11511.n4 535.449
R14184 a_48815_11511.t17 a_48815_11511.t13 437.233
R14185 a_48815_11511.t14 a_48815_11511.t10 437.233
R14186 a_48815_11511.t11 a_48815_11511.n2 313.873
R14187 a_48815_11511.n4 a_48815_11511.t8 294.986
R14188 a_48815_11511.n1 a_48815_11511.t16 272.288
R14189 a_48815_11511.n5 a_48815_11511.t5 245.184
R14190 a_48815_11511.n7 a_48815_11511.t14 218.628
R14191 a_48815_11511.n9 a_48815_11511.t17 217.024
R14192 a_48815_11511.n8 a_48815_11511.t7 214.686
R14193 a_48815_11511.t13 a_48815_11511.n8 214.686
R14194 a_48815_11511.n6 a_48815_11511.t4 214.686
R14195 a_48815_11511.t10 a_48815_11511.n6 214.686
R14196 a_48815_11511.n11 a_48815_11511.n0 192.754
R14197 a_48815_11511.n3 a_48815_11511.t11 190.152
R14198 a_48815_11511.n3 a_48815_11511.t6 190.152
R14199 a_48815_11511.n1 a_48815_11511.t9 160.666
R14200 a_48815_11511.n2 a_48815_11511.t19 160.666
R14201 a_48815_11511.n4 a_48815_11511.t12 110.859
R14202 a_48815_11511.n2 a_48815_11511.n1 96.129
R14203 a_48815_11511.n8 a_48815_11511.t18 80.333
R14204 a_48815_11511.t5 a_48815_11511.n3 80.333
R14205 a_48815_11511.n6 a_48815_11511.t15 80.333
R14206 a_48815_11511.t0 a_48815_11511.n11 28.568
R14207 a_48815_11511.n0 a_48815_11511.t3 28.565
R14208 a_48815_11511.n0 a_48815_11511.t2 28.565
R14209 a_48815_11511.n10 a_48815_11511.t1 20.07
R14210 a_48815_11511.n7 a_48815_11511.n5 14.9
R14211 a_48815_11511.n10 a_48815_11511.n9 3.139
R14212 a_48815_11511.n9 a_48815_11511.n7 2.599
R14213 a_48815_11511.n11 a_48815_11511.n10 1.101
R14214 a_51114_6548.n4 a_51114_6548.t9 214.335
R14215 a_51114_6548.t8 a_51114_6548.n4 214.335
R14216 a_51114_6548.n5 a_51114_6548.t8 143.851
R14217 a_51114_6548.n5 a_51114_6548.t10 135.658
R14218 a_51114_6548.n4 a_51114_6548.t7 80.333
R14219 a_51114_6548.n0 a_51114_6548.t4 28.565
R14220 a_51114_6548.n0 a_51114_6548.t6 28.565
R14221 a_51114_6548.n2 a_51114_6548.t1 28.565
R14222 a_51114_6548.n2 a_51114_6548.t5 28.565
R14223 a_51114_6548.n7 a_51114_6548.t0 28.565
R14224 a_51114_6548.t2 a_51114_6548.n7 28.565
R14225 a_51114_6548.n1 a_51114_6548.t3 9.714
R14226 a_51114_6548.n1 a_51114_6548.n0 1.003
R14227 a_51114_6548.n6 a_51114_6548.n3 0.833
R14228 a_51114_6548.n3 a_51114_6548.n2 0.653
R14229 a_51114_6548.n7 a_51114_6548.n6 0.653
R14230 a_51114_6548.n3 a_51114_6548.n1 0.341
R14231 a_51114_6548.n6 a_51114_6548.n5 0.032
R14232 a_63598_4278.n0 a_63598_4278.t9 214.335
R14233 a_63598_4278.t7 a_63598_4278.n0 214.335
R14234 a_63598_4278.n1 a_63598_4278.t7 143.851
R14235 a_63598_4278.n1 a_63598_4278.t8 135.658
R14236 a_63598_4278.n0 a_63598_4278.t10 80.333
R14237 a_63598_4278.n2 a_63598_4278.t4 28.565
R14238 a_63598_4278.n2 a_63598_4278.t6 28.565
R14239 a_63598_4278.n4 a_63598_4278.t5 28.565
R14240 a_63598_4278.n4 a_63598_4278.t2 28.565
R14241 a_63598_4278.n7 a_63598_4278.t1 28.565
R14242 a_63598_4278.t3 a_63598_4278.n7 28.565
R14243 a_63598_4278.n6 a_63598_4278.t0 9.714
R14244 a_63598_4278.n7 a_63598_4278.n6 1.003
R14245 a_63598_4278.n5 a_63598_4278.n3 0.833
R14246 a_63598_4278.n3 a_63598_4278.n2 0.653
R14247 a_63598_4278.n5 a_63598_4278.n4 0.653
R14248 a_63598_4278.n6 a_63598_4278.n5 0.341
R14249 a_63598_4278.n3 a_63598_4278.n1 0.032
R14250 a_61533_6910.n0 a_61533_6910.n8 122.999
R14251 a_61533_6910.n0 a_61533_6910.t3 14.282
R14252 a_61533_6910.t1 a_61533_6910.n0 14.282
R14253 a_61533_6910.n8 a_61533_6910.n6 50.575
R14254 a_61533_6910.n6 a_61533_6910.n4 74.302
R14255 a_61533_6910.n8 a_61533_6910.n7 157.665
R14256 a_61533_6910.n7 a_61533_6910.t4 8.7
R14257 a_61533_6910.n7 a_61533_6910.t0 8.7
R14258 a_61533_6910.n6 a_61533_6910.n5 90.416
R14259 a_61533_6910.n5 a_61533_6910.t2 14.282
R14260 a_61533_6910.n5 a_61533_6910.t6 14.282
R14261 a_61533_6910.n4 a_61533_6910.n3 90.436
R14262 a_61533_6910.n3 a_61533_6910.t7 14.282
R14263 a_61533_6910.n3 a_61533_6910.t5 14.282
R14264 a_61533_6910.n4 a_61533_6910.n1 670.272
R14265 a_61533_6910.n1 a_61533_6910.t9 408.806
R14266 a_61533_6910.t11 a_61533_6910.n2 160.666
R14267 a_61533_6910.n1 a_61533_6910.t11 989.744
R14268 a_61533_6910.n2 a_61533_6910.t10 287.241
R14269 a_61533_6910.n2 a_61533_6910.t8 287.241
R14270 a_61769_6178.t0 a_61769_6178.t1 17.4
R14271 A[5].n26 A[5].t33 3756.03
R14272 A[5].n12 A[5].n5 2643.13
R14273 A[5].n36 A[5].n26 2196.31
R14274 A[5].n15 A[5].t40 990.34
R14275 A[5].n17 A[5].t54 867.497
R14276 A[5].n17 A[5].t11 591.811
R14277 A[5].t51 A[5].t2 575.234
R14278 A[5].n31 A[5].n30 535.449
R14279 A[5].n37 A[5].n19 445.43
R14280 A[5].t43 A[5].t56 437.233
R14281 A[5].t17 A[5].t18 437.233
R14282 A[5].t33 A[5].t19 437.233
R14283 A[5].t25 A[5].t24 437.233
R14284 A[5].t0 A[5].t27 437.233
R14285 A[5].t13 A[5].t14 415.315
R14286 A[5].t58 A[5].t31 415.315
R14287 A[5].n11 A[5].n10 412.11
R14288 A[5].n15 A[5].t23 408.211
R14289 A[5].n8 A[5].t52 394.151
R14290 A[5].t30 A[5].n28 313.873
R14291 A[5].n30 A[5].t29 294.986
R14292 A[5].n10 A[5].t49 294.653
R14293 A[5].n14 A[5].t39 286.438
R14294 A[5].n14 A[5].t41 286.438
R14295 A[5].n16 A[5].t53 286.438
R14296 A[5].n16 A[5].t16 286.438
R14297 A[5].n1 A[5].t48 285.543
R14298 A[5].n27 A[5].t7 272.288
R14299 A[5].n7 A[5].t46 269.523
R14300 A[5].t52 A[5].n7 269.523
R14301 A[5].n25 A[5].t58 256.298
R14302 A[5].n31 A[5].t20 245.184
R14303 A[5].n11 A[5].n9 224.13
R14304 A[5].n3 A[5].t43 222.157
R14305 A[5].n23 A[5].t17 219.994
R14306 A[5].n33 A[5].t0 218.627
R14307 A[5].n23 A[5].t13 217.552
R14308 A[5].n35 A[5].t25 217.023
R14309 A[5].n0 A[5].t12 214.686
R14310 A[5].t56 A[5].n0 214.686
R14311 A[5].n21 A[5].t35 214.686
R14312 A[5].t18 A[5].n21 214.686
R14313 A[5].n20 A[5].t55 214.686
R14314 A[5].t19 A[5].n20 214.686
R14315 A[5].n34 A[5].t1 214.686
R14316 A[5].t24 A[5].n34 214.686
R14317 A[5].n32 A[5].t45 214.686
R14318 A[5].t27 A[5].n32 214.686
R14319 A[5].n22 A[5].t22 214.335
R14320 A[5].t14 A[5].n22 214.335
R14321 A[5].n24 A[5].t36 214.335
R14322 A[5].t31 A[5].n24 214.335
R14323 A[5].n6 A[5].t28 198.043
R14324 A[5].n29 A[5].t3 190.152
R14325 A[5].n29 A[5].t30 190.152
R14326 A[5].n4 A[5].t15 185.301
R14327 A[5].n4 A[5].t10 185.301
R14328 A[5].n3 A[5].n2 181.495
R14329 A[5].t40 A[5].n14 160.666
R14330 A[5].t54 A[5].n16 160.666
R14331 A[5].n1 A[5].t50 160.666
R14332 A[5].n2 A[5].t51 160.666
R14333 A[5].n7 A[5].t26 160.666
R14334 A[5].n27 A[5].t6 160.666
R14335 A[5].n28 A[5].t5 160.666
R14336 A[5].n12 A[5].n11 142.204
R14337 A[5].n5 A[5].t21 140.583
R14338 A[5] A[5].n37 138.722
R14339 A[5].n2 A[5].n1 114.089
R14340 A[5].n10 A[5].t4 111.663
R14341 A[5].n30 A[5].t8 110.859
R14342 A[5].n4 A[5].t32 107.646
R14343 A[5].n9 A[5].n8 97.816
R14344 A[5].n28 A[5].n27 96.129
R14345 A[5].n6 A[5].t47 93.989
R14346 A[5].n0 A[5].t59 80.333
R14347 A[5].n8 A[5].t9 80.333
R14348 A[5].n22 A[5].t42 80.333
R14349 A[5].n21 A[5].t37 80.333
R14350 A[5].n24 A[5].t34 80.333
R14351 A[5].n20 A[5].t57 80.333
R14352 A[5].n34 A[5].t38 80.333
R14353 A[5].t20 A[5].n29 80.333
R14354 A[5].n32 A[5].t44 80.333
R14355 A[5].n5 A[5].n4 61.856
R14356 A[5].n36 A[5].n35 45.674
R14357 A[5].n13 A[5].n3 40.051
R14358 A[5].n19 A[5].n18 28.418
R14359 A[5].n13 A[5].n12 27.336
R14360 A[5].n18 A[5].n17 24.266
R14361 A[5].n33 A[5].n31 14.9
R14362 A[5].n19 A[5].n13 11.117
R14363 A[5].n9 A[5].n6 6.615
R14364 A[5].n37 A[5].n36 3.545
R14365 A[5].n35 A[5].n33 2.599
R14366 A[5].n25 A[5].n23 0.426
R14367 A[5].n26 A[5].n25 0.09
R14368 A[5].n18 A[5].n15 0.004
R14369 a_55853_15446.n0 a_55853_15446.t9 214.335
R14370 a_55853_15446.t7 a_55853_15446.n0 214.335
R14371 a_55853_15446.n1 a_55853_15446.t7 143.851
R14372 a_55853_15446.n1 a_55853_15446.t8 135.658
R14373 a_55853_15446.n0 a_55853_15446.t10 80.333
R14374 a_55853_15446.n2 a_55853_15446.t3 28.565
R14375 a_55853_15446.n2 a_55853_15446.t4 28.565
R14376 a_55853_15446.n4 a_55853_15446.t5 28.565
R14377 a_55853_15446.n4 a_55853_15446.t0 28.565
R14378 a_55853_15446.n7 a_55853_15446.t1 28.565
R14379 a_55853_15446.t2 a_55853_15446.n7 28.565
R14380 a_55853_15446.n3 a_55853_15446.t6 9.714
R14381 a_55853_15446.n3 a_55853_15446.n2 1.003
R14382 a_55853_15446.n6 a_55853_15446.n5 0.833
R14383 a_55853_15446.n5 a_55853_15446.n4 0.653
R14384 a_55853_15446.n7 a_55853_15446.n6 0.653
R14385 a_55853_15446.n5 a_55853_15446.n3 0.341
R14386 a_55853_15446.n6 a_55853_15446.n1 0.032
R14387 opcode[3].n1 opcode[3].t9 1374.12
R14388 opcode[3].n8 opcode[3].t10 1374.12
R14389 opcode[3].n13 opcode[3].t25 1374.12
R14390 opcode[3].n18 opcode[3].t61 1374.12
R14391 opcode[3].n23 opcode[3].t32 1374.12
R14392 opcode[3].n28 opcode[3].t33 1374.12
R14393 opcode[3].n33 opcode[3].t47 1374.12
R14394 opcode[3].n38 opcode[3].t48 1374.12
R14395 opcode[3].n3 opcode[3].t26 623.291
R14396 opcode[3].n6 opcode[3].t52 623.291
R14397 opcode[3].n11 opcode[3].t45 623.291
R14398 opcode[3].n16 opcode[3].t49 623.291
R14399 opcode[3].n21 opcode[3].t19 623.291
R14400 opcode[3].n26 opcode[3].t60 623.291
R14401 opcode[3].n31 opcode[3].t40 623.291
R14402 opcode[3].n36 opcode[3].t63 623.291
R14403 opcode[3].n3 opcode[3].t1 610.283
R14404 opcode[3].n6 opcode[3].t3 610.283
R14405 opcode[3].n11 opcode[3].t12 610.283
R14406 opcode[3].n16 opcode[3].t7 610.283
R14407 opcode[3].n21 opcode[3].t38 610.283
R14408 opcode[3].n26 opcode[3].t16 610.283
R14409 opcode[3].n31 opcode[3].t39 610.283
R14410 opcode[3].n36 opcode[3].t42 610.283
R14411 opcode[3].n40 opcode[3].n39 490.381
R14412 opcode[3].n43 opcode[3].n42 333.112
R14413 opcode[3].n42 opcode[3].n41 327.388
R14414 opcode[3].n46 opcode[3].n45 327.18
R14415 opcode[3].n44 opcode[3].n43 327.076
R14416 opcode[3].n45 opcode[3].n44 326.139
R14417 opcode[3].n1 opcode[3].t23 326.034
R14418 opcode[3].n8 opcode[3].t46 326.034
R14419 opcode[3].n13 opcode[3].t54 326.034
R14420 opcode[3].n18 opcode[3].t35 326.034
R14421 opcode[3].n23 opcode[3].t20 326.034
R14422 opcode[3].n28 opcode[3].t11 326.034
R14423 opcode[3].n33 opcode[3].t2 326.034
R14424 opcode[3].n38 opcode[3].t57 326.034
R14425 opcode[3].n41 opcode[3].n40 325.931
R14426 opcode[3].n2 opcode[3].t5 286.438
R14427 opcode[3].n2 opcode[3].t28 286.438
R14428 opcode[3].n5 opcode[3].t51 286.438
R14429 opcode[3].n5 opcode[3].t53 286.438
R14430 opcode[3].n10 opcode[3].t44 286.438
R14431 opcode[3].n10 opcode[3].t55 286.438
R14432 opcode[3].n15 opcode[3].t29 286.438
R14433 opcode[3].n15 opcode[3].t50 286.438
R14434 opcode[3].n20 opcode[3].t17 286.438
R14435 opcode[3].n20 opcode[3].t36 286.438
R14436 opcode[3].n25 opcode[3].t59 286.438
R14437 opcode[3].n25 opcode[3].t22 286.438
R14438 opcode[3].n30 opcode[3].t14 286.438
R14439 opcode[3].n30 opcode[3].t43 286.438
R14440 opcode[3].n35 opcode[3].t62 286.438
R14441 opcode[3].n35 opcode[3].t18 286.438
R14442 opcode[3] opcode[3].n46 220.752
R14443 opcode[3].n0 opcode[3].t27 206.421
R14444 opcode[3].t23 opcode[3].n0 206.421
R14445 opcode[3].n7 opcode[3].t21 206.421
R14446 opcode[3].t46 opcode[3].n7 206.421
R14447 opcode[3].n12 opcode[3].t58 206.421
R14448 opcode[3].t54 opcode[3].n12 206.421
R14449 opcode[3].n17 opcode[3].t41 206.421
R14450 opcode[3].t35 opcode[3].n17 206.421
R14451 opcode[3].n22 opcode[3].t31 206.421
R14452 opcode[3].t20 opcode[3].n22 206.421
R14453 opcode[3].n27 opcode[3].t15 206.421
R14454 opcode[3].t11 opcode[3].n27 206.421
R14455 opcode[3].n32 opcode[3].t6 206.421
R14456 opcode[3].t2 opcode[3].n32 206.421
R14457 opcode[3].n37 opcode[3].t34 206.421
R14458 opcode[3].t57 opcode[3].n37 206.421
R14459 opcode[3].n46 opcode[3].n4 164.203
R14460 opcode[3].n45 opcode[3].n9 163.896
R14461 opcode[3].n43 opcode[3].n19 163.095
R14462 opcode[3].n41 opcode[3].n29 162.871
R14463 opcode[3].n44 opcode[3].n14 162.596
R14464 opcode[3].t26 opcode[3].n2 160.666
R14465 opcode[3].t52 opcode[3].n5 160.666
R14466 opcode[3].t45 opcode[3].n10 160.666
R14467 opcode[3].t49 opcode[3].n15 160.666
R14468 opcode[3].t19 opcode[3].n20 160.666
R14469 opcode[3].t60 opcode[3].n25 160.666
R14470 opcode[3].t40 opcode[3].n30 160.666
R14471 opcode[3].t63 opcode[3].n35 160.666
R14472 opcode[3].n42 opcode[3].n24 158.147
R14473 opcode[3].n40 opcode[3].n34 157.689
R14474 opcode[3].n0 opcode[3].t24 80.333
R14475 opcode[3].n7 opcode[3].t0 80.333
R14476 opcode[3].n12 opcode[3].t56 80.333
R14477 opcode[3].n17 opcode[3].t37 80.333
R14478 opcode[3].n22 opcode[3].t30 80.333
R14479 opcode[3].n27 opcode[3].t13 80.333
R14480 opcode[3].n32 opcode[3].t4 80.333
R14481 opcode[3].n37 opcode[3].t8 80.333
R14482 opcode[3] opcode[3].n47 14.9
R14483 opcode[3].n47 opcode[3] 14.601
R14484 opcode[3].n47 opcode[3] 1.772
R14485 opcode[3].n47 opcode[3] 1.736
R14486 opcode[3].n9 opcode[3].n6 1.617
R14487 opcode[3].n14 opcode[3].n11 1.617
R14488 opcode[3].n19 opcode[3].n16 1.617
R14489 opcode[3].n24 opcode[3].n21 1.617
R14490 opcode[3].n29 opcode[3].n26 1.617
R14491 opcode[3].n34 opcode[3].n31 1.617
R14492 opcode[3].n39 opcode[3].n36 1.617
R14493 opcode[3].n4 opcode[3].n3 1.616
R14494 opcode[3].n4 opcode[3].n1 0.003
R14495 opcode[3].n9 opcode[3].n8 0.003
R14496 opcode[3].n14 opcode[3].n13 0.003
R14497 opcode[3].n19 opcode[3].n18 0.003
R14498 opcode[3].n24 opcode[3].n23 0.003
R14499 opcode[3].n29 opcode[3].n28 0.003
R14500 opcode[3].n34 opcode[3].n33 0.003
R14501 opcode[3].n39 opcode[3].n38 0.003
R14502 a_3424_n2152.n2 a_3424_n2152.t6 448.382
R14503 a_3424_n2152.n1 a_3424_n2152.t5 286.438
R14504 a_3424_n2152.n1 a_3424_n2152.t7 286.438
R14505 a_3424_n2152.n0 a_3424_n2152.t4 247.69
R14506 a_3424_n2152.n4 a_3424_n2152.n3 182.117
R14507 a_3424_n2152.t6 a_3424_n2152.n1 160.666
R14508 a_3424_n2152.n3 a_3424_n2152.t0 28.568
R14509 a_3424_n2152.n4 a_3424_n2152.t1 28.565
R14510 a_3424_n2152.t2 a_3424_n2152.n4 28.565
R14511 a_3424_n2152.n0 a_3424_n2152.t3 18.127
R14512 a_3424_n2152.n2 a_3424_n2152.n0 4.039
R14513 a_3424_n2152.n3 a_3424_n2152.n2 0.937
R14514 a_37894_4002.n2 a_37894_4002.t10 214.335
R14515 a_37894_4002.t9 a_37894_4002.n2 214.335
R14516 a_37894_4002.n3 a_37894_4002.t9 143.851
R14517 a_37894_4002.n3 a_37894_4002.t7 135.658
R14518 a_37894_4002.n2 a_37894_4002.t8 80.333
R14519 a_37894_4002.n4 a_37894_4002.t4 28.565
R14520 a_37894_4002.n4 a_37894_4002.t6 28.565
R14521 a_37894_4002.n0 a_37894_4002.t5 28.565
R14522 a_37894_4002.n0 a_37894_4002.t2 28.565
R14523 a_37894_4002.n7 a_37894_4002.t3 28.565
R14524 a_37894_4002.t0 a_37894_4002.n7 28.565
R14525 a_37894_4002.n1 a_37894_4002.t1 9.714
R14526 a_37894_4002.n1 a_37894_4002.n0 1.003
R14527 a_37894_4002.n6 a_37894_4002.n5 0.833
R14528 a_37894_4002.n5 a_37894_4002.n4 0.653
R14529 a_37894_4002.n7 a_37894_4002.n6 0.653
R14530 a_37894_4002.n6 a_37894_4002.n1 0.341
R14531 a_37894_4002.n5 a_37894_4002.n3 0.032
R14532 a_38484_3565.t4 a_38484_3565.t6 800.071
R14533 a_38484_3565.n2 a_38484_3565.n1 659.097
R14534 a_38484_3565.n0 a_38484_3565.t5 285.109
R14535 a_38484_3565.n1 a_38484_3565.t4 193.602
R14536 a_38484_3565.n4 a_38484_3565.n3 192.754
R14537 a_38484_3565.n0 a_38484_3565.t7 160.666
R14538 a_38484_3565.n1 a_38484_3565.n0 91.507
R14539 a_38484_3565.n3 a_38484_3565.t0 28.568
R14540 a_38484_3565.t2 a_38484_3565.n4 28.565
R14541 a_38484_3565.n4 a_38484_3565.t1 28.565
R14542 a_38484_3565.n2 a_38484_3565.t3 19.061
R14543 a_38484_3565.n3 a_38484_3565.n2 1.005
R14544 a_11155_13581.n2 a_11155_13581.t6 448.381
R14545 a_11155_13581.n1 a_11155_13581.t5 286.438
R14546 a_11155_13581.n1 a_11155_13581.t4 286.438
R14547 a_11155_13581.n0 a_11155_13581.t7 247.69
R14548 a_11155_13581.n4 a_11155_13581.n3 182.117
R14549 a_11155_13581.t6 a_11155_13581.n1 160.666
R14550 a_11155_13581.n3 a_11155_13581.t0 28.568
R14551 a_11155_13581.n4 a_11155_13581.t1 28.565
R14552 a_11155_13581.t2 a_11155_13581.n4 28.565
R14553 a_11155_13581.n0 a_11155_13581.t3 18.127
R14554 a_11155_13581.n2 a_11155_13581.n0 4.036
R14555 a_11155_13581.n3 a_11155_13581.n2 0.937
R14556 a_10509_14454.n0 a_10509_14454.n9 167.433
R14557 a_10509_14454.t0 a_10509_14454.n0 14.282
R14558 a_10509_14454.n0 a_10509_14454.t1 14.282
R14559 a_10509_14454.n9 a_10509_14454.n8 77.784
R14560 a_10509_14454.n8 a_10509_14454.n6 77.456
R14561 a_10509_14454.n6 a_10509_14454.n4 77.456
R14562 a_10509_14454.n4 a_10509_14454.n2 75.815
R14563 a_10509_14454.n9 a_10509_14454.t2 104.259
R14564 a_10509_14454.n8 a_10509_14454.n7 89.977
R14565 a_10509_14454.n7 a_10509_14454.t4 14.282
R14566 a_10509_14454.n7 a_10509_14454.t5 14.282
R14567 a_10509_14454.n6 a_10509_14454.n5 89.977
R14568 a_10509_14454.n5 a_10509_14454.t3 14.282
R14569 a_10509_14454.n5 a_10509_14454.t7 14.282
R14570 a_10509_14454.n4 a_10509_14454.n3 89.977
R14571 a_10509_14454.n3 a_10509_14454.t6 14.282
R14572 a_10509_14454.n3 a_10509_14454.t8 14.282
R14573 a_10509_14454.n2 a_10509_14454.t10 104.259
R14574 a_10509_14454.n2 a_10509_14454.n1 167.433
R14575 a_10509_14454.n1 a_10509_14454.t11 14.282
R14576 a_10509_14454.n1 a_10509_14454.t9 14.282
R14577 a_9976_13724.t0 a_9976_13724.n0 14.283
R14578 a_9976_13724.n0 a_9976_13724.n5 0.852
R14579 a_9976_13724.n5 a_9976_13724.n6 4.366
R14580 a_9976_13724.n6 a_9976_13724.n7 258.161
R14581 a_9976_13724.n7 a_9976_13724.t6 14.282
R14582 a_9976_13724.n7 a_9976_13724.t5 14.282
R14583 a_9976_13724.n6 a_9976_13724.t7 14.283
R14584 a_9976_13724.n5 a_9976_13724.n4 97.614
R14585 a_9976_13724.n4 a_9976_13724.t9 200.029
R14586 a_9976_13724.t9 a_9976_13724.n3 206.421
R14587 a_9976_13724.n3 a_9976_13724.t11 80.333
R14588 a_9976_13724.n3 a_9976_13724.t8 206.421
R14589 a_9976_13724.n4 a_9976_13724.t10 1527.4
R14590 a_9976_13724.t10 a_9976_13724.n2 657.379
R14591 a_9976_13724.n2 a_9976_13724.t4 8.7
R14592 a_9976_13724.n2 a_9976_13724.t3 8.7
R14593 a_9976_13724.n0 a_9976_13724.n1 258.161
R14594 a_9976_13724.n1 a_9976_13724.t1 14.282
R14595 a_9976_13724.n1 a_9976_13724.t2 14.282
R14596 a_23787_8115.n2 a_23787_8115.t7 448.381
R14597 a_23787_8115.n1 a_23787_8115.t6 286.438
R14598 a_23787_8115.n1 a_23787_8115.t4 286.438
R14599 a_23787_8115.n0 a_23787_8115.t5 247.69
R14600 a_23787_8115.n4 a_23787_8115.n3 182.117
R14601 a_23787_8115.t7 a_23787_8115.n1 160.666
R14602 a_23787_8115.n3 a_23787_8115.t0 28.568
R14603 a_23787_8115.n4 a_23787_8115.t1 28.565
R14604 a_23787_8115.t2 a_23787_8115.n4 28.565
R14605 a_23787_8115.n0 a_23787_8115.t3 18.127
R14606 a_23787_8115.n2 a_23787_8115.n0 4.036
R14607 a_23787_8115.n3 a_23787_8115.n2 0.937
R14608 a_60201_9159.t5 a_60201_9159.t6 800.071
R14609 a_60201_9159.n3 a_60201_9159.n2 672.951
R14610 a_60201_9159.n1 a_60201_9159.t4 285.109
R14611 a_60201_9159.n2 a_60201_9159.t5 193.602
R14612 a_60201_9159.n1 a_60201_9159.t7 160.666
R14613 a_60201_9159.n2 a_60201_9159.n1 91.507
R14614 a_60201_9159.t0 a_60201_9159.n4 28.57
R14615 a_60201_9159.n0 a_60201_9159.t2 28.565
R14616 a_60201_9159.n0 a_60201_9159.t3 28.565
R14617 a_60201_9159.n4 a_60201_9159.t1 17.638
R14618 a_60201_9159.n3 a_60201_9159.n0 0.69
R14619 a_60201_9159.n4 a_60201_9159.n3 0.6
R14620 a_61197_9746.n0 a_61197_9746.t4 14.282
R14621 a_61197_9746.n0 a_61197_9746.t1 14.282
R14622 a_61197_9746.n1 a_61197_9746.t5 14.282
R14623 a_61197_9746.n1 a_61197_9746.t3 14.282
R14624 a_61197_9746.n3 a_61197_9746.t2 14.282
R14625 a_61197_9746.t0 a_61197_9746.n3 14.282
R14626 a_61197_9746.n3 a_61197_9746.n2 2.546
R14627 a_61197_9746.n2 a_61197_9746.n1 2.367
R14628 a_61197_9746.n2 a_61197_9746.n0 0.001
R14629 a_3700_13728.t1 a_3700_13728.n0 14.282
R14630 a_3700_13728.n0 a_3700_13728.t2 14.282
R14631 a_3700_13728.n0 a_3700_13728.n1 258.161
R14632 a_3700_13728.n1 a_3700_13728.t3 14.283
R14633 a_3700_13728.n1 a_3700_13728.n7 4.366
R14634 a_3700_13728.n7 a_3700_13728.n5 0.852
R14635 a_3700_13728.n5 a_3700_13728.n6 258.161
R14636 a_3700_13728.n6 a_3700_13728.t6 14.282
R14637 a_3700_13728.n6 a_3700_13728.t4 14.282
R14638 a_3700_13728.n5 a_3700_13728.t5 14.283
R14639 a_3700_13728.n7 a_3700_13728.n4 97.614
R14640 a_3700_13728.n4 a_3700_13728.t8 200.029
R14641 a_3700_13728.t8 a_3700_13728.n3 206.421
R14642 a_3700_13728.n3 a_3700_13728.t9 80.333
R14643 a_3700_13728.n3 a_3700_13728.t10 206.421
R14644 a_3700_13728.n4 a_3700_13728.t11 1527.4
R14645 a_3700_13728.t11 a_3700_13728.n2 657.379
R14646 a_3700_13728.n2 a_3700_13728.t0 8.7
R14647 a_3700_13728.n2 a_3700_13728.t7 8.7
R14648 a_3642_14458.n2 a_3642_14458.t7 867.497
R14649 a_3642_14458.n2 a_3642_14458.t5 591.811
R14650 a_3642_14458.n1 a_3642_14458.t6 286.438
R14651 a_3642_14458.n1 a_3642_14458.t4 286.438
R14652 a_3642_14458.n4 a_3642_14458.n0 185.55
R14653 a_3642_14458.t7 a_3642_14458.n1 160.666
R14654 a_3642_14458.t2 a_3642_14458.n4 28.568
R14655 a_3642_14458.n0 a_3642_14458.t0 28.565
R14656 a_3642_14458.n0 a_3642_14458.t1 28.565
R14657 a_3642_14458.n3 a_3642_14458.n2 25.354
R14658 a_3642_14458.n3 a_3642_14458.t3 21.376
R14659 a_3642_14458.n4 a_3642_14458.n3 1.638
R14660 a_8289_6359.n2 a_8289_6359.t4 990.34
R14661 a_8289_6359.n2 a_8289_6359.t6 408.211
R14662 a_8289_6359.n1 a_8289_6359.t5 286.438
R14663 a_8289_6359.n1 a_8289_6359.t7 286.438
R14664 a_8289_6359.n4 a_8289_6359.n0 197.272
R14665 a_8289_6359.t4 a_8289_6359.n1 160.666
R14666 a_8289_6359.n3 a_8289_6359.n2 50.288
R14667 a_8289_6359.t2 a_8289_6359.n4 28.568
R14668 a_8289_6359.n0 a_8289_6359.t1 28.565
R14669 a_8289_6359.n0 a_8289_6359.t0 28.565
R14670 a_8289_6359.n3 a_8289_6359.t3 18.144
R14671 a_8289_6359.n4 a_8289_6359.n3 0.52
R14672 a_67135_7303.n4 a_67135_7303.t8 214.335
R14673 a_67135_7303.t7 a_67135_7303.n4 214.335
R14674 a_67135_7303.n5 a_67135_7303.t7 143.851
R14675 a_67135_7303.n5 a_67135_7303.t9 135.658
R14676 a_67135_7303.n4 a_67135_7303.t10 80.333
R14677 a_67135_7303.n0 a_67135_7303.t5 28.565
R14678 a_67135_7303.n0 a_67135_7303.t4 28.565
R14679 a_67135_7303.n2 a_67135_7303.t1 28.565
R14680 a_67135_7303.n2 a_67135_7303.t3 28.565
R14681 a_67135_7303.n7 a_67135_7303.t2 28.565
R14682 a_67135_7303.t0 a_67135_7303.n7 28.565
R14683 a_67135_7303.n1 a_67135_7303.t6 9.714
R14684 a_67135_7303.n1 a_67135_7303.n0 1.003
R14685 a_67135_7303.n6 a_67135_7303.n3 0.833
R14686 a_67135_7303.n3 a_67135_7303.n2 0.653
R14687 a_67135_7303.n7 a_67135_7303.n6 0.653
R14688 a_67135_7303.n3 a_67135_7303.n1 0.341
R14689 a_67135_7303.n6 a_67135_7303.n5 0.032
R14690 a_67372_6666.t0 a_67372_6666.t1 17.4
R14691 a_16795_16385.n0 a_16795_16385.t7 214.335
R14692 a_16795_16385.t8 a_16795_16385.n0 214.335
R14693 a_16795_16385.n1 a_16795_16385.t8 143.851
R14694 a_16795_16385.n1 a_16795_16385.t10 135.658
R14695 a_16795_16385.n0 a_16795_16385.t9 80.333
R14696 a_16795_16385.n2 a_16795_16385.t6 28.565
R14697 a_16795_16385.n2 a_16795_16385.t4 28.565
R14698 a_16795_16385.n4 a_16795_16385.t5 28.565
R14699 a_16795_16385.n4 a_16795_16385.t0 28.565
R14700 a_16795_16385.n7 a_16795_16385.t1 28.565
R14701 a_16795_16385.t2 a_16795_16385.n7 28.565
R14702 a_16795_16385.n3 a_16795_16385.t3 9.714
R14703 a_16795_16385.n3 a_16795_16385.n2 1.003
R14704 a_16795_16385.n6 a_16795_16385.n5 0.833
R14705 a_16795_16385.n5 a_16795_16385.n4 0.653
R14706 a_16795_16385.n7 a_16795_16385.n6 0.653
R14707 a_16795_16385.n5 a_16795_16385.n3 0.341
R14708 a_16795_16385.n6 a_16795_16385.n1 0.032
R14709 a_7305_14428.n2 a_7305_14428.t5 867.497
R14710 a_7305_14428.n2 a_7305_14428.t7 591.811
R14711 a_7305_14428.n1 a_7305_14428.t4 286.438
R14712 a_7305_14428.n1 a_7305_14428.t6 286.438
R14713 a_7305_14428.n4 a_7305_14428.n0 192.754
R14714 a_7305_14428.t5 a_7305_14428.n1 160.666
R14715 a_7305_14428.n3 a_7305_14428.n2 31.175
R14716 a_7305_14428.t2 a_7305_14428.n4 28.568
R14717 a_7305_14428.n0 a_7305_14428.t1 28.565
R14718 a_7305_14428.n0 a_7305_14428.t0 28.565
R14719 a_7305_14428.n3 a_7305_14428.t3 18.726
R14720 a_7305_14428.n4 a_7305_14428.n3 1.123
R14721 a_1916_13125.t0 a_1916_13125.t1 17.4
R14722 a_35001_1426.n0 a_35001_1426.t7 214.335
R14723 a_35001_1426.t10 a_35001_1426.n0 214.335
R14724 a_35001_1426.n1 a_35001_1426.t10 143.851
R14725 a_35001_1426.n1 a_35001_1426.t8 135.658
R14726 a_35001_1426.n0 a_35001_1426.t9 80.333
R14727 a_35001_1426.n2 a_35001_1426.t1 28.565
R14728 a_35001_1426.n2 a_35001_1426.t0 28.565
R14729 a_35001_1426.n4 a_35001_1426.t2 28.565
R14730 a_35001_1426.n4 a_35001_1426.t4 28.565
R14731 a_35001_1426.t3 a_35001_1426.n7 28.565
R14732 a_35001_1426.n7 a_35001_1426.t5 28.565
R14733 a_35001_1426.n6 a_35001_1426.t6 9.714
R14734 a_35001_1426.n7 a_35001_1426.n6 1.003
R14735 a_35001_1426.n5 a_35001_1426.n3 0.833
R14736 a_35001_1426.n3 a_35001_1426.n2 0.653
R14737 a_35001_1426.n5 a_35001_1426.n4 0.653
R14738 a_35001_1426.n6 a_35001_1426.n5 0.341
R14739 a_35001_1426.n3 a_35001_1426.n1 0.032
R14740 a_35591_989.n8 a_35591_989.n7 861.987
R14741 a_35591_989.n7 a_35591_989.n6 560.726
R14742 a_35591_989.t11 a_35591_989.t5 415.315
R14743 a_35591_989.t12 a_35591_989.t13 415.315
R14744 a_35591_989.n3 a_35591_989.t17 394.151
R14745 a_35591_989.n6 a_35591_989.t16 294.653
R14746 a_35591_989.n2 a_35591_989.t6 269.523
R14747 a_35591_989.t17 a_35591_989.n2 269.523
R14748 a_35591_989.n10 a_35591_989.t11 217.716
R14749 a_35591_989.n9 a_35591_989.t7 214.335
R14750 a_35591_989.t5 a_35591_989.n9 214.335
R14751 a_35591_989.n1 a_35591_989.t14 214.335
R14752 a_35591_989.t13 a_35591_989.n1 214.335
R14753 a_35591_989.n8 a_35591_989.t12 198.921
R14754 a_35591_989.n4 a_35591_989.t8 198.043
R14755 a_35591_989.n12 a_35591_989.n0 192.754
R14756 a_35591_989.n2 a_35591_989.t9 160.666
R14757 a_35591_989.n6 a_35591_989.t19 111.663
R14758 a_35591_989.n5 a_35591_989.n3 97.816
R14759 a_35591_989.n4 a_35591_989.t18 93.989
R14760 a_35591_989.n9 a_35591_989.t15 80.333
R14761 a_35591_989.n3 a_35591_989.t10 80.333
R14762 a_35591_989.n1 a_35591_989.t4 80.333
R14763 a_35591_989.n7 a_35591_989.n5 65.07
R14764 a_35591_989.t2 a_35591_989.n12 28.568
R14765 a_35591_989.n0 a_35591_989.t1 28.565
R14766 a_35591_989.n0 a_35591_989.t0 28.565
R14767 a_35591_989.n11 a_35591_989.t3 18.825
R14768 a_35591_989.n10 a_35591_989.n8 16.411
R14769 a_35591_989.n5 a_35591_989.n4 6.615
R14770 a_35591_989.n11 a_35591_989.n10 2.988
R14771 a_35591_989.n12 a_35591_989.n11 1.105
R14772 a_39381_15765.t0 a_39381_15765.n0 14.282
R14773 a_39381_15765.n0 a_39381_15765.t1 14.282
R14774 a_39381_15765.n0 a_39381_15765.n8 122.747
R14775 a_39381_15765.n4 a_39381_15765.n6 74.302
R14776 a_39381_15765.n8 a_39381_15765.n4 50.575
R14777 a_39381_15765.n8 a_39381_15765.n7 157.665
R14778 a_39381_15765.n7 a_39381_15765.t4 8.7
R14779 a_39381_15765.n7 a_39381_15765.t2 8.7
R14780 a_39381_15765.n6 a_39381_15765.n5 90.436
R14781 a_39381_15765.n5 a_39381_15765.t5 14.282
R14782 a_39381_15765.n5 a_39381_15765.t6 14.282
R14783 a_39381_15765.n4 a_39381_15765.n3 90.416
R14784 a_39381_15765.n3 a_39381_15765.t7 14.282
R14785 a_39381_15765.n3 a_39381_15765.t3 14.282
R14786 a_39381_15765.n6 a_39381_15765.n1 293.294
R14787 a_39381_15765.t11 a_39381_15765.n2 160.666
R14788 a_39381_15765.n1 a_39381_15765.t11 867.393
R14789 a_39381_15765.n2 a_39381_15765.t8 287.241
R14790 a_39381_15765.n2 a_39381_15765.t10 287.241
R14791 a_39381_15765.n1 a_39381_15765.t9 545.094
R14792 a_70509_n2116.n0 a_70509_n2116.t2 14.282
R14793 a_70509_n2116.t0 a_70509_n2116.n0 14.282
R14794 a_70509_n2116.n0 a_70509_n2116.n1 258.161
R14795 a_70509_n2116.n1 a_70509_n2116.t1 14.283
R14796 a_70509_n2116.n1 a_70509_n2116.n5 0.852
R14797 a_70509_n2116.n5 a_70509_n2116.n6 4.366
R14798 a_70509_n2116.n6 a_70509_n2116.n7 258.161
R14799 a_70509_n2116.n7 a_70509_n2116.t4 14.282
R14800 a_70509_n2116.n7 a_70509_n2116.t5 14.282
R14801 a_70509_n2116.n6 a_70509_n2116.t6 14.283
R14802 a_70509_n2116.n5 a_70509_n2116.n4 73.514
R14803 a_70509_n2116.n4 a_70509_n2116.t9 1551.5
R14804 a_70509_n2116.t9 a_70509_n2116.n3 656.576
R14805 a_70509_n2116.n3 a_70509_n2116.t7 8.7
R14806 a_70509_n2116.n3 a_70509_n2116.t3 8.7
R14807 a_70509_n2116.n4 a_70509_n2116.t10 224.129
R14808 a_70509_n2116.t10 a_70509_n2116.n2 207.225
R14809 a_70509_n2116.n2 a_70509_n2116.t11 207.225
R14810 a_70509_n2116.n2 a_70509_n2116.t8 80.333
R14811 a_70509_n1998.t3 a_70509_n1998.n0 14.282
R14812 a_70509_n1998.n0 a_70509_n1998.t4 14.282
R14813 a_70509_n1998.n4 a_70509_n1998.n2 77.784
R14814 a_70509_n1998.n6 a_70509_n1998.n4 77.456
R14815 a_70509_n1998.n8 a_70509_n1998.n6 77.456
R14816 a_70509_n1998.n9 a_70509_n1998.n8 75.815
R14817 a_70509_n1998.n0 a_70509_n1998.n9 167.433
R14818 a_70509_n1998.n9 a_70509_n1998.t5 104.259
R14819 a_70509_n1998.n8 a_70509_n1998.n7 89.977
R14820 a_70509_n1998.n7 a_70509_n1998.t10 14.282
R14821 a_70509_n1998.n7 a_70509_n1998.t11 14.282
R14822 a_70509_n1998.n6 a_70509_n1998.n5 89.977
R14823 a_70509_n1998.n5 a_70509_n1998.t6 14.282
R14824 a_70509_n1998.n5 a_70509_n1998.t9 14.282
R14825 a_70509_n1998.n4 a_70509_n1998.n3 89.977
R14826 a_70509_n1998.n3 a_70509_n1998.t7 14.282
R14827 a_70509_n1998.n3 a_70509_n1998.t8 14.282
R14828 a_70509_n1998.n2 a_70509_n1998.t1 104.259
R14829 a_70509_n1998.n2 a_70509_n1998.n1 167.433
R14830 a_70509_n1998.n1 a_70509_n1998.t2 14.282
R14831 a_70509_n1998.n1 a_70509_n1998.t0 14.282
R14832 a_48248_308.t0 a_48248_308.t1 380.209
R14833 a_48855_n1313.n7 a_48855_n1313.n6 861.987
R14834 a_48855_n1313.n6 a_48855_n1313.n5 560.726
R14835 a_48855_n1313.t17 a_48855_n1313.t11 415.315
R14836 a_48855_n1313.t12 a_48855_n1313.t13 415.315
R14837 a_48855_n1313.n2 a_48855_n1313.t8 394.151
R14838 a_48855_n1313.n5 a_48855_n1313.t15 294.653
R14839 a_48855_n1313.n1 a_48855_n1313.t10 269.523
R14840 a_48855_n1313.t8 a_48855_n1313.n1 269.523
R14841 a_48855_n1313.n9 a_48855_n1313.t17 217.716
R14842 a_48855_n1313.n8 a_48855_n1313.t14 214.335
R14843 a_48855_n1313.t11 a_48855_n1313.n8 214.335
R14844 a_48855_n1313.n0 a_48855_n1313.t18 214.335
R14845 a_48855_n1313.t13 a_48855_n1313.n0 214.335
R14846 a_48855_n1313.n7 a_48855_n1313.t12 198.921
R14847 a_48855_n1313.n3 a_48855_n1313.t9 198.043
R14848 a_48855_n1313.n12 a_48855_n1313.n11 192.754
R14849 a_48855_n1313.n1 a_48855_n1313.t4 160.666
R14850 a_48855_n1313.n5 a_48855_n1313.t6 111.663
R14851 a_48855_n1313.n4 a_48855_n1313.n2 97.816
R14852 a_48855_n1313.n3 a_48855_n1313.t5 93.989
R14853 a_48855_n1313.n8 a_48855_n1313.t19 80.333
R14854 a_48855_n1313.n2 a_48855_n1313.t16 80.333
R14855 a_48855_n1313.n0 a_48855_n1313.t7 80.333
R14856 a_48855_n1313.n6 a_48855_n1313.n4 65.07
R14857 a_48855_n1313.n11 a_48855_n1313.t1 28.568
R14858 a_48855_n1313.n12 a_48855_n1313.t3 28.565
R14859 a_48855_n1313.t0 a_48855_n1313.n12 28.565
R14860 a_48855_n1313.n10 a_48855_n1313.t2 18.826
R14861 a_48855_n1313.n9 a_48855_n1313.n7 16.411
R14862 a_48855_n1313.n4 a_48855_n1313.n3 6.615
R14863 a_48855_n1313.n10 a_48855_n1313.n9 5.027
R14864 a_48855_n1313.n11 a_48855_n1313.n10 1.101
R14865 a_52887_1041.n0 a_52887_1041.t1 14.282
R14866 a_52887_1041.t0 a_52887_1041.n0 14.282
R14867 a_52887_1041.n1 a_52887_1041.n9 0.001
R14868 a_52887_1041.n0 a_52887_1041.n1 267.767
R14869 a_52887_1041.n9 a_52887_1041.t6 14.282
R14870 a_52887_1041.n9 a_52887_1041.t2 14.282
R14871 a_52887_1041.n1 a_52887_1041.n7 0.669
R14872 a_52887_1041.n7 a_52887_1041.n8 1.511
R14873 a_52887_1041.n8 a_52887_1041.t7 14.282
R14874 a_52887_1041.n8 a_52887_1041.t8 14.282
R14875 a_52887_1041.n7 a_52887_1041.n6 0.227
R14876 a_52887_1041.n6 a_52887_1041.n3 0.575
R14877 a_52887_1041.n6 a_52887_1041.n5 0.2
R14878 a_52887_1041.n5 a_52887_1041.t10 16.058
R14879 a_52887_1041.n5 a_52887_1041.n4 0.999
R14880 a_52887_1041.n4 a_52887_1041.t9 14.282
R14881 a_52887_1041.n4 a_52887_1041.t11 14.282
R14882 a_52887_1041.n3 a_52887_1041.n2 0.999
R14883 a_52887_1041.n2 a_52887_1041.t4 14.282
R14884 a_52887_1041.n2 a_52887_1041.t5 14.282
R14885 a_52887_1041.n3 a_52887_1041.t3 16.058
R14886 a_47709_7603.n1 a_47709_7603.t5 318.922
R14887 a_47709_7603.n0 a_47709_7603.t7 273.935
R14888 a_47709_7603.n0 a_47709_7603.t4 273.935
R14889 a_47709_7603.n1 a_47709_7603.t6 269.116
R14890 a_47709_7603.n4 a_47709_7603.n3 193.227
R14891 a_47709_7603.t5 a_47709_7603.n0 179.142
R14892 a_47709_7603.n2 a_47709_7603.n1 106.999
R14893 a_47709_7603.n3 a_47709_7603.t3 28.568
R14894 a_47709_7603.t0 a_47709_7603.n4 28.565
R14895 a_47709_7603.n4 a_47709_7603.t1 28.565
R14896 a_47709_7603.n2 a_47709_7603.t2 18.149
R14897 a_47709_7603.n3 a_47709_7603.n2 3.726
R14898 a_48136_6910.t0 a_48136_6910.n7 16.058
R14899 a_48136_6910.n7 a_48136_6910.n5 0.575
R14900 a_48136_6910.n5 a_48136_6910.n9 0.2
R14901 a_48136_6910.n9 a_48136_6910.t3 16.058
R14902 a_48136_6910.n9 a_48136_6910.n8 0.999
R14903 a_48136_6910.n8 a_48136_6910.t4 14.282
R14904 a_48136_6910.n8 a_48136_6910.t5 14.282
R14905 a_48136_6910.n7 a_48136_6910.n6 0.999
R14906 a_48136_6910.n6 a_48136_6910.t1 14.282
R14907 a_48136_6910.n6 a_48136_6910.t2 14.282
R14908 a_48136_6910.n5 a_48136_6910.n3 0.227
R14909 a_48136_6910.n3 a_48136_6910.n4 1.511
R14910 a_48136_6910.n4 a_48136_6910.t7 14.282
R14911 a_48136_6910.n4 a_48136_6910.t6 14.282
R14912 a_48136_6910.n3 a_48136_6910.n0 0.669
R14913 a_48136_6910.n0 a_48136_6910.n1 0.001
R14914 a_48136_6910.n0 a_48136_6910.n2 267.767
R14915 a_48136_6910.n2 a_48136_6910.t11 14.282
R14916 a_48136_6910.n2 a_48136_6910.t9 14.282
R14917 a_48136_6910.n1 a_48136_6910.t8 14.282
R14918 a_48136_6910.n1 a_48136_6910.t10 14.282
R14919 a_48254_6910.n8 a_48254_6910.n7 861.987
R14920 a_48254_6910.n7 a_48254_6910.n6 560.726
R14921 a_48254_6910.t12 a_48254_6910.t22 415.315
R14922 a_48254_6910.t13 a_48254_6910.t14 415.315
R14923 a_48254_6910.n3 a_48254_6910.t21 394.151
R14924 a_48254_6910.n6 a_48254_6910.t20 294.653
R14925 a_48254_6910.n2 a_48254_6910.t10 269.523
R14926 a_48254_6910.t21 a_48254_6910.n2 269.523
R14927 a_48254_6910.n10 a_48254_6910.t12 217.716
R14928 a_48254_6910.n11 a_48254_6910.n10 216.635
R14929 a_48254_6910.n9 a_48254_6910.t8 214.335
R14930 a_48254_6910.t22 a_48254_6910.n9 214.335
R14931 a_48254_6910.n1 a_48254_6910.t16 214.335
R14932 a_48254_6910.t14 a_48254_6910.n1 214.335
R14933 a_48254_6910.n8 a_48254_6910.t13 198.921
R14934 a_48254_6910.n4 a_48254_6910.t9 198.043
R14935 a_48254_6910.n2 a_48254_6910.t17 160.666
R14936 a_48254_6910.n14 a_48254_6910.n12 157.665
R14937 a_48254_6910.n14 a_48254_6910.n13 122.999
R14938 a_48254_6910.n6 a_48254_6910.t18 111.663
R14939 a_48254_6910.n5 a_48254_6910.n3 97.816
R14940 a_48254_6910.n4 a_48254_6910.t19 93.989
R14941 a_48254_6910.n11 a_48254_6910.n0 90.436
R14942 a_48254_6910.n16 a_48254_6910.n15 90.416
R14943 a_48254_6910.n9 a_48254_6910.t15 80.333
R14944 a_48254_6910.n3 a_48254_6910.t11 80.333
R14945 a_48254_6910.n1 a_48254_6910.t23 80.333
R14946 a_48254_6910.n15 a_48254_6910.n11 74.302
R14947 a_48254_6910.n7 a_48254_6910.n5 65.07
R14948 a_48254_6910.n15 a_48254_6910.n14 50.575
R14949 a_48254_6910.n10 a_48254_6910.n8 16.411
R14950 a_48254_6910.n0 a_48254_6910.t4 14.282
R14951 a_48254_6910.n0 a_48254_6910.t6 14.282
R14952 a_48254_6910.n13 a_48254_6910.t1 14.282
R14953 a_48254_6910.n13 a_48254_6910.t0 14.282
R14954 a_48254_6910.n16 a_48254_6910.t5 14.282
R14955 a_48254_6910.t2 a_48254_6910.n16 14.282
R14956 a_48254_6910.n12 a_48254_6910.t7 8.7
R14957 a_48254_6910.n12 a_48254_6910.t3 8.7
R14958 a_48254_6910.n5 a_48254_6910.n4 6.615
R14959 a_51119_8152.n0 a_51119_8152.t9 214.335
R14960 a_51119_8152.t8 a_51119_8152.n0 214.335
R14961 a_51119_8152.n1 a_51119_8152.t8 143.851
R14962 a_51119_8152.n1 a_51119_8152.t7 135.658
R14963 a_51119_8152.n0 a_51119_8152.t10 80.333
R14964 a_51119_8152.n2 a_51119_8152.t5 28.565
R14965 a_51119_8152.n2 a_51119_8152.t4 28.565
R14966 a_51119_8152.n4 a_51119_8152.t6 28.565
R14967 a_51119_8152.n4 a_51119_8152.t0 28.565
R14968 a_51119_8152.t2 a_51119_8152.n7 28.565
R14969 a_51119_8152.n7 a_51119_8152.t1 28.565
R14970 a_51119_8152.n6 a_51119_8152.t3 9.714
R14971 a_51119_8152.n7 a_51119_8152.n6 1.003
R14972 a_51119_8152.n5 a_51119_8152.n3 0.833
R14973 a_51119_8152.n3 a_51119_8152.n2 0.653
R14974 a_51119_8152.n5 a_51119_8152.n4 0.653
R14975 a_51119_8152.n6 a_51119_8152.n5 0.341
R14976 a_51119_8152.n3 a_51119_8152.n1 0.032
R14977 a_51709_7715.t6 a_51709_7715.t4 574.43
R14978 a_51709_7715.n0 a_51709_7715.t7 285.109
R14979 a_51709_7715.n2 a_51709_7715.n1 211.136
R14980 a_51709_7715.n4 a_51709_7715.n3 192.754
R14981 a_51709_7715.n0 a_51709_7715.t5 160.666
R14982 a_51709_7715.n1 a_51709_7715.t6 160.666
R14983 a_51709_7715.n1 a_51709_7715.n0 114.829
R14984 a_51709_7715.n3 a_51709_7715.t1 28.568
R14985 a_51709_7715.n4 a_51709_7715.t0 28.565
R14986 a_51709_7715.t2 a_51709_7715.n4 28.565
R14987 a_51709_7715.n2 a_51709_7715.t3 19.084
R14988 a_51709_7715.n3 a_51709_7715.n2 1.051
R14989 a_63595_1208.n2 a_63595_1208.t8 214.335
R14990 a_63595_1208.t7 a_63595_1208.n2 214.335
R14991 a_63595_1208.n3 a_63595_1208.t7 143.851
R14992 a_63595_1208.n3 a_63595_1208.t9 135.658
R14993 a_63595_1208.n2 a_63595_1208.t10 80.333
R14994 a_63595_1208.n4 a_63595_1208.t1 28.565
R14995 a_63595_1208.n4 a_63595_1208.t0 28.565
R14996 a_63595_1208.n0 a_63595_1208.t3 28.565
R14997 a_63595_1208.n0 a_63595_1208.t5 28.565
R14998 a_63595_1208.t2 a_63595_1208.n7 28.565
R14999 a_63595_1208.n7 a_63595_1208.t4 28.565
R15000 a_63595_1208.n1 a_63595_1208.t6 9.714
R15001 a_63595_1208.n1 a_63595_1208.n0 1.003
R15002 a_63595_1208.n6 a_63595_1208.n5 0.833
R15003 a_63595_1208.n5 a_63595_1208.n4 0.653
R15004 a_63595_1208.n7 a_63595_1208.n6 0.653
R15005 a_63595_1208.n6 a_63595_1208.n1 0.341
R15006 a_63595_1208.n5 a_63595_1208.n3 0.032
R15007 a_23700_6043.n1 a_23700_6043.t4 318.922
R15008 a_23700_6043.n0 a_23700_6043.t6 274.739
R15009 a_23700_6043.n0 a_23700_6043.t7 274.739
R15010 a_23700_6043.n1 a_23700_6043.t5 269.116
R15011 a_23700_6043.t4 a_23700_6043.n0 179.946
R15012 a_23700_6043.n2 a_23700_6043.n1 107.263
R15013 a_23700_6043.t2 a_23700_6043.n4 29.444
R15014 a_23700_6043.n3 a_23700_6043.t1 28.565
R15015 a_23700_6043.n3 a_23700_6043.t0 28.565
R15016 a_23700_6043.n2 a_23700_6043.t3 18.145
R15017 a_23700_6043.n4 a_23700_6043.n2 2.878
R15018 a_23700_6043.n4 a_23700_6043.n3 0.764
R15019 a_44702_7583.t0 a_44702_7583.t1 17.4
R15020 a_20054_1744.t1 a_20054_1744.n0 14.282
R15021 a_20054_1744.n0 a_20054_1744.t4 14.282
R15022 a_20054_1744.n0 a_20054_1744.n1 258.161
R15023 a_20054_1744.n1 a_20054_1744.n7 4.366
R15024 a_20054_1744.n7 a_20054_1744.n5 0.852
R15025 a_20054_1744.n5 a_20054_1744.n6 258.161
R15026 a_20054_1744.n6 a_20054_1744.t7 14.282
R15027 a_20054_1744.n6 a_20054_1744.t5 14.282
R15028 a_20054_1744.n5 a_20054_1744.t6 14.283
R15029 a_20054_1744.n7 a_20054_1744.n4 97.614
R15030 a_20054_1744.n4 a_20054_1744.t9 200.029
R15031 a_20054_1744.t9 a_20054_1744.n3 206.421
R15032 a_20054_1744.n3 a_20054_1744.t10 80.333
R15033 a_20054_1744.n3 a_20054_1744.t8 206.421
R15034 a_20054_1744.n4 a_20054_1744.t11 1527.4
R15035 a_20054_1744.t11 a_20054_1744.n2 657.379
R15036 a_20054_1744.n2 a_20054_1744.t0 8.7
R15037 a_20054_1744.n2 a_20054_1744.t2 8.7
R15038 a_20054_1744.n1 a_20054_1744.t3 14.283
R15039 a_20611_n2633.n1 a_20611_n2633.t6 867.497
R15040 a_20611_n2633.n1 a_20611_n2633.t4 615.911
R15041 a_20611_n2633.n0 a_20611_n2633.t5 286.438
R15042 a_20611_n2633.n0 a_20611_n2633.t7 286.438
R15043 a_20611_n2633.n4 a_20611_n2633.n3 185.55
R15044 a_20611_n2633.t6 a_20611_n2633.n0 160.666
R15045 a_20611_n2633.n3 a_20611_n2633.t1 28.568
R15046 a_20611_n2633.n4 a_20611_n2633.t0 28.565
R15047 a_20611_n2633.t2 a_20611_n2633.n4 28.565
R15048 a_20611_n2633.n2 a_20611_n2633.n1 22.948
R15049 a_20611_n2633.n2 a_20611_n2633.t3 20.412
R15050 a_20611_n2633.n3 a_20611_n2633.n2 1.813
R15051 a_1964_13805.n3 a_1964_13805.n2 1056.23
R15052 a_1964_13805.n2 a_1964_13805.t6 990.34
R15053 a_1964_13805.n2 a_1964_13805.t5 408.211
R15054 a_1964_13805.n1 a_1964_13805.t4 286.438
R15055 a_1964_13805.n1 a_1964_13805.t7 286.438
R15056 a_1964_13805.t6 a_1964_13805.n1 160.666
R15057 a_1964_13805.n3 a_1964_13805.n0 149.031
R15058 a_1964_13805.n4 a_1964_13805.n3 67.391
R15059 a_1964_13805.n0 a_1964_13805.t1 28.568
R15060 a_1964_13805.t0 a_1964_13805.n4 28.565
R15061 a_1964_13805.n4 a_1964_13805.t3 28.565
R15062 a_1964_13805.n0 a_1964_13805.t2 17.64
R15063 a_1089_14458.n0 a_1089_14458.n9 167.433
R15064 a_1089_14458.t3 a_1089_14458.n0 14.282
R15065 a_1089_14458.n0 a_1089_14458.t4 14.282
R15066 a_1089_14458.n9 a_1089_14458.n8 77.784
R15067 a_1089_14458.n8 a_1089_14458.n6 77.456
R15068 a_1089_14458.n6 a_1089_14458.n4 77.456
R15069 a_1089_14458.n4 a_1089_14458.n2 75.815
R15070 a_1089_14458.n9 a_1089_14458.t5 104.259
R15071 a_1089_14458.n8 a_1089_14458.n7 89.977
R15072 a_1089_14458.n7 a_1089_14458.t2 14.282
R15073 a_1089_14458.n7 a_1089_14458.t1 14.282
R15074 a_1089_14458.n6 a_1089_14458.n5 89.977
R15075 a_1089_14458.n5 a_1089_14458.t0 14.282
R15076 a_1089_14458.n5 a_1089_14458.t7 14.282
R15077 a_1089_14458.n4 a_1089_14458.n3 89.977
R15078 a_1089_14458.n3 a_1089_14458.t6 14.282
R15079 a_1089_14458.n3 a_1089_14458.t8 14.282
R15080 a_1089_14458.n2 a_1089_14458.t11 104.259
R15081 a_1089_14458.n2 a_1089_14458.n1 167.433
R15082 a_1089_14458.n1 a_1089_14458.t10 14.282
R15083 a_1089_14458.n1 a_1089_14458.t9 14.282
R15084 a_65651_3118.n0 a_65651_3118.n1 0.001
R15085 a_65651_3118.t0 a_65651_3118.n0 14.282
R15086 a_65651_3118.n0 a_65651_3118.t6 14.282
R15087 a_65651_3118.n1 a_65651_3118.n9 267.767
R15088 a_65651_3118.n9 a_65651_3118.t7 14.282
R15089 a_65651_3118.n9 a_65651_3118.t8 14.282
R15090 a_65651_3118.n1 a_65651_3118.n7 0.669
R15091 a_65651_3118.n7 a_65651_3118.n8 1.511
R15092 a_65651_3118.n8 a_65651_3118.t11 14.282
R15093 a_65651_3118.n8 a_65651_3118.t10 14.282
R15094 a_65651_3118.n7 a_65651_3118.n6 0.227
R15095 a_65651_3118.n6 a_65651_3118.n3 0.575
R15096 a_65651_3118.n6 a_65651_3118.n5 0.2
R15097 a_65651_3118.n5 a_65651_3118.t5 16.058
R15098 a_65651_3118.n5 a_65651_3118.n4 0.999
R15099 a_65651_3118.n4 a_65651_3118.t4 14.282
R15100 a_65651_3118.n4 a_65651_3118.t3 14.282
R15101 a_65651_3118.n3 a_65651_3118.n2 0.999
R15102 a_65651_3118.n2 a_65651_3118.t1 14.282
R15103 a_65651_3118.n2 a_65651_3118.t9 14.282
R15104 a_65651_3118.n3 a_65651_3118.t2 16.058
R15105 a_53312_9674.t5 a_53312_9674.n3 404.877
R15106 a_53312_9674.n2 a_53312_9674.t8 210.902
R15107 a_53312_9674.n4 a_53312_9674.t5 136.943
R15108 a_53312_9674.n3 a_53312_9674.n2 107.801
R15109 a_53312_9674.n2 a_53312_9674.t7 80.333
R15110 a_53312_9674.n3 a_53312_9674.t6 80.333
R15111 a_53312_9674.n1 a_53312_9674.t4 17.4
R15112 a_53312_9674.n1 a_53312_9674.t1 17.4
R15113 a_53312_9674.t0 a_53312_9674.n5 15.032
R15114 a_53312_9674.n0 a_53312_9674.t3 14.282
R15115 a_53312_9674.n0 a_53312_9674.t2 14.282
R15116 a_53312_9674.n5 a_53312_9674.n0 1.65
R15117 a_53312_9674.n4 a_53312_9674.n1 0.672
R15118 a_53312_9674.n5 a_53312_9674.n4 0.665
R15119 a_53576_9091.t6 a_53576_9091.t7 800.071
R15120 a_53576_9091.n3 a_53576_9091.n2 672.951
R15121 a_53576_9091.n1 a_53576_9091.t4 285.109
R15122 a_53576_9091.n2 a_53576_9091.t6 193.602
R15123 a_53576_9091.n1 a_53576_9091.t5 160.666
R15124 a_53576_9091.n2 a_53576_9091.n1 91.507
R15125 a_53576_9091.t2 a_53576_9091.n4 28.57
R15126 a_53576_9091.n0 a_53576_9091.t0 28.565
R15127 a_53576_9091.n0 a_53576_9091.t1 28.565
R15128 a_53576_9091.n4 a_53576_9091.t3 17.638
R15129 a_53576_9091.n3 a_53576_9091.n0 0.69
R15130 a_53576_9091.n4 a_53576_9091.n3 0.6
R15131 a_3923_n2178.n1 a_3923_n2178.t5 990.34
R15132 a_3923_n2178.n1 a_3923_n2178.t4 408.211
R15133 a_3923_n2178.n0 a_3923_n2178.t6 286.438
R15134 a_3923_n2178.n0 a_3923_n2178.t7 286.438
R15135 a_3923_n2178.n4 a_3923_n2178.n3 185.55
R15136 a_3923_n2178.t5 a_3923_n2178.n0 160.666
R15137 a_3923_n2178.n3 a_3923_n2178.t2 28.568
R15138 a_3923_n2178.t0 a_3923_n2178.n4 28.565
R15139 a_3923_n2178.n4 a_3923_n2178.t3 28.565
R15140 a_3923_n2178.n2 a_3923_n2178.n1 24.399
R15141 a_3923_n2178.n2 a_3923_n2178.t1 21.554
R15142 a_3923_n2178.n3 a_3923_n2178.n2 1.602
R15143 a_4568_n3485.t0 a_4568_n3485.t1 17.4
R15144 a_4300_1740.t5 a_4300_1740.n0 14.282
R15145 a_4300_1740.n0 a_4300_1740.t7 14.282
R15146 a_4300_1740.n0 a_4300_1740.n1 258.161
R15147 a_4300_1740.n1 a_4300_1740.t6 14.283
R15148 a_4300_1740.n1 a_4300_1740.n5 0.852
R15149 a_4300_1740.n5 a_4300_1740.n6 4.366
R15150 a_4300_1740.n6 a_4300_1740.n7 258.161
R15151 a_4300_1740.n7 a_4300_1740.t1 14.282
R15152 a_4300_1740.n7 a_4300_1740.t2 14.282
R15153 a_4300_1740.n6 a_4300_1740.t3 14.283
R15154 a_4300_1740.n5 a_4300_1740.n4 97.614
R15155 a_4300_1740.n4 a_4300_1740.t10 200.029
R15156 a_4300_1740.t10 a_4300_1740.n3 206.421
R15157 a_4300_1740.n3 a_4300_1740.t11 80.333
R15158 a_4300_1740.n3 a_4300_1740.t9 206.421
R15159 a_4300_1740.n4 a_4300_1740.t8 1527.4
R15160 a_4300_1740.t8 a_4300_1740.n2 657.379
R15161 a_4300_1740.n2 a_4300_1740.t0 8.7
R15162 a_4300_1740.n2 a_4300_1740.t4 8.7
R15163 a_21956_20862.t2 a_21956_20862.n0 14.282
R15164 a_21956_20862.n0 a_21956_20862.t3 14.282
R15165 a_21956_20862.n0 a_21956_20862.n1 258.161
R15166 a_21956_20862.n1 a_21956_20862.t4 14.283
R15167 a_21956_20862.n1 a_21956_20862.n7 4.366
R15168 a_21956_20862.n7 a_21956_20862.n5 0.852
R15169 a_21956_20862.n5 a_21956_20862.n6 258.161
R15170 a_21956_20862.n6 a_21956_20862.t6 14.282
R15171 a_21956_20862.n6 a_21956_20862.t5 14.282
R15172 a_21956_20862.n5 a_21956_20862.t7 14.283
R15173 a_21956_20862.n7 a_21956_20862.n4 97.614
R15174 a_21956_20862.n4 a_21956_20862.t11 200.029
R15175 a_21956_20862.t11 a_21956_20862.n3 206.421
R15176 a_21956_20862.n3 a_21956_20862.t9 80.333
R15177 a_21956_20862.n3 a_21956_20862.t10 206.421
R15178 a_21956_20862.n4 a_21956_20862.t8 1527.4
R15179 a_21956_20862.t8 a_21956_20862.n2 657.379
R15180 a_21956_20862.n2 a_21956_20862.t1 8.7
R15181 a_21956_20862.n2 a_21956_20862.t0 8.7
R15182 a_22489_21592.n0 a_22489_21592.t0 14.282
R15183 a_22489_21592.t6 a_22489_21592.n0 14.282
R15184 a_22489_21592.n0 a_22489_21592.n9 89.977
R15185 a_22489_21592.n6 a_22489_21592.n7 77.784
R15186 a_22489_21592.n9 a_22489_21592.n6 77.456
R15187 a_22489_21592.n9 a_22489_21592.n4 77.456
R15188 a_22489_21592.n4 a_22489_21592.n2 75.815
R15189 a_22489_21592.n7 a_22489_21592.n8 167.433
R15190 a_22489_21592.n8 a_22489_21592.t11 14.282
R15191 a_22489_21592.n8 a_22489_21592.t10 14.282
R15192 a_22489_21592.n7 a_22489_21592.t9 104.259
R15193 a_22489_21592.n6 a_22489_21592.n5 89.977
R15194 a_22489_21592.n5 a_22489_21592.t1 14.282
R15195 a_22489_21592.n5 a_22489_21592.t2 14.282
R15196 a_22489_21592.n4 a_22489_21592.n3 89.977
R15197 a_22489_21592.n3 a_22489_21592.t7 14.282
R15198 a_22489_21592.n3 a_22489_21592.t8 14.282
R15199 a_22489_21592.n2 a_22489_21592.t5 104.259
R15200 a_22489_21592.n2 a_22489_21592.n1 167.433
R15201 a_22489_21592.n1 a_22489_21592.t4 14.282
R15202 a_22489_21592.n1 a_22489_21592.t3 14.282
R15203 a_20103_5350.n0 a_20103_5350.n1 0.001
R15204 a_20103_5350.t0 a_20103_5350.n0 14.282
R15205 a_20103_5350.n0 a_20103_5350.t7 14.282
R15206 a_20103_5350.n1 a_20103_5350.n9 267.767
R15207 a_20103_5350.n9 a_20103_5350.t11 14.282
R15208 a_20103_5350.n9 a_20103_5350.t4 14.282
R15209 a_20103_5350.n1 a_20103_5350.n7 0.669
R15210 a_20103_5350.n7 a_20103_5350.n8 1.511
R15211 a_20103_5350.n8 a_20103_5350.t5 14.282
R15212 a_20103_5350.n8 a_20103_5350.t6 14.282
R15213 a_20103_5350.n7 a_20103_5350.n6 0.227
R15214 a_20103_5350.n6 a_20103_5350.n3 0.2
R15215 a_20103_5350.n6 a_20103_5350.n5 0.575
R15216 a_20103_5350.n5 a_20103_5350.t3 16.058
R15217 a_20103_5350.n5 a_20103_5350.n4 0.999
R15218 a_20103_5350.n4 a_20103_5350.t2 14.282
R15219 a_20103_5350.n4 a_20103_5350.t1 14.282
R15220 a_20103_5350.n3 a_20103_5350.n2 0.999
R15221 a_20103_5350.n2 a_20103_5350.t10 14.282
R15222 a_20103_5350.n2 a_20103_5350.t9 14.282
R15223 a_20103_5350.n3 a_20103_5350.t8 16.058
R15224 a_40296_23896.t5 a_40296_23896.t4 800.071
R15225 a_40296_23896.n2 a_40296_23896.n1 659.097
R15226 a_40296_23896.n0 a_40296_23896.t7 285.109
R15227 a_40296_23896.n1 a_40296_23896.t5 193.602
R15228 a_40296_23896.n4 a_40296_23896.n3 192.754
R15229 a_40296_23896.n0 a_40296_23896.t6 160.666
R15230 a_40296_23896.n1 a_40296_23896.n0 91.507
R15231 a_40296_23896.n3 a_40296_23896.t0 28.568
R15232 a_40296_23896.n4 a_40296_23896.t1 28.565
R15233 a_40296_23896.t2 a_40296_23896.n4 28.565
R15234 a_40296_23896.n2 a_40296_23896.t3 19.061
R15235 a_40296_23896.n3 a_40296_23896.n2 1.005
R15236 a_42756_17049.n0 a_42756_17049.t8 214.335
R15237 a_42756_17049.t10 a_42756_17049.n0 214.335
R15238 a_42756_17049.n1 a_42756_17049.t10 143.851
R15239 a_42756_17049.n1 a_42756_17049.t7 135.658
R15240 a_42756_17049.n0 a_42756_17049.t9 80.333
R15241 a_42756_17049.n2 a_42756_17049.t5 28.565
R15242 a_42756_17049.n2 a_42756_17049.t3 28.565
R15243 a_42756_17049.n4 a_42756_17049.t4 28.565
R15244 a_42756_17049.n4 a_42756_17049.t0 28.565
R15245 a_42756_17049.n7 a_42756_17049.t1 28.565
R15246 a_42756_17049.t2 a_42756_17049.n7 28.565
R15247 a_42756_17049.n3 a_42756_17049.t6 9.714
R15248 a_42756_17049.n3 a_42756_17049.n2 1.003
R15249 a_42756_17049.n6 a_42756_17049.n5 0.833
R15250 a_42756_17049.n5 a_42756_17049.n4 0.653
R15251 a_42756_17049.n7 a_42756_17049.n6 0.653
R15252 a_42756_17049.n5 a_42756_17049.n3 0.341
R15253 a_42756_17049.n6 a_42756_17049.n1 0.032
R15254 a_40011_18575.t6 a_40011_18575.t7 574.43
R15255 a_40011_18575.n1 a_40011_18575.t4 285.109
R15256 a_40011_18575.n3 a_40011_18575.n2 211.134
R15257 a_40011_18575.n4 a_40011_18575.n0 192.754
R15258 a_40011_18575.n1 a_40011_18575.t5 160.666
R15259 a_40011_18575.n2 a_40011_18575.t6 160.666
R15260 a_40011_18575.n2 a_40011_18575.n1 114.829
R15261 a_40011_18575.t2 a_40011_18575.n4 28.568
R15262 a_40011_18575.n0 a_40011_18575.t0 28.565
R15263 a_40011_18575.n0 a_40011_18575.t1 28.565
R15264 a_40011_18575.n3 a_40011_18575.t3 19.087
R15265 a_40011_18575.n4 a_40011_18575.n3 1.051
R15266 a_1681_1255.n1 a_1681_1255.t7 867.497
R15267 a_1681_1255.n1 a_1681_1255.t6 615.911
R15268 a_1681_1255.n0 a_1681_1255.t4 286.438
R15269 a_1681_1255.n0 a_1681_1255.t5 286.438
R15270 a_1681_1255.n4 a_1681_1255.n3 185.55
R15271 a_1681_1255.t7 a_1681_1255.n0 160.666
R15272 a_1681_1255.n2 a_1681_1255.n1 140.613
R15273 a_1681_1255.n3 a_1681_1255.t1 28.568
R15274 a_1681_1255.n4 a_1681_1255.t0 28.565
R15275 a_1681_1255.t2 a_1681_1255.n4 28.565
R15276 a_1681_1255.n2 a_1681_1255.t3 20.393
R15277 a_1681_1255.n3 a_1681_1255.n2 1.886
R15278 a_1156_1740.n0 a_1156_1740.t1 14.282
R15279 a_1156_1740.t0 a_1156_1740.n0 14.282
R15280 a_1156_1740.n0 a_1156_1740.n1 258.161
R15281 a_1156_1740.n1 a_1156_1740.n7 4.366
R15282 a_1156_1740.n7 a_1156_1740.n5 0.852
R15283 a_1156_1740.n5 a_1156_1740.n6 258.161
R15284 a_1156_1740.n6 a_1156_1740.t6 14.282
R15285 a_1156_1740.n6 a_1156_1740.t4 14.282
R15286 a_1156_1740.n5 a_1156_1740.t5 14.283
R15287 a_1156_1740.n7 a_1156_1740.n4 97.614
R15288 a_1156_1740.n4 a_1156_1740.t8 200.029
R15289 a_1156_1740.t8 a_1156_1740.n3 206.421
R15290 a_1156_1740.n3 a_1156_1740.t10 80.333
R15291 a_1156_1740.n3 a_1156_1740.t11 206.421
R15292 a_1156_1740.n4 a_1156_1740.t9 1527.4
R15293 a_1156_1740.t9 a_1156_1740.n2 657.379
R15294 a_1156_1740.n2 a_1156_1740.t7 8.7
R15295 a_1156_1740.n2 a_1156_1740.t2 8.7
R15296 a_1156_1740.n1 a_1156_1740.t3 14.283
R15297 a_70513_7422.t0 a_70513_7422.n9 104.259
R15298 a_70513_7422.n3 a_70513_7422.n1 77.784
R15299 a_70513_7422.n5 a_70513_7422.n3 77.456
R15300 a_70513_7422.n7 a_70513_7422.n5 77.456
R15301 a_70513_7422.n9 a_70513_7422.n7 75.815
R15302 a_70513_7422.n9 a_70513_7422.n8 167.433
R15303 a_70513_7422.n8 a_70513_7422.t4 14.282
R15304 a_70513_7422.n8 a_70513_7422.t5 14.282
R15305 a_70513_7422.n7 a_70513_7422.n6 89.977
R15306 a_70513_7422.n6 a_70513_7422.t8 14.282
R15307 a_70513_7422.n6 a_70513_7422.t6 14.282
R15308 a_70513_7422.n5 a_70513_7422.n4 89.977
R15309 a_70513_7422.n4 a_70513_7422.t10 14.282
R15310 a_70513_7422.n4 a_70513_7422.t7 14.282
R15311 a_70513_7422.n3 a_70513_7422.n2 89.977
R15312 a_70513_7422.n2 a_70513_7422.t9 14.282
R15313 a_70513_7422.n2 a_70513_7422.t11 14.282
R15314 a_70513_7422.n1 a_70513_7422.t3 104.259
R15315 a_70513_7422.n1 a_70513_7422.n0 167.433
R15316 a_70513_7422.n0 a_70513_7422.t1 14.282
R15317 a_70513_7422.n0 a_70513_7422.t2 14.282
R15318 a_55862_18700.n0 a_55862_18700.t8 214.335
R15319 a_55862_18700.t10 a_55862_18700.n0 214.335
R15320 a_55862_18700.n1 a_55862_18700.t10 143.851
R15321 a_55862_18700.n1 a_55862_18700.t7 135.658
R15322 a_55862_18700.n0 a_55862_18700.t9 80.333
R15323 a_55862_18700.n2 a_55862_18700.t5 28.565
R15324 a_55862_18700.n2 a_55862_18700.t3 28.565
R15325 a_55862_18700.n4 a_55862_18700.t4 28.565
R15326 a_55862_18700.n4 a_55862_18700.t2 28.565
R15327 a_55862_18700.n7 a_55862_18700.t1 28.565
R15328 a_55862_18700.t0 a_55862_18700.n7 28.565
R15329 a_55862_18700.n3 a_55862_18700.t6 9.714
R15330 a_55862_18700.n3 a_55862_18700.n2 1.003
R15331 a_55862_18700.n6 a_55862_18700.n5 0.833
R15332 a_55862_18700.n5 a_55862_18700.n4 0.653
R15333 a_55862_18700.n7 a_55862_18700.n6 0.653
R15334 a_55862_18700.n5 a_55862_18700.n3 0.341
R15335 a_55862_18700.n6 a_55862_18700.n1 0.032
R15336 a_508_8992.n1 a_508_8992.t7 990.34
R15337 a_508_8992.n1 a_508_8992.t4 408.211
R15338 a_508_8992.n0 a_508_8992.t6 286.438
R15339 a_508_8992.n0 a_508_8992.t5 286.438
R15340 a_508_8992.n4 a_508_8992.n3 185.55
R15341 a_508_8992.t7 a_508_8992.n0 160.666
R15342 a_508_8992.n3 a_508_8992.t1 28.568
R15343 a_508_8992.n4 a_508_8992.t0 28.565
R15344 a_508_8992.t2 a_508_8992.n4 28.565
R15345 a_508_8992.n2 a_508_8992.t3 23.417
R15346 a_508_8992.n2 a_508_8992.n1 12.315
R15347 a_508_8992.n3 a_508_8992.n2 0.002
R15348 a_67133_11394.n2 a_67133_11394.t7 214.335
R15349 a_67133_11394.t9 a_67133_11394.n2 214.335
R15350 a_67133_11394.n3 a_67133_11394.t9 143.851
R15351 a_67133_11394.n3 a_67133_11394.t8 135.658
R15352 a_67133_11394.n2 a_67133_11394.t10 80.333
R15353 a_67133_11394.n4 a_67133_11394.t4 28.565
R15354 a_67133_11394.n4 a_67133_11394.t3 28.565
R15355 a_67133_11394.n0 a_67133_11394.t6 28.565
R15356 a_67133_11394.n0 a_67133_11394.t5 28.565
R15357 a_67133_11394.n7 a_67133_11394.t2 28.565
R15358 a_67133_11394.t1 a_67133_11394.n7 28.565
R15359 a_67133_11394.n1 a_67133_11394.t0 9.714
R15360 a_67133_11394.n1 a_67133_11394.n0 1.003
R15361 a_67133_11394.n6 a_67133_11394.n5 0.833
R15362 a_67133_11394.n5 a_67133_11394.n4 0.653
R15363 a_67133_11394.n7 a_67133_11394.n6 0.653
R15364 a_67133_11394.n6 a_67133_11394.n1 0.341
R15365 a_67133_11394.n5 a_67133_11394.n3 0.032
R15366 a_44399_2324.n6 a_44399_2324.n5 501.28
R15367 a_44399_2324.t10 a_44399_2324.t11 437.233
R15368 a_44399_2324.t14 a_44399_2324.t8 415.315
R15369 a_44399_2324.t4 a_44399_2324.n3 313.873
R15370 a_44399_2324.n5 a_44399_2324.t6 294.986
R15371 a_44399_2324.n2 a_44399_2324.t16 272.288
R15372 a_44399_2324.n6 a_44399_2324.t12 236.01
R15373 a_44399_2324.n9 a_44399_2324.t10 216.627
R15374 a_44399_2324.n7 a_44399_2324.t14 216.111
R15375 a_44399_2324.n8 a_44399_2324.t7 214.686
R15376 a_44399_2324.t11 a_44399_2324.n8 214.686
R15377 a_44399_2324.n1 a_44399_2324.t18 214.335
R15378 a_44399_2324.t8 a_44399_2324.n1 214.335
R15379 a_44399_2324.n11 a_44399_2324.n0 192.754
R15380 a_44399_2324.n4 a_44399_2324.t4 190.152
R15381 a_44399_2324.n4 a_44399_2324.t17 190.152
R15382 a_44399_2324.n2 a_44399_2324.t9 160.666
R15383 a_44399_2324.n3 a_44399_2324.t19 160.666
R15384 a_44399_2324.n7 a_44399_2324.n6 148.428
R15385 a_44399_2324.n5 a_44399_2324.t15 110.859
R15386 a_44399_2324.n10 a_44399_2324.n9 102.569
R15387 a_44399_2324.n3 a_44399_2324.n2 96.129
R15388 a_44399_2324.n8 a_44399_2324.t13 80.333
R15389 a_44399_2324.n1 a_44399_2324.t5 80.333
R15390 a_44399_2324.t12 a_44399_2324.n4 80.333
R15391 a_44399_2324.t2 a_44399_2324.n11 28.568
R15392 a_44399_2324.n0 a_44399_2324.t0 28.565
R15393 a_44399_2324.n0 a_44399_2324.t1 28.565
R15394 a_44399_2324.n10 a_44399_2324.t3 18.523
R15395 a_44399_2324.n9 a_44399_2324.n7 2.923
R15396 a_44399_2324.n11 a_44399_2324.n10 1.167
R15397 a_41999_6796.n1 a_41999_6796.t7 318.922
R15398 a_41999_6796.n0 a_41999_6796.t4 274.739
R15399 a_41999_6796.n0 a_41999_6796.t5 274.739
R15400 a_41999_6796.n1 a_41999_6796.t6 269.116
R15401 a_41999_6796.t7 a_41999_6796.n0 179.946
R15402 a_41999_6796.n2 a_41999_6796.n1 105.178
R15403 a_41999_6796.n3 a_41999_6796.t2 29.444
R15404 a_41999_6796.n4 a_41999_6796.t1 28.565
R15405 a_41999_6796.t0 a_41999_6796.n4 28.565
R15406 a_41999_6796.n2 a_41999_6796.t3 18.145
R15407 a_41999_6796.n3 a_41999_6796.n2 2.878
R15408 a_41999_6796.n4 a_41999_6796.n3 0.764
R15409 a_41705_6822.t0 a_41705_6822.n0 14.282
R15410 a_41705_6822.n0 a_41705_6822.t1 14.282
R15411 a_41705_6822.n0 a_41705_6822.n14 90.436
R15412 a_41705_6822.n10 a_41705_6822.n13 50.575
R15413 a_41705_6822.n14 a_41705_6822.n10 74.302
R15414 a_41705_6822.n13 a_41705_6822.n12 157.665
R15415 a_41705_6822.n12 a_41705_6822.t6 8.7
R15416 a_41705_6822.n12 a_41705_6822.t3 8.7
R15417 a_41705_6822.n13 a_41705_6822.n11 122.999
R15418 a_41705_6822.n11 a_41705_6822.t4 14.282
R15419 a_41705_6822.n11 a_41705_6822.t7 14.282
R15420 a_41705_6822.n10 a_41705_6822.n9 90.416
R15421 a_41705_6822.n9 a_41705_6822.t5 14.282
R15422 a_41705_6822.n9 a_41705_6822.t2 14.282
R15423 a_41705_6822.n1 a_41705_6822.t12 220.285
R15424 a_41705_6822.n14 a_41705_6822.n1 3509.5
R15425 a_41705_6822.n1 a_41705_6822.n8 61.538
R15426 a_41705_6822.n8 a_41705_6822.n3 465.933
R15427 a_41705_6822.n8 a_41705_6822.n7 163.88
R15428 a_41705_6822.n7 a_41705_6822.n6 6.615
R15429 a_41705_6822.n6 a_41705_6822.t17 93.989
R15430 a_41705_6822.n7 a_41705_6822.n5 97.816
R15431 a_41705_6822.n5 a_41705_6822.t19 80.333
R15432 a_41705_6822.n5 a_41705_6822.t8 394.151
R15433 a_41705_6822.t8 a_41705_6822.n4 269.523
R15434 a_41705_6822.n4 a_41705_6822.t9 160.666
R15435 a_41705_6822.n4 a_41705_6822.t13 269.523
R15436 a_41705_6822.n6 a_41705_6822.t10 198.043
R15437 a_41705_6822.n3 a_41705_6822.t18 294.653
R15438 a_41705_6822.n3 a_41705_6822.t11 111.663
R15439 a_41705_6822.t12 a_41705_6822.t14 415.315
R15440 a_41705_6822.t14 a_41705_6822.n2 214.335
R15441 a_41705_6822.n2 a_41705_6822.t15 80.333
R15442 a_41705_6822.n2 a_41705_6822.t16 214.335
R15443 a_41587_6822.t0 a_41587_6822.n0 14.282
R15444 a_41587_6822.n0 a_41587_6822.t1 14.282
R15445 a_41587_6822.n1 a_41587_6822.n9 0.001
R15446 a_41587_6822.n0 a_41587_6822.n1 267.767
R15447 a_41587_6822.n9 a_41587_6822.t8 14.282
R15448 a_41587_6822.n9 a_41587_6822.t2 14.282
R15449 a_41587_6822.n1 a_41587_6822.n7 0.669
R15450 a_41587_6822.n7 a_41587_6822.n8 1.511
R15451 a_41587_6822.n8 a_41587_6822.t7 14.282
R15452 a_41587_6822.n8 a_41587_6822.t6 14.282
R15453 a_41587_6822.n7 a_41587_6822.n6 0.227
R15454 a_41587_6822.n6 a_41587_6822.n3 0.575
R15455 a_41587_6822.n6 a_41587_6822.n5 0.2
R15456 a_41587_6822.n5 a_41587_6822.t4 16.058
R15457 a_41587_6822.n5 a_41587_6822.n4 0.999
R15458 a_41587_6822.n4 a_41587_6822.t5 14.282
R15459 a_41587_6822.n4 a_41587_6822.t3 14.282
R15460 a_41587_6822.n3 a_41587_6822.n2 0.999
R15461 a_41587_6822.n2 a_41587_6822.t11 14.282
R15462 a_41587_6822.n2 a_41587_6822.t10 14.282
R15463 a_41587_6822.n3 a_41587_6822.t9 16.058
R15464 a_30645_3831.n0 a_30645_3831.t3 14.282
R15465 a_30645_3831.t1 a_30645_3831.n0 14.282
R15466 a_30645_3831.n0 a_30645_3831.n16 90.436
R15467 a_30645_3831.n16 a_30645_3831.n2 74.302
R15468 a_30645_3831.n2 a_30645_3831.n4 50.575
R15469 a_30645_3831.n4 a_30645_3831.n5 110.084
R15470 a_30645_3831.n16 a_30645_3831.n6 213.889
R15471 a_30645_3831.n6 a_30645_3831.n8 16.411
R15472 a_30645_3831.n8 a_30645_3831.t8 198.921
R15473 a_30645_3831.t8 a_30645_3831.t16 415.315
R15474 a_30645_3831.t16 a_30645_3831.n15 214.335
R15475 a_30645_3831.n15 a_30645_3831.t14 80.333
R15476 a_30645_3831.n15 a_30645_3831.t13 214.335
R15477 a_30645_3831.n8 a_30645_3831.n14 861.987
R15478 a_30645_3831.n14 a_30645_3831.n9 560.726
R15479 a_30645_3831.n14 a_30645_3831.n13 65.07
R15480 a_30645_3831.n13 a_30645_3831.n12 6.615
R15481 a_30645_3831.n12 a_30645_3831.t19 93.989
R15482 a_30645_3831.n12 a_30645_3831.t20 198.043
R15483 a_30645_3831.n13 a_30645_3831.n11 97.816
R15484 a_30645_3831.n11 a_30645_3831.t18 80.333
R15485 a_30645_3831.n11 a_30645_3831.t23 394.151
R15486 a_30645_3831.t23 a_30645_3831.n10 269.523
R15487 a_30645_3831.n10 a_30645_3831.t22 160.666
R15488 a_30645_3831.n10 a_30645_3831.t21 269.523
R15489 a_30645_3831.n9 a_30645_3831.t15 294.653
R15490 a_30645_3831.n9 a_30645_3831.t10 111.663
R15491 a_30645_3831.n6 a_30645_3831.t17 217.716
R15492 a_30645_3831.t17 a_30645_3831.t12 415.315
R15493 a_30645_3831.t12 a_30645_3831.n7 214.335
R15494 a_30645_3831.n7 a_30645_3831.t11 80.333
R15495 a_30645_3831.n7 a_30645_3831.t9 214.335
R15496 a_30645_3831.n5 a_30645_3831.t4 14.282
R15497 a_30645_3831.n5 a_30645_3831.t5 14.282
R15498 a_30645_3831.n4 a_30645_3831.n3 157.665
R15499 a_30645_3831.n3 a_30645_3831.t0 8.7
R15500 a_30645_3831.n3 a_30645_3831.t6 8.7
R15501 a_30645_3831.n2 a_30645_3831.n1 90.416
R15502 a_30645_3831.n1 a_30645_3831.t2 14.282
R15503 a_30645_3831.n1 a_30645_3831.t7 14.282
R15504 a_63010_16442.t0 a_63010_16442.t1 17.4
R15505 a_47282_17937.t8 a_47282_17937.n2 404.877
R15506 a_47282_17937.n1 a_47282_17937.t5 210.902
R15507 a_47282_17937.n3 a_47282_17937.t8 136.949
R15508 a_47282_17937.n2 a_47282_17937.n1 107.801
R15509 a_47282_17937.n1 a_47282_17937.t6 80.333
R15510 a_47282_17937.n2 a_47282_17937.t7 80.333
R15511 a_47282_17937.n0 a_47282_17937.t1 17.4
R15512 a_47282_17937.n0 a_47282_17937.t0 17.4
R15513 a_47282_17937.n4 a_47282_17937.t4 15.032
R15514 a_47282_17937.n5 a_47282_17937.t3 14.282
R15515 a_47282_17937.t2 a_47282_17937.n5 14.282
R15516 a_47282_17937.n5 a_47282_17937.n4 1.65
R15517 a_47282_17937.n3 a_47282_17937.n0 0.657
R15518 a_47282_17937.n4 a_47282_17937.n3 0.614
R15519 a_46215_18571.t6 a_46215_18571.t7 800.071
R15520 a_46215_18571.n3 a_46215_18571.n2 672.95
R15521 a_46215_18571.n1 a_46215_18571.t4 285.109
R15522 a_46215_18571.n2 a_46215_18571.t6 193.602
R15523 a_46215_18571.n1 a_46215_18571.t5 160.666
R15524 a_46215_18571.n2 a_46215_18571.n1 91.507
R15525 a_46215_18571.n0 a_46215_18571.t0 28.57
R15526 a_46215_18571.n4 a_46215_18571.t1 28.565
R15527 a_46215_18571.t2 a_46215_18571.n4 28.565
R15528 a_46215_18571.n0 a_46215_18571.t3 17.638
R15529 a_46215_18571.n4 a_46215_18571.n3 0.693
R15530 a_46215_18571.n3 a_46215_18571.n0 0.597
R15531 a_16859_20723.n2 a_16859_20723.t4 448.381
R15532 a_16859_20723.n1 a_16859_20723.t6 286.438
R15533 a_16859_20723.n1 a_16859_20723.t5 286.438
R15534 a_16859_20723.n0 a_16859_20723.t7 247.69
R15535 a_16859_20723.n4 a_16859_20723.n3 182.117
R15536 a_16859_20723.t4 a_16859_20723.n1 160.666
R15537 a_16859_20723.n3 a_16859_20723.t0 28.568
R15538 a_16859_20723.n4 a_16859_20723.t1 28.565
R15539 a_16859_20723.t2 a_16859_20723.n4 28.565
R15540 a_16859_20723.n0 a_16859_20723.t3 18.127
R15541 a_16859_20723.n2 a_16859_20723.n0 4.036
R15542 a_16859_20723.n3 a_16859_20723.n2 0.937
R15543 a_15680_20866.n0 a_15680_20866.t2 14.282
R15544 a_15680_20866.t1 a_15680_20866.n0 14.282
R15545 a_15680_20866.n0 a_15680_20866.n1 258.161
R15546 a_15680_20866.n1 a_15680_20866.n5 0.852
R15547 a_15680_20866.n5 a_15680_20866.n6 4.366
R15548 a_15680_20866.n6 a_15680_20866.n7 258.161
R15549 a_15680_20866.n7 a_15680_20866.t6 14.282
R15550 a_15680_20866.n7 a_15680_20866.t4 14.282
R15551 a_15680_20866.n6 a_15680_20866.t7 14.283
R15552 a_15680_20866.n5 a_15680_20866.n4 97.614
R15553 a_15680_20866.n4 a_15680_20866.t8 200.029
R15554 a_15680_20866.t8 a_15680_20866.n3 206.421
R15555 a_15680_20866.n3 a_15680_20866.t10 80.333
R15556 a_15680_20866.n3 a_15680_20866.t11 206.421
R15557 a_15680_20866.n4 a_15680_20866.t9 1527.4
R15558 a_15680_20866.t9 a_15680_20866.n2 657.379
R15559 a_15680_20866.n2 a_15680_20866.t5 8.7
R15560 a_15680_20866.n2 a_15680_20866.t0 8.7
R15561 a_15680_20866.n1 a_15680_20866.t3 14.283
R15562 a_16213_21596.n3 a_16213_21596.n2 167.433
R15563 a_16213_21596.n7 a_16213_21596.n6 167.433
R15564 a_16213_21596.n3 a_16213_21596.t8 104.259
R15565 a_16213_21596.n7 a_16213_21596.t3 104.259
R15566 a_16213_21596.n4 a_16213_21596.n1 89.977
R15567 a_16213_21596.n5 a_16213_21596.n0 89.977
R15568 a_16213_21596.n9 a_16213_21596.n8 89.977
R15569 a_16213_21596.n8 a_16213_21596.n7 77.784
R15570 a_16213_21596.n5 a_16213_21596.n4 77.456
R15571 a_16213_21596.n8 a_16213_21596.n5 77.456
R15572 a_16213_21596.n4 a_16213_21596.n3 75.815
R15573 a_16213_21596.n2 a_16213_21596.t6 14.282
R15574 a_16213_21596.n2 a_16213_21596.t7 14.282
R15575 a_16213_21596.n1 a_16213_21596.t10 14.282
R15576 a_16213_21596.n1 a_16213_21596.t11 14.282
R15577 a_16213_21596.n0 a_16213_21596.t9 14.282
R15578 a_16213_21596.n0 a_16213_21596.t0 14.282
R15579 a_16213_21596.n6 a_16213_21596.t4 14.282
R15580 a_16213_21596.n6 a_16213_21596.t5 14.282
R15581 a_16213_21596.n9 a_16213_21596.t1 14.282
R15582 a_16213_21596.t2 a_16213_21596.n9 14.282
R15583 a_20588_7655.t0 a_20588_7655.t1 17.4
R15584 a_19464_8258.n0 a_19464_8258.t2 14.282
R15585 a_19464_8258.t1 a_19464_8258.n0 14.282
R15586 a_19464_8258.n0 a_19464_8258.n1 258.161
R15587 a_19464_8258.n1 a_19464_8258.n5 0.852
R15588 a_19464_8258.n5 a_19464_8258.n6 4.366
R15589 a_19464_8258.n6 a_19464_8258.n7 258.161
R15590 a_19464_8258.n7 a_19464_8258.t5 14.282
R15591 a_19464_8258.n7 a_19464_8258.t6 14.282
R15592 a_19464_8258.n6 a_19464_8258.t7 14.283
R15593 a_19464_8258.n5 a_19464_8258.n4 97.614
R15594 a_19464_8258.n4 a_19464_8258.t10 200.029
R15595 a_19464_8258.t10 a_19464_8258.n3 206.421
R15596 a_19464_8258.n3 a_19464_8258.t8 80.333
R15597 a_19464_8258.n3 a_19464_8258.t11 206.421
R15598 a_19464_8258.n4 a_19464_8258.t9 1527.4
R15599 a_19464_8258.t9 a_19464_8258.n2 657.379
R15600 a_19464_8258.n2 a_19464_8258.t4 8.7
R15601 a_19464_8258.n2 a_19464_8258.t0 8.7
R15602 a_19464_8258.n1 a_19464_8258.t3 14.283
R15603 a_19357_21596.n0 a_19357_21596.t5 14.282
R15604 a_19357_21596.t0 a_19357_21596.n0 14.282
R15605 a_19357_21596.n0 a_19357_21596.n9 89.977
R15606 a_19357_21596.n6 a_19357_21596.n7 77.784
R15607 a_19357_21596.n9 a_19357_21596.n6 77.456
R15608 a_19357_21596.n9 a_19357_21596.n4 77.456
R15609 a_19357_21596.n4 a_19357_21596.n2 75.815
R15610 a_19357_21596.n7 a_19357_21596.n8 167.433
R15611 a_19357_21596.n8 a_19357_21596.t9 14.282
R15612 a_19357_21596.n8 a_19357_21596.t10 14.282
R15613 a_19357_21596.n7 a_19357_21596.t11 104.259
R15614 a_19357_21596.n6 a_19357_21596.n5 89.977
R15615 a_19357_21596.n5 a_19357_21596.t4 14.282
R15616 a_19357_21596.n5 a_19357_21596.t3 14.282
R15617 a_19357_21596.n4 a_19357_21596.n3 89.977
R15618 a_19357_21596.n3 a_19357_21596.t1 14.282
R15619 a_19357_21596.n3 a_19357_21596.t2 14.282
R15620 a_19357_21596.n2 a_19357_21596.t8 104.259
R15621 a_19357_21596.n2 a_19357_21596.n1 167.433
R15622 a_19357_21596.n1 a_19357_21596.t7 14.282
R15623 a_19357_21596.n1 a_19357_21596.t6 14.282
R15624 a_37848_2326.n6 a_37848_2326.n5 501.28
R15625 a_37848_2326.t16 a_37848_2326.t18 437.233
R15626 a_37848_2326.t7 a_37848_2326.t13 415.315
R15627 a_37848_2326.t19 a_37848_2326.n3 313.873
R15628 a_37848_2326.n5 a_37848_2326.t8 294.986
R15629 a_37848_2326.n2 a_37848_2326.t5 272.288
R15630 a_37848_2326.n6 a_37848_2326.t11 236.01
R15631 a_37848_2326.n9 a_37848_2326.t16 216.627
R15632 a_37848_2326.n7 a_37848_2326.t7 216.111
R15633 a_37848_2326.n8 a_37848_2326.t9 214.686
R15634 a_37848_2326.t18 a_37848_2326.n8 214.686
R15635 a_37848_2326.n1 a_37848_2326.t10 214.335
R15636 a_37848_2326.t13 a_37848_2326.n1 214.335
R15637 a_37848_2326.n4 a_37848_2326.t19 190.152
R15638 a_37848_2326.n4 a_37848_2326.t4 190.152
R15639 a_37848_2326.n2 a_37848_2326.t15 160.666
R15640 a_37848_2326.n3 a_37848_2326.t12 160.666
R15641 a_37848_2326.n7 a_37848_2326.n6 148.428
R15642 a_37848_2326.n5 a_37848_2326.t6 110.859
R15643 a_37848_2326.n3 a_37848_2326.n2 96.129
R15644 a_37848_2326.n8 a_37848_2326.t17 80.333
R15645 a_37848_2326.n1 a_37848_2326.t14 80.333
R15646 a_37848_2326.t11 a_37848_2326.n4 80.333
R15647 a_37848_2326.n0 a_37848_2326.t1 28.57
R15648 a_37848_2326.n11 a_37848_2326.t3 28.565
R15649 a_37848_2326.t0 a_37848_2326.n11 28.565
R15650 a_37848_2326.n0 a_37848_2326.t2 17.638
R15651 a_37848_2326.n10 a_37848_2326.n9 7.04
R15652 a_37848_2326.n9 a_37848_2326.n7 2.923
R15653 a_37848_2326.n11 a_37848_2326.n10 0.69
R15654 a_37848_2326.n10 a_37848_2326.n0 0.6
R15655 a_41991_1016.n1 a_41991_1016.t7 318.922
R15656 a_41991_1016.n0 a_41991_1016.t5 274.739
R15657 a_41991_1016.n0 a_41991_1016.t6 274.739
R15658 a_41991_1016.n1 a_41991_1016.t4 269.116
R15659 a_41991_1016.t7 a_41991_1016.n0 179.946
R15660 a_41991_1016.n2 a_41991_1016.n1 105.178
R15661 a_41991_1016.t2 a_41991_1016.n4 29.444
R15662 a_41991_1016.n3 a_41991_1016.t1 28.565
R15663 a_41991_1016.n3 a_41991_1016.t0 28.565
R15664 a_41991_1016.n2 a_41991_1016.t3 18.145
R15665 a_41991_1016.n4 a_41991_1016.n2 2.878
R15666 a_41991_1016.n4 a_41991_1016.n3 0.764
R15667 a_54903_1041.t0 a_54903_1041.n0 14.282
R15668 a_54903_1041.n0 a_54903_1041.t2 14.282
R15669 a_54903_1041.n0 a_54903_1041.n15 90.436
R15670 a_54903_1041.n11 a_54903_1041.n14 50.575
R15671 a_54903_1041.n15 a_54903_1041.n11 74.302
R15672 a_54903_1041.n14 a_54903_1041.n13 157.665
R15673 a_54903_1041.n13 a_54903_1041.t6 8.7
R15674 a_54903_1041.n13 a_54903_1041.t7 8.7
R15675 a_54903_1041.n14 a_54903_1041.n12 122.999
R15676 a_54903_1041.n12 a_54903_1041.t3 14.282
R15677 a_54903_1041.n12 a_54903_1041.t5 14.282
R15678 a_54903_1041.n11 a_54903_1041.n10 90.416
R15679 a_54903_1041.n10 a_54903_1041.t4 14.282
R15680 a_54903_1041.n10 a_54903_1041.t1 14.282
R15681 a_54903_1041.n15 a_54903_1041.n9 220.49
R15682 a_54903_1041.n9 a_54903_1041.n2 2.599
R15683 a_54903_1041.n2 a_54903_1041.t10 218.628
R15684 a_54903_1041.t10 a_54903_1041.t15 437.233
R15685 a_54903_1041.t15 a_54903_1041.n8 214.686
R15686 a_54903_1041.n8 a_54903_1041.t12 80.333
R15687 a_54903_1041.n8 a_54903_1041.t17 214.686
R15688 a_54903_1041.n2 a_54903_1041.n3 14.9
R15689 a_54903_1041.n3 a_54903_1041.n7 535.449
R15690 a_54903_1041.n7 a_54903_1041.t22 294.986
R15691 a_54903_1041.n7 a_54903_1041.t23 110.859
R15692 a_54903_1041.n3 a_54903_1041.t21 245.184
R15693 a_54903_1041.t21 a_54903_1041.n6 80.333
R15694 a_54903_1041.n6 a_54903_1041.t18 190.152
R15695 a_54903_1041.n6 a_54903_1041.t16 190.152
R15696 a_54903_1041.t16 a_54903_1041.n5 313.873
R15697 a_54903_1041.n5 a_54903_1041.t19 160.666
R15698 a_54903_1041.n5 a_54903_1041.n4 96.129
R15699 a_54903_1041.n4 a_54903_1041.t11 160.666
R15700 a_54903_1041.n4 a_54903_1041.t13 272.288
R15701 a_54903_1041.n9 a_54903_1041.t14 217.024
R15702 a_54903_1041.t14 a_54903_1041.t9 437.233
R15703 a_54903_1041.t9 a_54903_1041.n1 214.686
R15704 a_54903_1041.n1 a_54903_1041.t20 80.333
R15705 a_54903_1041.n1 a_54903_1041.t8 214.686
R15706 a_57722_4002.n4 a_57722_4002.t9 214.335
R15707 a_57722_4002.t10 a_57722_4002.n4 214.335
R15708 a_57722_4002.n5 a_57722_4002.t10 143.851
R15709 a_57722_4002.n5 a_57722_4002.t7 135.658
R15710 a_57722_4002.n4 a_57722_4002.t8 80.333
R15711 a_57722_4002.n0 a_57722_4002.t4 28.565
R15712 a_57722_4002.n0 a_57722_4002.t6 28.565
R15713 a_57722_4002.n2 a_57722_4002.t1 28.565
R15714 a_57722_4002.n2 a_57722_4002.t5 28.565
R15715 a_57722_4002.n7 a_57722_4002.t2 28.565
R15716 a_57722_4002.t0 a_57722_4002.n7 28.565
R15717 a_57722_4002.n1 a_57722_4002.t3 9.714
R15718 a_57722_4002.n1 a_57722_4002.n0 1.003
R15719 a_57722_4002.n6 a_57722_4002.n3 0.833
R15720 a_57722_4002.n3 a_57722_4002.n2 0.653
R15721 a_57722_4002.n7 a_57722_4002.n6 0.653
R15722 a_57722_4002.n3 a_57722_4002.n1 0.341
R15723 a_57722_4002.n6 a_57722_4002.n5 0.032
R15724 a_29954_7911.t0 a_29954_7911.n0 14.282
R15725 a_29954_7911.n0 a_29954_7911.t1 14.282
R15726 a_29954_7911.n1 a_29954_7911.n9 0.001
R15727 a_29954_7911.n0 a_29954_7911.n1 267.767
R15728 a_29954_7911.n9 a_29954_7911.t9 14.282
R15729 a_29954_7911.n9 a_29954_7911.t3 14.282
R15730 a_29954_7911.n1 a_29954_7911.n7 0.669
R15731 a_29954_7911.n7 a_29954_7911.n8 1.511
R15732 a_29954_7911.n8 a_29954_7911.t2 14.282
R15733 a_29954_7911.n8 a_29954_7911.t4 14.282
R15734 a_29954_7911.n7 a_29954_7911.n6 0.227
R15735 a_29954_7911.n6 a_29954_7911.n5 0.2
R15736 a_29954_7911.n6 a_29954_7911.n3 0.575
R15737 a_29954_7911.n5 a_29954_7911.t5 16.058
R15738 a_29954_7911.n5 a_29954_7911.n4 0.999
R15739 a_29954_7911.n4 a_29954_7911.t6 14.282
R15740 a_29954_7911.n4 a_29954_7911.t7 14.282
R15741 a_29954_7911.n3 a_29954_7911.n2 0.999
R15742 a_29954_7911.n2 a_29954_7911.t8 14.282
R15743 a_29954_7911.n2 a_29954_7911.t10 14.282
R15744 a_29954_7911.n3 a_29954_7911.t11 16.058
R15745 a_19563_6043.n1 a_19563_6043.t6 318.922
R15746 a_19563_6043.n0 a_19563_6043.t4 274.739
R15747 a_19563_6043.n0 a_19563_6043.t5 274.739
R15748 a_19563_6043.n1 a_19563_6043.t7 269.116
R15749 a_19563_6043.t6 a_19563_6043.n0 179.946
R15750 a_19563_6043.n2 a_19563_6043.n1 107.263
R15751 a_19563_6043.n3 a_19563_6043.t3 29.444
R15752 a_19563_6043.t0 a_19563_6043.n4 28.565
R15753 a_19563_6043.n4 a_19563_6043.t2 28.565
R15754 a_19563_6043.n2 a_19563_6043.t1 18.145
R15755 a_19563_6043.n3 a_19563_6043.n2 2.878
R15756 a_19563_6043.n4 a_19563_6043.n3 0.764
R15757 a_57730_9870.n4 a_57730_9870.t9 214.335
R15758 a_57730_9870.t8 a_57730_9870.n4 214.335
R15759 a_57730_9870.n5 a_57730_9870.t8 143.851
R15760 a_57730_9870.n5 a_57730_9870.t10 135.658
R15761 a_57730_9870.n4 a_57730_9870.t7 80.333
R15762 a_57730_9870.n0 a_57730_9870.t2 28.565
R15763 a_57730_9870.n0 a_57730_9870.t0 28.565
R15764 a_57730_9870.n2 a_57730_9870.t6 28.565
R15765 a_57730_9870.n2 a_57730_9870.t1 28.565
R15766 a_57730_9870.t4 a_57730_9870.n7 28.565
R15767 a_57730_9870.n7 a_57730_9870.t5 28.565
R15768 a_57730_9870.n1 a_57730_9870.t3 9.714
R15769 a_57730_9870.n1 a_57730_9870.n0 1.003
R15770 a_57730_9870.n6 a_57730_9870.n3 0.833
R15771 a_57730_9870.n3 a_57730_9870.n2 0.653
R15772 a_57730_9870.n7 a_57730_9870.n6 0.653
R15773 a_57730_9870.n3 a_57730_9870.n1 0.341
R15774 a_57730_9870.n6 a_57730_9870.n5 0.032
R15775 a_58320_9433.t6 a_58320_9433.t5 800.071
R15776 a_58320_9433.n2 a_58320_9433.n1 659.097
R15777 a_58320_9433.n0 a_58320_9433.t7 285.109
R15778 a_58320_9433.n1 a_58320_9433.t6 193.602
R15779 a_58320_9433.n4 a_58320_9433.n3 192.754
R15780 a_58320_9433.n0 a_58320_9433.t4 160.666
R15781 a_58320_9433.n1 a_58320_9433.n0 91.507
R15782 a_58320_9433.n3 a_58320_9433.t0 28.568
R15783 a_58320_9433.t2 a_58320_9433.n4 28.565
R15784 a_58320_9433.n4 a_58320_9433.t1 28.565
R15785 a_58320_9433.n2 a_58320_9433.t3 19.061
R15786 a_58320_9433.n3 a_58320_9433.n2 1.005
R15787 a_12478_20862.n0 a_12478_20862.t2 14.282
R15788 a_12478_20862.t1 a_12478_20862.n0 14.282
R15789 a_12478_20862.n0 a_12478_20862.n1 258.161
R15790 a_12478_20862.n1 a_12478_20862.n5 0.852
R15791 a_12478_20862.n5 a_12478_20862.n6 4.366
R15792 a_12478_20862.n6 a_12478_20862.n7 258.161
R15793 a_12478_20862.n7 a_12478_20862.t5 14.282
R15794 a_12478_20862.n7 a_12478_20862.t6 14.282
R15795 a_12478_20862.n6 a_12478_20862.t7 14.283
R15796 a_12478_20862.n5 a_12478_20862.n4 97.614
R15797 a_12478_20862.n4 a_12478_20862.t10 200.029
R15798 a_12478_20862.t10 a_12478_20862.n3 206.421
R15799 a_12478_20862.n3 a_12478_20862.t11 80.333
R15800 a_12478_20862.n3 a_12478_20862.t8 206.421
R15801 a_12478_20862.n4 a_12478_20862.t9 1527.4
R15802 a_12478_20862.t9 a_12478_20862.n2 657.379
R15803 a_12478_20862.n2 a_12478_20862.t4 8.7
R15804 a_12478_20862.n2 a_12478_20862.t0 8.7
R15805 a_12478_20862.n1 a_12478_20862.t3 14.283
R15806 a_13011_21592.n0 a_13011_21592.t0 14.282
R15807 a_13011_21592.t6 a_13011_21592.n0 14.282
R15808 a_13011_21592.n0 a_13011_21592.n9 89.977
R15809 a_13011_21592.n6 a_13011_21592.n7 77.784
R15810 a_13011_21592.n9 a_13011_21592.n6 77.456
R15811 a_13011_21592.n9 a_13011_21592.n4 77.456
R15812 a_13011_21592.n4 a_13011_21592.n2 75.815
R15813 a_13011_21592.n7 a_13011_21592.n8 167.433
R15814 a_13011_21592.n8 a_13011_21592.t5 14.282
R15815 a_13011_21592.n8 a_13011_21592.t4 14.282
R15816 a_13011_21592.n7 a_13011_21592.t3 104.259
R15817 a_13011_21592.n6 a_13011_21592.n5 89.977
R15818 a_13011_21592.n5 a_13011_21592.t2 14.282
R15819 a_13011_21592.n5 a_13011_21592.t1 14.282
R15820 a_13011_21592.n4 a_13011_21592.n3 89.977
R15821 a_13011_21592.n3 a_13011_21592.t7 14.282
R15822 a_13011_21592.n3 a_13011_21592.t8 14.282
R15823 a_13011_21592.n2 a_13011_21592.t11 104.259
R15824 a_13011_21592.n2 a_13011_21592.n1 167.433
R15825 a_13011_21592.n1 a_13011_21592.t10 14.282
R15826 a_13011_21592.n1 a_13011_21592.t9 14.282
R15827 a_40799_18571.t4 a_40799_18571.t6 800.071
R15828 a_40799_18571.n2 a_40799_18571.n1 659.095
R15829 a_40799_18571.n0 a_40799_18571.t7 285.109
R15830 a_40799_18571.n1 a_40799_18571.t4 193.602
R15831 a_40799_18571.n4 a_40799_18571.n3 192.754
R15832 a_40799_18571.n0 a_40799_18571.t5 160.666
R15833 a_40799_18571.n1 a_40799_18571.n0 91.507
R15834 a_40799_18571.n3 a_40799_18571.t0 28.568
R15835 a_40799_18571.n4 a_40799_18571.t1 28.565
R15836 a_40799_18571.t2 a_40799_18571.n4 28.565
R15837 a_40799_18571.n2 a_40799_18571.t3 19.063
R15838 a_40799_18571.n3 a_40799_18571.n2 1.005
R15839 a_30154_7310.n1 a_30154_7310.t7 318.119
R15840 a_30154_7310.n1 a_30154_7310.t5 269.919
R15841 a_30154_7310.n0 a_30154_7310.t4 267.853
R15842 a_30154_7310.n0 a_30154_7310.t6 267.853
R15843 a_30154_7310.t7 a_30154_7310.n0 160.666
R15844 a_30154_7310.n2 a_30154_7310.n1 107.263
R15845 a_30154_7310.n3 a_30154_7310.t2 29.444
R15846 a_30154_7310.t0 a_30154_7310.n4 28.565
R15847 a_30154_7310.n4 a_30154_7310.t3 28.565
R15848 a_30154_7310.n2 a_30154_7310.t1 18.145
R15849 a_30154_7310.n3 a_30154_7310.n2 2.878
R15850 a_30154_7310.n4 a_30154_7310.n3 0.764
R15851 a_30647_7968.n0 a_30647_7968.t5 14.282
R15852 a_30647_7968.t2 a_30647_7968.n0 14.282
R15853 a_30647_7968.n0 a_30647_7968.n16 90.416
R15854 a_30647_7968.n16 a_30647_7968.n2 74.302
R15855 a_30647_7968.n16 a_30647_7968.n4 50.575
R15856 a_30647_7968.n4 a_30647_7968.n5 110.084
R15857 a_30647_7968.n2 a_30647_7968.n6 210.799
R15858 a_30647_7968.n6 a_30647_7968.n8 16.411
R15859 a_30647_7968.n8 a_30647_7968.t14 198.921
R15860 a_30647_7968.t14 a_30647_7968.t15 415.315
R15861 a_30647_7968.t15 a_30647_7968.n15 214.335
R15862 a_30647_7968.n15 a_30647_7968.t22 80.333
R15863 a_30647_7968.n15 a_30647_7968.t23 214.335
R15864 a_30647_7968.n8 a_30647_7968.n14 861.987
R15865 a_30647_7968.n14 a_30647_7968.n9 560.726
R15866 a_30647_7968.n14 a_30647_7968.n13 65.07
R15867 a_30647_7968.n13 a_30647_7968.n12 6.615
R15868 a_30647_7968.n12 a_30647_7968.t8 93.989
R15869 a_30647_7968.n13 a_30647_7968.n11 97.816
R15870 a_30647_7968.n11 a_30647_7968.t9 80.333
R15871 a_30647_7968.n11 a_30647_7968.t12 394.151
R15872 a_30647_7968.t12 a_30647_7968.n10 269.523
R15873 a_30647_7968.n10 a_30647_7968.t13 160.666
R15874 a_30647_7968.n10 a_30647_7968.t16 269.523
R15875 a_30647_7968.n12 a_30647_7968.t20 198.043
R15876 a_30647_7968.n9 a_30647_7968.t11 294.653
R15877 a_30647_7968.n9 a_30647_7968.t10 111.663
R15878 a_30647_7968.n6 a_30647_7968.t21 217.716
R15879 a_30647_7968.t21 a_30647_7968.t17 415.315
R15880 a_30647_7968.t17 a_30647_7968.n7 214.335
R15881 a_30647_7968.n7 a_30647_7968.t18 80.333
R15882 a_30647_7968.n7 a_30647_7968.t19 214.335
R15883 a_30647_7968.n5 a_30647_7968.t6 14.282
R15884 a_30647_7968.n5 a_30647_7968.t7 14.282
R15885 a_30647_7968.n4 a_30647_7968.n3 157.665
R15886 a_30647_7968.n3 a_30647_7968.t0 8.7
R15887 a_30647_7968.n3 a_30647_7968.t1 8.7
R15888 a_30647_7968.n2 a_30647_7968.n1 90.436
R15889 a_30647_7968.n1 a_30647_7968.t4 14.282
R15890 a_30647_7968.n1 a_30647_7968.t3 14.282
R15891 a_30152_3173.n1 a_30152_3173.t4 318.119
R15892 a_30152_3173.n1 a_30152_3173.t6 269.919
R15893 a_30152_3173.n0 a_30152_3173.t5 267.853
R15894 a_30152_3173.n0 a_30152_3173.t7 267.853
R15895 a_30152_3173.t4 a_30152_3173.n0 160.666
R15896 a_30152_3173.n2 a_30152_3173.n1 107.263
R15897 a_30152_3173.t2 a_30152_3173.n4 29.444
R15898 a_30152_3173.n3 a_30152_3173.t0 28.565
R15899 a_30152_3173.n3 a_30152_3173.t1 28.565
R15900 a_30152_3173.n2 a_30152_3173.t3 18.145
R15901 a_30152_3173.n4 a_30152_3173.n2 2.878
R15902 a_30152_3173.n4 a_30152_3173.n3 0.764
R15903 a_29952_3774.n0 a_29952_3774.t11 14.282
R15904 a_29952_3774.t9 a_29952_3774.n0 14.282
R15905 a_29952_3774.n0 a_29952_3774.n9 0.999
R15906 a_29952_3774.n6 a_29952_3774.n8 0.2
R15907 a_29952_3774.n9 a_29952_3774.n6 0.575
R15908 a_29952_3774.n8 a_29952_3774.t3 16.058
R15909 a_29952_3774.n8 a_29952_3774.n7 0.999
R15910 a_29952_3774.n7 a_29952_3774.t5 14.282
R15911 a_29952_3774.n7 a_29952_3774.t4 14.282
R15912 a_29952_3774.n9 a_29952_3774.t10 16.058
R15913 a_29952_3774.n6 a_29952_3774.n4 0.227
R15914 a_29952_3774.n4 a_29952_3774.n5 1.511
R15915 a_29952_3774.n5 a_29952_3774.t8 14.282
R15916 a_29952_3774.n5 a_29952_3774.t7 14.282
R15917 a_29952_3774.n4 a_29952_3774.n1 0.669
R15918 a_29952_3774.n1 a_29952_3774.n2 0.001
R15919 a_29952_3774.n1 a_29952_3774.n3 267.767
R15920 a_29952_3774.n3 a_29952_3774.t0 14.282
R15921 a_29952_3774.n3 a_29952_3774.t2 14.282
R15922 a_29952_3774.n2 a_29952_3774.t1 14.282
R15923 a_29952_3774.n2 a_29952_3774.t6 14.282
R15924 a_37908_2352.n4 a_37908_2352.t9 214.335
R15925 a_37908_2352.t8 a_37908_2352.n4 214.335
R15926 a_37908_2352.n5 a_37908_2352.t8 143.851
R15927 a_37908_2352.n5 a_37908_2352.t7 135.658
R15928 a_37908_2352.n4 a_37908_2352.t10 80.333
R15929 a_37908_2352.n0 a_37908_2352.t4 28.565
R15930 a_37908_2352.n0 a_37908_2352.t5 28.565
R15931 a_37908_2352.n2 a_37908_2352.t1 28.565
R15932 a_37908_2352.n2 a_37908_2352.t3 28.565
R15933 a_37908_2352.n7 a_37908_2352.t0 28.565
R15934 a_37908_2352.t2 a_37908_2352.n7 28.565
R15935 a_37908_2352.n1 a_37908_2352.t6 9.714
R15936 a_37908_2352.n1 a_37908_2352.n0 1.003
R15937 a_37908_2352.n6 a_37908_2352.n3 0.833
R15938 a_37908_2352.n3 a_37908_2352.n2 0.653
R15939 a_37908_2352.n7 a_37908_2352.n6 0.653
R15940 a_37908_2352.n3 a_37908_2352.n1 0.341
R15941 a_37908_2352.n6 a_37908_2352.n5 0.032
R15942 a_39799_1042.n0 a_39799_1042.t5 14.282
R15943 a_39799_1042.t1 a_39799_1042.n0 14.282
R15944 a_39799_1042.n0 a_39799_1042.n12 90.416
R15945 a_39799_1042.n12 a_39799_1042.n11 50.575
R15946 a_39799_1042.n12 a_39799_1042.n8 74.302
R15947 a_39799_1042.n11 a_39799_1042.n10 157.665
R15948 a_39799_1042.n10 a_39799_1042.t4 8.7
R15949 a_39799_1042.n10 a_39799_1042.t0 8.7
R15950 a_39799_1042.n11 a_39799_1042.n9 122.999
R15951 a_39799_1042.n9 a_39799_1042.t3 14.282
R15952 a_39799_1042.n9 a_39799_1042.t2 14.282
R15953 a_39799_1042.n8 a_39799_1042.n7 90.436
R15954 a_39799_1042.n7 a_39799_1042.t6 14.282
R15955 a_39799_1042.n7 a_39799_1042.t7 14.282
R15956 a_39799_1042.n8 a_39799_1042.n1 342.688
R15957 a_39799_1042.n1 a_39799_1042.n6 126.566
R15958 a_39799_1042.n6 a_39799_1042.t11 294.653
R15959 a_39799_1042.n6 a_39799_1042.t13 111.663
R15960 a_39799_1042.n1 a_39799_1042.n5 552.333
R15961 a_39799_1042.n5 a_39799_1042.n4 6.615
R15962 a_39799_1042.n4 a_39799_1042.t8 93.989
R15963 a_39799_1042.n5 a_39799_1042.n3 97.816
R15964 a_39799_1042.n3 a_39799_1042.t15 80.333
R15965 a_39799_1042.n3 a_39799_1042.t9 394.151
R15966 a_39799_1042.t9 a_39799_1042.n2 269.523
R15967 a_39799_1042.n2 a_39799_1042.t14 160.666
R15968 a_39799_1042.n2 a_39799_1042.t10 269.523
R15969 a_39799_1042.n4 a_39799_1042.t12 198.043
R15970 a_41152_1735.n1 a_41152_1735.t7 318.922
R15971 a_41152_1735.n0 a_41152_1735.t4 273.935
R15972 a_41152_1735.n0 a_41152_1735.t5 273.935
R15973 a_41152_1735.n1 a_41152_1735.t6 269.116
R15974 a_41152_1735.n4 a_41152_1735.n3 193.227
R15975 a_41152_1735.t7 a_41152_1735.n0 179.142
R15976 a_41152_1735.n2 a_41152_1735.n1 106.999
R15977 a_41152_1735.n3 a_41152_1735.t1 28.568
R15978 a_41152_1735.n4 a_41152_1735.t0 28.565
R15979 a_41152_1735.t2 a_41152_1735.n4 28.565
R15980 a_41152_1735.n2 a_41152_1735.t3 18.149
R15981 a_41152_1735.n3 a_41152_1735.n2 3.726
R15982 a_13657_20719.n2 a_13657_20719.t6 448.381
R15983 a_13657_20719.n1 a_13657_20719.t5 286.438
R15984 a_13657_20719.n1 a_13657_20719.t7 286.438
R15985 a_13657_20719.n0 a_13657_20719.t4 247.69
R15986 a_13657_20719.n4 a_13657_20719.n3 182.117
R15987 a_13657_20719.t6 a_13657_20719.n1 160.666
R15988 a_13657_20719.n3 a_13657_20719.t0 28.568
R15989 a_13657_20719.n4 a_13657_20719.t1 28.565
R15990 a_13657_20719.t2 a_13657_20719.n4 28.565
R15991 a_13657_20719.n0 a_13657_20719.t3 18.127
R15992 a_13657_20719.n2 a_13657_20719.n0 4.036
R15993 a_13657_20719.n3 a_13657_20719.n2 0.937
R15994 a_30150_1105.n1 a_30150_1105.t6 318.119
R15995 a_30150_1105.n1 a_30150_1105.t4 269.919
R15996 a_30150_1105.n0 a_30150_1105.t7 267.853
R15997 a_30150_1105.n0 a_30150_1105.t5 267.853
R15998 a_30150_1105.t6 a_30150_1105.n0 160.666
R15999 a_30150_1105.n2 a_30150_1105.n1 107.263
R16000 a_30150_1105.t2 a_30150_1105.n4 29.444
R16001 a_30150_1105.n3 a_30150_1105.t0 28.565
R16002 a_30150_1105.n3 a_30150_1105.t1 28.565
R16003 a_30150_1105.n2 a_30150_1105.t3 18.145
R16004 a_30150_1105.n4 a_30150_1105.n2 2.878
R16005 a_30150_1105.n4 a_30150_1105.n3 0.764
R16006 a_9668_1744.n2 a_9668_1744.t4 448.382
R16007 a_9668_1744.n1 a_9668_1744.t6 286.438
R16008 a_9668_1744.n1 a_9668_1744.t7 286.438
R16009 a_9668_1744.n0 a_9668_1744.t5 247.69
R16010 a_9668_1744.n4 a_9668_1744.n3 182.117
R16011 a_9668_1744.t4 a_9668_1744.n1 160.666
R16012 a_9668_1744.n3 a_9668_1744.t1 28.568
R16013 a_9668_1744.n4 a_9668_1744.t0 28.565
R16014 a_9668_1744.t2 a_9668_1744.n4 28.565
R16015 a_9668_1744.n0 a_9668_1744.t3 18.127
R16016 a_9668_1744.n2 a_9668_1744.n0 4.039
R16017 a_9668_1744.n3 a_9668_1744.n2 0.937
R16018 a_9334_20862.n0 a_9334_20862.t7 14.282
R16019 a_9334_20862.t4 a_9334_20862.n0 14.282
R16020 a_9334_20862.n0 a_9334_20862.n1 258.161
R16021 a_9334_20862.n1 a_9334_20862.t5 14.283
R16022 a_9334_20862.n1 a_9334_20862.n7 4.366
R16023 a_9334_20862.n7 a_9334_20862.n5 0.852
R16024 a_9334_20862.n5 a_9334_20862.n6 258.161
R16025 a_9334_20862.n6 a_9334_20862.t2 14.282
R16026 a_9334_20862.n6 a_9334_20862.t1 14.282
R16027 a_9334_20862.n5 a_9334_20862.t3 14.283
R16028 a_9334_20862.n7 a_9334_20862.n4 97.614
R16029 a_9334_20862.n4 a_9334_20862.t8 200.029
R16030 a_9334_20862.t8 a_9334_20862.n3 206.421
R16031 a_9334_20862.n3 a_9334_20862.t9 80.333
R16032 a_9334_20862.n3 a_9334_20862.t10 206.421
R16033 a_9334_20862.n4 a_9334_20862.t11 1527.4
R16034 a_9334_20862.t11 a_9334_20862.n2 657.379
R16035 a_9334_20862.n2 a_9334_20862.t6 8.7
R16036 a_9334_20862.n2 a_9334_20862.t0 8.7
R16037 a_7055_n2174.n2 a_7055_n2174.t5 990.34
R16038 a_7055_n2174.n2 a_7055_n2174.t7 408.211
R16039 a_7055_n2174.n1 a_7055_n2174.t4 286.438
R16040 a_7055_n2174.n1 a_7055_n2174.t6 286.438
R16041 a_7055_n2174.n4 a_7055_n2174.n0 185.55
R16042 a_7055_n2174.t5 a_7055_n2174.n1 160.666
R16043 a_7055_n2174.t2 a_7055_n2174.n4 28.568
R16044 a_7055_n2174.n0 a_7055_n2174.t0 28.565
R16045 a_7055_n2174.n0 a_7055_n2174.t1 28.565
R16046 a_7055_n2174.n3 a_7055_n2174.n2 28.289
R16047 a_7055_n2174.n3 a_7055_n2174.t3 21.376
R16048 a_7055_n2174.n4 a_7055_n2174.n3 1.637
R16049 a_6813_6359.n1 a_6813_6359.t6 990.34
R16050 a_6813_6359.n1 a_6813_6359.t7 408.211
R16051 a_6813_6359.n0 a_6813_6359.t4 286.438
R16052 a_6813_6359.n0 a_6813_6359.t5 286.438
R16053 a_6813_6359.n4 a_6813_6359.n3 195.766
R16054 a_6813_6359.t6 a_6813_6359.n0 160.666
R16055 a_6813_6359.n2 a_6813_6359.n1 38.314
R16056 a_6813_6359.n3 a_6813_6359.t1 28.568
R16057 a_6813_6359.n4 a_6813_6359.t0 28.565
R16058 a_6813_6359.t2 a_6813_6359.n4 28.565
R16059 a_6813_6359.n2 a_6813_6359.t3 18.111
R16060 a_6813_6359.n3 a_6813_6359.n2 0.462
R16061 a_3700_10994.t0 a_3700_10994.n0 14.282
R16062 a_3700_10994.n0 a_3700_10994.t2 14.282
R16063 a_3700_10994.n0 a_3700_10994.n1 258.161
R16064 a_3700_10994.n1 a_3700_10994.t3 14.283
R16065 a_3700_10994.n1 a_3700_10994.n7 4.366
R16066 a_3700_10994.n7 a_3700_10994.n5 0.852
R16067 a_3700_10994.n5 a_3700_10994.n6 258.161
R16068 a_3700_10994.n6 a_3700_10994.t4 14.282
R16069 a_3700_10994.n6 a_3700_10994.t6 14.282
R16070 a_3700_10994.n5 a_3700_10994.t5 14.283
R16071 a_3700_10994.n7 a_3700_10994.n4 97.614
R16072 a_3700_10994.n4 a_3700_10994.t11 200.029
R16073 a_3700_10994.t11 a_3700_10994.n3 206.421
R16074 a_3700_10994.n3 a_3700_10994.t8 80.333
R16075 a_3700_10994.n3 a_3700_10994.t9 206.421
R16076 a_3700_10994.n4 a_3700_10994.t10 1527.4
R16077 a_3700_10994.t10 a_3700_10994.n2 657.379
R16078 a_3700_10994.n2 a_3700_10994.t1 8.7
R16079 a_3700_10994.n2 a_3700_10994.t7 8.7
R16080 a_58868_15769.n5 a_58868_15769.n7 0.2
R16081 a_58868_15769.n9 a_58868_15769.n5 0.575
R16082 a_58868_15769.t3 a_58868_15769.n9 16.058
R16083 a_58868_15769.n9 a_58868_15769.n8 0.999
R16084 a_58868_15769.n8 a_58868_15769.t5 14.282
R16085 a_58868_15769.n8 a_58868_15769.t4 14.282
R16086 a_58868_15769.n7 a_58868_15769.n6 0.999
R16087 a_58868_15769.n6 a_58868_15769.t9 14.282
R16088 a_58868_15769.n6 a_58868_15769.t10 14.282
R16089 a_58868_15769.n7 a_58868_15769.t11 16.058
R16090 a_58868_15769.n5 a_58868_15769.n3 0.227
R16091 a_58868_15769.n3 a_58868_15769.n4 1.511
R16092 a_58868_15769.n4 a_58868_15769.t1 14.282
R16093 a_58868_15769.n4 a_58868_15769.t0 14.282
R16094 a_58868_15769.n3 a_58868_15769.n0 0.669
R16095 a_58868_15769.n0 a_58868_15769.n1 0.001
R16096 a_58868_15769.n0 a_58868_15769.n2 267.767
R16097 a_58868_15769.n2 a_58868_15769.t8 14.282
R16098 a_58868_15769.n2 a_58868_15769.t7 14.282
R16099 a_58868_15769.n1 a_58868_15769.t6 14.282
R16100 a_58868_15769.n1 a_58868_15769.t2 14.282
R16101 a_70509_1146.t0 a_70509_1146.n0 14.282
R16102 a_70509_1146.n0 a_70509_1146.t2 14.282
R16103 a_70509_1146.n0 a_70509_1146.n1 167.433
R16104 a_70509_1146.n1 a_70509_1146.n3 77.784
R16105 a_70509_1146.n3 a_70509_1146.n5 77.456
R16106 a_70509_1146.n5 a_70509_1146.n7 77.456
R16107 a_70509_1146.n7 a_70509_1146.n8 75.815
R16108 a_70509_1146.n8 a_70509_1146.n9 167.433
R16109 a_70509_1146.n9 a_70509_1146.t3 14.282
R16110 a_70509_1146.n9 a_70509_1146.t5 14.282
R16111 a_70509_1146.n8 a_70509_1146.t4 104.259
R16112 a_70509_1146.n7 a_70509_1146.n6 89.977
R16113 a_70509_1146.n6 a_70509_1146.t7 14.282
R16114 a_70509_1146.n6 a_70509_1146.t6 14.282
R16115 a_70509_1146.n5 a_70509_1146.n4 89.977
R16116 a_70509_1146.n4 a_70509_1146.t11 14.282
R16117 a_70509_1146.n4 a_70509_1146.t8 14.282
R16118 a_70509_1146.n3 a_70509_1146.n2 89.977
R16119 a_70509_1146.n2 a_70509_1146.t10 14.282
R16120 a_70509_1146.n2 a_70509_1146.t9 14.282
R16121 a_70509_1146.n1 a_70509_1146.t1 104.259
R16122 a_70509_1028.n2 a_70509_1028.t11 1551.5
R16123 a_70509_1028.t11 a_70509_1028.n0 656.576
R16124 a_70509_1028.n4 a_70509_1028.n3 258.161
R16125 a_70509_1028.n7 a_70509_1028.n6 258.161
R16126 a_70509_1028.n2 a_70509_1028.t8 224.129
R16127 a_70509_1028.n1 a_70509_1028.t10 207.225
R16128 a_70509_1028.t8 a_70509_1028.n1 207.225
R16129 a_70509_1028.n1 a_70509_1028.t9 80.333
R16130 a_70509_1028.n5 a_70509_1028.n2 73.514
R16131 a_70509_1028.n4 a_70509_1028.t3 14.283
R16132 a_70509_1028.n6 a_70509_1028.t0 14.283
R16133 a_70509_1028.n3 a_70509_1028.t4 14.282
R16134 a_70509_1028.n3 a_70509_1028.t5 14.282
R16135 a_70509_1028.n7 a_70509_1028.t1 14.282
R16136 a_70509_1028.t2 a_70509_1028.n7 14.282
R16137 a_70509_1028.n0 a_70509_1028.t7 8.7
R16138 a_70509_1028.n0 a_70509_1028.t6 8.7
R16139 a_70509_1028.n5 a_70509_1028.n4 4.366
R16140 a_70509_1028.n6 a_70509_1028.n5 0.852
R16141 a_30152_4612.n1 a_30152_4612.t4 318.119
R16142 a_30152_4612.n1 a_30152_4612.t6 269.919
R16143 a_30152_4612.n0 a_30152_4612.t5 267.256
R16144 a_30152_4612.n0 a_30152_4612.t7 267.256
R16145 a_30152_4612.n4 a_30152_4612.n3 193.227
R16146 a_30152_4612.t4 a_30152_4612.n0 160.666
R16147 a_30152_4612.n2 a_30152_4612.n1 106.999
R16148 a_30152_4612.n3 a_30152_4612.t0 28.568
R16149 a_30152_4612.n4 a_30152_4612.t1 28.565
R16150 a_30152_4612.t2 a_30152_4612.n4 28.565
R16151 a_30152_4612.n2 a_30152_4612.t3 18.149
R16152 a_30152_4612.n3 a_30152_4612.n2 3.726
R16153 a_59627_1042.t0 a_59627_1042.n0 14.282
R16154 a_59627_1042.n0 a_59627_1042.t2 14.282
R16155 a_59627_1042.n0 a_59627_1042.n12 90.436
R16156 a_59627_1042.n8 a_59627_1042.n11 50.575
R16157 a_59627_1042.n12 a_59627_1042.n8 74.302
R16158 a_59627_1042.n11 a_59627_1042.n10 157.665
R16159 a_59627_1042.n10 a_59627_1042.t6 8.7
R16160 a_59627_1042.n10 a_59627_1042.t7 8.7
R16161 a_59627_1042.n11 a_59627_1042.n9 122.999
R16162 a_59627_1042.n9 a_59627_1042.t5 14.282
R16163 a_59627_1042.n9 a_59627_1042.t4 14.282
R16164 a_59627_1042.n8 a_59627_1042.n7 90.416
R16165 a_59627_1042.n7 a_59627_1042.t3 14.282
R16166 a_59627_1042.n7 a_59627_1042.t1 14.282
R16167 a_59627_1042.n12 a_59627_1042.n1 342.688
R16168 a_59627_1042.n1 a_59627_1042.n6 126.566
R16169 a_59627_1042.n6 a_59627_1042.t15 294.653
R16170 a_59627_1042.n6 a_59627_1042.t14 111.663
R16171 a_59627_1042.n1 a_59627_1042.n5 552.333
R16172 a_59627_1042.n5 a_59627_1042.n4 6.615
R16173 a_59627_1042.n4 a_59627_1042.t9 93.989
R16174 a_59627_1042.n5 a_59627_1042.n3 97.816
R16175 a_59627_1042.n3 a_59627_1042.t13 80.333
R16176 a_59627_1042.n3 a_59627_1042.t8 394.151
R16177 a_59627_1042.t8 a_59627_1042.n2 269.523
R16178 a_59627_1042.n2 a_59627_1042.t12 160.666
R16179 a_59627_1042.n2 a_59627_1042.t10 269.523
R16180 a_59627_1042.n4 a_59627_1042.t11 198.043
R16181 a_61407_1042.n0 a_61407_1042.t1 14.282
R16182 a_61407_1042.t0 a_61407_1042.n0 14.282
R16183 a_61407_1042.n1 a_61407_1042.n9 0.001
R16184 a_61407_1042.n0 a_61407_1042.n1 267.767
R16185 a_61407_1042.n9 a_61407_1042.t10 14.282
R16186 a_61407_1042.n9 a_61407_1042.t2 14.282
R16187 a_61407_1042.n1 a_61407_1042.n7 0.669
R16188 a_61407_1042.n7 a_61407_1042.n8 1.511
R16189 a_61407_1042.n8 a_61407_1042.t11 14.282
R16190 a_61407_1042.n8 a_61407_1042.t9 14.282
R16191 a_61407_1042.n7 a_61407_1042.n6 0.227
R16192 a_61407_1042.n6 a_61407_1042.n3 0.575
R16193 a_61407_1042.n6 a_61407_1042.n5 0.2
R16194 a_61407_1042.n5 a_61407_1042.t4 16.058
R16195 a_61407_1042.n5 a_61407_1042.n4 0.999
R16196 a_61407_1042.n4 a_61407_1042.t5 14.282
R16197 a_61407_1042.n4 a_61407_1042.t3 14.282
R16198 a_61407_1042.n3 a_61407_1042.n2 0.999
R16199 a_61407_1042.n2 a_61407_1042.t8 14.282
R16200 a_61407_1042.n2 a_61407_1042.t7 14.282
R16201 a_61407_1042.n3 a_61407_1042.t6 16.058
R16202 a_60671_22062.n2 a_60671_22062.t5 318.922
R16203 a_60671_22062.n1 a_60671_22062.t4 273.935
R16204 a_60671_22062.n1 a_60671_22062.t6 273.935
R16205 a_60671_22062.n2 a_60671_22062.t7 269.116
R16206 a_60671_22062.n4 a_60671_22062.n0 193.227
R16207 a_60671_22062.t5 a_60671_22062.n1 179.142
R16208 a_60671_22062.n3 a_60671_22062.n2 106.999
R16209 a_60671_22062.t2 a_60671_22062.n4 28.568
R16210 a_60671_22062.n0 a_60671_22062.t0 28.565
R16211 a_60671_22062.n0 a_60671_22062.t1 28.565
R16212 a_60671_22062.n3 a_60671_22062.t3 18.149
R16213 a_60671_22062.n4 a_60671_22062.n3 3.726
R16214 a_45939_15029.t0 a_45939_15029.t1 380.209
R16215 a_19178_n2148.n3 a_19178_n2148.t6 448.382
R16216 a_19178_n2148.n2 a_19178_n2148.t5 286.438
R16217 a_19178_n2148.n2 a_19178_n2148.t7 286.438
R16218 a_19178_n2148.n1 a_19178_n2148.t4 247.69
R16219 a_19178_n2148.n4 a_19178_n2148.n0 182.117
R16220 a_19178_n2148.t6 a_19178_n2148.n2 160.666
R16221 a_19178_n2148.t2 a_19178_n2148.n4 28.568
R16222 a_19178_n2148.n0 a_19178_n2148.t0 28.565
R16223 a_19178_n2148.n0 a_19178_n2148.t1 28.565
R16224 a_19178_n2148.n1 a_19178_n2148.t3 18.127
R16225 a_19178_n2148.n3 a_19178_n2148.n1 4.039
R16226 a_19178_n2148.n4 a_19178_n2148.n3 0.937
R16227 a_71842_1737.t0 a_71842_1737.t1 17.4
R16228 a_65769_n1230.n0 a_65769_n1230.t4 14.282
R16229 a_65769_n1230.t0 a_65769_n1230.n0 14.282
R16230 a_65769_n1230.n0 a_65769_n1230.n8 122.999
R16231 a_65769_n1230.n8 a_65769_n1230.n6 50.575
R16232 a_65769_n1230.n6 a_65769_n1230.n4 74.302
R16233 a_65769_n1230.n8 a_65769_n1230.n7 157.665
R16234 a_65769_n1230.n7 a_65769_n1230.t2 8.7
R16235 a_65769_n1230.n7 a_65769_n1230.t5 8.7
R16236 a_65769_n1230.n6 a_65769_n1230.n5 90.416
R16237 a_65769_n1230.n5 a_65769_n1230.t1 14.282
R16238 a_65769_n1230.n5 a_65769_n1230.t6 14.282
R16239 a_65769_n1230.n4 a_65769_n1230.n3 90.436
R16240 a_65769_n1230.n3 a_65769_n1230.t7 14.282
R16241 a_65769_n1230.n3 a_65769_n1230.t3 14.282
R16242 a_65769_n1230.n4 a_65769_n1230.n1 154.155
R16243 a_65769_n1230.n1 a_65769_n1230.t9 408.806
R16244 a_65769_n1230.t8 a_65769_n1230.n2 160.666
R16245 a_65769_n1230.n1 a_65769_n1230.t8 989.744
R16246 a_65769_n1230.n2 a_65769_n1230.t11 287.241
R16247 a_65769_n1230.n2 a_65769_n1230.t10 287.241
R16248 a_70509_10624.t3 a_70509_10624.n9 104.259
R16249 a_70509_10624.n9 a_70509_10624.n2 77.784
R16250 a_70509_10624.n2 a_70509_10624.n4 77.456
R16251 a_70509_10624.n4 a_70509_10624.n6 77.456
R16252 a_70509_10624.n6 a_70509_10624.n7 75.815
R16253 a_70509_10624.n7 a_70509_10624.n8 167.433
R16254 a_70509_10624.n8 a_70509_10624.t2 14.282
R16255 a_70509_10624.n8 a_70509_10624.t1 14.282
R16256 a_70509_10624.n7 a_70509_10624.t0 104.259
R16257 a_70509_10624.n6 a_70509_10624.n5 89.977
R16258 a_70509_10624.n5 a_70509_10624.t5 14.282
R16259 a_70509_10624.n5 a_70509_10624.t7 14.282
R16260 a_70509_10624.n4 a_70509_10624.n3 89.977
R16261 a_70509_10624.n3 a_70509_10624.t11 14.282
R16262 a_70509_10624.n3 a_70509_10624.t6 14.282
R16263 a_70509_10624.n2 a_70509_10624.n1 89.977
R16264 a_70509_10624.n1 a_70509_10624.t10 14.282
R16265 a_70509_10624.n1 a_70509_10624.t9 14.282
R16266 a_70509_10624.n9 a_70509_10624.n0 167.433
R16267 a_70509_10624.n0 a_70509_10624.t4 14.282
R16268 a_70509_10624.n0 a_70509_10624.t8 14.282
R16269 a_40859_18597.n0 a_40859_18597.t5 14.282
R16270 a_40859_18597.n0 a_40859_18597.t4 14.282
R16271 a_40859_18597.n1 a_40859_18597.t1 14.282
R16272 a_40859_18597.n1 a_40859_18597.t0 14.282
R16273 a_40859_18597.t3 a_40859_18597.n3 14.282
R16274 a_40859_18597.n3 a_40859_18597.t2 14.282
R16275 a_40859_18597.n2 a_40859_18597.n0 2.546
R16276 a_40859_18597.n2 a_40859_18597.n1 2.367
R16277 a_40859_18597.n3 a_40859_18597.n2 0.001
R16278 a_11165_8115.n2 a_11165_8115.t5 448.381
R16279 a_11165_8115.n1 a_11165_8115.t6 286.438
R16280 a_11165_8115.n1 a_11165_8115.t7 286.438
R16281 a_11165_8115.n0 a_11165_8115.t4 247.69
R16282 a_11165_8115.n4 a_11165_8115.n3 182.117
R16283 a_11165_8115.t5 a_11165_8115.n1 160.666
R16284 a_11165_8115.n3 a_11165_8115.t1 28.568
R16285 a_11165_8115.n4 a_11165_8115.t0 28.565
R16286 a_11165_8115.t2 a_11165_8115.n4 28.565
R16287 a_11165_8115.n0 a_11165_8115.t3 18.127
R16288 a_11165_8115.n2 a_11165_8115.n0 4.036
R16289 a_11165_8115.n3 a_11165_8115.n2 0.937
R16290 a_30152_n964.n1 a_30152_n964.t7 318.119
R16291 a_30152_n964.n1 a_30152_n964.t5 269.919
R16292 a_30152_n964.n0 a_30152_n964.t6 267.853
R16293 a_30152_n964.n0 a_30152_n964.t4 267.853
R16294 a_30152_n964.t7 a_30152_n964.n0 160.666
R16295 a_30152_n964.n2 a_30152_n964.n1 107.263
R16296 a_30152_n964.n3 a_30152_n964.t0 29.444
R16297 a_30152_n964.t2 a_30152_n964.n4 28.565
R16298 a_30152_n964.n4 a_30152_n964.t1 28.565
R16299 a_30152_n964.n2 a_30152_n964.t3 18.145
R16300 a_30152_n964.n3 a_30152_n964.n2 2.878
R16301 a_30152_n964.n4 a_30152_n964.n3 0.764
R16302 a_29952_n363.t3 a_29952_n363.n0 14.282
R16303 a_29952_n363.n0 a_29952_n363.t4 14.282
R16304 a_29952_n363.n0 a_29952_n363.n9 0.999
R16305 a_29952_n363.n9 a_29952_n363.n6 0.2
R16306 a_29952_n363.n6 a_29952_n363.n8 0.575
R16307 a_29952_n363.n9 a_29952_n363.t5 16.058
R16308 a_29952_n363.n8 a_29952_n363.n7 0.999
R16309 a_29952_n363.n7 a_29952_n363.t6 14.282
R16310 a_29952_n363.n7 a_29952_n363.t11 14.282
R16311 a_29952_n363.n8 a_29952_n363.t7 16.058
R16312 a_29952_n363.n6 a_29952_n363.n4 0.227
R16313 a_29952_n363.n4 a_29952_n363.n5 1.511
R16314 a_29952_n363.n5 a_29952_n363.t9 14.282
R16315 a_29952_n363.n5 a_29952_n363.t8 14.282
R16316 a_29952_n363.n4 a_29952_n363.n1 0.669
R16317 a_29952_n363.n1 a_29952_n363.n2 0.001
R16318 a_29952_n363.n1 a_29952_n363.n3 267.767
R16319 a_29952_n363.n3 a_29952_n363.t0 14.282
R16320 a_29952_n363.n3 a_29952_n363.t1 14.282
R16321 a_29952_n363.n2 a_29952_n363.t2 14.282
R16322 a_29952_n363.n2 a_29952_n363.t10 14.282
R16323 a_30645_n306.n0 a_30645_n306.t1 14.282
R16324 a_30645_n306.t3 a_30645_n306.n0 14.282
R16325 a_30645_n306.n0 a_30645_n306.n16 90.416
R16326 a_30645_n306.n16 a_30645_n306.n2 74.302
R16327 a_30645_n306.n16 a_30645_n306.n4 50.575
R16328 a_30645_n306.n4 a_30645_n306.n5 110.084
R16329 a_30645_n306.n2 a_30645_n306.n6 691.471
R16330 a_30645_n306.n6 a_30645_n306.n8 16.411
R16331 a_30645_n306.n8 a_30645_n306.t17 198.921
R16332 a_30645_n306.t17 a_30645_n306.t10 415.315
R16333 a_30645_n306.t10 a_30645_n306.n15 214.335
R16334 a_30645_n306.n15 a_30645_n306.t22 80.333
R16335 a_30645_n306.n15 a_30645_n306.t20 214.335
R16336 a_30645_n306.n8 a_30645_n306.n14 861.987
R16337 a_30645_n306.n14 a_30645_n306.n9 560.726
R16338 a_30645_n306.n14 a_30645_n306.n13 65.07
R16339 a_30645_n306.n13 a_30645_n306.n12 6.615
R16340 a_30645_n306.n12 a_30645_n306.t14 93.989
R16341 a_30645_n306.n12 a_30645_n306.t16 198.043
R16342 a_30645_n306.n13 a_30645_n306.n11 97.816
R16343 a_30645_n306.n11 a_30645_n306.t13 80.333
R16344 a_30645_n306.n11 a_30645_n306.t9 394.151
R16345 a_30645_n306.t9 a_30645_n306.n10 269.523
R16346 a_30645_n306.n10 a_30645_n306.t19 160.666
R16347 a_30645_n306.n10 a_30645_n306.t18 269.523
R16348 a_30645_n306.n9 a_30645_n306.t15 294.653
R16349 a_30645_n306.n9 a_30645_n306.t11 111.663
R16350 a_30645_n306.n6 a_30645_n306.t23 217.716
R16351 a_30645_n306.t23 a_30645_n306.t8 415.315
R16352 a_30645_n306.t8 a_30645_n306.n7 214.335
R16353 a_30645_n306.n7 a_30645_n306.t21 80.333
R16354 a_30645_n306.n7 a_30645_n306.t12 214.335
R16355 a_30645_n306.n5 a_30645_n306.t7 14.282
R16356 a_30645_n306.n5 a_30645_n306.t4 14.282
R16357 a_30645_n306.n4 a_30645_n306.n3 157.665
R16358 a_30645_n306.n3 a_30645_n306.t6 8.7
R16359 a_30645_n306.n3 a_30645_n306.t5 8.7
R16360 a_30645_n306.n2 a_30645_n306.n1 90.436
R16361 a_30645_n306.n1 a_30645_n306.t2 14.282
R16362 a_30645_n306.n1 a_30645_n306.t0 14.282
R16363 a_44696_1713.t0 a_44696_1713.t1 17.4
R16364 a_63527_9231.n2 a_63527_9231.t9 214.335
R16365 a_63527_9231.t8 a_63527_9231.n2 214.335
R16366 a_63527_9231.n3 a_63527_9231.t8 143.851
R16367 a_63527_9231.n3 a_63527_9231.t10 135.658
R16368 a_63527_9231.n2 a_63527_9231.t7 80.333
R16369 a_63527_9231.n4 a_63527_9231.t0 28.565
R16370 a_63527_9231.n4 a_63527_9231.t1 28.565
R16371 a_63527_9231.n0 a_63527_9231.t6 28.565
R16372 a_63527_9231.n0 a_63527_9231.t5 28.565
R16373 a_63527_9231.t2 a_63527_9231.n7 28.565
R16374 a_63527_9231.n7 a_63527_9231.t4 28.565
R16375 a_63527_9231.n1 a_63527_9231.t3 9.714
R16376 a_63527_9231.n1 a_63527_9231.n0 1.003
R16377 a_63527_9231.n6 a_63527_9231.n5 0.833
R16378 a_63527_9231.n5 a_63527_9231.n4 0.653
R16379 a_63527_9231.n7 a_63527_9231.n6 0.653
R16380 a_63527_9231.n6 a_63527_9231.n1 0.341
R16381 a_63527_9231.n5 a_63527_9231.n3 0.032
R16382 a_64117_8794.n4 a_64117_8794.n3 563.136
R16383 a_64117_8794.t4 a_64117_8794.t5 437.233
R16384 a_64117_8794.t6 a_64117_8794.n1 313.873
R16385 a_64117_8794.n3 a_64117_8794.t15 294.986
R16386 a_64117_8794.n0 a_64117_8794.t8 272.288
R16387 a_64117_8794.n6 a_64117_8794.t4 217.824
R16388 a_64117_8794.n5 a_64117_8794.t11 214.686
R16389 a_64117_8794.t5 a_64117_8794.n5 214.686
R16390 a_64117_8794.n9 a_64117_8794.n8 192.754
R16391 a_64117_8794.n2 a_64117_8794.t6 190.152
R16392 a_64117_8794.n2 a_64117_8794.t14 190.152
R16393 a_64117_8794.n4 a_64117_8794.t13 178.973
R16394 a_64117_8794.n0 a_64117_8794.t9 160.666
R16395 a_64117_8794.n1 a_64117_8794.t10 160.666
R16396 a_64117_8794.n6 a_64117_8794.n4 133.838
R16397 a_64117_8794.n3 a_64117_8794.t7 110.859
R16398 a_64117_8794.n1 a_64117_8794.n0 96.129
R16399 a_64117_8794.t13 a_64117_8794.n2 80.333
R16400 a_64117_8794.n5 a_64117_8794.t12 80.333
R16401 a_64117_8794.n8 a_64117_8794.t0 28.568
R16402 a_64117_8794.t2 a_64117_8794.n9 28.565
R16403 a_64117_8794.n9 a_64117_8794.t1 28.565
R16404 a_64117_8794.n7 a_64117_8794.t3 18.822
R16405 a_64117_8794.n7 a_64117_8794.n6 5.647
R16406 a_64117_8794.n8 a_64117_8794.n7 1.105
R16407 a_66063_6587.n1 a_66063_6587.t4 318.922
R16408 a_66063_6587.n0 a_66063_6587.t5 274.739
R16409 a_66063_6587.n0 a_66063_6587.t6 274.739
R16410 a_66063_6587.n1 a_66063_6587.t7 269.116
R16411 a_66063_6587.t4 a_66063_6587.n0 179.946
R16412 a_66063_6587.n2 a_66063_6587.n1 107.263
R16413 a_66063_6587.t2 a_66063_6587.n4 29.444
R16414 a_66063_6587.n3 a_66063_6587.t1 28.565
R16415 a_66063_6587.n3 a_66063_6587.t0 28.565
R16416 a_66063_6587.n2 a_66063_6587.t3 18.145
R16417 a_66063_6587.n4 a_66063_6587.n2 2.878
R16418 a_66063_6587.n4 a_66063_6587.n3 0.764
R16419 a_59082_1735.n1 a_59082_1735.t5 318.922
R16420 a_59082_1735.n0 a_59082_1735.t6 273.935
R16421 a_59082_1735.n0 a_59082_1735.t7 273.935
R16422 a_59082_1735.n1 a_59082_1735.t4 269.116
R16423 a_59082_1735.n4 a_59082_1735.n3 193.227
R16424 a_59082_1735.t5 a_59082_1735.n0 179.142
R16425 a_59082_1735.n2 a_59082_1735.n1 106.999
R16426 a_59082_1735.n3 a_59082_1735.t2 28.568
R16427 a_59082_1735.n4 a_59082_1735.t3 28.565
R16428 a_59082_1735.t0 a_59082_1735.n4 28.565
R16429 a_59082_1735.n2 a_59082_1735.t1 18.149
R16430 a_59082_1735.n3 a_59082_1735.n2 3.726
R16431 a_59627_310.t0 a_59627_310.t1 380.209
R16432 a_35575_3749.n4 a_35575_3749.n3 535.449
R16433 a_35575_3749.t17 a_35575_3749.t13 437.233
R16434 a_35575_3749.t7 a_35575_3749.t11 437.233
R16435 a_35575_3749.t8 a_35575_3749.n1 313.873
R16436 a_35575_3749.n3 a_35575_3749.t10 294.986
R16437 a_35575_3749.n0 a_35575_3749.t15 272.288
R16438 a_35575_3749.n4 a_35575_3749.t4 245.184
R16439 a_35575_3749.n6 a_35575_3749.t7 218.628
R16440 a_35575_3749.n8 a_35575_3749.t17 217.026
R16441 a_35575_3749.n7 a_35575_3749.t18 214.686
R16442 a_35575_3749.t13 a_35575_3749.n7 214.686
R16443 a_35575_3749.n5 a_35575_3749.t5 214.686
R16444 a_35575_3749.t11 a_35575_3749.n5 214.686
R16445 a_35575_3749.n11 a_35575_3749.n10 192.754
R16446 a_35575_3749.n2 a_35575_3749.t8 190.152
R16447 a_35575_3749.n2 a_35575_3749.t9 190.152
R16448 a_35575_3749.n0 a_35575_3749.t6 160.666
R16449 a_35575_3749.n1 a_35575_3749.t16 160.666
R16450 a_35575_3749.n3 a_35575_3749.t14 110.859
R16451 a_35575_3749.n1 a_35575_3749.n0 96.129
R16452 a_35575_3749.n7 a_35575_3749.t12 80.333
R16453 a_35575_3749.t4 a_35575_3749.n2 80.333
R16454 a_35575_3749.n5 a_35575_3749.t19 80.333
R16455 a_35575_3749.n10 a_35575_3749.t2 28.568
R16456 a_35575_3749.n11 a_35575_3749.t3 28.565
R16457 a_35575_3749.t1 a_35575_3749.n11 28.565
R16458 a_35575_3749.n9 a_35575_3749.t0 18.722
R16459 a_35575_3749.n6 a_35575_3749.n4 14.9
R16460 a_35575_3749.n8 a_35575_3749.n6 2.603
R16461 a_35575_3749.n9 a_35575_3749.n8 2.382
R16462 a_35575_3749.n10 a_35575_3749.n9 1.281
R16463 a_40093_1016.n1 a_40093_1016.t4 318.922
R16464 a_40093_1016.n0 a_40093_1016.t7 274.739
R16465 a_40093_1016.n0 a_40093_1016.t6 274.739
R16466 a_40093_1016.n1 a_40093_1016.t5 269.116
R16467 a_40093_1016.t4 a_40093_1016.n0 179.946
R16468 a_40093_1016.n2 a_40093_1016.n1 107.263
R16469 a_40093_1016.n3 a_40093_1016.t0 29.444
R16470 a_40093_1016.t2 a_40093_1016.n4 28.565
R16471 a_40093_1016.n4 a_40093_1016.t1 28.565
R16472 a_40093_1016.n2 a_40093_1016.t3 18.145
R16473 a_40093_1016.n3 a_40093_1016.n2 2.878
R16474 a_40093_1016.n4 a_40093_1016.n3 0.764
R16475 A[1].n8 A[1].n7 3623.58
R16476 A[1].n15 A[1].t11 990.34
R16477 A[1].n17 A[1].t21 867.497
R16478 A[1].n17 A[1].t28 591.811
R16479 A[1].t14 A[1].t26 575.234
R16480 A[1].n29 A[1].n19 553.37
R16481 A[1].n24 A[1].n23 535.449
R16482 A[1].t33 A[1].t41 437.233
R16483 A[1].t38 A[1].t31 437.233
R16484 A[1].t37 A[1].t40 437.233
R16485 A[1].n5 A[1].n4 412.11
R16486 A[1].n15 A[1].t8 408.211
R16487 A[1].n2 A[1].t36 394.151
R16488 A[1].t9 A[1].n21 313.873
R16489 A[1].n23 A[1].t32 294.986
R16490 A[1].n4 A[1].t35 294.653
R16491 A[1].n14 A[1].t10 286.438
R16492 A[1].n14 A[1].t22 286.438
R16493 A[1].n16 A[1].t4 286.438
R16494 A[1].n16 A[1].t25 286.438
R16495 A[1].n10 A[1].t16 284.688
R16496 A[1].n20 A[1].t0 272.288
R16497 A[1].n1 A[1].t19 269.523
R16498 A[1].t36 A[1].n1 269.523
R16499 A[1].n24 A[1].t3 245.184
R16500 A[1].n5 A[1].n3 224.13
R16501 A[1].n12 A[1].t33 220.332
R16502 A[1].n26 A[1].t37 218.628
R16503 A[1].n28 A[1].t38 217.024
R16504 A[1].n9 A[1].t43 214.686
R16505 A[1].t41 A[1].n9 214.686
R16506 A[1].n27 A[1].t29 214.686
R16507 A[1].t31 A[1].n27 214.686
R16508 A[1].n25 A[1].t20 214.686
R16509 A[1].t40 A[1].n25 214.686
R16510 A[1].n0 A[1].t23 198.043
R16511 A[1].n22 A[1].t9 190.152
R16512 A[1].n22 A[1].t6 190.152
R16513 A[1].n6 A[1].t1 190.121
R16514 A[1].n6 A[1].t34 190.121
R16515 A[1].n12 A[1].n11 183.203
R16516 A[1].n10 A[1].t12 160.666
R16517 A[1].n11 A[1].t14 160.666
R16518 A[1].n1 A[1].t5 160.666
R16519 A[1].t11 A[1].n14 160.666
R16520 A[1].t21 A[1].n16 160.666
R16521 A[1].n20 A[1].t2 160.666
R16522 A[1].n21 A[1].t18 160.666
R16523 A[1].n8 A[1].n5 140.87
R16524 A[1].n7 A[1].t7 137.369
R16525 A[1].n11 A[1].n10 115.593
R16526 A[1].n6 A[1].t17 112.466
R16527 A[1].n4 A[1].t13 111.663
R16528 A[1].n23 A[1].t27 110.859
R16529 A[1].n3 A[1].n2 97.816
R16530 A[1].n21 A[1].n20 96.129
R16531 A[1].n0 A[1].t39 93.989
R16532 A[1].n9 A[1].t42 80.333
R16533 A[1].n2 A[1].t15 80.333
R16534 A[1].n27 A[1].t30 80.333
R16535 A[1].t3 A[1].n22 80.333
R16536 A[1].n25 A[1].t24 80.333
R16537 A[1].n7 A[1].n6 61.856
R16538 A[1] A[1].n29 45.279
R16539 A[1].n29 A[1].n28 26.946
R16540 A[1].n13 A[1].n12 26.822
R16541 A[1].n18 A[1].n17 25.214
R16542 A[1].n26 A[1].n24 14.9
R16543 A[1].n19 A[1].n13 14.192
R16544 A[1].n13 A[1].n8 8.399
R16545 A[1].n3 A[1].n0 6.615
R16546 A[1].n28 A[1].n26 2.599
R16547 A[1].n19 A[1].n18 2.07
R16548 A[1].n18 A[1].n15 0.004
R16549 a_59187_17949.t5 a_59187_17949.n3 404.877
R16550 a_59187_17949.n2 a_59187_17949.t6 210.902
R16551 a_59187_17949.n4 a_59187_17949.t5 136.949
R16552 a_59187_17949.n3 a_59187_17949.n2 107.801
R16553 a_59187_17949.n2 a_59187_17949.t7 80.333
R16554 a_59187_17949.n3 a_59187_17949.t8 80.333
R16555 a_59187_17949.n1 a_59187_17949.t2 17.4
R16556 a_59187_17949.n1 a_59187_17949.t1 17.4
R16557 a_59187_17949.t0 a_59187_17949.n5 15.032
R16558 a_59187_17949.n0 a_59187_17949.t4 14.282
R16559 a_59187_17949.n0 a_59187_17949.t3 14.282
R16560 a_59187_17949.n5 a_59187_17949.n0 1.65
R16561 a_59187_17949.n4 a_59187_17949.n1 0.657
R16562 a_59187_17949.n5 a_59187_17949.n4 0.614
R16563 a_54713_3294.n8 a_54713_3294.n7 861.987
R16564 a_54713_3294.n7 a_54713_3294.n6 560.726
R16565 a_54713_3294.t13 a_54713_3294.t12 415.315
R16566 a_54713_3294.t18 a_54713_3294.t14 415.315
R16567 a_54713_3294.n3 a_54713_3294.t5 394.151
R16568 a_54713_3294.n6 a_54713_3294.t16 294.653
R16569 a_54713_3294.n2 a_54713_3294.t7 269.523
R16570 a_54713_3294.t5 a_54713_3294.n2 269.523
R16571 a_54713_3294.n10 a_54713_3294.t13 217.716
R16572 a_54713_3294.n9 a_54713_3294.t19 214.335
R16573 a_54713_3294.t12 a_54713_3294.n9 214.335
R16574 a_54713_3294.n1 a_54713_3294.t4 214.335
R16575 a_54713_3294.t14 a_54713_3294.n1 214.335
R16576 a_54713_3294.n8 a_54713_3294.t18 198.921
R16577 a_54713_3294.n4 a_54713_3294.t11 198.043
R16578 a_54713_3294.n2 a_54713_3294.t15 160.666
R16579 a_54713_3294.n6 a_54713_3294.t9 111.663
R16580 a_54713_3294.n5 a_54713_3294.n3 97.816
R16581 a_54713_3294.n4 a_54713_3294.t6 93.989
R16582 a_54713_3294.n9 a_54713_3294.t8 80.333
R16583 a_54713_3294.n3 a_54713_3294.t17 80.333
R16584 a_54713_3294.n1 a_54713_3294.t10 80.333
R16585 a_54713_3294.n7 a_54713_3294.n5 65.07
R16586 a_54713_3294.n0 a_54713_3294.t1 28.57
R16587 a_54713_3294.t0 a_54713_3294.n12 28.565
R16588 a_54713_3294.n12 a_54713_3294.t2 28.565
R16589 a_54713_3294.n0 a_54713_3294.t3 17.638
R16590 a_54713_3294.n10 a_54713_3294.n8 16.411
R16591 a_54713_3294.n11 a_54713_3294.n10 7.315
R16592 a_54713_3294.n5 a_54713_3294.n4 6.615
R16593 a_54713_3294.n12 a_54713_3294.n11 0.69
R16594 a_54713_3294.n11 a_54713_3294.n0 0.6
R16595 a_57744_8220.n0 a_57744_8220.t8 214.335
R16596 a_57744_8220.t9 a_57744_8220.n0 214.335
R16597 a_57744_8220.n1 a_57744_8220.t9 143.851
R16598 a_57744_8220.n1 a_57744_8220.t10 135.658
R16599 a_57744_8220.n0 a_57744_8220.t7 80.333
R16600 a_57744_8220.n2 a_57744_8220.t2 28.565
R16601 a_57744_8220.n2 a_57744_8220.t1 28.565
R16602 a_57744_8220.n4 a_57744_8220.t0 28.565
R16603 a_57744_8220.n4 a_57744_8220.t4 28.565
R16604 a_57744_8220.n7 a_57744_8220.t6 28.565
R16605 a_57744_8220.t3 a_57744_8220.n7 28.565
R16606 a_57744_8220.n6 a_57744_8220.t5 9.714
R16607 a_57744_8220.n7 a_57744_8220.n6 1.003
R16608 a_57744_8220.n5 a_57744_8220.n3 0.833
R16609 a_57744_8220.n3 a_57744_8220.n2 0.653
R16610 a_57744_8220.n5 a_57744_8220.n4 0.653
R16611 a_57744_8220.n6 a_57744_8220.n5 0.341
R16612 a_57744_8220.n3 a_57744_8220.n1 0.032
R16613 a_39807_6090.t0 a_39807_6090.t1 380.209
R16614 a_53010_6842.t1 a_53010_6842.n0 14.282
R16615 a_53010_6842.n0 a_53010_6842.t3 14.282
R16616 a_53010_6842.n0 a_53010_6842.n12 90.436
R16617 a_53010_6842.n8 a_53010_6842.n11 50.575
R16618 a_53010_6842.n12 a_53010_6842.n8 74.302
R16619 a_53010_6842.n11 a_53010_6842.n10 157.665
R16620 a_53010_6842.n10 a_53010_6842.t4 8.7
R16621 a_53010_6842.n10 a_53010_6842.t0 8.7
R16622 a_53010_6842.n11 a_53010_6842.n9 122.999
R16623 a_53010_6842.n9 a_53010_6842.t7 14.282
R16624 a_53010_6842.n9 a_53010_6842.t6 14.282
R16625 a_53010_6842.n8 a_53010_6842.n7 90.416
R16626 a_53010_6842.n7 a_53010_6842.t5 14.282
R16627 a_53010_6842.n7 a_53010_6842.t2 14.282
R16628 a_53010_6842.n12 a_53010_6842.n1 342.688
R16629 a_53010_6842.n1 a_53010_6842.n6 126.566
R16630 a_53010_6842.n6 a_53010_6842.t12 294.653
R16631 a_53010_6842.n6 a_53010_6842.t11 111.663
R16632 a_53010_6842.n1 a_53010_6842.n5 552.333
R16633 a_53010_6842.n5 a_53010_6842.n4 6.615
R16634 a_53010_6842.n4 a_53010_6842.t10 93.989
R16635 a_53010_6842.n5 a_53010_6842.n3 97.816
R16636 a_53010_6842.n3 a_53010_6842.t15 80.333
R16637 a_53010_6842.n3 a_53010_6842.t8 394.151
R16638 a_53010_6842.t8 a_53010_6842.n2 269.523
R16639 a_53010_6842.n2 a_53010_6842.t9 160.666
R16640 a_53010_6842.n2 a_53010_6842.t14 269.523
R16641 a_53010_6842.n4 a_53010_6842.t13 198.043
R16642 a_54790_6842.t3 a_54790_6842.n7 16.058
R16643 a_54790_6842.n7 a_54790_6842.n5 0.575
R16644 a_54790_6842.n5 a_54790_6842.n9 0.2
R16645 a_54790_6842.n9 a_54790_6842.t1 16.058
R16646 a_54790_6842.n9 a_54790_6842.n8 0.999
R16647 a_54790_6842.n8 a_54790_6842.t2 14.282
R16648 a_54790_6842.n8 a_54790_6842.t0 14.282
R16649 a_54790_6842.n7 a_54790_6842.n6 0.999
R16650 a_54790_6842.n6 a_54790_6842.t4 14.282
R16651 a_54790_6842.n6 a_54790_6842.t5 14.282
R16652 a_54790_6842.n5 a_54790_6842.n3 0.227
R16653 a_54790_6842.n3 a_54790_6842.n4 1.511
R16654 a_54790_6842.n4 a_54790_6842.t11 14.282
R16655 a_54790_6842.n4 a_54790_6842.t10 14.282
R16656 a_54790_6842.n3 a_54790_6842.n0 0.669
R16657 a_54790_6842.n0 a_54790_6842.n1 0.001
R16658 a_54790_6842.n0 a_54790_6842.n2 267.767
R16659 a_54790_6842.n2 a_54790_6842.t6 14.282
R16660 a_54790_6842.n2 a_54790_6842.t7 14.282
R16661 a_54790_6842.n1 a_54790_6842.t9 14.282
R16662 a_54790_6842.n1 a_54790_6842.t8 14.282
R16663 a_53891_18572.t5 a_53891_18572.t6 800.071
R16664 a_53891_18572.n3 a_53891_18572.n2 659.095
R16665 a_53891_18572.n1 a_53891_18572.t7 285.109
R16666 a_53891_18572.n2 a_53891_18572.t5 193.602
R16667 a_53891_18572.n4 a_53891_18572.n0 192.754
R16668 a_53891_18572.n1 a_53891_18572.t4 160.666
R16669 a_53891_18572.n2 a_53891_18572.n1 91.507
R16670 a_53891_18572.t2 a_53891_18572.n4 28.568
R16671 a_53891_18572.n0 a_53891_18572.t0 28.565
R16672 a_53891_18572.n0 a_53891_18572.t1 28.565
R16673 a_53891_18572.n3 a_53891_18572.t3 19.063
R16674 a_53891_18572.n4 a_53891_18572.n3 1.005
R16675 a_53951_18598.n0 a_53951_18598.t2 14.282
R16676 a_53951_18598.n0 a_53951_18598.t1 14.282
R16677 a_53951_18598.n1 a_53951_18598.t5 14.282
R16678 a_53951_18598.n1 a_53951_18598.t3 14.282
R16679 a_53951_18598.t0 a_53951_18598.n3 14.282
R16680 a_53951_18598.n3 a_53951_18598.t4 14.282
R16681 a_53951_18598.n2 a_53951_18598.n0 2.546
R16682 a_53951_18598.n2 a_53951_18598.n1 2.367
R16683 a_53951_18598.n3 a_53951_18598.n2 0.001
R16684 a_10227_1744.n0 a_10227_1744.n9 167.433
R16685 a_10227_1744.t0 a_10227_1744.n0 14.282
R16686 a_10227_1744.n0 a_10227_1744.t2 14.282
R16687 a_10227_1744.n9 a_10227_1744.n8 75.815
R16688 a_10227_1744.n8 a_10227_1744.n6 77.456
R16689 a_10227_1744.n6 a_10227_1744.n4 77.456
R16690 a_10227_1744.n4 a_10227_1744.n2 77.784
R16691 a_10227_1744.n9 a_10227_1744.t1 104.259
R16692 a_10227_1744.n8 a_10227_1744.n7 89.977
R16693 a_10227_1744.n7 a_10227_1744.t4 14.282
R16694 a_10227_1744.n7 a_10227_1744.t5 14.282
R16695 a_10227_1744.n6 a_10227_1744.n5 89.977
R16696 a_10227_1744.n5 a_10227_1744.t3 14.282
R16697 a_10227_1744.n5 a_10227_1744.t7 14.282
R16698 a_10227_1744.n4 a_10227_1744.n3 89.977
R16699 a_10227_1744.n3 a_10227_1744.t8 14.282
R16700 a_10227_1744.n3 a_10227_1744.t6 14.282
R16701 a_10227_1744.n2 a_10227_1744.t10 104.259
R16702 a_10227_1744.n2 a_10227_1744.n1 167.433
R16703 a_10227_1744.n1 a_10227_1744.t11 14.282
R16704 a_10227_1744.n1 a_10227_1744.t9 14.282
R16705 a_30154_11447.n1 a_30154_11447.t5 318.119
R16706 a_30154_11447.n1 a_30154_11447.t6 269.919
R16707 a_30154_11447.n0 a_30154_11447.t7 267.853
R16708 a_30154_11447.n0 a_30154_11447.t4 267.853
R16709 a_30154_11447.t5 a_30154_11447.n0 160.666
R16710 a_30154_11447.n2 a_30154_11447.n1 107.263
R16711 a_30154_11447.n3 a_30154_11447.t0 29.444
R16712 a_30154_11447.n4 a_30154_11447.t1 28.565
R16713 a_30154_11447.t2 a_30154_11447.n4 28.565
R16714 a_30154_11447.n2 a_30154_11447.t3 18.145
R16715 a_30154_11447.n3 a_30154_11447.n2 2.878
R16716 a_30154_11447.n4 a_30154_11447.n3 0.764
R16717 a_53357_22238.t7 a_53357_22238.t6 574.43
R16718 a_53357_22238.n1 a_53357_22238.t5 285.109
R16719 a_53357_22238.n3 a_53357_22238.n2 211.136
R16720 a_53357_22238.n4 a_53357_22238.n0 192.754
R16721 a_53357_22238.n1 a_53357_22238.t4 160.666
R16722 a_53357_22238.n2 a_53357_22238.t7 160.666
R16723 a_53357_22238.n2 a_53357_22238.n1 114.829
R16724 a_53357_22238.t0 a_53357_22238.n4 28.568
R16725 a_53357_22238.n0 a_53357_22238.t3 28.565
R16726 a_53357_22238.n0 a_53357_22238.t2 28.565
R16727 a_53357_22238.n3 a_53357_22238.t1 19.084
R16728 a_53357_22238.n4 a_53357_22238.n3 1.051
R16729 a_56220_24201.n0 a_56220_24201.t5 14.282
R16730 a_56220_24201.n0 a_56220_24201.t3 14.282
R16731 a_56220_24201.n1 a_56220_24201.t2 14.282
R16732 a_56220_24201.n1 a_56220_24201.t1 14.282
R16733 a_56220_24201.t0 a_56220_24201.n3 14.282
R16734 a_56220_24201.n3 a_56220_24201.t4 14.282
R16735 a_56220_24201.n2 a_56220_24201.n0 2.546
R16736 a_56220_24201.n2 a_56220_24201.n1 2.367
R16737 a_56220_24201.n3 a_56220_24201.n2 0.001
R16738 a_56102_24201.t6 a_56102_24201.n2 404.877
R16739 a_56102_24201.n1 a_56102_24201.t8 210.902
R16740 a_56102_24201.n3 a_56102_24201.t6 136.943
R16741 a_56102_24201.n2 a_56102_24201.n1 107.801
R16742 a_56102_24201.n1 a_56102_24201.t7 80.333
R16743 a_56102_24201.n2 a_56102_24201.t5 80.333
R16744 a_56102_24201.n0 a_56102_24201.t0 17.4
R16745 a_56102_24201.n0 a_56102_24201.t4 17.4
R16746 a_56102_24201.n4 a_56102_24201.t1 15.032
R16747 a_56102_24201.n5 a_56102_24201.t2 14.282
R16748 a_56102_24201.t3 a_56102_24201.n5 14.282
R16749 a_56102_24201.n5 a_56102_24201.n4 1.65
R16750 a_56102_24201.n3 a_56102_24201.n0 0.672
R16751 a_56102_24201.n4 a_56102_24201.n3 0.665
R16752 a_4879_10851.n2 a_4879_10851.t6 448.381
R16753 a_4879_10851.n1 a_4879_10851.t4 286.438
R16754 a_4879_10851.n1 a_4879_10851.t7 286.438
R16755 a_4879_10851.n0 a_4879_10851.t5 247.69
R16756 a_4879_10851.n4 a_4879_10851.n3 182.117
R16757 a_4879_10851.t6 a_4879_10851.n1 160.666
R16758 a_4879_10851.n3 a_4879_10851.t1 28.568
R16759 a_4879_10851.t2 a_4879_10851.n4 28.565
R16760 a_4879_10851.n4 a_4879_10851.t0 28.565
R16761 a_4879_10851.n0 a_4879_10851.t3 18.127
R16762 a_4879_10851.n2 a_4879_10851.n0 4.036
R16763 a_4879_10851.n3 a_4879_10851.n2 0.937
R16764 a_70459_8189.n2 a_70459_8189.t7 448.381
R16765 a_70459_8189.n1 a_70459_8189.t4 287.241
R16766 a_70459_8189.n1 a_70459_8189.t6 287.241
R16767 a_70459_8189.n0 a_70459_8189.t5 247.733
R16768 a_70459_8189.n4 a_70459_8189.n3 182.117
R16769 a_70459_8189.t7 a_70459_8189.n1 160.666
R16770 a_70459_8189.n3 a_70459_8189.t0 28.568
R16771 a_70459_8189.n4 a_70459_8189.t1 28.565
R16772 a_70459_8189.t2 a_70459_8189.n4 28.565
R16773 a_70459_8189.n0 a_70459_8189.t3 18.127
R16774 a_70459_8189.n2 a_70459_8189.n0 4.036
R16775 a_70459_8189.n3 a_70459_8189.n2 0.937
R16776 a_35004_7464.n2 a_35004_7464.t9 214.335
R16777 a_35004_7464.t7 a_35004_7464.n2 214.335
R16778 a_35004_7464.n3 a_35004_7464.t7 143.851
R16779 a_35004_7464.n3 a_35004_7464.t8 135.658
R16780 a_35004_7464.n2 a_35004_7464.t10 80.333
R16781 a_35004_7464.n4 a_35004_7464.t5 28.565
R16782 a_35004_7464.n4 a_35004_7464.t4 28.565
R16783 a_35004_7464.n0 a_35004_7464.t2 28.565
R16784 a_35004_7464.n0 a_35004_7464.t3 28.565
R16785 a_35004_7464.n7 a_35004_7464.t6 28.565
R16786 a_35004_7464.t1 a_35004_7464.n7 28.565
R16787 a_35004_7464.n1 a_35004_7464.t0 9.714
R16788 a_35004_7464.n1 a_35004_7464.n0 1.003
R16789 a_35004_7464.n6 a_35004_7464.n5 0.833
R16790 a_35004_7464.n5 a_35004_7464.n4 0.653
R16791 a_35004_7464.n7 a_35004_7464.n6 0.653
R16792 a_35004_7464.n6 a_35004_7464.n1 0.341
R16793 a_35004_7464.n5 a_35004_7464.n3 0.032
R16794 a_43055_24209.t7 a_43055_24209.n3 404.877
R16795 a_43055_24209.n2 a_43055_24209.t8 210.902
R16796 a_43055_24209.n4 a_43055_24209.t7 136.943
R16797 a_43055_24209.n3 a_43055_24209.n2 107.801
R16798 a_43055_24209.n2 a_43055_24209.t6 80.333
R16799 a_43055_24209.n3 a_43055_24209.t5 80.333
R16800 a_43055_24209.n1 a_43055_24209.t4 17.4
R16801 a_43055_24209.n1 a_43055_24209.t2 17.4
R16802 a_43055_24209.t0 a_43055_24209.n5 15.032
R16803 a_43055_24209.n0 a_43055_24209.t3 14.282
R16804 a_43055_24209.n0 a_43055_24209.t1 14.282
R16805 a_43055_24209.n5 a_43055_24209.n0 1.65
R16806 a_43055_24209.n4 a_43055_24209.n1 0.672
R16807 a_43055_24209.n5 a_43055_24209.n4 0.665
R16808 a_43319_23626.n6 a_43319_23626.n5 501.28
R16809 a_43319_23626.t16 a_43319_23626.t4 437.233
R16810 a_43319_23626.t15 a_43319_23626.t17 415.315
R16811 a_43319_23626.t9 a_43319_23626.n3 313.873
R16812 a_43319_23626.n5 a_43319_23626.t13 294.986
R16813 a_43319_23626.n2 a_43319_23626.t5 272.288
R16814 a_43319_23626.n6 a_43319_23626.t10 236.01
R16815 a_43319_23626.n9 a_43319_23626.t16 216.627
R16816 a_43319_23626.n7 a_43319_23626.t15 216.111
R16817 a_43319_23626.n8 a_43319_23626.t11 214.686
R16818 a_43319_23626.t4 a_43319_23626.n8 214.686
R16819 a_43319_23626.n1 a_43319_23626.t7 214.335
R16820 a_43319_23626.t17 a_43319_23626.n1 214.335
R16821 a_43319_23626.n4 a_43319_23626.t9 190.152
R16822 a_43319_23626.n4 a_43319_23626.t8 190.152
R16823 a_43319_23626.n2 a_43319_23626.t6 160.666
R16824 a_43319_23626.n3 a_43319_23626.t14 160.666
R16825 a_43319_23626.n7 a_43319_23626.n6 148.428
R16826 a_43319_23626.n5 a_43319_23626.t19 110.859
R16827 a_43319_23626.n3 a_43319_23626.n2 96.129
R16828 a_43319_23626.n8 a_43319_23626.t12 80.333
R16829 a_43319_23626.n1 a_43319_23626.t18 80.333
R16830 a_43319_23626.t10 a_43319_23626.n4 80.333
R16831 a_43319_23626.t2 a_43319_23626.n11 28.57
R16832 a_43319_23626.n0 a_43319_23626.t0 28.565
R16833 a_43319_23626.n0 a_43319_23626.t1 28.565
R16834 a_43319_23626.n11 a_43319_23626.t3 17.638
R16835 a_43319_23626.n10 a_43319_23626.n9 5.375
R16836 a_43319_23626.n9 a_43319_23626.n7 2.923
R16837 a_43319_23626.n10 a_43319_23626.n0 0.69
R16838 a_43319_23626.n11 a_43319_23626.n10 0.6
R16839 a_5659_15753.t8 a_5659_15753.n2 406.978
R16840 a_5659_15753.n1 a_5659_15753.t5 207.38
R16841 a_5659_15753.n3 a_5659_15753.t8 136.949
R16842 a_5659_15753.n2 a_5659_15753.n1 112.003
R16843 a_5659_15753.n1 a_5659_15753.t6 80.333
R16844 a_5659_15753.n2 a_5659_15753.t7 80.333
R16845 a_5659_15753.n0 a_5659_15753.t2 17.4
R16846 a_5659_15753.n0 a_5659_15753.t0 17.4
R16847 a_5659_15753.n4 a_5659_15753.t3 15.036
R16848 a_5659_15753.n5 a_5659_15753.t4 14.282
R16849 a_5659_15753.t1 a_5659_15753.n5 14.282
R16850 a_5659_15753.n5 a_5659_15753.n4 1.654
R16851 a_5659_15753.n3 a_5659_15753.n0 0.657
R16852 a_5659_15753.n4 a_5659_15753.n3 0.614
R16853 a_5794_16410.n1 a_5794_16410.t3 14.282
R16854 a_5794_16410.n1 a_5794_16410.t0 14.282
R16855 a_5794_16410.n0 a_5794_16410.t4 14.282
R16856 a_5794_16410.n0 a_5794_16410.t5 14.282
R16857 a_5794_16410.n3 a_5794_16410.t1 14.282
R16858 a_5794_16410.t2 a_5794_16410.n3 14.282
R16859 a_5794_16410.n2 a_5794_16410.n0 2.538
R16860 a_5794_16410.n3 a_5794_16410.n2 2.375
R16861 a_5794_16410.n2 a_5794_16410.n1 0.001
R16862 a_54245_18572.t6 a_54245_18572.t7 574.43
R16863 a_54245_18572.n0 a_54245_18572.t4 285.109
R16864 a_54245_18572.n2 a_54245_18572.n1 197.215
R16865 a_54245_18572.n4 a_54245_18572.n3 192.754
R16866 a_54245_18572.n0 a_54245_18572.t5 160.666
R16867 a_54245_18572.n1 a_54245_18572.t6 160.666
R16868 a_54245_18572.n1 a_54245_18572.n0 114.829
R16869 a_54245_18572.n3 a_54245_18572.t1 28.568
R16870 a_54245_18572.t2 a_54245_18572.n4 28.565
R16871 a_54245_18572.n4 a_54245_18572.t0 28.565
R16872 a_54245_18572.n2 a_54245_18572.t3 18.838
R16873 a_54245_18572.n3 a_54245_18572.n2 1.129
R16874 a_70513_16900.t0 a_70513_16900.n9 104.259
R16875 a_70513_16900.n9 a_70513_16900.n2 77.784
R16876 a_70513_16900.n2 a_70513_16900.n4 77.456
R16877 a_70513_16900.n4 a_70513_16900.n6 77.456
R16878 a_70513_16900.n6 a_70513_16900.n7 75.815
R16879 a_70513_16900.n7 a_70513_16900.n8 167.433
R16880 a_70513_16900.n8 a_70513_16900.t5 14.282
R16881 a_70513_16900.n8 a_70513_16900.t3 14.282
R16882 a_70513_16900.n7 a_70513_16900.t4 104.259
R16883 a_70513_16900.n6 a_70513_16900.n5 89.977
R16884 a_70513_16900.n5 a_70513_16900.t7 14.282
R16885 a_70513_16900.n5 a_70513_16900.t8 14.282
R16886 a_70513_16900.n4 a_70513_16900.n3 89.977
R16887 a_70513_16900.n3 a_70513_16900.t9 14.282
R16888 a_70513_16900.n3 a_70513_16900.t6 14.282
R16889 a_70513_16900.n2 a_70513_16900.n1 89.977
R16890 a_70513_16900.n1 a_70513_16900.t11 14.282
R16891 a_70513_16900.n1 a_70513_16900.t10 14.282
R16892 a_70513_16900.n9 a_70513_16900.n0 167.433
R16893 a_70513_16900.n0 a_70513_16900.t1 14.282
R16894 a_70513_16900.n0 a_70513_16900.t2 14.282
R16895 a_9918_14454.n1 a_9918_14454.t5 867.497
R16896 a_9918_14454.n1 a_9918_14454.t6 591.811
R16897 a_9918_14454.n0 a_9918_14454.t4 286.438
R16898 a_9918_14454.n0 a_9918_14454.t7 286.438
R16899 a_9918_14454.n4 a_9918_14454.n3 185.55
R16900 a_9918_14454.t5 a_9918_14454.n0 160.666
R16901 a_9918_14454.n3 a_9918_14454.t1 28.568
R16902 a_9918_14454.t2 a_9918_14454.n4 28.565
R16903 a_9918_14454.n4 a_9918_14454.t0 28.565
R16904 a_9918_14454.n2 a_9918_14454.n1 25.445
R16905 a_9918_14454.n2 a_9918_14454.t3 21.376
R16906 a_9918_14454.n3 a_9918_14454.n2 1.637
R16907 a_9976_10990.n0 a_9976_10990.t1 14.282
R16908 a_9976_10990.t0 a_9976_10990.n0 14.282
R16909 a_9976_10990.n0 a_9976_10990.n1 258.161
R16910 a_9976_10990.n1 a_9976_10990.n5 0.852
R16911 a_9976_10990.n5 a_9976_10990.n6 4.366
R16912 a_9976_10990.n6 a_9976_10990.n7 258.161
R16913 a_9976_10990.n7 a_9976_10990.t4 14.282
R16914 a_9976_10990.n7 a_9976_10990.t5 14.282
R16915 a_9976_10990.n6 a_9976_10990.t6 14.283
R16916 a_9976_10990.n5 a_9976_10990.n4 97.614
R16917 a_9976_10990.n4 a_9976_10990.t10 200.029
R16918 a_9976_10990.t10 a_9976_10990.n3 206.421
R16919 a_9976_10990.n3 a_9976_10990.t11 80.333
R16920 a_9976_10990.n3 a_9976_10990.t8 206.421
R16921 a_9976_10990.n4 a_9976_10990.t9 1527.4
R16922 a_9976_10990.t9 a_9976_10990.n2 657.379
R16923 a_9976_10990.n2 a_9976_10990.t7 8.7
R16924 a_9976_10990.n2 a_9976_10990.t3 8.7
R16925 a_9976_10990.n1 a_9976_10990.t2 14.283
R16926 a_10509_11720.t3 a_10509_11720.n9 104.259
R16927 a_10509_11720.n6 a_10509_11720.n7 77.784
R16928 a_10509_11720.n4 a_10509_11720.n6 77.456
R16929 a_10509_11720.n2 a_10509_11720.n4 77.456
R16930 a_10509_11720.n9 a_10509_11720.n2 75.815
R16931 a_10509_11720.n7 a_10509_11720.n8 167.433
R16932 a_10509_11720.n8 a_10509_11720.t2 14.282
R16933 a_10509_11720.n8 a_10509_11720.t1 14.282
R16934 a_10509_11720.n7 a_10509_11720.t0 104.259
R16935 a_10509_11720.n6 a_10509_11720.n5 89.977
R16936 a_10509_11720.n5 a_10509_11720.t7 14.282
R16937 a_10509_11720.n5 a_10509_11720.t8 14.282
R16938 a_10509_11720.n4 a_10509_11720.n3 89.977
R16939 a_10509_11720.n3 a_10509_11720.t6 14.282
R16940 a_10509_11720.n3 a_10509_11720.t9 14.282
R16941 a_10509_11720.n2 a_10509_11720.n1 89.977
R16942 a_10509_11720.n1 a_10509_11720.t10 14.282
R16943 a_10509_11720.n1 a_10509_11720.t11 14.282
R16944 a_10509_11720.n9 a_10509_11720.n0 167.433
R16945 a_10509_11720.n0 a_10509_11720.t4 14.282
R16946 a_10509_11720.n0 a_10509_11720.t5 14.282
R16947 a_49904_21370.t0 a_49904_21370.n0 14.282
R16948 a_49904_21370.n0 a_49904_21370.t1 14.282
R16949 a_49904_21370.n0 a_49904_21370.n9 0.999
R16950 a_49904_21370.n6 a_49904_21370.n8 0.575
R16951 a_49904_21370.n9 a_49904_21370.n6 0.2
R16952 a_49904_21370.n9 a_49904_21370.t2 16.058
R16953 a_49904_21370.n8 a_49904_21370.n7 0.999
R16954 a_49904_21370.n7 a_49904_21370.t9 14.282
R16955 a_49904_21370.n7 a_49904_21370.t11 14.282
R16956 a_49904_21370.n8 a_49904_21370.t10 16.058
R16957 a_49904_21370.n6 a_49904_21370.n4 0.227
R16958 a_49904_21370.n4 a_49904_21370.n5 1.511
R16959 a_49904_21370.n5 a_49904_21370.t5 14.282
R16960 a_49904_21370.n5 a_49904_21370.t4 14.282
R16961 a_49904_21370.n4 a_49904_21370.n1 0.669
R16962 a_49904_21370.n1 a_49904_21370.n2 0.001
R16963 a_49904_21370.n1 a_49904_21370.n3 267.767
R16964 a_49904_21370.n3 a_49904_21370.t7 14.282
R16965 a_49904_21370.n3 a_49904_21370.t6 14.282
R16966 a_49904_21370.n2 a_49904_21370.t3 14.282
R16967 a_49904_21370.n2 a_49904_21370.t8 14.282
R16968 a_55848_17050.n0 a_55848_17050.t9 214.335
R16969 a_55848_17050.t8 a_55848_17050.n0 214.335
R16970 a_55848_17050.n1 a_55848_17050.t8 143.851
R16971 a_55848_17050.n1 a_55848_17050.t7 135.658
R16972 a_55848_17050.n0 a_55848_17050.t10 80.333
R16973 a_55848_17050.n2 a_55848_17050.t0 28.565
R16974 a_55848_17050.n2 a_55848_17050.t1 28.565
R16975 a_55848_17050.n4 a_55848_17050.t2 28.565
R16976 a_55848_17050.n4 a_55848_17050.t6 28.565
R16977 a_55848_17050.n7 a_55848_17050.t5 28.565
R16978 a_55848_17050.t4 a_55848_17050.n7 28.565
R16979 a_55848_17050.n3 a_55848_17050.t3 9.714
R16980 a_55848_17050.n3 a_55848_17050.n2 1.003
R16981 a_55848_17050.n6 a_55848_17050.n5 0.833
R16982 a_55848_17050.n5 a_55848_17050.n4 0.653
R16983 a_55848_17050.n7 a_55848_17050.n6 0.653
R16984 a_55848_17050.n5 a_55848_17050.n3 0.341
R16985 a_55848_17050.n6 a_55848_17050.n1 0.032
R16986 a_53103_18576.t6 a_53103_18576.t7 574.43
R16987 a_53103_18576.n0 a_53103_18576.t4 285.109
R16988 a_53103_18576.n2 a_53103_18576.n1 211.134
R16989 a_53103_18576.n4 a_53103_18576.n3 192.754
R16990 a_53103_18576.n0 a_53103_18576.t5 160.666
R16991 a_53103_18576.n1 a_53103_18576.t6 160.666
R16992 a_53103_18576.n1 a_53103_18576.n0 114.829
R16993 a_53103_18576.n3 a_53103_18576.t1 28.568
R16994 a_53103_18576.t2 a_53103_18576.n4 28.565
R16995 a_53103_18576.n4 a_53103_18576.t0 28.565
R16996 a_53103_18576.n2 a_53103_18576.t3 19.087
R16997 a_53103_18576.n3 a_53103_18576.n2 1.051
R16998 a_46652_3872.t7 a_46652_3872.n3 404.877
R16999 a_46652_3872.n2 a_46652_3872.t5 210.902
R17000 a_46652_3872.n4 a_46652_3872.t7 136.943
R17001 a_46652_3872.n3 a_46652_3872.n2 107.801
R17002 a_46652_3872.n2 a_46652_3872.t6 80.333
R17003 a_46652_3872.n3 a_46652_3872.t8 80.333
R17004 a_46652_3872.n1 a_46652_3872.t4 17.4
R17005 a_46652_3872.n1 a_46652_3872.t1 17.4
R17006 a_46652_3872.t0 a_46652_3872.n5 15.032
R17007 a_46652_3872.n0 a_46652_3872.t2 14.282
R17008 a_46652_3872.n0 a_46652_3872.t3 14.282
R17009 a_46652_3872.n5 a_46652_3872.n0 1.65
R17010 a_46652_3872.n4 a_46652_3872.n1 0.672
R17011 a_46652_3872.n5 a_46652_3872.n4 0.665
R17012 a_46916_3289.t5 a_46916_3289.t6 800.071
R17013 a_46916_3289.n3 a_46916_3289.n2 672.951
R17014 a_46916_3289.n1 a_46916_3289.t7 285.109
R17015 a_46916_3289.n2 a_46916_3289.t5 193.602
R17016 a_46916_3289.n1 a_46916_3289.t4 160.666
R17017 a_46916_3289.n2 a_46916_3289.n1 91.507
R17018 a_46916_3289.n0 a_46916_3289.t0 28.57
R17019 a_46916_3289.t2 a_46916_3289.n4 28.565
R17020 a_46916_3289.n4 a_46916_3289.t1 28.565
R17021 a_46916_3289.n0 a_46916_3289.t3 17.638
R17022 a_46916_3289.n4 a_46916_3289.n3 0.69
R17023 a_46916_3289.n3 a_46916_3289.n0 0.6
R17024 a_31379_7968.t0 a_31379_7968.t1 379.845
R17025 a_70455_14535.n2 a_70455_14535.t5 448.381
R17026 a_70455_14535.n1 a_70455_14535.t7 287.241
R17027 a_70455_14535.n1 a_70455_14535.t4 287.241
R17028 a_70455_14535.n0 a_70455_14535.t6 247.733
R17029 a_70455_14535.n4 a_70455_14535.n3 182.117
R17030 a_70455_14535.t5 a_70455_14535.n1 160.666
R17031 a_70455_14535.n3 a_70455_14535.t0 28.568
R17032 a_70455_14535.n4 a_70455_14535.t1 28.565
R17033 a_70455_14535.t2 a_70455_14535.n4 28.565
R17034 a_70455_14535.n0 a_70455_14535.t3 18.127
R17035 a_70455_14535.n2 a_70455_14535.n0 4.036
R17036 a_70455_14535.n3 a_70455_14535.n2 0.937
R17037 a_70509_13768.t0 a_70509_13768.n9 104.259
R17038 a_70509_13768.n9 a_70509_13768.n2 77.784
R17039 a_70509_13768.n2 a_70509_13768.n4 77.456
R17040 a_70509_13768.n4 a_70509_13768.n6 77.456
R17041 a_70509_13768.n6 a_70509_13768.n7 75.815
R17042 a_70509_13768.n7 a_70509_13768.n8 167.433
R17043 a_70509_13768.n8 a_70509_13768.t4 14.282
R17044 a_70509_13768.n8 a_70509_13768.t5 14.282
R17045 a_70509_13768.n7 a_70509_13768.t3 104.259
R17046 a_70509_13768.n6 a_70509_13768.n5 89.977
R17047 a_70509_13768.n5 a_70509_13768.t7 14.282
R17048 a_70509_13768.n5 a_70509_13768.t6 14.282
R17049 a_70509_13768.n4 a_70509_13768.n3 89.977
R17050 a_70509_13768.n3 a_70509_13768.t9 14.282
R17051 a_70509_13768.n3 a_70509_13768.t8 14.282
R17052 a_70509_13768.n2 a_70509_13768.n1 89.977
R17053 a_70509_13768.n1 a_70509_13768.t11 14.282
R17054 a_70509_13768.n1 a_70509_13768.t10 14.282
R17055 a_70509_13768.n9 a_70509_13768.n0 167.433
R17056 a_70509_13768.n0 a_70509_13768.t1 14.282
R17057 a_70509_13768.n0 a_70509_13768.t2 14.282
R17058 a_70509_13650.n0 a_70509_13650.t2 14.282
R17059 a_70509_13650.t0 a_70509_13650.n0 14.282
R17060 a_70509_13650.n0 a_70509_13650.n1 258.161
R17061 a_70509_13650.n1 a_70509_13650.t1 14.283
R17062 a_70509_13650.n1 a_70509_13650.n5 0.852
R17063 a_70509_13650.n5 a_70509_13650.n6 4.366
R17064 a_70509_13650.n6 a_70509_13650.n7 258.161
R17065 a_70509_13650.n7 a_70509_13650.t6 14.282
R17066 a_70509_13650.n7 a_70509_13650.t5 14.282
R17067 a_70509_13650.n6 a_70509_13650.t4 14.283
R17068 a_70509_13650.n5 a_70509_13650.n4 73.514
R17069 a_70509_13650.n4 a_70509_13650.t9 1551.5
R17070 a_70509_13650.t9 a_70509_13650.n3 656.576
R17071 a_70509_13650.n3 a_70509_13650.t3 8.7
R17072 a_70509_13650.n3 a_70509_13650.t7 8.7
R17073 a_70509_13650.n4 a_70509_13650.t11 224.129
R17074 a_70509_13650.t11 a_70509_13650.n2 207.225
R17075 a_70509_13650.n2 a_70509_13650.t10 207.225
R17076 a_70509_13650.n2 a_70509_13650.t8 80.333
R17077 a_14357_10851.n2 a_14357_10851.t6 448.381
R17078 a_14357_10851.n1 a_14357_10851.t5 286.438
R17079 a_14357_10851.n1 a_14357_10851.t4 286.438
R17080 a_14357_10851.n0 a_14357_10851.t7 247.69
R17081 a_14357_10851.n4 a_14357_10851.n3 182.117
R17082 a_14357_10851.t6 a_14357_10851.n1 160.666
R17083 a_14357_10851.n3 a_14357_10851.t0 28.568
R17084 a_14357_10851.n4 a_14357_10851.t1 28.565
R17085 a_14357_10851.t2 a_14357_10851.n4 28.565
R17086 a_14357_10851.n0 a_14357_10851.t3 18.127
R17087 a_14357_10851.n2 a_14357_10851.n0 4.036
R17088 a_14357_10851.n3 a_14357_10851.n2 0.937
R17089 a_29952_9980.t6 a_29952_9980.n9 16.058
R17090 a_29952_9980.n9 a_29952_9980.n5 0.2
R17091 a_29952_9980.n5 a_29952_9980.n7 0.575
R17092 a_29952_9980.n9 a_29952_9980.n8 0.999
R17093 a_29952_9980.n8 a_29952_9980.t7 14.282
R17094 a_29952_9980.n8 a_29952_9980.t8 14.282
R17095 a_29952_9980.n7 a_29952_9980.n6 0.999
R17096 a_29952_9980.n6 a_29952_9980.t10 14.282
R17097 a_29952_9980.n6 a_29952_9980.t9 14.282
R17098 a_29952_9980.n7 a_29952_9980.t11 16.058
R17099 a_29952_9980.n5 a_29952_9980.n3 0.227
R17100 a_29952_9980.n3 a_29952_9980.n4 1.511
R17101 a_29952_9980.n4 a_29952_9980.t5 14.282
R17102 a_29952_9980.n4 a_29952_9980.t4 14.282
R17103 a_29952_9980.n3 a_29952_9980.n0 0.669
R17104 a_29952_9980.n0 a_29952_9980.n1 0.001
R17105 a_29952_9980.n0 a_29952_9980.n2 267.767
R17106 a_29952_9980.n2 a_29952_9980.t1 14.282
R17107 a_29952_9980.n2 a_29952_9980.t2 14.282
R17108 a_29952_9980.n1 a_29952_9980.t0 14.282
R17109 a_29952_9980.n1 a_29952_9980.t3 14.282
R17110 a_57676_2326.n4 a_57676_2326.n3 501.28
R17111 a_57676_2326.t7 a_57676_2326.t8 437.233
R17112 a_57676_2326.t14 a_57676_2326.t18 415.315
R17113 a_57676_2326.t13 a_57676_2326.n1 313.873
R17114 a_57676_2326.n3 a_57676_2326.t16 294.986
R17115 a_57676_2326.n0 a_57676_2326.t15 272.288
R17116 a_57676_2326.n4 a_57676_2326.t9 236.01
R17117 a_57676_2326.n8 a_57676_2326.t7 216.627
R17118 a_57676_2326.n6 a_57676_2326.t14 216.069
R17119 a_57676_2326.n7 a_57676_2326.t6 214.686
R17120 a_57676_2326.t8 a_57676_2326.n7 214.686
R17121 a_57676_2326.n5 a_57676_2326.t12 214.335
R17122 a_57676_2326.t18 a_57676_2326.n5 214.335
R17123 a_57676_2326.n11 a_57676_2326.n10 192.754
R17124 a_57676_2326.n2 a_57676_2326.t13 190.152
R17125 a_57676_2326.n2 a_57676_2326.t4 190.152
R17126 a_57676_2326.n0 a_57676_2326.t11 160.666
R17127 a_57676_2326.n1 a_57676_2326.t5 160.666
R17128 a_57676_2326.n6 a_57676_2326.n4 148.384
R17129 a_57676_2326.n3 a_57676_2326.t10 110.859
R17130 a_57676_2326.n1 a_57676_2326.n0 96.129
R17131 a_57676_2326.n7 a_57676_2326.t19 80.333
R17132 a_57676_2326.n5 a_57676_2326.t17 80.333
R17133 a_57676_2326.t9 a_57676_2326.n2 80.333
R17134 a_57676_2326.n9 a_57676_2326.n8 47.31
R17135 a_57676_2326.n10 a_57676_2326.t1 28.568
R17136 a_57676_2326.n11 a_57676_2326.t0 28.565
R17137 a_57676_2326.t2 a_57676_2326.n11 28.565
R17138 a_57676_2326.n9 a_57676_2326.t3 18.466
R17139 a_57676_2326.n8 a_57676_2326.n6 2.697
R17140 a_57676_2326.n10 a_57676_2326.n9 1.161
R17141 a_51100_4001.n0 a_51100_4001.t8 214.335
R17142 a_51100_4001.t7 a_51100_4001.n0 214.335
R17143 a_51100_4001.n1 a_51100_4001.t7 143.851
R17144 a_51100_4001.n1 a_51100_4001.t9 135.658
R17145 a_51100_4001.n0 a_51100_4001.t10 80.333
R17146 a_51100_4001.n2 a_51100_4001.t5 28.565
R17147 a_51100_4001.n2 a_51100_4001.t4 28.565
R17148 a_51100_4001.n4 a_51100_4001.t6 28.565
R17149 a_51100_4001.n4 a_51100_4001.t1 28.565
R17150 a_51100_4001.n7 a_51100_4001.t2 28.565
R17151 a_51100_4001.t0 a_51100_4001.n7 28.565
R17152 a_51100_4001.n6 a_51100_4001.t3 9.714
R17153 a_51100_4001.n7 a_51100_4001.n6 1.003
R17154 a_51100_4001.n5 a_51100_4001.n3 0.833
R17155 a_51100_4001.n3 a_51100_4001.n2 0.653
R17156 a_51100_4001.n5 a_51100_4001.n4 0.653
R17157 a_51100_4001.n6 a_51100_4001.n5 0.341
R17158 a_51100_4001.n3 a_51100_4001.n1 0.032
R17159 a_51690_3564.t6 a_51690_3564.t4 800.071
R17160 a_51690_3564.n2 a_51690_3564.n1 659.097
R17161 a_51690_3564.n0 a_51690_3564.t7 285.109
R17162 a_51690_3564.n1 a_51690_3564.t6 193.602
R17163 a_51690_3564.n4 a_51690_3564.n3 192.754
R17164 a_51690_3564.n0 a_51690_3564.t5 160.666
R17165 a_51690_3564.n1 a_51690_3564.n0 91.507
R17166 a_51690_3564.n3 a_51690_3564.t1 28.568
R17167 a_51690_3564.n4 a_51690_3564.t0 28.565
R17168 a_51690_3564.t2 a_51690_3564.n4 28.565
R17169 a_51690_3564.n2 a_51690_3564.t3 19.061
R17170 a_51690_3564.n3 a_51690_3564.n2 1.005
R17171 a_70459_17667.n2 a_70459_17667.t4 448.381
R17172 a_70459_17667.n1 a_70459_17667.t5 287.241
R17173 a_70459_17667.n1 a_70459_17667.t7 287.241
R17174 a_70459_17667.n0 a_70459_17667.t6 247.733
R17175 a_70459_17667.n4 a_70459_17667.n3 182.117
R17176 a_70459_17667.t4 a_70459_17667.n1 160.666
R17177 a_70459_17667.n3 a_70459_17667.t0 28.568
R17178 a_70459_17667.n4 a_70459_17667.t1 28.565
R17179 a_70459_17667.t2 a_70459_17667.n4 28.565
R17180 a_70459_17667.n0 a_70459_17667.t3 18.127
R17181 a_70459_17667.n2 a_70459_17667.n0 4.036
R17182 a_70459_17667.n3 a_70459_17667.n2 0.937
R17183 a_19937_8962.t0 a_19937_8962.n0 14.282
R17184 a_19937_8962.n0 a_19937_8962.t7 14.282
R17185 a_19937_8962.n0 a_19937_8962.n8 90.436
R17186 a_19937_8962.n8 a_19937_8962.n5 74.302
R17187 a_19937_8962.n5 a_19937_8962.n7 50.575
R17188 a_19937_8962.n7 a_19937_8962.n6 157.665
R17189 a_19937_8962.n6 a_19937_8962.t1 8.7
R17190 a_19937_8962.n6 a_19937_8962.t2 8.7
R17191 a_19937_8962.n5 a_19937_8962.n4 90.416
R17192 a_19937_8962.n4 a_19937_8962.t6 14.282
R17193 a_19937_8962.n4 a_19937_8962.t3 14.282
R17194 a_19937_8962.n7 a_19937_8962.n3 122.746
R17195 a_19937_8962.n3 a_19937_8962.t5 14.282
R17196 a_19937_8962.n3 a_19937_8962.t4 14.282
R17197 a_19937_8962.n8 a_19937_8962.n1 1100.5
R17198 a_19937_8962.n1 a_19937_8962.t9 591.811
R17199 a_19937_8962.n1 a_19937_8962.t10 867.497
R17200 a_19937_8962.t10 a_19937_8962.n2 160.666
R17201 a_19937_8962.n2 a_19937_8962.t8 286.438
R17202 a_19937_8962.n2 a_19937_8962.t11 286.438
R17203 a_19997_8988.t9 a_19997_8988.n9 104.259
R17204 a_19997_8988.n6 a_19997_8988.n7 77.784
R17205 a_19997_8988.n4 a_19997_8988.n6 77.456
R17206 a_19997_8988.n2 a_19997_8988.n4 77.456
R17207 a_19997_8988.n9 a_19997_8988.n2 75.815
R17208 a_19997_8988.n7 a_19997_8988.n8 167.433
R17209 a_19997_8988.n8 a_19997_8988.t6 14.282
R17210 a_19997_8988.n8 a_19997_8988.t7 14.282
R17211 a_19997_8988.n7 a_19997_8988.t8 104.259
R17212 a_19997_8988.n6 a_19997_8988.n5 89.977
R17213 a_19997_8988.n5 a_19997_8988.t1 14.282
R17214 a_19997_8988.n5 a_19997_8988.t2 14.282
R17215 a_19997_8988.n4 a_19997_8988.n3 89.977
R17216 a_19997_8988.n3 a_19997_8988.t0 14.282
R17217 a_19997_8988.n3 a_19997_8988.t3 14.282
R17218 a_19997_8988.n2 a_19997_8988.n1 89.977
R17219 a_19997_8988.n1 a_19997_8988.t4 14.282
R17220 a_19997_8988.n1 a_19997_8988.t5 14.282
R17221 a_19997_8988.n9 a_19997_8988.n0 167.433
R17222 a_19997_8988.n0 a_19997_8988.t11 14.282
R17223 a_19997_8988.n0 a_19997_8988.t10 14.282
R17224 a_7432_1744.n0 a_7432_1744.t7 14.282
R17225 a_7432_1744.t4 a_7432_1744.n0 14.282
R17226 a_7432_1744.n0 a_7432_1744.n1 258.161
R17227 a_7432_1744.n1 a_7432_1744.n7 4.366
R17228 a_7432_1744.n7 a_7432_1744.n5 0.852
R17229 a_7432_1744.n5 a_7432_1744.n6 258.161
R17230 a_7432_1744.n6 a_7432_1744.t2 14.282
R17231 a_7432_1744.n6 a_7432_1744.t3 14.282
R17232 a_7432_1744.n5 a_7432_1744.t1 14.283
R17233 a_7432_1744.n7 a_7432_1744.n4 97.614
R17234 a_7432_1744.n4 a_7432_1744.t9 200.029
R17235 a_7432_1744.t9 a_7432_1744.n3 206.421
R17236 a_7432_1744.n3 a_7432_1744.t8 80.333
R17237 a_7432_1744.n3 a_7432_1744.t11 206.421
R17238 a_7432_1744.n4 a_7432_1744.t10 1527.4
R17239 a_7432_1744.t10 a_7432_1744.n2 657.379
R17240 a_7432_1744.n2 a_7432_1744.t0 8.7
R17241 a_7432_1744.n2 a_7432_1744.t5 8.7
R17242 a_7432_1744.n1 a_7432_1744.t6 14.283
R17243 a_7989_n2633.n1 a_7989_n2633.t6 867.497
R17244 a_7989_n2633.n1 a_7989_n2633.t4 615.911
R17245 a_7989_n2633.n0 a_7989_n2633.t5 286.438
R17246 a_7989_n2633.n0 a_7989_n2633.t7 286.438
R17247 a_7989_n2633.n4 a_7989_n2633.n3 185.55
R17248 a_7989_n2633.t6 a_7989_n2633.n0 160.666
R17249 a_7989_n2633.n3 a_7989_n2633.t1 28.568
R17250 a_7989_n2633.t2 a_7989_n2633.n4 28.565
R17251 a_7989_n2633.n4 a_7989_n2633.t0 28.565
R17252 a_7989_n2633.n2 a_7989_n2633.n1 22.152
R17253 a_7989_n2633.n2 a_7989_n2633.t3 20.4
R17254 a_7989_n2633.n3 a_7989_n2633.n2 1.828
R17255 a_54952_21339.n1 a_54952_21339.t7 318.922
R17256 a_54952_21339.n0 a_54952_21339.t4 274.739
R17257 a_54952_21339.n0 a_54952_21339.t5 274.739
R17258 a_54952_21339.n1 a_54952_21339.t6 269.116
R17259 a_54952_21339.t7 a_54952_21339.n0 179.946
R17260 a_54952_21339.n2 a_54952_21339.n1 107.263
R17261 a_54952_21339.n3 a_54952_21339.t1 29.444
R17262 a_54952_21339.t2 a_54952_21339.n4 28.565
R17263 a_54952_21339.n4 a_54952_21339.t0 28.565
R17264 a_54952_21339.n2 a_54952_21339.t3 18.145
R17265 a_54952_21339.n3 a_54952_21339.n2 2.878
R17266 a_54952_21339.n4 a_54952_21339.n3 0.764
R17267 a_44459_2350.n0 a_44459_2350.t7 214.335
R17268 a_44459_2350.t10 a_44459_2350.n0 214.335
R17269 a_44459_2350.n1 a_44459_2350.t10 143.851
R17270 a_44459_2350.n1 a_44459_2350.t9 135.658
R17271 a_44459_2350.n0 a_44459_2350.t8 80.333
R17272 a_44459_2350.n2 a_44459_2350.t5 28.565
R17273 a_44459_2350.n2 a_44459_2350.t4 28.565
R17274 a_44459_2350.n4 a_44459_2350.t6 28.565
R17275 a_44459_2350.n4 a_44459_2350.t1 28.565
R17276 a_44459_2350.n7 a_44459_2350.t0 28.565
R17277 a_44459_2350.t2 a_44459_2350.n7 28.565
R17278 a_44459_2350.n6 a_44459_2350.t3 9.714
R17279 a_44459_2350.n7 a_44459_2350.n6 1.003
R17280 a_44459_2350.n5 a_44459_2350.n3 0.833
R17281 a_44459_2350.n3 a_44459_2350.n2 0.653
R17282 a_44459_2350.n5 a_44459_2350.n4 0.653
R17283 a_44459_2350.n6 a_44459_2350.n5 0.341
R17284 a_44459_2350.n3 a_44459_2350.n1 0.032
R17285 a_15946_15776.t0 a_15946_15776.t1 17.4
R17286 a_42761_15445.n0 a_42761_15445.t10 214.335
R17287 a_42761_15445.t9 a_42761_15445.n0 214.335
R17288 a_42761_15445.n1 a_42761_15445.t9 143.851
R17289 a_42761_15445.n1 a_42761_15445.t7 135.658
R17290 a_42761_15445.n0 a_42761_15445.t8 80.333
R17291 a_42761_15445.n2 a_42761_15445.t6 28.565
R17292 a_42761_15445.n2 a_42761_15445.t4 28.565
R17293 a_42761_15445.n4 a_42761_15445.t5 28.565
R17294 a_42761_15445.n4 a_42761_15445.t0 28.565
R17295 a_42761_15445.n7 a_42761_15445.t1 28.565
R17296 a_42761_15445.t2 a_42761_15445.n7 28.565
R17297 a_42761_15445.n3 a_42761_15445.t3 9.714
R17298 a_42761_15445.n3 a_42761_15445.n2 1.003
R17299 a_42761_15445.n6 a_42761_15445.n5 0.833
R17300 a_42761_15445.n5 a_42761_15445.n4 0.653
R17301 a_42761_15445.n7 a_42761_15445.n6 0.653
R17302 a_42761_15445.n5 a_42761_15445.n3 0.341
R17303 a_42761_15445.n6 a_42761_15445.n1 0.032
R17304 a_41153_18571.t6 a_41153_18571.t7 574.43
R17305 a_41153_18571.n0 a_41153_18571.t4 285.109
R17306 a_41153_18571.n2 a_41153_18571.n1 197.215
R17307 a_41153_18571.n4 a_41153_18571.n3 192.754
R17308 a_41153_18571.n0 a_41153_18571.t5 160.666
R17309 a_41153_18571.n1 a_41153_18571.t6 160.666
R17310 a_41153_18571.n1 a_41153_18571.n0 114.829
R17311 a_41153_18571.n3 a_41153_18571.t0 28.568
R17312 a_41153_18571.n4 a_41153_18571.t1 28.565
R17313 a_41153_18571.t2 a_41153_18571.n4 28.565
R17314 a_41153_18571.n2 a_41153_18571.t3 18.838
R17315 a_41153_18571.n3 a_41153_18571.n2 1.129
R17316 a_13188_8262.t0 a_13188_8262.n0 14.282
R17317 a_13188_8262.n0 a_13188_8262.t7 14.282
R17318 a_13188_8262.n0 a_13188_8262.n1 258.161
R17319 a_13188_8262.n1 a_13188_8262.t5 14.283
R17320 a_13188_8262.n1 a_13188_8262.n7 4.366
R17321 a_13188_8262.n7 a_13188_8262.n5 0.852
R17322 a_13188_8262.n5 a_13188_8262.n6 258.161
R17323 a_13188_8262.n6 a_13188_8262.t2 14.282
R17324 a_13188_8262.n6 a_13188_8262.t3 14.282
R17325 a_13188_8262.n5 a_13188_8262.t4 14.283
R17326 a_13188_8262.n7 a_13188_8262.n4 97.614
R17327 a_13188_8262.n4 a_13188_8262.t10 200.029
R17328 a_13188_8262.t10 a_13188_8262.n3 206.421
R17329 a_13188_8262.n3 a_13188_8262.t8 80.333
R17330 a_13188_8262.n3 a_13188_8262.t11 206.421
R17331 a_13188_8262.n4 a_13188_8262.t9 1527.4
R17332 a_13188_8262.t9 a_13188_8262.n2 657.379
R17333 a_13188_8262.n2 a_13188_8262.t6 8.7
R17334 a_13188_8262.n2 a_13188_8262.t1 8.7
R17335 a_13721_8992.n0 a_13721_8992.t2 14.282
R17336 a_13721_8992.t0 a_13721_8992.n0 14.282
R17337 a_13721_8992.n0 a_13721_8992.n9 89.977
R17338 a_13721_8992.n6 a_13721_8992.n7 77.784
R17339 a_13721_8992.n9 a_13721_8992.n6 77.456
R17340 a_13721_8992.n9 a_13721_8992.n4 77.456
R17341 a_13721_8992.n4 a_13721_8992.n2 75.815
R17342 a_13721_8992.n7 a_13721_8992.n8 167.433
R17343 a_13721_8992.n8 a_13721_8992.t6 14.282
R17344 a_13721_8992.n8 a_13721_8992.t4 14.282
R17345 a_13721_8992.n7 a_13721_8992.t5 104.259
R17346 a_13721_8992.n6 a_13721_8992.n5 89.977
R17347 a_13721_8992.n5 a_13721_8992.t3 14.282
R17348 a_13721_8992.n5 a_13721_8992.t1 14.282
R17349 a_13721_8992.n4 a_13721_8992.n3 89.977
R17350 a_13721_8992.n3 a_13721_8992.t8 14.282
R17351 a_13721_8992.n3 a_13721_8992.t7 14.282
R17352 a_13721_8992.n2 a_13721_8992.t10 104.259
R17353 a_13721_8992.n2 a_13721_8992.n1 167.433
R17354 a_13721_8992.n1 a_13721_8992.t11 14.282
R17355 a_13721_8992.n1 a_13721_8992.t9 14.282
R17356 a_61343_9163.n2 a_61343_9163.t4 989.744
R17357 a_61343_9163.n3 a_61343_9163.n2 494.286
R17358 a_61343_9163.n2 a_61343_9163.t5 408.806
R17359 a_61343_9163.n1 a_61343_9163.t7 287.241
R17360 a_61343_9163.n1 a_61343_9163.t6 287.241
R17361 a_61343_9163.t4 a_61343_9163.n1 160.666
R17362 a_61343_9163.n0 a_61343_9163.t1 28.57
R17363 a_61343_9163.n4 a_61343_9163.t2 28.565
R17364 a_61343_9163.t0 a_61343_9163.n4 28.565
R17365 a_61343_9163.n0 a_61343_9163.t3 17.638
R17366 a_61343_9163.n4 a_61343_9163.n3 0.69
R17367 a_61343_9163.n3 a_61343_9163.n0 0.6
R17368 a_38723_16458.n1 a_38723_16458.t6 318.922
R17369 a_38723_16458.n0 a_38723_16458.t5 274.739
R17370 a_38723_16458.n0 a_38723_16458.t7 274.739
R17371 a_38723_16458.n1 a_38723_16458.t4 269.116
R17372 a_38723_16458.t6 a_38723_16458.n0 179.946
R17373 a_38723_16458.n2 a_38723_16458.n1 105.178
R17374 a_38723_16458.n3 a_38723_16458.t0 29.444
R17375 a_38723_16458.n4 a_38723_16458.t1 28.565
R17376 a_38723_16458.t2 a_38723_16458.n4 28.565
R17377 a_38723_16458.n2 a_38723_16458.t3 18.145
R17378 a_38723_16458.n3 a_38723_16458.n2 2.878
R17379 a_38723_16458.n4 a_38723_16458.n3 0.764
R17380 a_9918_11720.n1 a_9918_11720.t7 990.34
R17381 a_9918_11720.n1 a_9918_11720.t6 408.211
R17382 a_9918_11720.n0 a_9918_11720.t4 286.438
R17383 a_9918_11720.n0 a_9918_11720.t5 286.438
R17384 a_9918_11720.n2 a_9918_11720.n1 216.826
R17385 a_9918_11720.n4 a_9918_11720.n3 185.55
R17386 a_9918_11720.t7 a_9918_11720.n0 160.666
R17387 a_9918_11720.n3 a_9918_11720.t1 28.568
R17388 a_9918_11720.t2 a_9918_11720.n4 28.565
R17389 a_9918_11720.n4 a_9918_11720.t0 28.565
R17390 a_9918_11720.n2 a_9918_11720.t3 21.562
R17391 a_9918_11720.n3 a_9918_11720.n2 1.603
R17392 a_51105_9802.n4 a_51105_9802.t9 214.335
R17393 a_51105_9802.t8 a_51105_9802.n4 214.335
R17394 a_51105_9802.n5 a_51105_9802.t8 143.851
R17395 a_51105_9802.n5 a_51105_9802.t10 135.658
R17396 a_51105_9802.n4 a_51105_9802.t7 80.333
R17397 a_51105_9802.n0 a_51105_9802.t3 28.565
R17398 a_51105_9802.n0 a_51105_9802.t5 28.565
R17399 a_51105_9802.n2 a_51105_9802.t0 28.565
R17400 a_51105_9802.n2 a_51105_9802.t4 28.565
R17401 a_51105_9802.t2 a_51105_9802.n7 28.565
R17402 a_51105_9802.n7 a_51105_9802.t1 28.565
R17403 a_51105_9802.n1 a_51105_9802.t6 9.714
R17404 a_51105_9802.n1 a_51105_9802.n0 1.003
R17405 a_51105_9802.n6 a_51105_9802.n3 0.833
R17406 a_51105_9802.n3 a_51105_9802.n2 0.653
R17407 a_51105_9802.n7 a_51105_9802.n6 0.653
R17408 a_51105_9802.n3 a_51105_9802.n1 0.341
R17409 a_51105_9802.n6 a_51105_9802.n5 0.032
R17410 a_42964_22066.n2 a_42964_22066.t6 318.922
R17411 a_42964_22066.n1 a_42964_22066.t5 273.935
R17412 a_42964_22066.n1 a_42964_22066.t7 273.935
R17413 a_42964_22066.n2 a_42964_22066.t4 269.116
R17414 a_42964_22066.n4 a_42964_22066.n0 193.227
R17415 a_42964_22066.t6 a_42964_22066.n1 179.142
R17416 a_42964_22066.n3 a_42964_22066.n2 106.999
R17417 a_42964_22066.t0 a_42964_22066.n4 28.568
R17418 a_42964_22066.n0 a_42964_22066.t2 28.565
R17419 a_42964_22066.n0 a_42964_22066.t1 28.565
R17420 a_42964_22066.n3 a_42964_22066.t3 18.149
R17421 a_42964_22066.n4 a_42964_22066.n3 3.726
R17422 a_43509_20641.t0 a_43509_20641.t1 380.209
R17423 a_43509_21373.t0 a_43509_21373.n0 14.282
R17424 a_43509_21373.n0 a_43509_21373.t5 14.282
R17425 a_43509_21373.n0 a_43509_21373.n8 90.436
R17426 a_43509_21373.n4 a_43509_21373.n7 50.575
R17427 a_43509_21373.n8 a_43509_21373.n4 74.302
R17428 a_43509_21373.n7 a_43509_21373.n6 157.665
R17429 a_43509_21373.n6 a_43509_21373.t4 8.7
R17430 a_43509_21373.n6 a_43509_21373.t7 8.7
R17431 a_43509_21373.n7 a_43509_21373.n5 122.999
R17432 a_43509_21373.n5 a_43509_21373.t3 14.282
R17433 a_43509_21373.n5 a_43509_21373.t2 14.282
R17434 a_43509_21373.n4 a_43509_21373.n3 90.416
R17435 a_43509_21373.n3 a_43509_21373.t1 14.282
R17436 a_43509_21373.n3 a_43509_21373.t6 14.282
R17437 a_43509_21373.n8 a_43509_21373.n1 3155.65
R17438 a_43509_21373.t8 a_43509_21373.n2 160.666
R17439 a_43509_21373.n1 a_43509_21373.t8 867.393
R17440 a_43509_21373.n2 a_43509_21373.t9 287.241
R17441 a_43509_21373.n2 a_43509_21373.t10 287.241
R17442 a_43509_21373.n1 a_43509_21373.t11 545.094
R17443 a_14498_15776.t0 a_14498_15776.t1 17.4
R17444 a_70459_5045.n2 a_70459_5045.t5 448.381
R17445 a_70459_5045.n1 a_70459_5045.t6 287.241
R17446 a_70459_5045.n1 a_70459_5045.t7 287.241
R17447 a_70459_5045.n0 a_70459_5045.t4 247.733
R17448 a_70459_5045.n4 a_70459_5045.n3 182.117
R17449 a_70459_5045.t5 a_70459_5045.n1 160.666
R17450 a_70459_5045.n3 a_70459_5045.t1 28.568
R17451 a_70459_5045.t2 a_70459_5045.n4 28.565
R17452 a_70459_5045.n4 a_70459_5045.t0 28.565
R17453 a_70459_5045.n0 a_70459_5045.t3 18.127
R17454 a_70459_5045.n2 a_70459_5045.n0 4.036
R17455 a_70459_5045.n3 a_70459_5045.n2 0.937
R17456 a_1089_11724.n0 a_1089_11724.n9 167.433
R17457 a_1089_11724.t0 a_1089_11724.n0 14.282
R17458 a_1089_11724.n0 a_1089_11724.t1 14.282
R17459 a_1089_11724.n9 a_1089_11724.n8 77.784
R17460 a_1089_11724.n8 a_1089_11724.n6 77.456
R17461 a_1089_11724.n6 a_1089_11724.n4 77.456
R17462 a_1089_11724.n4 a_1089_11724.n2 75.815
R17463 a_1089_11724.n9 a_1089_11724.t2 104.259
R17464 a_1089_11724.n8 a_1089_11724.n7 89.977
R17465 a_1089_11724.n7 a_1089_11724.t10 14.282
R17466 a_1089_11724.n7 a_1089_11724.t9 14.282
R17467 a_1089_11724.n6 a_1089_11724.n5 89.977
R17468 a_1089_11724.n5 a_1089_11724.t8 14.282
R17469 a_1089_11724.n5 a_1089_11724.t11 14.282
R17470 a_1089_11724.n4 a_1089_11724.n3 89.977
R17471 a_1089_11724.n3 a_1089_11724.t6 14.282
R17472 a_1089_11724.n3 a_1089_11724.t7 14.282
R17473 a_1089_11724.n2 a_1089_11724.t4 104.259
R17474 a_1089_11724.n2 a_1089_11724.n1 167.433
R17475 a_1089_11724.n1 a_1089_11724.t3 14.282
R17476 a_1089_11724.n1 a_1089_11724.t5 14.282
R17477 a_61189_3878.n0 a_61189_3878.t3 14.282
R17478 a_61189_3878.n0 a_61189_3878.t2 14.282
R17479 a_61189_3878.n1 a_61189_3878.t4 14.282
R17480 a_61189_3878.n1 a_61189_3878.t5 14.282
R17481 a_61189_3878.t0 a_61189_3878.n3 14.282
R17482 a_61189_3878.n3 a_61189_3878.t1 14.282
R17483 a_61189_3878.n3 a_61189_3878.n2 2.546
R17484 a_61189_3878.n2 a_61189_3878.n1 2.367
R17485 a_61189_3878.n2 a_61189_3878.n0 0.001
R17486 a_65224_7306.n1 a_65224_7306.t7 318.922
R17487 a_65224_7306.n0 a_65224_7306.t4 273.935
R17488 a_65224_7306.n0 a_65224_7306.t5 273.935
R17489 a_65224_7306.n1 a_65224_7306.t6 269.116
R17490 a_65224_7306.n4 a_65224_7306.n3 193.227
R17491 a_65224_7306.t7 a_65224_7306.n0 179.142
R17492 a_65224_7306.n2 a_65224_7306.n1 106.999
R17493 a_65224_7306.n3 a_65224_7306.t1 28.568
R17494 a_65224_7306.t0 a_65224_7306.n4 28.565
R17495 a_65224_7306.n4 a_65224_7306.t2 28.565
R17496 a_65224_7306.n2 a_65224_7306.t3 18.149
R17497 a_65224_7306.n3 a_65224_7306.n2 3.726
R17498 a_65651_6613.n0 a_65651_6613.n1 0.001
R17499 a_65651_6613.t0 a_65651_6613.n0 14.282
R17500 a_65651_6613.n0 a_65651_6613.t8 14.282
R17501 a_65651_6613.n1 a_65651_6613.n9 267.767
R17502 a_65651_6613.n9 a_65651_6613.t6 14.282
R17503 a_65651_6613.n9 a_65651_6613.t7 14.282
R17504 a_65651_6613.n1 a_65651_6613.n7 0.669
R17505 a_65651_6613.n7 a_65651_6613.n8 1.511
R17506 a_65651_6613.n8 a_65651_6613.t5 14.282
R17507 a_65651_6613.n8 a_65651_6613.t1 14.282
R17508 a_65651_6613.n7 a_65651_6613.n6 0.227
R17509 a_65651_6613.n6 a_65651_6613.n3 0.575
R17510 a_65651_6613.n6 a_65651_6613.n5 0.2
R17511 a_65651_6613.n5 a_65651_6613.t2 16.058
R17512 a_65651_6613.n5 a_65651_6613.n4 0.999
R17513 a_65651_6613.n4 a_65651_6613.t3 14.282
R17514 a_65651_6613.n4 a_65651_6613.t4 14.282
R17515 a_65651_6613.n3 a_65651_6613.n2 0.999
R17516 a_65651_6613.n2 a_65651_6613.t9 14.282
R17517 a_65651_6613.n2 a_65651_6613.t10 14.282
R17518 a_65651_6613.n3 a_65651_6613.t11 16.058
R17519 a_65769_6613.n1 a_65769_6613.t11 989.744
R17520 a_65769_6613.n7 a_65769_6613.n1 653.122
R17521 a_65769_6613.n1 a_65769_6613.t10 408.806
R17522 a_65769_6613.n0 a_65769_6613.t8 287.241
R17523 a_65769_6613.n0 a_65769_6613.t9 287.241
R17524 a_65769_6613.t11 a_65769_6613.n0 160.666
R17525 a_65769_6613.n5 a_65769_6613.n3 157.665
R17526 a_65769_6613.n5 a_65769_6613.n4 122.999
R17527 a_65769_6613.n8 a_65769_6613.n7 90.436
R17528 a_65769_6613.n6 a_65769_6613.n2 90.416
R17529 a_65769_6613.n7 a_65769_6613.n6 74.302
R17530 a_65769_6613.n6 a_65769_6613.n5 50.575
R17531 a_65769_6613.n2 a_65769_6613.t1 14.282
R17532 a_65769_6613.n2 a_65769_6613.t6 14.282
R17533 a_65769_6613.n4 a_65769_6613.t5 14.282
R17534 a_65769_6613.n4 a_65769_6613.t7 14.282
R17535 a_65769_6613.n8 a_65769_6613.t0 14.282
R17536 a_65769_6613.t2 a_65769_6613.n8 14.282
R17537 a_65769_6613.n3 a_65769_6613.t3 8.7
R17538 a_65769_6613.n3 a_65769_6613.t4 8.7
R17539 a_56366_23618.n6 a_56366_23618.n5 501.28
R17540 a_56366_23618.t6 a_56366_23618.t18 437.233
R17541 a_56366_23618.t5 a_56366_23618.t7 415.315
R17542 a_56366_23618.t16 a_56366_23618.n3 313.873
R17543 a_56366_23618.n5 a_56366_23618.t4 294.986
R17544 a_56366_23618.n2 a_56366_23618.t10 272.288
R17545 a_56366_23618.n6 a_56366_23618.t12 236.01
R17546 a_56366_23618.n9 a_56366_23618.t6 216.627
R17547 a_56366_23618.n7 a_56366_23618.t5 216.111
R17548 a_56366_23618.n8 a_56366_23618.t13 214.686
R17549 a_56366_23618.t18 a_56366_23618.n8 214.686
R17550 a_56366_23618.n1 a_56366_23618.t9 214.335
R17551 a_56366_23618.t7 a_56366_23618.n1 214.335
R17552 a_56366_23618.n4 a_56366_23618.t16 190.152
R17553 a_56366_23618.n4 a_56366_23618.t14 190.152
R17554 a_56366_23618.n2 a_56366_23618.t11 160.666
R17555 a_56366_23618.n3 a_56366_23618.t17 160.666
R17556 a_56366_23618.n7 a_56366_23618.n6 148.428
R17557 a_56366_23618.n5 a_56366_23618.t19 110.859
R17558 a_56366_23618.n3 a_56366_23618.n2 96.129
R17559 a_56366_23618.n8 a_56366_23618.t15 80.333
R17560 a_56366_23618.n1 a_56366_23618.t8 80.333
R17561 a_56366_23618.t12 a_56366_23618.n4 80.333
R17562 a_56366_23618.t2 a_56366_23618.n11 28.57
R17563 a_56366_23618.n0 a_56366_23618.t0 28.565
R17564 a_56366_23618.n0 a_56366_23618.t1 28.565
R17565 a_56366_23618.n11 a_56366_23618.t3 17.638
R17566 a_56366_23618.n10 a_56366_23618.n9 5.767
R17567 a_56366_23618.n9 a_56366_23618.n7 2.923
R17568 a_56366_23618.n10 a_56366_23618.n0 0.69
R17569 a_56366_23618.n11 a_56366_23618.n10 0.6
R17570 a_63350_20637.t0 a_63350_20637.t1 17.4
R17571 a_31377_4067.t0 a_31377_4067.t1 17.4
R17572 a_64192_n2074.n6 a_64192_n2074.n5 465.933
R17573 a_64192_n2074.t12 a_64192_n2074.t4 415.315
R17574 a_64192_n2074.n2 a_64192_n2074.t5 394.151
R17575 a_64192_n2074.n5 a_64192_n2074.t11 294.653
R17576 a_64192_n2074.n1 a_64192_n2074.t9 269.523
R17577 a_64192_n2074.t5 a_64192_n2074.n1 269.523
R17578 a_64192_n2074.n8 a_64192_n2074.t12 220.285
R17579 a_64192_n2074.n7 a_64192_n2074.t8 214.335
R17580 a_64192_n2074.t4 a_64192_n2074.n7 214.335
R17581 a_64192_n2074.n3 a_64192_n2074.t13 198.043
R17582 a_64192_n2074.n10 a_64192_n2074.n0 192.754
R17583 a_64192_n2074.n6 a_64192_n2074.n4 163.88
R17584 a_64192_n2074.n1 a_64192_n2074.t15 160.666
R17585 a_64192_n2074.n5 a_64192_n2074.t6 111.663
R17586 a_64192_n2074.n4 a_64192_n2074.n2 97.816
R17587 a_64192_n2074.n3 a_64192_n2074.t7 93.989
R17588 a_64192_n2074.n7 a_64192_n2074.t14 80.333
R17589 a_64192_n2074.n2 a_64192_n2074.t10 80.333
R17590 a_64192_n2074.n8 a_64192_n2074.n6 61.538
R17591 a_64192_n2074.t0 a_64192_n2074.n10 28.568
R17592 a_64192_n2074.n0 a_64192_n2074.t3 28.565
R17593 a_64192_n2074.n0 a_64192_n2074.t2 28.565
R17594 a_64192_n2074.n9 a_64192_n2074.t1 18.824
R17595 a_64192_n2074.n4 a_64192_n2074.n3 6.615
R17596 a_64192_n2074.n9 a_64192_n2074.n8 2.736
R17597 a_64192_n2074.n10 a_64192_n2074.n9 1.105
R17598 a_67135_n540.n0 a_67135_n540.t9 214.335
R17599 a_67135_n540.t7 a_67135_n540.n0 214.335
R17600 a_67135_n540.n1 a_67135_n540.t7 143.851
R17601 a_67135_n540.n1 a_67135_n540.t8 135.658
R17602 a_67135_n540.n0 a_67135_n540.t10 80.333
R17603 a_67135_n540.n2 a_67135_n540.t5 28.565
R17604 a_67135_n540.n2 a_67135_n540.t4 28.565
R17605 a_67135_n540.n4 a_67135_n540.t6 28.565
R17606 a_67135_n540.n4 a_67135_n540.t0 28.565
R17607 a_67135_n540.t2 a_67135_n540.n7 28.565
R17608 a_67135_n540.n7 a_67135_n540.t1 28.565
R17609 a_67135_n540.n6 a_67135_n540.t3 9.714
R17610 a_67135_n540.n7 a_67135_n540.n6 1.003
R17611 a_67135_n540.n5 a_67135_n540.n3 0.833
R17612 a_67135_n540.n3 a_67135_n540.n2 0.653
R17613 a_67135_n540.n5 a_67135_n540.n4 0.653
R17614 a_67135_n540.n6 a_67135_n540.n5 0.341
R17615 a_67135_n540.n3 a_67135_n540.n1 0.032
R17616 a_52674_17946.t6 a_52674_17946.n2 404.877
R17617 a_52674_17946.n1 a_52674_17946.t7 210.902
R17618 a_52674_17946.n3 a_52674_17946.t6 136.949
R17619 a_52674_17946.n2 a_52674_17946.n1 107.801
R17620 a_52674_17946.n1 a_52674_17946.t8 80.333
R17621 a_52674_17946.n2 a_52674_17946.t5 80.333
R17622 a_52674_17946.n0 a_52674_17946.t1 17.4
R17623 a_52674_17946.n0 a_52674_17946.t4 17.4
R17624 a_52674_17946.n4 a_52674_17946.t2 15.032
R17625 a_52674_17946.t0 a_52674_17946.n5 14.282
R17626 a_52674_17946.n5 a_52674_17946.t3 14.282
R17627 a_52674_17946.n5 a_52674_17946.n4 1.65
R17628 a_52674_17946.n3 a_52674_17946.n0 0.657
R17629 a_52674_17946.n4 a_52674_17946.n3 0.614
R17630 a_8011_13581.n2 a_8011_13581.t6 448.381
R17631 a_8011_13581.n1 a_8011_13581.t5 286.438
R17632 a_8011_13581.n1 a_8011_13581.t4 286.438
R17633 a_8011_13581.n0 a_8011_13581.t7 247.69
R17634 a_8011_13581.n4 a_8011_13581.n3 182.117
R17635 a_8011_13581.t6 a_8011_13581.n1 160.666
R17636 a_8011_13581.n3 a_8011_13581.t0 28.568
R17637 a_8011_13581.n4 a_8011_13581.t1 28.565
R17638 a_8011_13581.t2 a_8011_13581.n4 28.565
R17639 a_8011_13581.n0 a_8011_13581.t3 18.127
R17640 a_8011_13581.n2 a_8011_13581.n0 4.036
R17641 a_8011_13581.n3 a_8011_13581.n2 0.937
R17642 a_7365_14454.n4 a_7365_14454.n3 167.433
R17643 a_7365_14454.n9 a_7365_14454.n8 167.433
R17644 a_7365_14454.n8 a_7365_14454.t0 104.259
R17645 a_7365_14454.n4 a_7365_14454.t9 104.259
R17646 a_7365_14454.n7 a_7365_14454.n0 89.977
R17647 a_7365_14454.n6 a_7365_14454.n1 89.977
R17648 a_7365_14454.n5 a_7365_14454.n2 89.977
R17649 a_7365_14454.n5 a_7365_14454.n4 77.784
R17650 a_7365_14454.n7 a_7365_14454.n6 77.456
R17651 a_7365_14454.n6 a_7365_14454.n5 77.456
R17652 a_7365_14454.n8 a_7365_14454.n7 75.815
R17653 a_7365_14454.n0 a_7365_14454.t8 14.282
R17654 a_7365_14454.n0 a_7365_14454.t6 14.282
R17655 a_7365_14454.n1 a_7365_14454.t7 14.282
R17656 a_7365_14454.n1 a_7365_14454.t3 14.282
R17657 a_7365_14454.n2 a_7365_14454.t4 14.282
R17658 a_7365_14454.n2 a_7365_14454.t5 14.282
R17659 a_7365_14454.n3 a_7365_14454.t10 14.282
R17660 a_7365_14454.n3 a_7365_14454.t11 14.282
R17661 a_7365_14454.n9 a_7365_14454.t1 14.282
R17662 a_7365_14454.t2 a_7365_14454.n9 14.282
R17663 a_40724_17941.t5 a_40724_17941.n2 404.877
R17664 a_40724_17941.n1 a_40724_17941.t6 210.902
R17665 a_40724_17941.n3 a_40724_17941.t5 136.949
R17666 a_40724_17941.n2 a_40724_17941.n1 107.801
R17667 a_40724_17941.n1 a_40724_17941.t7 80.333
R17668 a_40724_17941.n2 a_40724_17941.t8 80.333
R17669 a_40724_17941.n0 a_40724_17941.t4 17.4
R17670 a_40724_17941.n0 a_40724_17941.t0 17.4
R17671 a_40724_17941.n4 a_40724_17941.t1 15.032
R17672 a_40724_17941.n5 a_40724_17941.t2 14.282
R17673 a_40724_17941.t3 a_40724_17941.n5 14.282
R17674 a_40724_17941.n5 a_40724_17941.n4 1.65
R17675 a_40724_17941.n3 a_40724_17941.n0 0.657
R17676 a_40724_17941.n4 a_40724_17941.n3 0.614
R17677 a_37903_748.n4 a_37903_748.t10 214.335
R17678 a_37903_748.t8 a_37903_748.n4 214.335
R17679 a_37903_748.n5 a_37903_748.t8 143.851
R17680 a_37903_748.n5 a_37903_748.t9 135.658
R17681 a_37903_748.n4 a_37903_748.t7 80.333
R17682 a_37903_748.n0 a_37903_748.t4 28.565
R17683 a_37903_748.n0 a_37903_748.t6 28.565
R17684 a_37903_748.n2 a_37903_748.t1 28.565
R17685 a_37903_748.n2 a_37903_748.t5 28.565
R17686 a_37903_748.t2 a_37903_748.n7 28.565
R17687 a_37903_748.n7 a_37903_748.t0 28.565
R17688 a_37903_748.n1 a_37903_748.t3 9.714
R17689 a_37903_748.n1 a_37903_748.n0 1.003
R17690 a_37903_748.n6 a_37903_748.n3 0.833
R17691 a_37903_748.n3 a_37903_748.n2 0.653
R17692 a_37903_748.n7 a_37903_748.n6 0.653
R17693 a_37903_748.n3 a_37903_748.n1 0.341
R17694 a_37903_748.n6 a_37903_748.n5 0.032
R17695 a_38493_311.t5 a_38493_311.t7 574.43
R17696 a_38493_311.n0 a_38493_311.t6 285.109
R17697 a_38493_311.n2 a_38493_311.n1 197.217
R17698 a_38493_311.n4 a_38493_311.n3 192.754
R17699 a_38493_311.n0 a_38493_311.t4 160.666
R17700 a_38493_311.n1 a_38493_311.t5 160.666
R17701 a_38493_311.n1 a_38493_311.n0 114.829
R17702 a_38493_311.n3 a_38493_311.t0 28.568
R17703 a_38493_311.t2 a_38493_311.n4 28.565
R17704 a_38493_311.n4 a_38493_311.t1 28.565
R17705 a_38493_311.n2 a_38493_311.t3 18.838
R17706 a_38493_311.n3 a_38493_311.n2 1.129
R17707 a_47912_3876.n1 a_47912_3876.t1 14.282
R17708 a_47912_3876.n1 a_47912_3876.t5 14.282
R17709 a_47912_3876.n0 a_47912_3876.t4 14.282
R17710 a_47912_3876.n0 a_47912_3876.t3 14.282
R17711 a_47912_3876.n3 a_47912_3876.t0 14.282
R17712 a_47912_3876.t2 a_47912_3876.n3 14.282
R17713 a_47912_3876.n2 a_47912_3876.n0 2.546
R17714 a_47912_3876.n3 a_47912_3876.n2 2.367
R17715 a_47912_3876.n2 a_47912_3876.n1 0.001
R17716 a_14367_8119.n2 a_14367_8119.t7 448.381
R17717 a_14367_8119.n1 a_14367_8119.t4 286.438
R17718 a_14367_8119.n1 a_14367_8119.t5 286.438
R17719 a_14367_8119.n0 a_14367_8119.t6 247.69
R17720 a_14367_8119.n4 a_14367_8119.n3 182.117
R17721 a_14367_8119.t7 a_14367_8119.n1 160.666
R17722 a_14367_8119.n3 a_14367_8119.t1 28.568
R17723 a_14367_8119.n4 a_14367_8119.t0 28.565
R17724 a_14367_8119.t2 a_14367_8119.n4 28.565
R17725 a_14367_8119.n0 a_14367_8119.t3 18.127
R17726 a_14367_8119.n2 a_14367_8119.n0 4.036
R17727 a_14367_8119.n3 a_14367_8119.n2 0.937
R17728 a_60758_18575.t7 a_60758_18575.t4 574.43
R17729 a_60758_18575.n1 a_60758_18575.t5 285.109
R17730 a_60758_18575.n3 a_60758_18575.n2 197.215
R17731 a_60758_18575.n4 a_60758_18575.n0 192.754
R17732 a_60758_18575.n1 a_60758_18575.t6 160.666
R17733 a_60758_18575.n2 a_60758_18575.t7 160.666
R17734 a_60758_18575.n2 a_60758_18575.n1 114.829
R17735 a_60758_18575.t0 a_60758_18575.n4 28.568
R17736 a_60758_18575.n0 a_60758_18575.t3 28.565
R17737 a_60758_18575.n0 a_60758_18575.t1 28.565
R17738 a_60758_18575.n3 a_60758_18575.t2 18.838
R17739 a_60758_18575.n4 a_60758_18575.n3 1.129
R17740 a_60329_17945.t5 a_60329_17945.n3 404.877
R17741 a_60329_17945.n2 a_60329_17945.t6 210.902
R17742 a_60329_17945.n4 a_60329_17945.t5 136.949
R17743 a_60329_17945.n3 a_60329_17945.n2 107.801
R17744 a_60329_17945.n2 a_60329_17945.t7 80.333
R17745 a_60329_17945.n3 a_60329_17945.t8 80.333
R17746 a_60329_17945.n1 a_60329_17945.t0 17.4
R17747 a_60329_17945.n1 a_60329_17945.t4 17.4
R17748 a_60329_17945.t1 a_60329_17945.n5 15.032
R17749 a_60329_17945.n0 a_60329_17945.t2 14.282
R17750 a_60329_17945.n0 a_60329_17945.t3 14.282
R17751 a_60329_17945.n5 a_60329_17945.n0 1.65
R17752 a_60329_17945.n4 a_60329_17945.n1 0.657
R17753 a_60329_17945.n5 a_60329_17945.n4 0.614
R17754 a_20515_5324.n2 a_20515_5324.t4 318.922
R17755 a_20515_5324.n1 a_20515_5324.t6 273.935
R17756 a_20515_5324.n1 a_20515_5324.t7 273.935
R17757 a_20515_5324.n2 a_20515_5324.t5 269.116
R17758 a_20515_5324.n4 a_20515_5324.n0 193.227
R17759 a_20515_5324.t4 a_20515_5324.n1 179.142
R17760 a_20515_5324.n3 a_20515_5324.n2 106.999
R17761 a_20515_5324.t2 a_20515_5324.n4 28.568
R17762 a_20515_5324.n0 a_20515_5324.t0 28.565
R17763 a_20515_5324.n0 a_20515_5324.t1 28.565
R17764 a_20515_5324.n3 a_20515_5324.t3 18.149
R17765 a_20515_5324.n4 a_20515_5324.n3 3.726
R17766 a_52460_1734.n1 a_52460_1734.t5 318.922
R17767 a_52460_1734.n0 a_52460_1734.t4 273.935
R17768 a_52460_1734.n0 a_52460_1734.t6 273.935
R17769 a_52460_1734.n1 a_52460_1734.t7 269.116
R17770 a_52460_1734.n4 a_52460_1734.n3 193.227
R17771 a_52460_1734.t5 a_52460_1734.n0 179.142
R17772 a_52460_1734.n2 a_52460_1734.n1 106.999
R17773 a_52460_1734.n3 a_52460_1734.t1 28.568
R17774 a_52460_1734.n4 a_52460_1734.t0 28.565
R17775 a_52460_1734.t2 a_52460_1734.n4 28.565
R17776 a_52460_1734.n2 a_52460_1734.t3 18.149
R17777 a_52460_1734.n3 a_52460_1734.n2 3.726
R17778 a_22526_4620.t0 a_22526_4620.t1 17.4
R17779 a_37902_9782.n0 a_37902_9782.t9 214.335
R17780 a_37902_9782.t7 a_37902_9782.n0 214.335
R17781 a_37902_9782.n1 a_37902_9782.t7 143.851
R17782 a_37902_9782.n1 a_37902_9782.t8 135.658
R17783 a_37902_9782.n0 a_37902_9782.t10 80.333
R17784 a_37902_9782.n2 a_37902_9782.t5 28.565
R17785 a_37902_9782.n2 a_37902_9782.t4 28.565
R17786 a_37902_9782.n4 a_37902_9782.t6 28.565
R17787 a_37902_9782.n4 a_37902_9782.t1 28.565
R17788 a_37902_9782.t3 a_37902_9782.n7 28.565
R17789 a_37902_9782.n7 a_37902_9782.t2 28.565
R17790 a_37902_9782.n6 a_37902_9782.t0 9.714
R17791 a_37902_9782.n7 a_37902_9782.n6 1.003
R17792 a_37902_9782.n5 a_37902_9782.n3 0.833
R17793 a_37902_9782.n3 a_37902_9782.n2 0.653
R17794 a_37902_9782.n5 a_37902_9782.n4 0.653
R17795 a_37902_9782.n6 a_37902_9782.n5 0.341
R17796 a_37902_9782.n3 a_37902_9782.n1 0.032
R17797 a_7551_6363.n1 a_7551_6363.t7 990.34
R17798 a_7551_6363.n1 a_7551_6363.t4 408.211
R17799 a_7551_6363.n0 a_7551_6363.t5 286.438
R17800 a_7551_6363.n0 a_7551_6363.t6 286.438
R17801 a_7551_6363.n4 a_7551_6363.n3 192.754
R17802 a_7551_6363.t7 a_7551_6363.n0 160.666
R17803 a_7551_6363.n2 a_7551_6363.n1 44.149
R17804 a_7551_6363.n3 a_7551_6363.t0 28.568
R17805 a_7551_6363.t2 a_7551_6363.n4 28.565
R17806 a_7551_6363.n4 a_7551_6363.t1 28.565
R17807 a_7551_6363.n2 a_7551_6363.t3 18.09
R17808 a_7551_6363.n3 a_7551_6363.n2 0.478
R17809 a_11110_7655.t0 a_11110_7655.t1 17.4
R17810 a_9986_8258.t5 a_9986_8258.n0 14.282
R17811 a_9986_8258.n0 a_9986_8258.t7 14.282
R17812 a_9986_8258.n0 a_9986_8258.n1 258.161
R17813 a_9986_8258.n1 a_9986_8258.n5 0.852
R17814 a_9986_8258.n5 a_9986_8258.n6 4.366
R17815 a_9986_8258.n6 a_9986_8258.n7 258.161
R17816 a_9986_8258.n7 a_9986_8258.t1 14.282
R17817 a_9986_8258.n7 a_9986_8258.t2 14.282
R17818 a_9986_8258.n6 a_9986_8258.t0 14.283
R17819 a_9986_8258.n5 a_9986_8258.n4 97.614
R17820 a_9986_8258.n4 a_9986_8258.t9 200.029
R17821 a_9986_8258.t9 a_9986_8258.n3 206.421
R17822 a_9986_8258.n3 a_9986_8258.t11 80.333
R17823 a_9986_8258.n3 a_9986_8258.t10 206.421
R17824 a_9986_8258.n4 a_9986_8258.t8 1527.4
R17825 a_9986_8258.t8 a_9986_8258.n2 657.379
R17826 a_9986_8258.n2 a_9986_8258.t3 8.7
R17827 a_9986_8258.n2 a_9986_8258.t4 8.7
R17828 a_9986_8258.n1 a_9986_8258.t6 14.283
R17829 a_4233_11724.t3 a_4233_11724.n9 104.259
R17830 a_4233_11724.n6 a_4233_11724.n7 77.784
R17831 a_4233_11724.n4 a_4233_11724.n6 77.456
R17832 a_4233_11724.n2 a_4233_11724.n4 77.456
R17833 a_4233_11724.n9 a_4233_11724.n2 75.815
R17834 a_4233_11724.n7 a_4233_11724.n8 167.433
R17835 a_4233_11724.n8 a_4233_11724.t1 14.282
R17836 a_4233_11724.n8 a_4233_11724.t0 14.282
R17837 a_4233_11724.n7 a_4233_11724.t2 104.259
R17838 a_4233_11724.n6 a_4233_11724.n5 89.977
R17839 a_4233_11724.n5 a_4233_11724.t11 14.282
R17840 a_4233_11724.n5 a_4233_11724.t10 14.282
R17841 a_4233_11724.n4 a_4233_11724.n3 89.977
R17842 a_4233_11724.n3 a_4233_11724.t9 14.282
R17843 a_4233_11724.n3 a_4233_11724.t6 14.282
R17844 a_4233_11724.n2 a_4233_11724.n1 89.977
R17845 a_4233_11724.n1 a_4233_11724.t5 14.282
R17846 a_4233_11724.n1 a_4233_11724.t4 14.282
R17847 a_4233_11724.n9 a_4233_11724.n0 167.433
R17848 a_4233_11724.n0 a_4233_11724.t7 14.282
R17849 a_4233_11724.n0 a_4233_11724.t8 14.282
R17850 a_41161_15765.t0 a_41161_15765.n0 14.282
R17851 a_41161_15765.n0 a_41161_15765.t1 14.282
R17852 a_41161_15765.n0 a_41161_15765.n9 0.999
R17853 a_41161_15765.n9 a_41161_15765.n6 0.2
R17854 a_41161_15765.n6 a_41161_15765.n8 0.575
R17855 a_41161_15765.n8 a_41161_15765.t5 16.058
R17856 a_41161_15765.n8 a_41161_15765.n7 0.999
R17857 a_41161_15765.n7 a_41161_15765.t6 14.282
R17858 a_41161_15765.n7 a_41161_15765.t11 14.282
R17859 a_41161_15765.n9 a_41161_15765.t7 16.058
R17860 a_41161_15765.n6 a_41161_15765.n4 0.227
R17861 a_41161_15765.n4 a_41161_15765.n5 1.511
R17862 a_41161_15765.n5 a_41161_15765.t3 14.282
R17863 a_41161_15765.n5 a_41161_15765.t2 14.282
R17864 a_41161_15765.n4 a_41161_15765.n1 0.669
R17865 a_41161_15765.n1 a_41161_15765.n2 0.001
R17866 a_41161_15765.n1 a_41161_15765.n3 267.767
R17867 a_41161_15765.n3 a_41161_15765.t10 14.282
R17868 a_41161_15765.n3 a_41161_15765.t9 14.282
R17869 a_41161_15765.n2 a_41161_15765.t8 14.282
R17870 a_41161_15765.n2 a_41161_15765.t4 14.282
R17871 a_70459_20811.n2 a_70459_20811.t5 448.381
R17872 a_70459_20811.n1 a_70459_20811.t7 287.241
R17873 a_70459_20811.n1 a_70459_20811.t4 287.241
R17874 a_70459_20811.n0 a_70459_20811.t6 247.733
R17875 a_70459_20811.n4 a_70459_20811.n3 182.117
R17876 a_70459_20811.t5 a_70459_20811.n1 160.666
R17877 a_70459_20811.n3 a_70459_20811.t0 28.568
R17878 a_70459_20811.n4 a_70459_20811.t1 28.565
R17879 a_70459_20811.t2 a_70459_20811.n4 28.565
R17880 a_70459_20811.n0 a_70459_20811.t3 18.127
R17881 a_70459_20811.n2 a_70459_20811.n0 4.036
R17882 a_70459_20811.n3 a_70459_20811.n2 0.937
R17883 a_61178_15743.n1 a_61178_15743.t6 318.922
R17884 a_61178_15743.n0 a_61178_15743.t5 273.935
R17885 a_61178_15743.n0 a_61178_15743.t7 273.935
R17886 a_61178_15743.n1 a_61178_15743.t4 269.116
R17887 a_61178_15743.n4 a_61178_15743.n3 193.227
R17888 a_61178_15743.t6 a_61178_15743.n0 179.142
R17889 a_61178_15743.n2 a_61178_15743.n1 106.999
R17890 a_61178_15743.n3 a_61178_15743.t0 28.568
R17891 a_61178_15743.n4 a_61178_15743.t1 28.565
R17892 a_61178_15743.t2 a_61178_15743.n4 28.565
R17893 a_61178_15743.n2 a_61178_15743.t3 18.149
R17894 a_61178_15743.n3 a_61178_15743.n2 3.726
R17895 a_65651_n1230.t0 a_65651_n1230.n0 14.282
R17896 a_65651_n1230.n0 a_65651_n1230.t1 14.282
R17897 a_65651_n1230.n0 a_65651_n1230.n9 0.999
R17898 a_65651_n1230.n9 a_65651_n1230.n6 0.575
R17899 a_65651_n1230.n6 a_65651_n1230.n8 0.2
R17900 a_65651_n1230.n8 a_65651_n1230.t2 16.058
R17901 a_65651_n1230.n8 a_65651_n1230.n7 0.999
R17902 a_65651_n1230.n7 a_65651_n1230.t7 14.282
R17903 a_65651_n1230.n7 a_65651_n1230.t8 14.282
R17904 a_65651_n1230.n9 a_65651_n1230.t3 16.058
R17905 a_65651_n1230.n6 a_65651_n1230.n4 0.227
R17906 a_65651_n1230.n4 a_65651_n1230.n5 1.511
R17907 a_65651_n1230.n5 a_65651_n1230.t11 14.282
R17908 a_65651_n1230.n5 a_65651_n1230.t9 14.282
R17909 a_65651_n1230.n4 a_65651_n1230.n1 0.669
R17910 a_65651_n1230.n1 a_65651_n1230.n2 0.001
R17911 a_65651_n1230.n1 a_65651_n1230.n3 267.767
R17912 a_65651_n1230.n3 a_65651_n1230.t4 14.282
R17913 a_65651_n1230.n3 a_65651_n1230.t5 14.282
R17914 a_65651_n1230.n2 a_65651_n1230.t10 14.282
R17915 a_65651_n1230.n2 a_65651_n1230.t6 14.282
R17916 a_31377_n306.t0 a_31377_n306.t1 379.845
R17917 a_9700_n2148.n3 a_9700_n2148.t6 448.382
R17918 a_9700_n2148.n2 a_9700_n2148.t5 286.438
R17919 a_9700_n2148.n2 a_9700_n2148.t7 286.438
R17920 a_9700_n2148.n1 a_9700_n2148.t4 247.69
R17921 a_9700_n2148.n4 a_9700_n2148.n0 182.117
R17922 a_9700_n2148.t6 a_9700_n2148.n2 160.666
R17923 a_9700_n2148.t2 a_9700_n2148.n4 28.568
R17924 a_9700_n2148.n0 a_9700_n2148.t0 28.565
R17925 a_9700_n2148.n0 a_9700_n2148.t1 28.565
R17926 a_9700_n2148.n1 a_9700_n2148.t3 18.127
R17927 a_9700_n2148.n3 a_9700_n2148.n1 4.039
R17928 a_9700_n2148.n4 a_9700_n2148.n3 0.937
R17929 a_10608_n2148.t0 a_10608_n2148.n0 14.283
R17930 a_10608_n2148.n0 a_10608_n2148.n7 258.161
R17931 a_10608_n2148.n7 a_10608_n2148.t1 14.282
R17932 a_10608_n2148.n7 a_10608_n2148.t2 14.282
R17933 a_10608_n2148.n0 a_10608_n2148.n4 0.852
R17934 a_10608_n2148.n4 a_10608_n2148.n5 4.366
R17935 a_10608_n2148.n5 a_10608_n2148.n6 258.161
R17936 a_10608_n2148.n6 a_10608_n2148.t5 14.282
R17937 a_10608_n2148.n6 a_10608_n2148.t4 14.282
R17938 a_10608_n2148.n5 a_10608_n2148.t6 14.283
R17939 a_10608_n2148.n4 a_10608_n2148.n3 97.614
R17940 a_10608_n2148.n3 a_10608_n2148.t8 200.029
R17941 a_10608_n2148.t8 a_10608_n2148.n2 206.421
R17942 a_10608_n2148.n2 a_10608_n2148.t9 80.333
R17943 a_10608_n2148.n2 a_10608_n2148.t10 206.421
R17944 a_10608_n2148.n3 a_10608_n2148.t11 1527.4
R17945 a_10608_n2148.t11 a_10608_n2148.n1 657.379
R17946 a_10608_n2148.n1 a_10608_n2148.t7 8.7
R17947 a_10608_n2148.n1 a_10608_n2148.t3 8.7
R17948 a_11080_n3481.t0 a_11080_n3481.t1 17.4
R17949 a_4804_n3485.t0 a_4804_n3485.t1 17.4
R17950 a_59262_18579.t5 a_59262_18579.t4 800.071
R17951 a_59262_18579.n3 a_59262_18579.n2 672.95
R17952 a_59262_18579.n1 a_59262_18579.t6 285.109
R17953 a_59262_18579.n2 a_59262_18579.t5 193.602
R17954 a_59262_18579.n1 a_59262_18579.t7 160.666
R17955 a_59262_18579.n2 a_59262_18579.n1 91.507
R17956 a_59262_18579.n0 a_59262_18579.t0 28.57
R17957 a_59262_18579.n4 a_59262_18579.t1 28.565
R17958 a_59262_18579.t2 a_59262_18579.n4 28.565
R17959 a_59262_18579.n0 a_59262_18579.t3 17.638
R17960 a_59262_18579.n4 a_59262_18579.n3 0.693
R17961 a_59262_18579.n3 a_59262_18579.n0 0.597
R17962 a_47800_9746.t8 a_47800_9746.n3 404.877
R17963 a_47800_9746.n2 a_47800_9746.t6 210.902
R17964 a_47800_9746.n4 a_47800_9746.t8 136.943
R17965 a_47800_9746.n3 a_47800_9746.n2 107.801
R17966 a_47800_9746.n2 a_47800_9746.t7 80.333
R17967 a_47800_9746.n3 a_47800_9746.t5 80.333
R17968 a_47800_9746.n1 a_47800_9746.t0 17.4
R17969 a_47800_9746.n1 a_47800_9746.t2 17.4
R17970 a_47800_9746.t1 a_47800_9746.n5 15.032
R17971 a_47800_9746.n0 a_47800_9746.t4 14.282
R17972 a_47800_9746.n0 a_47800_9746.t3 14.282
R17973 a_47800_9746.n5 a_47800_9746.n0 1.65
R17974 a_47800_9746.n4 a_47800_9746.n1 0.672
R17975 a_47800_9746.n5 a_47800_9746.n4 0.665
R17976 a_48064_9163.n5 a_48064_9163.n4 535.449
R17977 a_48064_9163.t5 a_48064_9163.t18 437.233
R17978 a_48064_9163.t19 a_48064_9163.t6 437.233
R17979 a_48064_9163.t15 a_48064_9163.n2 313.873
R17980 a_48064_9163.n4 a_48064_9163.t12 294.986
R17981 a_48064_9163.n1 a_48064_9163.t4 272.288
R17982 a_48064_9163.n5 a_48064_9163.t9 245.184
R17983 a_48064_9163.n7 a_48064_9163.t19 218.628
R17984 a_48064_9163.n9 a_48064_9163.t5 217.024
R17985 a_48064_9163.n8 a_48064_9163.t17 214.686
R17986 a_48064_9163.t18 a_48064_9163.n8 214.686
R17987 a_48064_9163.n6 a_48064_9163.t13 214.686
R17988 a_48064_9163.t6 a_48064_9163.n6 214.686
R17989 a_48064_9163.n3 a_48064_9163.t15 190.152
R17990 a_48064_9163.n3 a_48064_9163.t10 190.152
R17991 a_48064_9163.n1 a_48064_9163.t16 160.666
R17992 a_48064_9163.n2 a_48064_9163.t11 160.666
R17993 a_48064_9163.n4 a_48064_9163.t14 110.859
R17994 a_48064_9163.n2 a_48064_9163.n1 96.129
R17995 a_48064_9163.n8 a_48064_9163.t7 80.333
R17996 a_48064_9163.t9 a_48064_9163.n3 80.333
R17997 a_48064_9163.n6 a_48064_9163.t8 80.333
R17998 a_48064_9163.t2 a_48064_9163.n11 28.57
R17999 a_48064_9163.n0 a_48064_9163.t1 28.565
R18000 a_48064_9163.n0 a_48064_9163.t0 28.565
R18001 a_48064_9163.n11 a_48064_9163.t3 17.638
R18002 a_48064_9163.n7 a_48064_9163.n5 14.9
R18003 a_48064_9163.n10 a_48064_9163.n9 8.819
R18004 a_48064_9163.n9 a_48064_9163.n7 2.599
R18005 a_48064_9163.n10 a_48064_9163.n0 0.69
R18006 a_48064_9163.n11 a_48064_9163.n10 0.6
R18007 a_38498_1915.t6 a_38498_1915.t4 574.43
R18008 a_38498_1915.n0 a_38498_1915.t7 285.109
R18009 a_38498_1915.n2 a_38498_1915.n1 211.136
R18010 a_38498_1915.n4 a_38498_1915.n3 192.754
R18011 a_38498_1915.n0 a_38498_1915.t5 160.666
R18012 a_38498_1915.n1 a_38498_1915.t6 160.666
R18013 a_38498_1915.n1 a_38498_1915.n0 114.829
R18014 a_38498_1915.n3 a_38498_1915.t1 28.568
R18015 a_38498_1915.n4 a_38498_1915.t0 28.565
R18016 a_38498_1915.t2 a_38498_1915.n4 28.565
R18017 a_38498_1915.n2 a_38498_1915.t3 19.084
R18018 a_38498_1915.n3 a_38498_1915.n2 1.051
R18019 a_3058_20866.t5 a_3058_20866.n0 14.282
R18020 a_3058_20866.n0 a_3058_20866.t6 14.282
R18021 a_3058_20866.n0 a_3058_20866.n1 258.161
R18022 a_3058_20866.n1 a_3058_20866.t7 14.283
R18023 a_3058_20866.n1 a_3058_20866.n7 4.366
R18024 a_3058_20866.n7 a_3058_20866.n5 0.852
R18025 a_3058_20866.n5 a_3058_20866.n6 258.161
R18026 a_3058_20866.n6 a_3058_20866.t2 14.282
R18027 a_3058_20866.n6 a_3058_20866.t1 14.282
R18028 a_3058_20866.n5 a_3058_20866.t3 14.283
R18029 a_3058_20866.n7 a_3058_20866.n4 97.614
R18030 a_3058_20866.n4 a_3058_20866.t9 200.029
R18031 a_3058_20866.t9 a_3058_20866.n3 206.421
R18032 a_3058_20866.n3 a_3058_20866.t10 80.333
R18033 a_3058_20866.n3 a_3058_20866.t11 206.421
R18034 a_3058_20866.n4 a_3058_20866.t8 1527.4
R18035 a_3058_20866.t8 a_3058_20866.n2 657.379
R18036 a_3058_20866.n2 a_3058_20866.t4 8.7
R18037 a_3058_20866.n2 a_3058_20866.t0 8.7
R18038 a_55197_1015.n1 a_55197_1015.t5 318.922
R18039 a_55197_1015.n0 a_55197_1015.t6 274.739
R18040 a_55197_1015.n0 a_55197_1015.t7 274.739
R18041 a_55197_1015.n1 a_55197_1015.t4 269.116
R18042 a_55197_1015.t5 a_55197_1015.n0 179.946
R18043 a_55197_1015.n2 a_55197_1015.n1 105.178
R18044 a_55197_1015.n3 a_55197_1015.t1 29.444
R18045 a_55197_1015.n4 a_55197_1015.t0 28.565
R18046 a_55197_1015.t2 a_55197_1015.n4 28.565
R18047 a_55197_1015.n2 a_55197_1015.t3 18.145
R18048 a_55197_1015.n3 a_55197_1015.n2 2.878
R18049 a_55197_1015.n4 a_55197_1015.n3 0.764
R18050 a_54903_309.t0 a_54903_309.t1 380.209
R18051 a_45805_1733.n1 a_45805_1733.t5 318.922
R18052 a_45805_1733.n0 a_45805_1733.t7 273.935
R18053 a_45805_1733.n0 a_45805_1733.t6 273.935
R18054 a_45805_1733.n1 a_45805_1733.t4 269.116
R18055 a_45805_1733.n4 a_45805_1733.n3 193.227
R18056 a_45805_1733.t5 a_45805_1733.n0 179.142
R18057 a_45805_1733.n2 a_45805_1733.n1 106.999
R18058 a_45805_1733.n3 a_45805_1733.t0 28.568
R18059 a_45805_1733.t2 a_45805_1733.n4 28.565
R18060 a_45805_1733.n4 a_45805_1733.t1 28.565
R18061 a_45805_1733.n2 a_45805_1733.t3 18.149
R18062 a_45805_1733.n3 a_45805_1733.n2 3.726
R18063 a_46350_308.t0 a_46350_308.t1 380.209
R18064 a_46350_1040.n0 a_46350_1040.n12 122.999
R18065 a_46350_1040.t0 a_46350_1040.n0 14.282
R18066 a_46350_1040.n0 a_46350_1040.t2 14.282
R18067 a_46350_1040.n12 a_46350_1040.n10 50.575
R18068 a_46350_1040.n10 a_46350_1040.n8 74.302
R18069 a_46350_1040.n12 a_46350_1040.n11 157.665
R18070 a_46350_1040.n11 a_46350_1040.t3 8.7
R18071 a_46350_1040.n11 a_46350_1040.t4 8.7
R18072 a_46350_1040.n10 a_46350_1040.n9 90.416
R18073 a_46350_1040.n9 a_46350_1040.t1 14.282
R18074 a_46350_1040.n9 a_46350_1040.t5 14.282
R18075 a_46350_1040.n8 a_46350_1040.n7 90.436
R18076 a_46350_1040.n7 a_46350_1040.t7 14.282
R18077 a_46350_1040.n7 a_46350_1040.t6 14.282
R18078 a_46350_1040.n8 a_46350_1040.n1 342.688
R18079 a_46350_1040.n1 a_46350_1040.n6 126.566
R18080 a_46350_1040.n6 a_46350_1040.t9 294.653
R18081 a_46350_1040.n6 a_46350_1040.t13 111.663
R18082 a_46350_1040.n1 a_46350_1040.n5 552.333
R18083 a_46350_1040.n5 a_46350_1040.n4 6.615
R18084 a_46350_1040.n4 a_46350_1040.t15 93.989
R18085 a_46350_1040.n5 a_46350_1040.n3 97.816
R18086 a_46350_1040.n3 a_46350_1040.t12 80.333
R18087 a_46350_1040.n3 a_46350_1040.t8 394.151
R18088 a_46350_1040.t8 a_46350_1040.n2 269.523
R18089 a_46350_1040.n2 a_46350_1040.t14 160.666
R18090 a_46350_1040.n2 a_46350_1040.t11 269.523
R18091 a_46350_1040.n4 a_46350_1040.t10 198.043
R18092 a_46650_6884.n1 a_46650_6884.t7 318.922
R18093 a_46650_6884.n0 a_46650_6884.t5 274.739
R18094 a_46650_6884.n0 a_46650_6884.t6 274.739
R18095 a_46650_6884.n1 a_46650_6884.t4 269.116
R18096 a_46650_6884.t7 a_46650_6884.n0 179.946
R18097 a_46650_6884.n2 a_46650_6884.n1 107.263
R18098 a_46650_6884.t0 a_46650_6884.n4 29.444
R18099 a_46650_6884.n3 a_46650_6884.t3 28.565
R18100 a_46650_6884.n3 a_46650_6884.t2 28.565
R18101 a_46650_6884.n2 a_46650_6884.t1 18.145
R18102 a_46650_6884.n4 a_46650_6884.n2 2.878
R18103 a_46650_6884.n4 a_46650_6884.n3 0.764
R18104 a_46356_6178.t0 a_46356_6178.t1 380.209
R18105 a_62361_17053.n0 a_62361_17053.t8 214.335
R18106 a_62361_17053.t10 a_62361_17053.n0 214.335
R18107 a_62361_17053.n1 a_62361_17053.t10 143.851
R18108 a_62361_17053.n1 a_62361_17053.t7 135.658
R18109 a_62361_17053.n0 a_62361_17053.t9 80.333
R18110 a_62361_17053.n2 a_62361_17053.t4 28.565
R18111 a_62361_17053.n2 a_62361_17053.t5 28.565
R18112 a_62361_17053.n4 a_62361_17053.t6 28.565
R18113 a_62361_17053.n4 a_62361_17053.t0 28.565
R18114 a_62361_17053.n7 a_62361_17053.t1 28.565
R18115 a_62361_17053.t2 a_62361_17053.n7 28.565
R18116 a_62361_17053.n3 a_62361_17053.t3 9.714
R18117 a_62361_17053.n3 a_62361_17053.n2 1.003
R18118 a_62361_17053.n6 a_62361_17053.n5 0.833
R18119 a_62361_17053.n5 a_62361_17053.n4 0.653
R18120 a_62361_17053.n7 a_62361_17053.n6 0.653
R18121 a_62361_17053.n5 a_62361_17053.n3 0.341
R18122 a_62361_17053.n6 a_62361_17053.n1 0.032
R18123 a_59616_18579.t7 a_59616_18579.t4 574.43
R18124 a_59616_18579.n1 a_59616_18579.t5 285.109
R18125 a_59616_18579.n3 a_59616_18579.n2 211.134
R18126 a_59616_18579.n4 a_59616_18579.n0 192.754
R18127 a_59616_18579.n1 a_59616_18579.t6 160.666
R18128 a_59616_18579.n2 a_59616_18579.t7 160.666
R18129 a_59616_18579.n2 a_59616_18579.n1 114.829
R18130 a_59616_18579.t2 a_59616_18579.n4 28.568
R18131 a_59616_18579.n0 a_59616_18579.t0 28.565
R18132 a_59616_18579.n0 a_59616_18579.t1 28.565
R18133 a_59616_18579.n3 a_59616_18579.t3 19.087
R18134 a_59616_18579.n4 a_59616_18579.n3 1.051
R18135 a_23081_8962.n0 a_23081_8962.t1 14.282
R18136 a_23081_8962.t0 a_23081_8962.n0 14.282
R18137 a_23081_8962.n0 a_23081_8962.n8 122.747
R18138 a_23081_8962.n4 a_23081_8962.n6 74.302
R18139 a_23081_8962.n8 a_23081_8962.n4 50.575
R18140 a_23081_8962.n8 a_23081_8962.n7 157.665
R18141 a_23081_8962.n7 a_23081_8962.t4 8.7
R18142 a_23081_8962.n7 a_23081_8962.t2 8.7
R18143 a_23081_8962.n6 a_23081_8962.n5 90.436
R18144 a_23081_8962.n5 a_23081_8962.t6 14.282
R18145 a_23081_8962.n5 a_23081_8962.t7 14.282
R18146 a_23081_8962.n4 a_23081_8962.n3 90.416
R18147 a_23081_8962.n3 a_23081_8962.t5 14.282
R18148 a_23081_8962.n3 a_23081_8962.t3 14.282
R18149 a_23081_8962.n6 a_23081_8962.n1 1297.45
R18150 a_23081_8962.n1 a_23081_8962.t11 591.811
R18151 a_23081_8962.n1 a_23081_8962.t10 867.497
R18152 a_23081_8962.t10 a_23081_8962.n2 160.666
R18153 a_23081_8962.n2 a_23081_8962.t8 286.438
R18154 a_23081_8962.n2 a_23081_8962.t9 286.438
R18155 a_22608_8258.n0 a_22608_8258.t2 14.282
R18156 a_22608_8258.t1 a_22608_8258.n0 14.282
R18157 a_22608_8258.n0 a_22608_8258.n1 258.161
R18158 a_22608_8258.n1 a_22608_8258.t3 14.283
R18159 a_22608_8258.n1 a_22608_8258.n7 4.366
R18160 a_22608_8258.n7 a_22608_8258.n5 0.852
R18161 a_22608_8258.n5 a_22608_8258.n6 258.161
R18162 a_22608_8258.n6 a_22608_8258.t5 14.282
R18163 a_22608_8258.n6 a_22608_8258.t7 14.282
R18164 a_22608_8258.n5 a_22608_8258.t6 14.283
R18165 a_22608_8258.n7 a_22608_8258.n4 97.614
R18166 a_22608_8258.n4 a_22608_8258.t9 200.029
R18167 a_22608_8258.t9 a_22608_8258.n3 206.421
R18168 a_22608_8258.n3 a_22608_8258.t8 80.333
R18169 a_22608_8258.n3 a_22608_8258.t11 206.421
R18170 a_22608_8258.n4 a_22608_8258.t10 1527.4
R18171 a_22608_8258.t10 a_22608_8258.n2 657.379
R18172 a_22608_8258.n2 a_22608_8258.t4 8.7
R18173 a_22608_8258.n2 a_22608_8258.t0 8.7
R18174 a_23141_8988.n3 a_23141_8988.n2 167.433
R18175 a_23141_8988.n7 a_23141_8988.n6 167.433
R18176 a_23141_8988.n3 a_23141_8988.t7 104.259
R18177 a_23141_8988.n7 a_23141_8988.t11 104.259
R18178 a_23141_8988.n4 a_23141_8988.n1 89.977
R18179 a_23141_8988.n5 a_23141_8988.n0 89.977
R18180 a_23141_8988.n9 a_23141_8988.n8 89.977
R18181 a_23141_8988.n8 a_23141_8988.n7 77.784
R18182 a_23141_8988.n5 a_23141_8988.n4 77.456
R18183 a_23141_8988.n8 a_23141_8988.n5 77.456
R18184 a_23141_8988.n4 a_23141_8988.n3 75.815
R18185 a_23141_8988.n2 a_23141_8988.t6 14.282
R18186 a_23141_8988.n2 a_23141_8988.t8 14.282
R18187 a_23141_8988.n1 a_23141_8988.t5 14.282
R18188 a_23141_8988.n1 a_23141_8988.t3 14.282
R18189 a_23141_8988.n0 a_23141_8988.t4 14.282
R18190 a_23141_8988.n0 a_23141_8988.t1 14.282
R18191 a_23141_8988.n6 a_23141_8988.t9 14.282
R18192 a_23141_8988.n6 a_23141_8988.t10 14.282
R18193 a_23141_8988.n9 a_23141_8988.t0 14.282
R18194 a_23141_8988.t2 a_23141_8988.n9 14.282
R18195 a_46140_17941.t8 a_46140_17941.n2 404.877
R18196 a_46140_17941.n1 a_46140_17941.t5 210.902
R18197 a_46140_17941.n3 a_46140_17941.t8 136.949
R18198 a_46140_17941.n2 a_46140_17941.n1 107.801
R18199 a_46140_17941.n1 a_46140_17941.t6 80.333
R18200 a_46140_17941.n2 a_46140_17941.t7 80.333
R18201 a_46140_17941.n0 a_46140_17941.t3 17.4
R18202 a_46140_17941.n0 a_46140_17941.t2 17.4
R18203 a_46140_17941.n4 a_46140_17941.t4 15.032
R18204 a_46140_17941.n5 a_46140_17941.t1 14.282
R18205 a_46140_17941.t0 a_46140_17941.n5 14.282
R18206 a_46140_17941.n5 a_46140_17941.n4 1.65
R18207 a_46140_17941.n3 a_46140_17941.n0 0.657
R18208 a_46140_17941.n4 a_46140_17941.n3 0.614
R18209 a_39689_6822.n0 a_39689_6822.t4 14.282
R18210 a_39689_6822.t3 a_39689_6822.n0 14.282
R18211 a_39689_6822.n0 a_39689_6822.n9 0.999
R18212 a_39689_6822.n9 a_39689_6822.n6 0.575
R18213 a_39689_6822.n6 a_39689_6822.n8 0.2
R18214 a_39689_6822.n8 a_39689_6822.t9 16.058
R18215 a_39689_6822.n8 a_39689_6822.n7 0.999
R18216 a_39689_6822.n7 a_39689_6822.t10 14.282
R18217 a_39689_6822.n7 a_39689_6822.t11 14.282
R18218 a_39689_6822.n9 a_39689_6822.t5 16.058
R18219 a_39689_6822.n6 a_39689_6822.n4 0.227
R18220 a_39689_6822.n4 a_39689_6822.n5 1.511
R18221 a_39689_6822.n5 a_39689_6822.t6 14.282
R18222 a_39689_6822.n5 a_39689_6822.t7 14.282
R18223 a_39689_6822.n4 a_39689_6822.n1 0.669
R18224 a_39689_6822.n1 a_39689_6822.n2 0.001
R18225 a_39689_6822.n1 a_39689_6822.n3 267.767
R18226 a_39689_6822.n3 a_39689_6822.t1 14.282
R18227 a_39689_6822.n3 a_39689_6822.t2 14.282
R18228 a_39689_6822.n2 a_39689_6822.t8 14.282
R18229 a_39689_6822.n2 a_39689_6822.t0 14.282
R18230 a_45281_16454.n1 a_45281_16454.t5 318.922
R18231 a_45281_16454.n0 a_45281_16454.t4 274.739
R18232 a_45281_16454.n0 a_45281_16454.t6 274.739
R18233 a_45281_16454.n1 a_45281_16454.t7 269.116
R18234 a_45281_16454.t5 a_45281_16454.n0 179.946
R18235 a_45281_16454.n2 a_45281_16454.n1 105.178
R18236 a_45281_16454.t2 a_45281_16454.n4 29.444
R18237 a_45281_16454.n3 a_45281_16454.t0 28.565
R18238 a_45281_16454.n3 a_45281_16454.t1 28.565
R18239 a_45281_16454.n2 a_45281_16454.t3 18.145
R18240 a_45281_16454.n4 a_45281_16454.n2 2.878
R18241 a_45281_16454.n4 a_45281_16454.n3 0.764
R18242 a_24594_4618.t0 a_24594_4618.t1 17.4
R18243 a_14357_13585.n2 a_14357_13585.t5 448.381
R18244 a_14357_13585.n1 a_14357_13585.t4 286.438
R18245 a_14357_13585.n1 a_14357_13585.t6 286.438
R18246 a_14357_13585.n0 a_14357_13585.t7 247.69
R18247 a_14357_13585.n4 a_14357_13585.n3 182.117
R18248 a_14357_13585.t5 a_14357_13585.n1 160.666
R18249 a_14357_13585.n3 a_14357_13585.t0 28.568
R18250 a_14357_13585.n4 a_14357_13585.t1 28.565
R18251 a_14357_13585.t2 a_14357_13585.n4 28.565
R18252 a_14357_13585.n0 a_14357_13585.t3 18.127
R18253 a_14357_13585.n2 a_14357_13585.n0 4.036
R18254 a_14357_13585.n3 a_14357_13585.n2 0.937
R18255 a_47179_16454.n1 a_47179_16454.t5 318.922
R18256 a_47179_16454.n0 a_47179_16454.t4 274.739
R18257 a_47179_16454.n0 a_47179_16454.t6 274.739
R18258 a_47179_16454.n1 a_47179_16454.t7 269.116
R18259 a_47179_16454.t5 a_47179_16454.n0 179.946
R18260 a_47179_16454.n2 a_47179_16454.n1 107.263
R18261 a_47179_16454.t2 a_47179_16454.n4 29.444
R18262 a_47179_16454.n3 a_47179_16454.t0 28.565
R18263 a_47179_16454.n3 a_47179_16454.t1 28.565
R18264 a_47179_16454.n2 a_47179_16454.t3 18.145
R18265 a_47179_16454.n4 a_47179_16454.n2 2.878
R18266 a_47179_16454.n4 a_47179_16454.n3 0.764
R18267 a_47719_15761.t0 a_47719_15761.n0 14.282
R18268 a_47719_15761.n0 a_47719_15761.t1 14.282
R18269 a_47719_15761.n0 a_47719_15761.n9 0.999
R18270 a_47719_15761.n6 a_47719_15761.n8 0.2
R18271 a_47719_15761.n9 a_47719_15761.n6 0.575
R18272 a_47719_15761.n9 a_47719_15761.t5 16.058
R18273 a_47719_15761.n8 a_47719_15761.n7 0.999
R18274 a_47719_15761.n7 a_47719_15761.t7 14.282
R18275 a_47719_15761.n7 a_47719_15761.t6 14.282
R18276 a_47719_15761.n8 a_47719_15761.t8 16.058
R18277 a_47719_15761.n6 a_47719_15761.n4 0.227
R18278 a_47719_15761.n4 a_47719_15761.n5 1.511
R18279 a_47719_15761.n5 a_47719_15761.t9 14.282
R18280 a_47719_15761.n5 a_47719_15761.t11 14.282
R18281 a_47719_15761.n4 a_47719_15761.n1 0.669
R18282 a_47719_15761.n1 a_47719_15761.n2 0.001
R18283 a_47719_15761.n1 a_47719_15761.n3 267.767
R18284 a_47719_15761.n3 a_47719_15761.t4 14.282
R18285 a_47719_15761.n3 a_47719_15761.t3 14.282
R18286 a_47719_15761.n2 a_47719_15761.t2 14.282
R18287 a_47719_15761.n2 a_47719_15761.t10 14.282
R18288 a_51346_110.t0 a_51346_110.t1 17.4
R18289 a_41579_1042.n2 a_41579_1042.n0 267.767
R18290 a_41579_1042.n6 a_41579_1042.t5 16.058
R18291 a_41579_1042.n4 a_41579_1042.t10 16.058
R18292 a_41579_1042.n5 a_41579_1042.t4 14.282
R18293 a_41579_1042.n5 a_41579_1042.t3 14.282
R18294 a_41579_1042.n3 a_41579_1042.t9 14.282
R18295 a_41579_1042.n3 a_41579_1042.t11 14.282
R18296 a_41579_1042.n1 a_41579_1042.t8 14.282
R18297 a_41579_1042.n1 a_41579_1042.t1 14.282
R18298 a_41579_1042.n0 a_41579_1042.t7 14.282
R18299 a_41579_1042.n0 a_41579_1042.t6 14.282
R18300 a_41579_1042.n9 a_41579_1042.t0 14.282
R18301 a_41579_1042.t2 a_41579_1042.n9 14.282
R18302 a_41579_1042.n9 a_41579_1042.n8 1.511
R18303 a_41579_1042.n6 a_41579_1042.n5 0.999
R18304 a_41579_1042.n4 a_41579_1042.n3 0.999
R18305 a_41579_1042.n8 a_41579_1042.n2 0.669
R18306 a_41579_1042.n7 a_41579_1042.n6 0.575
R18307 a_41579_1042.n8 a_41579_1042.n7 0.227
R18308 a_41579_1042.n7 a_41579_1042.n4 0.2
R18309 a_41579_1042.n2 a_41579_1042.n1 0.001
R18310 a_15426_6045.n1 a_15426_6045.t6 318.922
R18311 a_15426_6045.n0 a_15426_6045.t7 274.739
R18312 a_15426_6045.n0 a_15426_6045.t5 274.739
R18313 a_15426_6045.n1 a_15426_6045.t4 269.116
R18314 a_15426_6045.t6 a_15426_6045.n0 179.946
R18315 a_15426_6045.n2 a_15426_6045.n1 107.263
R18316 a_15426_6045.t2 a_15426_6045.n4 29.444
R18317 a_15426_6045.n3 a_15426_6045.t1 28.565
R18318 a_15426_6045.n3 a_15426_6045.t0 28.565
R18319 a_15426_6045.n2 a_15426_6045.t3 18.145
R18320 a_15426_6045.n4 a_15426_6045.n2 2.878
R18321 a_15426_6045.n4 a_15426_6045.n3 0.764
R18322 a_16084_4620.t0 a_16084_4620.t1 380.209
R18323 a_19927_14428.n2 a_19927_14428.t4 867.497
R18324 a_19927_14428.n2 a_19927_14428.t6 591.811
R18325 a_19927_14428.n1 a_19927_14428.t7 286.438
R18326 a_19927_14428.n1 a_19927_14428.t5 286.438
R18327 a_19927_14428.n4 a_19927_14428.n0 192.754
R18328 a_19927_14428.t4 a_19927_14428.n1 160.666
R18329 a_19927_14428.t0 a_19927_14428.n4 28.568
R18330 a_19927_14428.n0 a_19927_14428.t2 28.565
R18331 a_19927_14428.n0 a_19927_14428.t1 28.565
R18332 a_19927_14428.n3 a_19927_14428.n2 19.25
R18333 a_19927_14428.n3 a_19927_14428.t3 18.726
R18334 a_19927_14428.n4 a_19927_14428.n3 1.123
R18335 a_19987_14454.n0 a_19987_14454.t0 14.282
R18336 a_19987_14454.t3 a_19987_14454.n0 14.282
R18337 a_19987_14454.n0 a_19987_14454.n9 89.977
R18338 a_19987_14454.n6 a_19987_14454.n7 77.784
R18339 a_19987_14454.n9 a_19987_14454.n6 77.456
R18340 a_19987_14454.n9 a_19987_14454.n4 77.456
R18341 a_19987_14454.n4 a_19987_14454.n2 75.815
R18342 a_19987_14454.n7 a_19987_14454.n8 167.433
R18343 a_19987_14454.n8 a_19987_14454.t9 14.282
R18344 a_19987_14454.n8 a_19987_14454.t11 14.282
R18345 a_19987_14454.n7 a_19987_14454.t10 104.259
R18346 a_19987_14454.n6 a_19987_14454.n5 89.977
R18347 a_19987_14454.n5 a_19987_14454.t2 14.282
R18348 a_19987_14454.n5 a_19987_14454.t1 14.282
R18349 a_19987_14454.n4 a_19987_14454.n3 89.977
R18350 a_19987_14454.n3 a_19987_14454.t4 14.282
R18351 a_19987_14454.n3 a_19987_14454.t5 14.282
R18352 a_19987_14454.n2 a_19987_14454.t8 104.259
R18353 a_19987_14454.n2 a_19987_14454.n1 167.433
R18354 a_19987_14454.n1 a_19987_14454.t7 14.282
R18355 a_19987_14454.n1 a_19987_14454.t6 14.282
R18356 a_19454_13724.t1 a_19454_13724.n0 14.282
R18357 a_19454_13724.n0 a_19454_13724.t2 14.282
R18358 a_19454_13724.n0 a_19454_13724.n1 258.161
R18359 a_19454_13724.n1 a_19454_13724.t4 14.283
R18360 a_19454_13724.n1 a_19454_13724.n7 4.366
R18361 a_19454_13724.n7 a_19454_13724.n5 0.852
R18362 a_19454_13724.n5 a_19454_13724.n6 258.161
R18363 a_19454_13724.n6 a_19454_13724.t7 14.282
R18364 a_19454_13724.n6 a_19454_13724.t6 14.282
R18365 a_19454_13724.n5 a_19454_13724.t5 14.283
R18366 a_19454_13724.n7 a_19454_13724.n4 97.614
R18367 a_19454_13724.n4 a_19454_13724.t8 200.029
R18368 a_19454_13724.t8 a_19454_13724.n3 206.421
R18369 a_19454_13724.n3 a_19454_13724.t9 80.333
R18370 a_19454_13724.n3 a_19454_13724.t10 206.421
R18371 a_19454_13724.n4 a_19454_13724.t11 1527.4
R18372 a_19454_13724.t11 a_19454_13724.n2 657.379
R18373 a_19454_13724.n2 a_19454_13724.t3 8.7
R18374 a_19454_13724.n2 a_19454_13724.t0 8.7
R18375 B[2].t14 B[2].t11 799.268
R18376 B[2].n9 B[2].n8 650.893
R18377 B[2].n5 B[2].n4 618.566
R18378 B[2].n14 B[2].n10 592.056
R18379 B[2].t1 B[2].t6 415.315
R18380 B[2].t12 B[2].n2 313.873
R18381 B[2].t9 B[2].n12 313.069
R18382 B[2].n10 B[2].t10 294.986
R18383 B[2].n7 B[2].t3 285.543
R18384 B[2].n4 B[2].t7 273.077
R18385 B[2].n1 B[2].t15 272.288
R18386 B[2].n11 B[2].t0 271.484
R18387 B[2].n6 B[2].t1 217.526
R18388 B[2].n0 B[2].t21 214.335
R18389 B[2].t6 B[2].n0 214.335
R18390 B[2].n5 B[2].t19 204.679
R18391 B[2].n14 B[2].t4 204.672
R18392 B[2].n8 B[2].t14 194.406
R18393 B[2].n13 B[2].t9 190.955
R18394 B[2].n13 B[2].t20 190.955
R18395 B[2].n3 B[2].t8 190.152
R18396 B[2].n3 B[2].t12 190.152
R18397 B[2].n1 B[2].t22 160.666
R18398 B[2].n2 B[2].t2 160.666
R18399 B[2].n7 B[2].t5 160.666
R18400 B[2].n12 B[2].t13 160.666
R18401 B[2].n11 B[2].t16 160.666
R18402 B[2].n4 B[2].t17 137.369
R18403 B[2].n10 B[2].t18 110.859
R18404 B[2].n2 B[2].n1 96.129
R18405 B[2].n12 B[2].n11 96.129
R18406 B[2].n8 B[2].n7 91.137
R18407 B[2].n0 B[2].t23 80.333
R18408 B[2].t19 B[2].n3 80.333
R18409 B[2].t4 B[2].n13 80.333
R18410 B[2].n15 B[2].n14 61.78
R18411 B[2].n6 B[2].n5 50.417
R18412 B[2] B[2].n15 48.774
R18413 B[2].n15 B[2].n9 9.758
R18414 B[2].n9 B[2].n6 4.527
R18415 a_58312_3565.t4 a_58312_3565.t5 800.071
R18416 a_58312_3565.n2 a_58312_3565.n1 659.097
R18417 a_58312_3565.n0 a_58312_3565.t6 285.109
R18418 a_58312_3565.n1 a_58312_3565.t4 193.602
R18419 a_58312_3565.n4 a_58312_3565.n3 192.754
R18420 a_58312_3565.n0 a_58312_3565.t7 160.666
R18421 a_58312_3565.n1 a_58312_3565.n0 91.507
R18422 a_58312_3565.n3 a_58312_3565.t1 28.568
R18423 a_58312_3565.t2 a_58312_3565.n4 28.565
R18424 a_58312_3565.n4 a_58312_3565.t0 28.565
R18425 a_58312_3565.n2 a_58312_3565.t3 19.061
R18426 a_58312_3565.n3 a_58312_3565.n2 1.005
R18427 a_53713_16459.n1 a_53713_16459.t6 318.922
R18428 a_53713_16459.n0 a_53713_16459.t5 274.739
R18429 a_53713_16459.n0 a_53713_16459.t7 274.739
R18430 a_53713_16459.n1 a_53713_16459.t4 269.116
R18431 a_53713_16459.t6 a_53713_16459.n0 179.946
R18432 a_53713_16459.n2 a_53713_16459.n1 107.263
R18433 a_53713_16459.t2 a_53713_16459.n4 29.444
R18434 a_53713_16459.n3 a_53713_16459.t0 28.565
R18435 a_53713_16459.n3 a_53713_16459.t1 28.565
R18436 a_53713_16459.n2 a_53713_16459.t3 18.145
R18437 a_53713_16459.n4 a_53713_16459.n2 2.878
R18438 a_53713_16459.n4 a_53713_16459.n3 0.764
R18439 a_59910_20638.t6 a_59910_20638.t5 574.43
R18440 a_59910_20638.n1 a_59910_20638.t4 285.109
R18441 a_59910_20638.n3 a_59910_20638.n2 197.217
R18442 a_59910_20638.n4 a_59910_20638.n0 192.754
R18443 a_59910_20638.n1 a_59910_20638.t7 160.666
R18444 a_59910_20638.n2 a_59910_20638.t6 160.666
R18445 a_59910_20638.n2 a_59910_20638.n1 114.829
R18446 a_59910_20638.t0 a_59910_20638.n4 28.568
R18447 a_59910_20638.n0 a_59910_20638.t2 28.565
R18448 a_59910_20638.n0 a_59910_20638.t1 28.565
R18449 a_59910_20638.n3 a_59910_20638.t3 18.838
R18450 a_59910_20638.n4 a_59910_20638.n3 1.129
R18451 a_61636_24201.n0 a_61636_24201.t3 14.282
R18452 a_61636_24201.n0 a_61636_24201.t4 14.282
R18453 a_61636_24201.n1 a_61636_24201.t2 14.282
R18454 a_61636_24201.n1 a_61636_24201.t1 14.282
R18455 a_61636_24201.t0 a_61636_24201.n3 14.282
R18456 a_61636_24201.n3 a_61636_24201.t5 14.282
R18457 a_61636_24201.n2 a_61636_24201.n0 2.546
R18458 a_61636_24201.n2 a_61636_24201.n1 2.367
R18459 a_61636_24201.n3 a_61636_24201.n2 0.001
R18460 a_13602_20259.t0 a_13602_20259.t1 17.4
R18461 a_3652_8992.n1 a_3652_8992.t5 990.34
R18462 a_3652_8992.n1 a_3652_8992.t7 408.211
R18463 a_3652_8992.n0 a_3652_8992.t4 286.438
R18464 a_3652_8992.n0 a_3652_8992.t6 286.438
R18465 a_3652_8992.n4 a_3652_8992.n3 185.55
R18466 a_3652_8992.t5 a_3652_8992.n0 160.666
R18467 a_3652_8992.n3 a_3652_8992.t1 28.568
R18468 a_3652_8992.n4 a_3652_8992.t0 28.565
R18469 a_3652_8992.t2 a_3652_8992.n4 28.565
R18470 a_3652_8992.n2 a_3652_8992.t3 21.476
R18471 a_3652_8992.n2 a_3652_8992.n1 11.714
R18472 a_3652_8992.n3 a_3652_8992.n2 1.537
R18473 a_17501_10851.n2 a_17501_10851.t5 448.381
R18474 a_17501_10851.n1 a_17501_10851.t4 286.438
R18475 a_17501_10851.n1 a_17501_10851.t7 286.438
R18476 a_17501_10851.n0 a_17501_10851.t6 247.69
R18477 a_17501_10851.n4 a_17501_10851.n3 182.117
R18478 a_17501_10851.t5 a_17501_10851.n1 160.666
R18479 a_17501_10851.n3 a_17501_10851.t0 28.568
R18480 a_17501_10851.n4 a_17501_10851.t1 28.565
R18481 a_17501_10851.t2 a_17501_10851.n4 28.565
R18482 a_17501_10851.n0 a_17501_10851.t3 18.127
R18483 a_17501_10851.n2 a_17501_10851.n0 4.036
R18484 a_17501_10851.n3 a_17501_10851.n2 0.937
R18485 a_43803_21347.n1 a_43803_21347.t7 318.922
R18486 a_43803_21347.n0 a_43803_21347.t6 274.739
R18487 a_43803_21347.n0 a_43803_21347.t4 274.739
R18488 a_43803_21347.n1 a_43803_21347.t5 269.116
R18489 a_43803_21347.t7 a_43803_21347.n0 179.946
R18490 a_43803_21347.n2 a_43803_21347.n1 105.178
R18491 a_43803_21347.n3 a_43803_21347.t0 29.444
R18492 a_43803_21347.n4 a_43803_21347.t1 28.565
R18493 a_43803_21347.t2 a_43803_21347.n4 28.565
R18494 a_43803_21347.n2 a_43803_21347.t3 18.145
R18495 a_43803_21347.n3 a_43803_21347.n2 2.878
R18496 a_43803_21347.n4 a_43803_21347.n3 0.764
R18497 a_43391_21373.n0 a_43391_21373.n9 1.511
R18498 a_43391_21373.t3 a_43391_21373.n0 14.282
R18499 a_43391_21373.n0 a_43391_21373.t4 14.282
R18500 a_43391_21373.n9 a_43391_21373.n5 0.227
R18501 a_43391_21373.n9 a_43391_21373.n6 0.669
R18502 a_43391_21373.n6 a_43391_21373.n7 0.001
R18503 a_43391_21373.n6 a_43391_21373.n8 267.767
R18504 a_43391_21373.n8 a_43391_21373.t6 14.282
R18505 a_43391_21373.n8 a_43391_21373.t7 14.282
R18506 a_43391_21373.n7 a_43391_21373.t5 14.282
R18507 a_43391_21373.n7 a_43391_21373.t8 14.282
R18508 a_43391_21373.n5 a_43391_21373.n2 0.575
R18509 a_43391_21373.n5 a_43391_21373.n4 0.2
R18510 a_43391_21373.n4 a_43391_21373.t11 16.058
R18511 a_43391_21373.n4 a_43391_21373.n3 0.999
R18512 a_43391_21373.n3 a_43391_21373.t10 14.282
R18513 a_43391_21373.n3 a_43391_21373.t9 14.282
R18514 a_43391_21373.n2 a_43391_21373.n1 0.999
R18515 a_43391_21373.n1 a_43391_21373.t1 14.282
R18516 a_43391_21373.n1 a_43391_21373.t0 14.282
R18517 a_43391_21373.n2 a_43391_21373.t2 16.058
R18518 a_50022_20638.t0 a_50022_20638.t1 380.209
R18519 a_50022_21370.n0 a_50022_21370.t7 14.282
R18520 a_50022_21370.t0 a_50022_21370.n0 14.282
R18521 a_50022_21370.n0 a_50022_21370.n8 90.416
R18522 a_50022_21370.n8 a_50022_21370.n7 50.575
R18523 a_50022_21370.n8 a_50022_21370.n4 74.302
R18524 a_50022_21370.n7 a_50022_21370.n6 157.665
R18525 a_50022_21370.n6 a_50022_21370.t4 8.7
R18526 a_50022_21370.n6 a_50022_21370.t3 8.7
R18527 a_50022_21370.n7 a_50022_21370.n5 122.999
R18528 a_50022_21370.n5 a_50022_21370.t6 14.282
R18529 a_50022_21370.n5 a_50022_21370.t5 14.282
R18530 a_50022_21370.n4 a_50022_21370.n3 90.436
R18531 a_50022_21370.n3 a_50022_21370.t1 14.282
R18532 a_50022_21370.n3 a_50022_21370.t2 14.282
R18533 a_50022_21370.n4 a_50022_21370.n1 2011.09
R18534 a_50022_21370.t10 a_50022_21370.n2 160.666
R18535 a_50022_21370.n1 a_50022_21370.t10 867.393
R18536 a_50022_21370.n2 a_50022_21370.t9 287.241
R18537 a_50022_21370.n2 a_50022_21370.t8 287.241
R18538 a_50022_21370.n1 a_50022_21370.t11 545.094
R18539 a_71842_14595.t0 a_71842_14595.t1 17.4
R18540 a_30154_12886.n1 a_30154_12886.t4 318.119
R18541 a_30154_12886.n1 a_30154_12886.t5 269.919
R18542 a_30154_12886.n0 a_30154_12886.t6 267.256
R18543 a_30154_12886.n0 a_30154_12886.t7 267.256
R18544 a_30154_12886.n4 a_30154_12886.n3 193.227
R18545 a_30154_12886.t4 a_30154_12886.n0 160.666
R18546 a_30154_12886.n2 a_30154_12886.n1 106.999
R18547 a_30154_12886.n3 a_30154_12886.t1 28.568
R18548 a_30154_12886.t2 a_30154_12886.n4 28.565
R18549 a_30154_12886.n4 a_30154_12886.t0 28.565
R18550 a_30154_12886.n2 a_30154_12886.t3 18.149
R18551 a_30154_12886.n3 a_30154_12886.n2 3.726
R18552 a_5108_13805.n2 a_5108_13805.t6 990.34
R18553 a_5108_13805.n3 a_5108_13805.n2 566.592
R18554 a_5108_13805.n2 a_5108_13805.t7 408.211
R18555 a_5108_13805.n1 a_5108_13805.t5 286.438
R18556 a_5108_13805.n1 a_5108_13805.t4 286.438
R18557 a_5108_13805.t6 a_5108_13805.n1 160.666
R18558 a_5108_13805.n3 a_5108_13805.n0 100.603
R18559 a_5108_13805.n4 a_5108_13805.n3 100.24
R18560 a_5108_13805.n0 a_5108_13805.t0 28.568
R18561 a_5108_13805.n4 a_5108_13805.t1 28.565
R18562 a_5108_13805.t2 a_5108_13805.n4 28.565
R18563 a_5108_13805.n0 a_5108_13805.t3 17.64
R18564 a_4233_14458.n0 a_4233_14458.t6 14.282
R18565 a_4233_14458.t0 a_4233_14458.n0 14.282
R18566 a_4233_14458.n0 a_4233_14458.n9 89.977
R18567 a_4233_14458.n6 a_4233_14458.n7 77.784
R18568 a_4233_14458.n9 a_4233_14458.n6 77.456
R18569 a_4233_14458.n9 a_4233_14458.n4 77.456
R18570 a_4233_14458.n4 a_4233_14458.n2 75.815
R18571 a_4233_14458.n7 a_4233_14458.n8 167.433
R18572 a_4233_14458.n8 a_4233_14458.t4 14.282
R18573 a_4233_14458.n8 a_4233_14458.t5 14.282
R18574 a_4233_14458.n7 a_4233_14458.t3 104.259
R18575 a_4233_14458.n6 a_4233_14458.n5 89.977
R18576 a_4233_14458.n5 a_4233_14458.t8 14.282
R18577 a_4233_14458.n5 a_4233_14458.t7 14.282
R18578 a_4233_14458.n4 a_4233_14458.n3 89.977
R18579 a_4233_14458.n3 a_4233_14458.t1 14.282
R18580 a_4233_14458.n3 a_4233_14458.t2 14.282
R18581 a_4233_14458.n2 a_4233_14458.t10 104.259
R18582 a_4233_14458.n2 a_4233_14458.n1 167.433
R18583 a_4233_14458.n1 a_4233_14458.t9 14.282
R18584 a_4233_14458.n1 a_4233_14458.t11 14.282
R18585 a_65224_3811.n1 a_65224_3811.t4 318.922
R18586 a_65224_3811.n0 a_65224_3811.t5 273.935
R18587 a_65224_3811.n0 a_65224_3811.t6 273.935
R18588 a_65224_3811.n1 a_65224_3811.t7 269.116
R18589 a_65224_3811.n4 a_65224_3811.n3 193.227
R18590 a_65224_3811.t4 a_65224_3811.n0 179.142
R18591 a_65224_3811.n2 a_65224_3811.n1 106.999
R18592 a_65224_3811.n3 a_65224_3811.t1 28.568
R18593 a_65224_3811.t0 a_65224_3811.n4 28.565
R18594 a_65224_3811.n4 a_65224_3811.t3 28.565
R18595 a_65224_3811.n2 a_65224_3811.t2 18.149
R18596 a_65224_3811.n3 a_65224_3811.n2 3.726
R18597 a_65769_3118.t0 a_65769_3118.n0 14.282
R18598 a_65769_3118.n0 a_65769_3118.t2 14.282
R18599 a_65769_3118.n0 a_65769_3118.n8 90.436
R18600 a_65769_3118.n4 a_65769_3118.n7 50.575
R18601 a_65769_3118.n8 a_65769_3118.n4 74.302
R18602 a_65769_3118.n7 a_65769_3118.n6 157.665
R18603 a_65769_3118.n6 a_65769_3118.t6 8.7
R18604 a_65769_3118.n6 a_65769_3118.t7 8.7
R18605 a_65769_3118.n7 a_65769_3118.n5 122.999
R18606 a_65769_3118.n5 a_65769_3118.t4 14.282
R18607 a_65769_3118.n5 a_65769_3118.t5 14.282
R18608 a_65769_3118.n4 a_65769_3118.n3 90.416
R18609 a_65769_3118.n3 a_65769_3118.t3 14.282
R18610 a_65769_3118.n3 a_65769_3118.t1 14.282
R18611 a_65769_3118.n8 a_65769_3118.n1 1255.94
R18612 a_65769_3118.n1 a_65769_3118.t9 408.806
R18613 a_65769_3118.t8 a_65769_3118.n2 160.666
R18614 a_65769_3118.n1 a_65769_3118.t8 989.744
R18615 a_65769_3118.n2 a_65769_3118.t11 287.241
R18616 a_65769_3118.n2 a_65769_3118.t10 287.241
R18617 a_24240_5350.n5 a_24240_5350.n7 0.2
R18618 a_24240_5350.n9 a_24240_5350.n5 0.575
R18619 a_24240_5350.t0 a_24240_5350.n9 16.058
R18620 a_24240_5350.n9 a_24240_5350.n8 0.999
R18621 a_24240_5350.n8 a_24240_5350.t5 14.282
R18622 a_24240_5350.n8 a_24240_5350.t4 14.282
R18623 a_24240_5350.n7 a_24240_5350.n6 0.999
R18624 a_24240_5350.n6 a_24240_5350.t11 14.282
R18625 a_24240_5350.n6 a_24240_5350.t9 14.282
R18626 a_24240_5350.n7 a_24240_5350.t10 16.058
R18627 a_24240_5350.n5 a_24240_5350.n3 0.227
R18628 a_24240_5350.n3 a_24240_5350.n4 1.511
R18629 a_24240_5350.n4 a_24240_5350.t7 14.282
R18630 a_24240_5350.n4 a_24240_5350.t8 14.282
R18631 a_24240_5350.n3 a_24240_5350.n0 0.669
R18632 a_24240_5350.n0 a_24240_5350.n1 0.001
R18633 a_24240_5350.n0 a_24240_5350.n2 267.767
R18634 a_24240_5350.n2 a_24240_5350.t3 14.282
R18635 a_24240_5350.n2 a_24240_5350.t1 14.282
R18636 a_24240_5350.n1 a_24240_5350.t2 14.282
R18637 a_24240_5350.n1 a_24240_5350.t6 14.282
R18638 a_25100_20862.t1 a_25100_20862.n0 14.282
R18639 a_25100_20862.n0 a_25100_20862.t2 14.282
R18640 a_25100_20862.n0 a_25100_20862.n1 258.161
R18641 a_25100_20862.n1 a_25100_20862.t3 14.283
R18642 a_25100_20862.n1 a_25100_20862.n7 4.366
R18643 a_25100_20862.n7 a_25100_20862.n5 0.852
R18644 a_25100_20862.n5 a_25100_20862.n6 258.161
R18645 a_25100_20862.n6 a_25100_20862.t5 14.282
R18646 a_25100_20862.n6 a_25100_20862.t7 14.282
R18647 a_25100_20862.n5 a_25100_20862.t6 14.283
R18648 a_25100_20862.n7 a_25100_20862.n4 97.614
R18649 a_25100_20862.n4 a_25100_20862.t8 200.029
R18650 a_25100_20862.t8 a_25100_20862.n3 206.421
R18651 a_25100_20862.n3 a_25100_20862.t9 80.333
R18652 a_25100_20862.n3 a_25100_20862.t10 206.421
R18653 a_25100_20862.n4 a_25100_20862.t11 1527.4
R18654 a_25100_20862.t11 a_25100_20862.n2 657.379
R18655 a_25100_20862.n2 a_25100_20862.t4 8.7
R18656 a_25100_20862.n2 a_25100_20862.t0 8.7
R18657 a_25633_21592.n0 a_25633_21592.t0 14.282
R18658 a_25633_21592.t6 a_25633_21592.n0 14.282
R18659 a_25633_21592.n0 a_25633_21592.n9 89.977
R18660 a_25633_21592.n6 a_25633_21592.n7 77.784
R18661 a_25633_21592.n9 a_25633_21592.n6 77.456
R18662 a_25633_21592.n9 a_25633_21592.n4 77.456
R18663 a_25633_21592.n4 a_25633_21592.n2 75.815
R18664 a_25633_21592.n7 a_25633_21592.n8 167.433
R18665 a_25633_21592.n8 a_25633_21592.t10 14.282
R18666 a_25633_21592.n8 a_25633_21592.t9 14.282
R18667 a_25633_21592.n7 a_25633_21592.t11 104.259
R18668 a_25633_21592.n6 a_25633_21592.n5 89.977
R18669 a_25633_21592.n5 a_25633_21592.t2 14.282
R18670 a_25633_21592.n5 a_25633_21592.t1 14.282
R18671 a_25633_21592.n4 a_25633_21592.n3 89.977
R18672 a_25633_21592.n3 a_25633_21592.t7 14.282
R18673 a_25633_21592.n3 a_25633_21592.t8 14.282
R18674 a_25633_21592.n2 a_25633_21592.t5 104.259
R18675 a_25633_21592.n2 a_25633_21592.n1 167.433
R18676 a_25633_21592.n1 a_25633_21592.t4 14.282
R18677 a_25633_21592.n1 a_25633_21592.t3 14.282
R18678 a_16014_1740.n2 a_16014_1740.t4 448.382
R18679 a_16014_1740.n1 a_16014_1740.t6 286.438
R18680 a_16014_1740.n1 a_16014_1740.t7 286.438
R18681 a_16014_1740.n0 a_16014_1740.t5 247.69
R18682 a_16014_1740.n4 a_16014_1740.n3 182.117
R18683 a_16014_1740.t4 a_16014_1740.n1 160.666
R18684 a_16014_1740.n3 a_16014_1740.t0 28.568
R18685 a_16014_1740.n4 a_16014_1740.t1 28.565
R18686 a_16014_1740.t2 a_16014_1740.n4 28.565
R18687 a_16014_1740.n0 a_16014_1740.t3 18.127
R18688 a_16014_1740.n2 a_16014_1740.n0 4.039
R18689 a_16014_1740.n3 a_16014_1740.n2 0.937
R18690 a_30152_6681.n1 a_30152_6681.t5 318.119
R18691 a_30152_6681.n1 a_30152_6681.t7 269.919
R18692 a_30152_6681.n0 a_30152_6681.t6 267.256
R18693 a_30152_6681.n0 a_30152_6681.t4 267.256
R18694 a_30152_6681.n4 a_30152_6681.n3 193.227
R18695 a_30152_6681.t5 a_30152_6681.n0 160.666
R18696 a_30152_6681.n2 a_30152_6681.n1 106.999
R18697 a_30152_6681.n3 a_30152_6681.t0 28.568
R18698 a_30152_6681.n4 a_30152_6681.t1 28.565
R18699 a_30152_6681.t2 a_30152_6681.n4 28.565
R18700 a_30152_6681.n2 a_30152_6681.t3 18.149
R18701 a_30152_6681.n3 a_30152_6681.n2 3.726
R18702 a_29952_5843.t0 a_29952_5843.n9 16.058
R18703 a_29952_5843.n9 a_29952_5843.n5 0.2
R18704 a_29952_5843.n5 a_29952_5843.n7 0.575
R18705 a_29952_5843.n9 a_29952_5843.n8 0.999
R18706 a_29952_5843.n8 a_29952_5843.t9 14.282
R18707 a_29952_5843.n8 a_29952_5843.t10 14.282
R18708 a_29952_5843.n7 a_29952_5843.n6 0.999
R18709 a_29952_5843.n6 a_29952_5843.t6 14.282
R18710 a_29952_5843.n6 a_29952_5843.t5 14.282
R18711 a_29952_5843.n7 a_29952_5843.t4 16.058
R18712 a_29952_5843.n5 a_29952_5843.n3 0.227
R18713 a_29952_5843.n3 a_29952_5843.n4 1.511
R18714 a_29952_5843.n4 a_29952_5843.t3 14.282
R18715 a_29952_5843.n4 a_29952_5843.t2 14.282
R18716 a_29952_5843.n3 a_29952_5843.n0 0.669
R18717 a_29952_5843.n0 a_29952_5843.n1 0.001
R18718 a_29952_5843.n0 a_29952_5843.n2 267.767
R18719 a_29952_5843.n2 a_29952_5843.t11 14.282
R18720 a_29952_5843.n2 a_29952_5843.t7 14.282
R18721 a_29952_5843.n1 a_29952_5843.t8 14.282
R18722 a_29952_5843.n1 a_29952_5843.t1 14.282
R18723 a_41251_9658.t7 a_41251_9658.n3 404.877
R18724 a_41251_9658.n2 a_41251_9658.t8 210.902
R18725 a_41251_9658.n4 a_41251_9658.t7 136.943
R18726 a_41251_9658.n3 a_41251_9658.n2 107.801
R18727 a_41251_9658.n2 a_41251_9658.t5 80.333
R18728 a_41251_9658.n3 a_41251_9658.t6 80.333
R18729 a_41251_9658.n1 a_41251_9658.t0 17.4
R18730 a_41251_9658.n1 a_41251_9658.t2 17.4
R18731 a_41251_9658.t1 a_41251_9658.n5 15.032
R18732 a_41251_9658.n0 a_41251_9658.t3 14.282
R18733 a_41251_9658.n0 a_41251_9658.t4 14.282
R18734 a_41251_9658.n5 a_41251_9658.n0 1.65
R18735 a_41251_9658.n4 a_41251_9658.n1 0.672
R18736 a_41251_9658.n5 a_41251_9658.n4 0.665
R18737 B[3].t28 B[3].t19 800.875
R18738 B[3].n9 B[3].n8 650.874
R18739 B[3].n4 B[3].n3 618.566
R18740 B[3].n21 B[3].n17 592.056
R18741 B[3].t11 B[3].t39 437.233
R18742 B[3].t5 B[3].t20 437.233
R18743 B[3].t34 B[3].t35 437.233
R18744 B[3].t31 B[3].t38 415.315
R18745 B[3].t21 B[3].t12 415.315
R18746 B[3].t8 B[3].n1 313.873
R18747 B[3].t1 B[3].n19 313.069
R18748 B[3].n17 B[3].t3 294.986
R18749 B[3].n7 B[3].t23 284.688
R18750 B[3].n3 B[3].t10 273.077
R18751 B[3].n0 B[3].t16 272.288
R18752 B[3].n18 B[3].t18 271.484
R18753 B[3].n12 B[3].t21 225.375
R18754 B[3].n15 B[3].t34 223.992
R18755 B[3].n15 B[3].t5 217.885
R18756 B[3].n6 B[3].t31 217.532
R18757 B[3].n12 B[3].t11 216.848
R18758 B[3].n11 B[3].t14 214.686
R18759 B[3].t39 B[3].n11 214.686
R18760 B[3].n13 B[3].t2 214.686
R18761 B[3].t20 B[3].n13 214.686
R18762 B[3].n14 B[3].t7 214.686
R18763 B[3].t35 B[3].n14 214.686
R18764 B[3].n5 B[3].t36 214.335
R18765 B[3].t38 B[3].n5 214.335
R18766 B[3].n10 B[3].t25 214.335
R18767 B[3].t12 B[3].n10 214.335
R18768 B[3].n4 B[3].t32 204.679
R18769 B[3].n21 B[3].t29 204.672
R18770 B[3].n8 B[3].t28 192.799
R18771 B[3].n20 B[3].t1 190.955
R18772 B[3].n20 B[3].t22 190.955
R18773 B[3].n2 B[3].t4 190.152
R18774 B[3].n2 B[3].t8 190.152
R18775 B[3].n0 B[3].t30 160.666
R18776 B[3].n1 B[3].t0 160.666
R18777 B[3].n7 B[3].t26 160.666
R18778 B[3].n19 B[3].t6 160.666
R18779 B[3].n18 B[3].t13 160.666
R18780 B[3].n3 B[3].t27 137.369
R18781 B[3].n17 B[3].t17 110.859
R18782 B[3].n1 B[3].n0 96.129
R18783 B[3].n19 B[3].n18 96.129
R18784 B[3].n8 B[3].n7 91.889
R18785 B[3].n5 B[3].t37 80.333
R18786 B[3].t32 B[3].n2 80.333
R18787 B[3].n11 B[3].t15 80.333
R18788 B[3].n10 B[3].t24 80.333
R18789 B[3].n13 B[3].t33 80.333
R18790 B[3].n14 B[3].t9 80.333
R18791 B[3].t29 B[3].n20 80.333
R18792 B[3].n16 B[3].n12 62.924
R18793 B[3].n6 B[3].n4 50.557
R18794 B[3] B[3].n23 48.773
R18795 B[3].n22 B[3].n21 45.981
R18796 B[3].n23 B[3].n22 28.632
R18797 B[3].n23 B[3].n9 14.285
R18798 B[3].n22 B[3].n16 13.481
R18799 B[3].n9 B[3].n6 4.969
R18800 B[3].n16 B[3].n15 0.469
R18801 a_62366_15449.n0 a_62366_15449.t7 214.335
R18802 a_62366_15449.t10 a_62366_15449.n0 214.335
R18803 a_62366_15449.n1 a_62366_15449.t10 143.851
R18804 a_62366_15449.n1 a_62366_15449.t9 135.658
R18805 a_62366_15449.n0 a_62366_15449.t8 80.333
R18806 a_62366_15449.n4 a_62366_15449.t1 28.565
R18807 a_62366_15449.n4 a_62366_15449.t2 28.565
R18808 a_62366_15449.n2 a_62366_15449.t6 28.565
R18809 a_62366_15449.n2 a_62366_15449.t4 28.565
R18810 a_62366_15449.t3 a_62366_15449.n7 28.565
R18811 a_62366_15449.n7 a_62366_15449.t5 28.565
R18812 a_62366_15449.n5 a_62366_15449.t0 9.714
R18813 a_62366_15449.n5 a_62366_15449.n4 1.003
R18814 a_62366_15449.n6 a_62366_15449.n3 0.833
R18815 a_62366_15449.n3 a_62366_15449.n2 0.653
R18816 a_62366_15449.n7 a_62366_15449.n6 0.653
R18817 a_62366_15449.n6 a_62366_15449.n5 0.341
R18818 a_62366_15449.n3 a_62366_15449.n1 0.032
R18819 a_14310_5328.n1 a_14310_5328.t7 318.922
R18820 a_14310_5328.n0 a_14310_5328.t5 273.935
R18821 a_14310_5328.n0 a_14310_5328.t6 273.935
R18822 a_14310_5328.n1 a_14310_5328.t4 269.116
R18823 a_14310_5328.n4 a_14310_5328.n3 193.227
R18824 a_14310_5328.t7 a_14310_5328.n0 179.142
R18825 a_14310_5328.n2 a_14310_5328.n1 106.999
R18826 a_14310_5328.n3 a_14310_5328.t1 28.568
R18827 a_14310_5328.n4 a_14310_5328.t0 28.565
R18828 a_14310_5328.t2 a_14310_5328.n4 28.565
R18829 a_14310_5328.n2 a_14310_5328.t3 18.149
R18830 a_14310_5328.n3 a_14310_5328.n2 3.726
R18831 a_41611_21373.t1 a_41611_21373.n0 14.282
R18832 a_41611_21373.n0 a_41611_21373.t6 14.282
R18833 a_41611_21373.n0 a_41611_21373.n12 90.416
R18834 a_41611_21373.n12 a_41611_21373.n11 50.575
R18835 a_41611_21373.n12 a_41611_21373.n8 74.302
R18836 a_41611_21373.n11 a_41611_21373.n10 157.665
R18837 a_41611_21373.n10 a_41611_21373.t0 8.7
R18838 a_41611_21373.n10 a_41611_21373.t7 8.7
R18839 a_41611_21373.n11 a_41611_21373.n9 122.999
R18840 a_41611_21373.n9 a_41611_21373.t3 14.282
R18841 a_41611_21373.n9 a_41611_21373.t2 14.282
R18842 a_41611_21373.n8 a_41611_21373.n7 90.436
R18843 a_41611_21373.n7 a_41611_21373.t4 14.282
R18844 a_41611_21373.n7 a_41611_21373.t5 14.282
R18845 a_41611_21373.n8 a_41611_21373.n1 342.688
R18846 a_41611_21373.n1 a_41611_21373.n6 126.566
R18847 a_41611_21373.n6 a_41611_21373.t8 294.653
R18848 a_41611_21373.n6 a_41611_21373.t9 111.663
R18849 a_41611_21373.n1 a_41611_21373.n5 552.333
R18850 a_41611_21373.n5 a_41611_21373.n4 6.615
R18851 a_41611_21373.n4 a_41611_21373.t14 93.989
R18852 a_41611_21373.n5 a_41611_21373.n3 97.816
R18853 a_41611_21373.n3 a_41611_21373.t15 80.333
R18854 a_41611_21373.n3 a_41611_21373.t10 394.151
R18855 a_41611_21373.t10 a_41611_21373.n2 269.523
R18856 a_41611_21373.n2 a_41611_21373.t11 160.666
R18857 a_41611_21373.n2 a_41611_21373.t12 269.523
R18858 a_41611_21373.n4 a_41611_21373.t13 198.043
R18859 a_43745_20641.t0 a_43745_20641.t1 17.4
R18860 a_54572_9678.n0 a_54572_9678.t0 14.282
R18861 a_54572_9678.n0 a_54572_9678.t4 14.282
R18862 a_54572_9678.n1 a_54572_9678.t2 14.282
R18863 a_54572_9678.n1 a_54572_9678.t1 14.282
R18864 a_54572_9678.t3 a_54572_9678.n3 14.282
R18865 a_54572_9678.n3 a_54572_9678.t5 14.282
R18866 a_54572_9678.n3 a_54572_9678.n2 2.546
R18867 a_54572_9678.n2 a_54572_9678.n1 2.367
R18868 a_54572_9678.n2 a_54572_9678.n0 0.001
R18869 a_63408_21343.n1 a_63408_21343.t6 318.922
R18870 a_63408_21343.n0 a_63408_21343.t5 274.739
R18871 a_63408_21343.n0 a_63408_21343.t7 274.739
R18872 a_63408_21343.n1 a_63408_21343.t4 269.116
R18873 a_63408_21343.t6 a_63408_21343.n0 179.946
R18874 a_63408_21343.n2 a_63408_21343.n1 105.178
R18875 a_63408_21343.n3 a_63408_21343.t1 29.444
R18876 a_63408_21343.t2 a_63408_21343.n4 28.565
R18877 a_63408_21343.n4 a_63408_21343.t0 28.565
R18878 a_63408_21343.n2 a_63408_21343.t3 18.145
R18879 a_63408_21343.n3 a_63408_21343.n2 2.878
R18880 a_63408_21343.n4 a_63408_21343.n3 0.764
R18881 a_63114_20637.t0 a_63114_20637.t1 380.209
R18882 a_22290_1744.n2 a_22290_1744.t7 448.382
R18883 a_22290_1744.n1 a_22290_1744.t4 286.438
R18884 a_22290_1744.n1 a_22290_1744.t5 286.438
R18885 a_22290_1744.n0 a_22290_1744.t6 247.69
R18886 a_22290_1744.n4 a_22290_1744.n3 182.117
R18887 a_22290_1744.t7 a_22290_1744.n1 160.666
R18888 a_22290_1744.n3 a_22290_1744.t0 28.568
R18889 a_22290_1744.t2 a_22290_1744.n4 28.565
R18890 a_22290_1744.n4 a_22290_1744.t1 28.565
R18891 a_22290_1744.n0 a_22290_1744.t3 18.127
R18892 a_22290_1744.n2 a_22290_1744.n0 4.039
R18893 a_22290_1744.n3 a_22290_1744.n2 0.937
R18894 a_10459_8962.t1 a_10459_8962.n0 14.282
R18895 a_10459_8962.n0 a_10459_8962.t6 14.282
R18896 a_10459_8962.n0 a_10459_8962.n8 122.747
R18897 a_10459_8962.n4 a_10459_8962.n6 74.302
R18898 a_10459_8962.n8 a_10459_8962.n4 50.575
R18899 a_10459_8962.n8 a_10459_8962.n7 157.665
R18900 a_10459_8962.n7 a_10459_8962.t0 8.7
R18901 a_10459_8962.n7 a_10459_8962.t7 8.7
R18902 a_10459_8962.n6 a_10459_8962.n5 90.436
R18903 a_10459_8962.n5 a_10459_8962.t3 14.282
R18904 a_10459_8962.n5 a_10459_8962.t4 14.282
R18905 a_10459_8962.n4 a_10459_8962.n3 90.416
R18906 a_10459_8962.n3 a_10459_8962.t5 14.282
R18907 a_10459_8962.n3 a_10459_8962.t2 14.282
R18908 a_10459_8962.n6 a_10459_8962.n1 1401.44
R18909 a_10459_8962.n1 a_10459_8962.t10 591.811
R18910 a_10459_8962.n1 a_10459_8962.t8 867.497
R18911 a_10459_8962.t8 a_10459_8962.n2 160.666
R18912 a_10459_8962.n2 a_10459_8962.t11 286.438
R18913 a_10459_8962.n2 a_10459_8962.t9 286.438
R18914 a_6784_8988.n2 a_6784_8988.t6 990.34
R18915 a_6784_8988.n2 a_6784_8988.t4 408.211
R18916 a_6784_8988.n1 a_6784_8988.t5 286.438
R18917 a_6784_8988.n1 a_6784_8988.t7 286.438
R18918 a_6784_8988.n4 a_6784_8988.n0 185.55
R18919 a_6784_8988.t6 a_6784_8988.n1 160.666
R18920 a_6784_8988.t2 a_6784_8988.n4 28.568
R18921 a_6784_8988.n0 a_6784_8988.t1 28.565
R18922 a_6784_8988.n0 a_6784_8988.t0 28.565
R18923 a_6784_8988.n3 a_6784_8988.t3 21.476
R18924 a_6784_8988.n3 a_6784_8988.n2 12.479
R18925 a_6784_8988.n4 a_6784_8988.n3 1.537
R18926 a_61819_1016.n1 a_61819_1016.t4 318.922
R18927 a_61819_1016.n0 a_61819_1016.t7 274.739
R18928 a_61819_1016.n0 a_61819_1016.t5 274.739
R18929 a_61819_1016.n1 a_61819_1016.t6 269.116
R18930 a_61819_1016.t4 a_61819_1016.n0 179.946
R18931 a_61819_1016.n2 a_61819_1016.n1 105.178
R18932 a_61819_1016.t2 a_61819_1016.n4 29.444
R18933 a_61819_1016.n3 a_61819_1016.t1 28.565
R18934 a_61819_1016.n3 a_61819_1016.t0 28.565
R18935 a_61819_1016.n2 a_61819_1016.t3 18.145
R18936 a_61819_1016.n4 a_61819_1016.n2 2.878
R18937 a_61819_1016.n4 a_61819_1016.n3 0.764
R18938 a_30152_5242.n1 a_30152_5242.t5 318.119
R18939 a_30152_5242.n1 a_30152_5242.t6 269.919
R18940 a_30152_5242.n0 a_30152_5242.t7 267.853
R18941 a_30152_5242.n0 a_30152_5242.t4 267.853
R18942 a_30152_5242.t5 a_30152_5242.n0 160.666
R18943 a_30152_5242.n2 a_30152_5242.n1 107.263
R18944 a_30152_5242.n3 a_30152_5242.t1 29.444
R18945 a_30152_5242.t2 a_30152_5242.n4 28.565
R18946 a_30152_5242.n4 a_30152_5242.t0 28.565
R18947 a_30152_5242.n2 a_30152_5242.t3 18.145
R18948 a_30152_5242.n3 a_30152_5242.n2 2.878
R18949 a_30152_5242.n4 a_30152_5242.n3 0.764
R18950 a_29954_12048.n8 a_29954_12048.n7 267.767
R18951 a_29954_12048.n1 a_29954_12048.t7 16.058
R18952 a_29954_12048.n3 a_29954_12048.t11 16.058
R18953 a_29954_12048.n0 a_29954_12048.t8 14.282
R18954 a_29954_12048.n0 a_29954_12048.t6 14.282
R18955 a_29954_12048.n2 a_29954_12048.t9 14.282
R18956 a_29954_12048.n2 a_29954_12048.t10 14.282
R18957 a_29954_12048.n5 a_29954_12048.t0 14.282
R18958 a_29954_12048.n5 a_29954_12048.t1 14.282
R18959 a_29954_12048.n7 a_29954_12048.t4 14.282
R18960 a_29954_12048.n7 a_29954_12048.t5 14.282
R18961 a_29954_12048.t2 a_29954_12048.n9 14.282
R18962 a_29954_12048.n9 a_29954_12048.t3 14.282
R18963 a_29954_12048.n6 a_29954_12048.n5 1.511
R18964 a_29954_12048.n1 a_29954_12048.n0 0.999
R18965 a_29954_12048.n3 a_29954_12048.n2 0.999
R18966 a_29954_12048.n8 a_29954_12048.n6 0.669
R18967 a_29954_12048.n4 a_29954_12048.n1 0.575
R18968 a_29954_12048.n6 a_29954_12048.n4 0.227
R18969 a_29954_12048.n4 a_29954_12048.n3 0.2
R18970 a_29954_12048.n9 a_29954_12048.n8 0.001
R18971 a_30150_2544.n2 a_30150_2544.t7 318.119
R18972 a_30150_2544.n2 a_30150_2544.t5 269.919
R18973 a_30150_2544.n1 a_30150_2544.t4 267.256
R18974 a_30150_2544.n1 a_30150_2544.t6 267.256
R18975 a_30150_2544.n4 a_30150_2544.n0 193.227
R18976 a_30150_2544.t7 a_30150_2544.n1 160.666
R18977 a_30150_2544.n3 a_30150_2544.n2 106.999
R18978 a_30150_2544.t2 a_30150_2544.n4 28.568
R18979 a_30150_2544.n0 a_30150_2544.t0 28.565
R18980 a_30150_2544.n0 a_30150_2544.t1 28.565
R18981 a_30150_2544.n3 a_30150_2544.t3 18.149
R18982 a_30150_2544.n4 a_30150_2544.n3 3.726
R18983 a_30643_1763.t1 a_30643_1763.n0 14.282
R18984 a_30643_1763.n0 a_30643_1763.t6 14.282
R18985 a_30643_1763.n0 a_30643_1763.n16 90.416
R18986 a_30643_1763.n16 a_30643_1763.n2 74.302
R18987 a_30643_1763.n16 a_30643_1763.n4 50.575
R18988 a_30643_1763.n4 a_30643_1763.n5 110.084
R18989 a_30643_1763.n2 a_30643_1763.n6 670.431
R18990 a_30643_1763.n6 a_30643_1763.n8 16.411
R18991 a_30643_1763.n8 a_30643_1763.t10 198.921
R18992 a_30643_1763.t10 a_30643_1763.t19 415.315
R18993 a_30643_1763.t19 a_30643_1763.n15 214.335
R18994 a_30643_1763.n15 a_30643_1763.t16 80.333
R18995 a_30643_1763.n15 a_30643_1763.t15 214.335
R18996 a_30643_1763.n8 a_30643_1763.n14 861.987
R18997 a_30643_1763.n14 a_30643_1763.n9 560.726
R18998 a_30643_1763.n14 a_30643_1763.n13 65.07
R18999 a_30643_1763.n13 a_30643_1763.n12 6.615
R19000 a_30643_1763.n12 a_30643_1763.t9 93.989
R19001 a_30643_1763.n12 a_30643_1763.t17 198.043
R19002 a_30643_1763.n13 a_30643_1763.n11 97.816
R19003 a_30643_1763.n11 a_30643_1763.t23 80.333
R19004 a_30643_1763.n11 a_30643_1763.t22 394.151
R19005 a_30643_1763.t22 a_30643_1763.n10 269.523
R19006 a_30643_1763.n10 a_30643_1763.t21 160.666
R19007 a_30643_1763.n10 a_30643_1763.t20 269.523
R19008 a_30643_1763.n9 a_30643_1763.t18 294.653
R19009 a_30643_1763.n9 a_30643_1763.t12 111.663
R19010 a_30643_1763.n6 a_30643_1763.t8 217.716
R19011 a_30643_1763.t8 a_30643_1763.t14 415.315
R19012 a_30643_1763.t14 a_30643_1763.n7 214.335
R19013 a_30643_1763.n7 a_30643_1763.t13 80.333
R19014 a_30643_1763.n7 a_30643_1763.t11 214.335
R19015 a_30643_1763.n5 a_30643_1763.t4 14.282
R19016 a_30643_1763.n5 a_30643_1763.t7 14.282
R19017 a_30643_1763.n4 a_30643_1763.n3 157.665
R19018 a_30643_1763.n3 a_30643_1763.t0 8.7
R19019 a_30643_1763.n3 a_30643_1763.t5 8.7
R19020 a_30643_1763.n2 a_30643_1763.n1 90.436
R19021 a_30643_1763.n1 a_30643_1763.t3 14.282
R19022 a_30643_1763.n1 a_30643_1763.t2 14.282
R19023 a_29950_1706.n8 a_29950_1706.n7 267.767
R19024 a_29950_1706.n1 a_29950_1706.t11 16.058
R19025 a_29950_1706.n3 a_29950_1706.t8 16.058
R19026 a_29950_1706.n0 a_29950_1706.t9 14.282
R19027 a_29950_1706.n0 a_29950_1706.t10 14.282
R19028 a_29950_1706.n2 a_29950_1706.t6 14.282
R19029 a_29950_1706.n2 a_29950_1706.t7 14.282
R19030 a_29950_1706.n5 a_29950_1706.t3 14.282
R19031 a_29950_1706.n5 a_29950_1706.t4 14.282
R19032 a_29950_1706.n7 a_29950_1706.t0 14.282
R19033 a_29950_1706.n7 a_29950_1706.t1 14.282
R19034 a_29950_1706.n9 a_29950_1706.t5 14.282
R19035 a_29950_1706.t2 a_29950_1706.n9 14.282
R19036 a_29950_1706.n6 a_29950_1706.n5 1.511
R19037 a_29950_1706.n1 a_29950_1706.n0 0.999
R19038 a_29950_1706.n3 a_29950_1706.n2 0.999
R19039 a_29950_1706.n8 a_29950_1706.n6 0.669
R19040 a_29950_1706.n4 a_29950_1706.n1 0.575
R19041 a_29950_1706.n6 a_29950_1706.n4 0.227
R19042 a_29950_1706.n4 a_29950_1706.n3 0.2
R19043 a_29950_1706.n9 a_29950_1706.n8 0.001
R19044 a_17040_20263.t0 a_17040_20263.t1 17.4
R19045 a_49968_14830.t0 a_49968_14830.t1 17.4
R19046 a_49319_15441.n0 a_49319_15441.t7 214.335
R19047 a_49319_15441.t10 a_49319_15441.n0 214.335
R19048 a_49319_15441.n1 a_49319_15441.t10 143.851
R19049 a_49319_15441.n1 a_49319_15441.t9 135.658
R19050 a_49319_15441.n0 a_49319_15441.t8 80.333
R19051 a_49319_15441.n4 a_49319_15441.t0 28.565
R19052 a_49319_15441.n4 a_49319_15441.t1 28.565
R19053 a_49319_15441.n2 a_49319_15441.t5 28.565
R19054 a_49319_15441.n2 a_49319_15441.t6 28.565
R19055 a_49319_15441.t2 a_49319_15441.n7 28.565
R19056 a_49319_15441.n7 a_49319_15441.t4 28.565
R19057 a_49319_15441.n5 a_49319_15441.t3 9.714
R19058 a_49319_15441.n5 a_49319_15441.n4 1.003
R19059 a_49319_15441.n6 a_49319_15441.n3 0.833
R19060 a_49319_15441.n3 a_49319_15441.n2 0.653
R19061 a_49319_15441.n7 a_49319_15441.n6 0.653
R19062 a_49319_15441.n6 a_49319_15441.n5 0.341
R19063 a_49319_15441.n3 a_49319_15441.n1 0.032
R19064 a_11100_10387.t0 a_11100_10387.t1 17.4
R19065 a_45035_3563.t5 a_45035_3563.t7 800.071
R19066 a_45035_3563.n2 a_45035_3563.n1 659.097
R19067 a_45035_3563.n0 a_45035_3563.t6 285.109
R19068 a_45035_3563.n1 a_45035_3563.t5 193.602
R19069 a_45035_3563.n4 a_45035_3563.n3 192.754
R19070 a_45035_3563.n0 a_45035_3563.t4 160.666
R19071 a_45035_3563.n1 a_45035_3563.n0 91.507
R19072 a_45035_3563.n3 a_45035_3563.t1 28.568
R19073 a_45035_3563.t2 a_45035_3563.n4 28.565
R19074 a_45035_3563.n4 a_45035_3563.t0 28.565
R19075 a_45035_3563.n2 a_45035_3563.t3 19.061
R19076 a_45035_3563.n3 a_45035_3563.n2 1.005
R19077 a_46770_3872.n0 a_46770_3872.t4 14.282
R19078 a_46770_3872.n0 a_46770_3872.t1 14.282
R19079 a_46770_3872.n1 a_46770_3872.t3 14.282
R19080 a_46770_3872.n1 a_46770_3872.t5 14.282
R19081 a_46770_3872.n3 a_46770_3872.t2 14.282
R19082 a_46770_3872.t0 a_46770_3872.n3 14.282
R19083 a_46770_3872.n3 a_46770_3872.n2 2.546
R19084 a_46770_3872.n2 a_46770_3872.n1 2.367
R19085 a_46770_3872.n2 a_46770_3872.n0 0.001
R19086 a_59921_1016.n1 a_59921_1016.t4 318.922
R19087 a_59921_1016.n0 a_59921_1016.t5 274.739
R19088 a_59921_1016.n0 a_59921_1016.t6 274.739
R19089 a_59921_1016.n1 a_59921_1016.t7 269.116
R19090 a_59921_1016.t4 a_59921_1016.n0 179.946
R19091 a_59921_1016.n2 a_59921_1016.n1 107.263
R19092 a_59921_1016.n3 a_59921_1016.t1 29.444
R19093 a_59921_1016.n4 a_59921_1016.t0 28.565
R19094 a_59921_1016.t2 a_59921_1016.n4 28.565
R19095 a_59921_1016.n2 a_59921_1016.t3 18.145
R19096 a_59921_1016.n3 a_59921_1016.n2 2.878
R19097 a_59921_1016.n4 a_59921_1016.n3 0.764
R19098 a_59509_1042.n0 a_59509_1042.n9 1.511
R19099 a_59509_1042.t0 a_59509_1042.n0 14.282
R19100 a_59509_1042.n0 a_59509_1042.t8 14.282
R19101 a_59509_1042.n9 a_59509_1042.n5 0.227
R19102 a_59509_1042.n9 a_59509_1042.n6 0.669
R19103 a_59509_1042.n6 a_59509_1042.n7 0.001
R19104 a_59509_1042.n6 a_59509_1042.n8 267.767
R19105 a_59509_1042.n8 a_59509_1042.t11 14.282
R19106 a_59509_1042.n8 a_59509_1042.t9 14.282
R19107 a_59509_1042.n7 a_59509_1042.t4 14.282
R19108 a_59509_1042.n7 a_59509_1042.t10 14.282
R19109 a_59509_1042.n5 a_59509_1042.n2 0.575
R19110 a_59509_1042.n5 a_59509_1042.n4 0.2
R19111 a_59509_1042.n4 a_59509_1042.t5 16.058
R19112 a_59509_1042.n4 a_59509_1042.n3 0.999
R19113 a_59509_1042.n3 a_59509_1042.t6 14.282
R19114 a_59509_1042.n3 a_59509_1042.t7 14.282
R19115 a_59509_1042.n2 a_59509_1042.n1 0.999
R19116 a_59509_1042.n1 a_59509_1042.t3 14.282
R19117 a_59509_1042.n1 a_59509_1042.t1 14.282
R19118 a_59509_1042.n2 a_59509_1042.t2 16.058
R19119 a_41493_21373.n0 a_41493_21373.t5 14.282
R19120 a_41493_21373.t3 a_41493_21373.n0 14.282
R19121 a_41493_21373.n0 a_41493_21373.n9 0.999
R19122 a_41493_21373.n6 a_41493_21373.n8 0.575
R19123 a_41493_21373.n9 a_41493_21373.n6 0.2
R19124 a_41493_21373.n9 a_41493_21373.t4 16.058
R19125 a_41493_21373.n8 a_41493_21373.n7 0.999
R19126 a_41493_21373.n7 a_41493_21373.t1 14.282
R19127 a_41493_21373.n7 a_41493_21373.t0 14.282
R19128 a_41493_21373.n8 a_41493_21373.t2 16.058
R19129 a_41493_21373.n6 a_41493_21373.n4 0.227
R19130 a_41493_21373.n4 a_41493_21373.n5 1.511
R19131 a_41493_21373.n5 a_41493_21373.t8 14.282
R19132 a_41493_21373.n5 a_41493_21373.t7 14.282
R19133 a_41493_21373.n4 a_41493_21373.n1 0.669
R19134 a_41493_21373.n1 a_41493_21373.n2 0.001
R19135 a_41493_21373.n1 a_41493_21373.n3 267.767
R19136 a_41493_21373.n3 a_41493_21373.t10 14.282
R19137 a_41493_21373.n3 a_41493_21373.t11 14.282
R19138 a_41493_21373.n2 a_41493_21373.t6 14.282
R19139 a_41493_21373.n2 a_41493_21373.t9 14.282
R19140 a_48418_21344.n1 a_48418_21344.t5 318.922
R19141 a_48418_21344.n0 a_48418_21344.t4 274.739
R19142 a_48418_21344.n0 a_48418_21344.t6 274.739
R19143 a_48418_21344.n1 a_48418_21344.t7 269.116
R19144 a_48418_21344.t5 a_48418_21344.n0 179.946
R19145 a_48418_21344.n2 a_48418_21344.n1 107.263
R19146 a_48418_21344.n3 a_48418_21344.t1 29.444
R19147 a_48418_21344.t2 a_48418_21344.n4 28.565
R19148 a_48418_21344.n4 a_48418_21344.t0 28.565
R19149 a_48418_21344.n2 a_48418_21344.t3 18.145
R19150 a_48418_21344.n3 a_48418_21344.n2 2.878
R19151 a_48418_21344.n4 a_48418_21344.n3 0.764
R19152 a_60980_1735.n1 a_60980_1735.t6 318.922
R19153 a_60980_1735.n0 a_60980_1735.t4 273.935
R19154 a_60980_1735.n0 a_60980_1735.t5 273.935
R19155 a_60980_1735.n1 a_60980_1735.t7 269.116
R19156 a_60980_1735.n4 a_60980_1735.n3 193.227
R19157 a_60980_1735.t6 a_60980_1735.n0 179.142
R19158 a_60980_1735.n2 a_60980_1735.n1 106.999
R19159 a_60980_1735.n3 a_60980_1735.t1 28.568
R19160 a_60980_1735.n4 a_60980_1735.t0 28.565
R19161 a_60980_1735.t2 a_60980_1735.n4 28.565
R19162 a_60980_1735.n2 a_60980_1735.t3 18.149
R19163 a_60980_1735.n3 a_60980_1735.n2 3.726
R19164 a_39681_1042.t6 a_39681_1042.n0 14.282
R19165 a_39681_1042.n0 a_39681_1042.t11 14.282
R19166 a_39681_1042.n0 a_39681_1042.n9 0.999
R19167 a_39681_1042.n9 a_39681_1042.n6 0.575
R19168 a_39681_1042.n6 a_39681_1042.n8 0.2
R19169 a_39681_1042.n8 a_39681_1042.t4 16.058
R19170 a_39681_1042.n8 a_39681_1042.n7 0.999
R19171 a_39681_1042.n7 a_39681_1042.t3 14.282
R19172 a_39681_1042.n7 a_39681_1042.t5 14.282
R19173 a_39681_1042.n9 a_39681_1042.t7 16.058
R19174 a_39681_1042.n6 a_39681_1042.n4 0.227
R19175 a_39681_1042.n4 a_39681_1042.n5 1.511
R19176 a_39681_1042.n5 a_39681_1042.t0 14.282
R19177 a_39681_1042.n5 a_39681_1042.t1 14.282
R19178 a_39681_1042.n4 a_39681_1042.n1 0.669
R19179 a_39681_1042.n1 a_39681_1042.n2 0.001
R19180 a_39681_1042.n1 a_39681_1042.n3 267.767
R19181 a_39681_1042.n3 a_39681_1042.t10 14.282
R19182 a_39681_1042.n3 a_39681_1042.t8 14.282
R19183 a_39681_1042.n2 a_39681_1042.t2 14.282
R19184 a_39681_1042.n2 a_39681_1042.t9 14.282
R19185 a_46232_1040.t6 a_46232_1040.n0 14.282
R19186 a_46232_1040.n0 a_46232_1040.t8 14.282
R19187 a_46232_1040.n0 a_46232_1040.n9 0.999
R19188 a_46232_1040.n6 a_46232_1040.n8 0.575
R19189 a_46232_1040.n9 a_46232_1040.n6 0.2
R19190 a_46232_1040.n9 a_46232_1040.t7 16.058
R19191 a_46232_1040.n8 a_46232_1040.n7 0.999
R19192 a_46232_1040.n7 a_46232_1040.t2 14.282
R19193 a_46232_1040.n7 a_46232_1040.t1 14.282
R19194 a_46232_1040.n8 a_46232_1040.t0 16.058
R19195 a_46232_1040.n6 a_46232_1040.n4 0.227
R19196 a_46232_1040.n4 a_46232_1040.n5 1.511
R19197 a_46232_1040.n5 a_46232_1040.t4 14.282
R19198 a_46232_1040.n5 a_46232_1040.t5 14.282
R19199 a_46232_1040.n4 a_46232_1040.n1 0.669
R19200 a_46232_1040.n1 a_46232_1040.n2 0.001
R19201 a_46232_1040.n1 a_46232_1040.n3 267.767
R19202 a_46232_1040.n3 a_46232_1040.t9 14.282
R19203 a_46232_1040.n3 a_46232_1040.t10 14.282
R19204 a_46232_1040.n2 a_46232_1040.t3 14.282
R19205 a_46232_1040.n2 a_46232_1040.t11 14.282
R19206 a_21860_15776.t0 a_21860_15776.t1 17.4
R19207 a_23135_20719.n3 a_23135_20719.t6 448.381
R19208 a_23135_20719.n2 a_23135_20719.t5 286.438
R19209 a_23135_20719.n2 a_23135_20719.t7 286.438
R19210 a_23135_20719.n1 a_23135_20719.t4 247.69
R19211 a_23135_20719.n4 a_23135_20719.n0 182.117
R19212 a_23135_20719.t6 a_23135_20719.n2 160.666
R19213 a_23135_20719.t2 a_23135_20719.n4 28.568
R19214 a_23135_20719.n0 a_23135_20719.t0 28.565
R19215 a_23135_20719.n0 a_23135_20719.t1 28.565
R19216 a_23135_20719.n1 a_23135_20719.t3 18.127
R19217 a_23135_20719.n3 a_23135_20719.n1 4.036
R19218 a_23135_20719.n4 a_23135_20719.n3 0.937
R19219 a_23080_20259.t0 a_23080_20259.t1 17.4
R19220 a_56011_22058.n1 a_56011_22058.t6 318.922
R19221 a_56011_22058.n0 a_56011_22058.t5 273.935
R19222 a_56011_22058.n0 a_56011_22058.t7 273.935
R19223 a_56011_22058.n1 a_56011_22058.t4 269.116
R19224 a_56011_22058.n4 a_56011_22058.n3 193.227
R19225 a_56011_22058.t6 a_56011_22058.n0 179.142
R19226 a_56011_22058.n2 a_56011_22058.n1 106.999
R19227 a_56011_22058.n3 a_56011_22058.t1 28.568
R19228 a_56011_22058.t2 a_56011_22058.n4 28.565
R19229 a_56011_22058.n4 a_56011_22058.t0 28.565
R19230 a_56011_22058.n2 a_56011_22058.t3 18.149
R19231 a_56011_22058.n3 a_56011_22058.n2 3.726
R19232 a_13429_1740.n0 a_13429_1740.t2 14.282
R19233 a_13429_1740.t0 a_13429_1740.n0 14.282
R19234 a_13429_1740.n0 a_13429_1740.n9 89.977
R19235 a_13429_1740.n9 a_13429_1740.n7 75.815
R19236 a_13429_1740.n9 a_13429_1740.n6 77.456
R19237 a_13429_1740.n6 a_13429_1740.n4 77.456
R19238 a_13429_1740.n4 a_13429_1740.n2 77.784
R19239 a_13429_1740.n7 a_13429_1740.n8 167.433
R19240 a_13429_1740.n8 a_13429_1740.t7 14.282
R19241 a_13429_1740.n8 a_13429_1740.t6 14.282
R19242 a_13429_1740.n7 a_13429_1740.t8 104.259
R19243 a_13429_1740.n6 a_13429_1740.n5 89.977
R19244 a_13429_1740.n5 a_13429_1740.t1 14.282
R19245 a_13429_1740.n5 a_13429_1740.t4 14.282
R19246 a_13429_1740.n4 a_13429_1740.n3 89.977
R19247 a_13429_1740.n3 a_13429_1740.t3 14.282
R19248 a_13429_1740.n3 a_13429_1740.t5 14.282
R19249 a_13429_1740.n2 a_13429_1740.t9 104.259
R19250 a_13429_1740.n2 a_13429_1740.n1 167.433
R19251 a_13429_1740.n1 a_13429_1740.t11 14.282
R19252 a_13429_1740.n1 a_13429_1740.t10 14.282
R19253 a_51114_2351.n0 a_51114_2351.t10 214.335
R19254 a_51114_2351.t9 a_51114_2351.n0 214.335
R19255 a_51114_2351.n1 a_51114_2351.t9 143.851
R19256 a_51114_2351.n1 a_51114_2351.t8 135.658
R19257 a_51114_2351.n0 a_51114_2351.t7 80.333
R19258 a_51114_2351.n2 a_51114_2351.t4 28.565
R19259 a_51114_2351.n2 a_51114_2351.t6 28.565
R19260 a_51114_2351.n4 a_51114_2351.t5 28.565
R19261 a_51114_2351.n4 a_51114_2351.t1 28.565
R19262 a_51114_2351.n7 a_51114_2351.t0 28.565
R19263 a_51114_2351.t2 a_51114_2351.n7 28.565
R19264 a_51114_2351.n6 a_51114_2351.t3 9.714
R19265 a_51114_2351.n7 a_51114_2351.n6 1.003
R19266 a_51114_2351.n5 a_51114_2351.n3 0.833
R19267 a_51114_2351.n3 a_51114_2351.n2 0.653
R19268 a_51114_2351.n5 a_51114_2351.n4 0.653
R19269 a_51114_2351.n6 a_51114_2351.n5 0.341
R19270 a_51114_2351.n3 a_51114_2351.n1 0.032
R19271 a_42266_11512.n5 a_42266_11512.n4 535.449
R19272 a_42266_11512.t18 a_42266_11512.t16 437.233
R19273 a_42266_11512.t13 a_42266_11512.t10 437.233
R19274 a_42266_11512.t9 a_42266_11512.n2 313.873
R19275 a_42266_11512.n4 a_42266_11512.t14 294.986
R19276 a_42266_11512.n1 a_42266_11512.t17 272.288
R19277 a_42266_11512.n5 a_42266_11512.t11 245.184
R19278 a_42266_11512.n7 a_42266_11512.t13 218.628
R19279 a_42266_11512.n9 a_42266_11512.t18 217.024
R19280 a_42266_11512.n8 a_42266_11512.t19 214.686
R19281 a_42266_11512.t16 a_42266_11512.n8 214.686
R19282 a_42266_11512.n6 a_42266_11512.t8 214.686
R19283 a_42266_11512.t10 a_42266_11512.n6 214.686
R19284 a_42266_11512.n11 a_42266_11512.n0 192.754
R19285 a_42266_11512.n3 a_42266_11512.t9 190.152
R19286 a_42266_11512.n3 a_42266_11512.t4 190.152
R19287 a_42266_11512.n1 a_42266_11512.t12 160.666
R19288 a_42266_11512.n2 a_42266_11512.t6 160.666
R19289 a_42266_11512.n4 a_42266_11512.t7 110.859
R19290 a_42266_11512.n2 a_42266_11512.n1 96.129
R19291 a_42266_11512.n8 a_42266_11512.t5 80.333
R19292 a_42266_11512.t11 a_42266_11512.n3 80.333
R19293 a_42266_11512.n6 a_42266_11512.t15 80.333
R19294 a_42266_11512.t0 a_42266_11512.n11 28.568
R19295 a_42266_11512.n0 a_42266_11512.t3 28.565
R19296 a_42266_11512.n0 a_42266_11512.t2 28.565
R19297 a_42266_11512.n10 a_42266_11512.t1 18.819
R19298 a_42266_11512.n7 a_42266_11512.n5 14.9
R19299 a_42266_11512.n10 a_42266_11512.n9 2.96
R19300 a_42266_11512.n9 a_42266_11512.n7 2.599
R19301 a_42266_11512.n11 a_42266_11512.n10 1.098
R19302 a_41697_310.t0 a_41697_310.t1 380.209
R19303 a_55504_n1325.n7 a_55504_n1325.n6 861.987
R19304 a_55504_n1325.n6 a_55504_n1325.n5 560.726
R19305 a_55504_n1325.t4 a_55504_n1325.t18 415.315
R19306 a_55504_n1325.t11 a_55504_n1325.t12 415.315
R19307 a_55504_n1325.n2 a_55504_n1325.t15 394.151
R19308 a_55504_n1325.n5 a_55504_n1325.t6 294.653
R19309 a_55504_n1325.n1 a_55504_n1325.t19 269.523
R19310 a_55504_n1325.t15 a_55504_n1325.n1 269.523
R19311 a_55504_n1325.n9 a_55504_n1325.t4 217.716
R19312 a_55504_n1325.n8 a_55504_n1325.t7 214.335
R19313 a_55504_n1325.t18 a_55504_n1325.n8 214.335
R19314 a_55504_n1325.n0 a_55504_n1325.t13 214.335
R19315 a_55504_n1325.t12 a_55504_n1325.n0 214.335
R19316 a_55504_n1325.n7 a_55504_n1325.t11 198.921
R19317 a_55504_n1325.n3 a_55504_n1325.t8 198.043
R19318 a_55504_n1325.n12 a_55504_n1325.n11 192.754
R19319 a_55504_n1325.n1 a_55504_n1325.t9 160.666
R19320 a_55504_n1325.n5 a_55504_n1325.t5 111.663
R19321 a_55504_n1325.n4 a_55504_n1325.n2 97.816
R19322 a_55504_n1325.n3 a_55504_n1325.t16 93.989
R19323 a_55504_n1325.n8 a_55504_n1325.t14 80.333
R19324 a_55504_n1325.n2 a_55504_n1325.t10 80.333
R19325 a_55504_n1325.n0 a_55504_n1325.t17 80.333
R19326 a_55504_n1325.n6 a_55504_n1325.n4 65.07
R19327 a_55504_n1325.n11 a_55504_n1325.t0 28.568
R19328 a_55504_n1325.n12 a_55504_n1325.t1 28.565
R19329 a_55504_n1325.t2 a_55504_n1325.n12 28.565
R19330 a_55504_n1325.n10 a_55504_n1325.t3 18.827
R19331 a_55504_n1325.n9 a_55504_n1325.n7 16.411
R19332 a_55504_n1325.n4 a_55504_n1325.n3 6.615
R19333 a_55504_n1325.n10 a_55504_n1325.n9 4.58
R19334 a_55504_n1325.n11 a_55504_n1325.n10 1.105
R19335 a_57959_3365.t0 a_57959_3365.t1 17.4
R19336 a_17692_7659.t0 a_17692_7659.t1 17.4
R19337 a_498_14458.n2 a_498_14458.t5 867.497
R19338 a_498_14458.n2 a_498_14458.t7 591.811
R19339 a_498_14458.n1 a_498_14458.t4 286.438
R19340 a_498_14458.n1 a_498_14458.t6 286.438
R19341 a_498_14458.n4 a_498_14458.n0 185.55
R19342 a_498_14458.t5 a_498_14458.n1 160.666
R19343 a_498_14458.t2 a_498_14458.n4 28.568
R19344 a_498_14458.n0 a_498_14458.t0 28.565
R19345 a_498_14458.n0 a_498_14458.t1 28.565
R19346 a_498_14458.n3 a_498_14458.n2 25.537
R19347 a_498_14458.n3 a_498_14458.t3 21.376
R19348 a_498_14458.n4 a_498_14458.n3 1.637
R19349 a_6071_6357.n2 a_6071_6357.t7 990.34
R19350 a_6071_6357.n2 a_6071_6357.t5 408.211
R19351 a_6071_6357.n1 a_6071_6357.t6 286.438
R19352 a_6071_6357.n1 a_6071_6357.t4 286.438
R19353 a_6071_6357.n4 a_6071_6357.n0 197.272
R19354 a_6071_6357.t7 a_6071_6357.n1 160.666
R19355 a_6071_6357.n3 a_6071_6357.n2 32.172
R19356 a_6071_6357.t2 a_6071_6357.n4 28.568
R19357 a_6071_6357.n0 a_6071_6357.t1 28.565
R19358 a_6071_6357.n0 a_6071_6357.t0 28.565
R19359 a_6071_6357.n3 a_6071_6357.t3 18.103
R19360 a_6071_6357.n4 a_6071_6357.n3 0.459
R19361 a_57684_8194.n6 a_57684_8194.n5 501.28
R19362 a_57684_8194.t6 a_57684_8194.t18 437.233
R19363 a_57684_8194.t13 a_57684_8194.t5 415.315
R19364 a_57684_8194.t10 a_57684_8194.n3 313.873
R19365 a_57684_8194.n5 a_57684_8194.t14 294.986
R19366 a_57684_8194.n2 a_57684_8194.t11 272.288
R19367 a_57684_8194.n6 a_57684_8194.t19 236.01
R19368 a_57684_8194.n9 a_57684_8194.t6 216.627
R19369 a_57684_8194.n7 a_57684_8194.t13 216.111
R19370 a_57684_8194.n8 a_57684_8194.t17 214.686
R19371 a_57684_8194.t18 a_57684_8194.n8 214.686
R19372 a_57684_8194.n1 a_57684_8194.t8 214.335
R19373 a_57684_8194.t5 a_57684_8194.n1 214.335
R19374 a_57684_8194.n4 a_57684_8194.t10 190.152
R19375 a_57684_8194.n4 a_57684_8194.t12 190.152
R19376 a_57684_8194.n2 a_57684_8194.t4 160.666
R19377 a_57684_8194.n3 a_57684_8194.t15 160.666
R19378 a_57684_8194.n7 a_57684_8194.n6 148.428
R19379 a_57684_8194.n5 a_57684_8194.t7 110.859
R19380 a_57684_8194.n3 a_57684_8194.n2 96.129
R19381 a_57684_8194.n8 a_57684_8194.t9 80.333
R19382 a_57684_8194.n1 a_57684_8194.t16 80.333
R19383 a_57684_8194.t19 a_57684_8194.n4 80.333
R19384 a_57684_8194.n0 a_57684_8194.t1 28.57
R19385 a_57684_8194.n11 a_57684_8194.t3 28.565
R19386 a_57684_8194.t0 a_57684_8194.n11 28.565
R19387 a_57684_8194.n0 a_57684_8194.t2 17.638
R19388 a_57684_8194.n10 a_57684_8194.n9 11.942
R19389 a_57684_8194.n9 a_57684_8194.n7 2.923
R19390 a_57684_8194.n11 a_57684_8194.n10 0.69
R19391 a_57684_8194.n10 a_57684_8194.n0 0.6
R19392 a_59901_23892.t4 a_59901_23892.t7 800.071
R19393 a_59901_23892.n2 a_59901_23892.n1 659.097
R19394 a_59901_23892.n0 a_59901_23892.t6 285.109
R19395 a_59901_23892.n1 a_59901_23892.t4 193.602
R19396 a_59901_23892.n4 a_59901_23892.n3 192.754
R19397 a_59901_23892.n0 a_59901_23892.t5 160.666
R19398 a_59901_23892.n1 a_59901_23892.n0 91.507
R19399 a_59901_23892.n3 a_59901_23892.t0 28.568
R19400 a_59901_23892.n4 a_59901_23892.t1 28.565
R19401 a_59901_23892.t2 a_59901_23892.n4 28.565
R19402 a_59901_23892.n2 a_59901_23892.t3 19.061
R19403 a_59901_23892.n3 a_59901_23892.n2 1.005
R19404 a_38501_6091.t6 a_38501_6091.t4 574.43
R19405 a_38501_6091.n0 a_38501_6091.t7 285.109
R19406 a_38501_6091.n2 a_38501_6091.n1 197.217
R19407 a_38501_6091.n4 a_38501_6091.n3 192.754
R19408 a_38501_6091.n0 a_38501_6091.t5 160.666
R19409 a_38501_6091.n1 a_38501_6091.t6 160.666
R19410 a_38501_6091.n1 a_38501_6091.n0 114.829
R19411 a_38501_6091.n3 a_38501_6091.t3 28.568
R19412 a_38501_6091.t0 a_38501_6091.n4 28.565
R19413 a_38501_6091.n4 a_38501_6091.t2 28.565
R19414 a_38501_6091.n2 a_38501_6091.t1 18.838
R19415 a_38501_6091.n3 a_38501_6091.n2 1.129
R19416 a_40109_9654.t5 a_40109_9654.n2 404.877
R19417 a_40109_9654.n1 a_40109_9654.t7 210.902
R19418 a_40109_9654.n3 a_40109_9654.t5 136.943
R19419 a_40109_9654.n2 a_40109_9654.n1 107.801
R19420 a_40109_9654.n1 a_40109_9654.t8 80.333
R19421 a_40109_9654.n2 a_40109_9654.t6 80.333
R19422 a_40109_9654.n0 a_40109_9654.t0 17.4
R19423 a_40109_9654.n0 a_40109_9654.t1 17.4
R19424 a_40109_9654.n4 a_40109_9654.t3 15.032
R19425 a_40109_9654.t2 a_40109_9654.n5 14.282
R19426 a_40109_9654.n5 a_40109_9654.t4 14.282
R19427 a_40109_9654.n5 a_40109_9654.n4 1.65
R19428 a_40109_9654.n3 a_40109_9654.n0 0.672
R19429 a_40109_9654.n4 a_40109_9654.n3 0.665
R19430 a_44451_9870.n0 a_44451_9870.t9 214.335
R19431 a_44451_9870.t8 a_44451_9870.n0 214.335
R19432 a_44451_9870.n1 a_44451_9870.t8 143.851
R19433 a_44451_9870.n1 a_44451_9870.t7 135.658
R19434 a_44451_9870.n0 a_44451_9870.t10 80.333
R19435 a_44451_9870.n2 a_44451_9870.t4 28.565
R19436 a_44451_9870.n2 a_44451_9870.t6 28.565
R19437 a_44451_9870.n4 a_44451_9870.t5 28.565
R19438 a_44451_9870.n4 a_44451_9870.t1 28.565
R19439 a_44451_9870.t2 a_44451_9870.n7 28.565
R19440 a_44451_9870.n7 a_44451_9870.t0 28.565
R19441 a_44451_9870.n6 a_44451_9870.t3 9.714
R19442 a_44451_9870.n7 a_44451_9870.n6 1.003
R19443 a_44451_9870.n5 a_44451_9870.n3 0.833
R19444 a_44451_9870.n3 a_44451_9870.n2 0.653
R19445 a_44451_9870.n5 a_44451_9870.n4 0.653
R19446 a_44451_9870.n6 a_44451_9870.n5 0.341
R19447 a_44451_9870.n3 a_44451_9870.n1 0.032
R19448 a_64188_3841.n5 a_64188_3841.n4 465.933
R19449 a_64188_3841.t11 a_64188_3841.t5 415.315
R19450 a_64188_3841.n1 a_64188_3841.t6 394.151
R19451 a_64188_3841.n4 a_64188_3841.t4 294.653
R19452 a_64188_3841.n0 a_64188_3841.t10 269.523
R19453 a_64188_3841.t6 a_64188_3841.n0 269.523
R19454 a_64188_3841.n7 a_64188_3841.t11 220.285
R19455 a_64188_3841.n6 a_64188_3841.t9 214.335
R19456 a_64188_3841.t5 a_64188_3841.n6 214.335
R19457 a_64188_3841.n2 a_64188_3841.t14 198.043
R19458 a_64188_3841.n10 a_64188_3841.n9 192.754
R19459 a_64188_3841.n5 a_64188_3841.n3 163.88
R19460 a_64188_3841.n0 a_64188_3841.t15 160.666
R19461 a_64188_3841.n4 a_64188_3841.t8 111.663
R19462 a_64188_3841.n3 a_64188_3841.n1 97.816
R19463 a_64188_3841.n2 a_64188_3841.t7 93.989
R19464 a_64188_3841.n6 a_64188_3841.t13 80.333
R19465 a_64188_3841.n1 a_64188_3841.t12 80.333
R19466 a_64188_3841.n7 a_64188_3841.n5 61.538
R19467 a_64188_3841.n9 a_64188_3841.t1 28.568
R19468 a_64188_3841.n10 a_64188_3841.t0 28.565
R19469 a_64188_3841.t2 a_64188_3841.n10 28.565
R19470 a_64188_3841.n8 a_64188_3841.t3 18.824
R19471 a_64188_3841.n3 a_64188_3841.n2 6.615
R19472 a_64188_3841.n8 a_64188_3841.n7 5.5
R19473 a_64188_3841.n9 a_64188_3841.n8 1.105
R19474 a_46644_1014.n1 a_46644_1014.t4 318.922
R19475 a_46644_1014.n0 a_46644_1014.t5 274.739
R19476 a_46644_1014.n0 a_46644_1014.t7 274.739
R19477 a_46644_1014.n1 a_46644_1014.t6 269.116
R19478 a_46644_1014.t4 a_46644_1014.n0 179.946
R19479 a_46644_1014.n2 a_46644_1014.n1 107.263
R19480 a_46644_1014.n3 a_46644_1014.t1 29.444
R19481 a_46644_1014.n4 a_46644_1014.t0 28.565
R19482 a_46644_1014.t2 a_46644_1014.n4 28.565
R19483 a_46644_1014.n2 a_46644_1014.t3 18.145
R19484 a_46644_1014.n3 a_46644_1014.n2 2.878
R19485 a_46644_1014.n4 a_46644_1014.n3 0.764
R19486 a_17447_1255.n1 a_17447_1255.t6 867.497
R19487 a_17447_1255.n1 a_17447_1255.t4 615.911
R19488 a_17447_1255.n0 a_17447_1255.t5 286.438
R19489 a_17447_1255.n0 a_17447_1255.t7 286.438
R19490 a_17447_1255.n4 a_17447_1255.n3 185.55
R19491 a_17447_1255.t6 a_17447_1255.n0 160.666
R19492 a_17447_1255.n2 a_17447_1255.n1 128.838
R19493 a_17447_1255.n3 a_17447_1255.t0 28.568
R19494 a_17447_1255.n4 a_17447_1255.t1 28.565
R19495 a_17447_1255.t2 a_17447_1255.n4 28.565
R19496 a_17447_1255.n2 a_17447_1255.t3 20.393
R19497 a_17447_1255.n3 a_17447_1255.n2 1.834
R19498 a_17394_407.t0 a_17394_407.t1 17.4
R19499 a_248_1740.n2 a_248_1740.t5 448.382
R19500 a_248_1740.n1 a_248_1740.t7 286.438
R19501 a_248_1740.n1 a_248_1740.t4 286.438
R19502 a_248_1740.n0 a_248_1740.t6 247.69
R19503 a_248_1740.n4 a_248_1740.n3 182.117
R19504 a_248_1740.t5 a_248_1740.n1 160.666
R19505 a_248_1740.n3 a_248_1740.t0 28.568
R19506 a_248_1740.t2 a_248_1740.n4 28.565
R19507 a_248_1740.n4 a_248_1740.t1 28.565
R19508 a_248_1740.n0 a_248_1740.t3 18.127
R19509 a_248_1740.n2 a_248_1740.n0 4.039
R19510 a_248_1740.n3 a_248_1740.n2 0.937
R19511 a_54363_7535.n1 a_54363_7535.t6 318.922
R19512 a_54363_7535.n0 a_54363_7535.t4 273.935
R19513 a_54363_7535.n0 a_54363_7535.t7 273.935
R19514 a_54363_7535.n1 a_54363_7535.t5 269.116
R19515 a_54363_7535.n4 a_54363_7535.n3 193.227
R19516 a_54363_7535.t6 a_54363_7535.n0 179.142
R19517 a_54363_7535.n2 a_54363_7535.n1 106.999
R19518 a_54363_7535.n3 a_54363_7535.t1 28.568
R19519 a_54363_7535.n4 a_54363_7535.t0 28.565
R19520 a_54363_7535.t2 a_54363_7535.n4 28.565
R19521 a_54363_7535.n2 a_54363_7535.t3 18.149
R19522 a_54363_7535.n3 a_54363_7535.n2 3.726
R19523 a_47711_18567.t7 a_47711_18567.t4 574.43
R19524 a_47711_18567.n1 a_47711_18567.t5 285.109
R19525 a_47711_18567.n3 a_47711_18567.n2 197.215
R19526 a_47711_18567.n4 a_47711_18567.n0 192.754
R19527 a_47711_18567.n1 a_47711_18567.t6 160.666
R19528 a_47711_18567.n2 a_47711_18567.t7 160.666
R19529 a_47711_18567.n2 a_47711_18567.n1 114.829
R19530 a_47711_18567.t2 a_47711_18567.n4 28.568
R19531 a_47711_18567.n0 a_47711_18567.t0 28.565
R19532 a_47711_18567.n0 a_47711_18567.t1 28.565
R19533 a_47711_18567.n3 a_47711_18567.t3 18.838
R19534 a_47711_18567.n4 a_47711_18567.n3 1.129
R19535 a_13778_1740.t1 a_13778_1740.n0 14.282
R19536 a_13778_1740.n0 a_13778_1740.t2 14.282
R19537 a_13778_1740.n0 a_13778_1740.n1 258.161
R19538 a_13778_1740.n1 a_13778_1740.n7 4.366
R19539 a_13778_1740.n7 a_13778_1740.n5 0.852
R19540 a_13778_1740.n5 a_13778_1740.n6 258.161
R19541 a_13778_1740.n6 a_13778_1740.t5 14.282
R19542 a_13778_1740.n6 a_13778_1740.t7 14.282
R19543 a_13778_1740.n5 a_13778_1740.t6 14.283
R19544 a_13778_1740.n7 a_13778_1740.n4 97.614
R19545 a_13778_1740.n4 a_13778_1740.t11 200.029
R19546 a_13778_1740.t11 a_13778_1740.n3 206.421
R19547 a_13778_1740.n3 a_13778_1740.t8 80.333
R19548 a_13778_1740.n3 a_13778_1740.t9 206.421
R19549 a_13778_1740.n4 a_13778_1740.t10 1527.4
R19550 a_13778_1740.t10 a_13778_1740.n2 657.379
R19551 a_13778_1740.n2 a_13778_1740.t4 8.7
R19552 a_13778_1740.n2 a_13778_1740.t0 8.7
R19553 a_13778_1740.n1 a_13778_1740.t3 14.283
R19554 a_14335_n2637.n1 a_14335_n2637.t6 867.497
R19555 a_14335_n2637.n1 a_14335_n2637.t5 615.911
R19556 a_14335_n2637.n0 a_14335_n2637.t4 286.438
R19557 a_14335_n2637.n0 a_14335_n2637.t7 286.438
R19558 a_14335_n2637.n4 a_14335_n2637.n3 185.55
R19559 a_14335_n2637.t6 a_14335_n2637.n0 160.666
R19560 a_14335_n2637.n3 a_14335_n2637.t0 28.568
R19561 a_14335_n2637.t2 a_14335_n2637.n4 28.565
R19562 a_14335_n2637.n4 a_14335_n2637.t1 28.565
R19563 a_14335_n2637.n2 a_14335_n2637.n1 22.12
R19564 a_14335_n2637.n2 a_14335_n2637.t3 20.393
R19565 a_14335_n2637.n3 a_14335_n2637.n2 1.842
R19566 a_18824_20866.t0 a_18824_20866.n0 14.282
R19567 a_18824_20866.n0 a_18824_20866.t1 14.282
R19568 a_18824_20866.n0 a_18824_20866.n1 258.161
R19569 a_18824_20866.n1 a_18824_20866.t3 14.283
R19570 a_18824_20866.n1 a_18824_20866.n7 4.366
R19571 a_18824_20866.n7 a_18824_20866.n5 0.852
R19572 a_18824_20866.n5 a_18824_20866.n6 258.161
R19573 a_18824_20866.n6 a_18824_20866.t6 14.282
R19574 a_18824_20866.n6 a_18824_20866.t5 14.282
R19575 a_18824_20866.n5 a_18824_20866.t7 14.283
R19576 a_18824_20866.n7 a_18824_20866.n4 97.614
R19577 a_18824_20866.n4 a_18824_20866.t9 200.029
R19578 a_18824_20866.t9 a_18824_20866.n3 206.421
R19579 a_18824_20866.n3 a_18824_20866.t10 80.333
R19580 a_18824_20866.n3 a_18824_20866.t8 206.421
R19581 a_18824_20866.n4 a_18824_20866.t11 1527.4
R19582 a_18824_20866.t11 a_18824_20866.n2 657.379
R19583 a_18824_20866.n2 a_18824_20866.t2 8.7
R19584 a_18824_20866.n2 a_18824_20866.t4 8.7
R19585 a_6832_10990.n0 a_6832_10990.t1 14.282
R19586 a_6832_10990.t0 a_6832_10990.n0 14.282
R19587 a_6832_10990.n0 a_6832_10990.n1 258.161
R19588 a_6832_10990.n1 a_6832_10990.n5 0.852
R19589 a_6832_10990.n5 a_6832_10990.n6 4.366
R19590 a_6832_10990.n6 a_6832_10990.n7 258.161
R19591 a_6832_10990.n7 a_6832_10990.t5 14.282
R19592 a_6832_10990.n7 a_6832_10990.t6 14.282
R19593 a_6832_10990.n6 a_6832_10990.t3 14.283
R19594 a_6832_10990.n5 a_6832_10990.n4 97.614
R19595 a_6832_10990.n4 a_6832_10990.t10 200.029
R19596 a_6832_10990.t10 a_6832_10990.n3 206.421
R19597 a_6832_10990.n3 a_6832_10990.t11 80.333
R19598 a_6832_10990.n3 a_6832_10990.t8 206.421
R19599 a_6832_10990.n4 a_6832_10990.t9 1527.4
R19600 a_6832_10990.t9 a_6832_10990.n2 657.379
R19601 a_6832_10990.n2 a_6832_10990.t4 8.7
R19602 a_6832_10990.n2 a_6832_10990.t7 8.7
R19603 a_6832_10990.n1 a_6832_10990.t2 14.283
R19604 a_22172_5352.t3 a_22172_5352.n7 16.058
R19605 a_22172_5352.n7 a_22172_5352.n5 0.2
R19606 a_22172_5352.n5 a_22172_5352.n9 0.575
R19607 a_22172_5352.n9 a_22172_5352.t8 16.058
R19608 a_22172_5352.n9 a_22172_5352.n8 0.999
R19609 a_22172_5352.n8 a_22172_5352.t7 14.282
R19610 a_22172_5352.n8 a_22172_5352.t9 14.282
R19611 a_22172_5352.n7 a_22172_5352.n6 0.999
R19612 a_22172_5352.n6 a_22172_5352.t11 14.282
R19613 a_22172_5352.n6 a_22172_5352.t10 14.282
R19614 a_22172_5352.n5 a_22172_5352.n3 0.227
R19615 a_22172_5352.n3 a_22172_5352.n4 1.511
R19616 a_22172_5352.n4 a_22172_5352.t6 14.282
R19617 a_22172_5352.n4 a_22172_5352.t4 14.282
R19618 a_22172_5352.n3 a_22172_5352.n0 0.669
R19619 a_22172_5352.n0 a_22172_5352.n1 0.001
R19620 a_22172_5352.n0 a_22172_5352.n2 267.767
R19621 a_22172_5352.n2 a_22172_5352.t0 14.282
R19622 a_22172_5352.n2 a_22172_5352.t2 14.282
R19623 a_22172_5352.n1 a_22172_5352.t1 14.282
R19624 a_22172_5352.n1 a_22172_5352.t5 14.282
R19625 a_49963_16434.t0 a_49963_16434.t1 17.4
R19626 a_49314_17045.n0 a_49314_17045.t8 214.335
R19627 a_49314_17045.t10 a_49314_17045.n0 214.335
R19628 a_49314_17045.n1 a_49314_17045.t10 143.851
R19629 a_49314_17045.n1 a_49314_17045.t7 135.658
R19630 a_49314_17045.n0 a_49314_17045.t9 80.333
R19631 a_49314_17045.n4 a_49314_17045.t0 28.565
R19632 a_49314_17045.n4 a_49314_17045.t1 28.565
R19633 a_49314_17045.n2 a_49314_17045.t4 28.565
R19634 a_49314_17045.n2 a_49314_17045.t5 28.565
R19635 a_49314_17045.t2 a_49314_17045.n7 28.565
R19636 a_49314_17045.n7 a_49314_17045.t6 28.565
R19637 a_49314_17045.n5 a_49314_17045.t3 9.714
R19638 a_49314_17045.n5 a_49314_17045.n4 1.003
R19639 a_49314_17045.n6 a_49314_17045.n3 0.833
R19640 a_49314_17045.n3 a_49314_17045.n2 0.653
R19641 a_49314_17045.n7 a_49314_17045.n6 0.653
R19642 a_49314_17045.n6 a_49314_17045.n5 0.341
R19643 a_49314_17045.n3 a_49314_17045.n1 0.032
R19644 a_8056_15820.n2 a_8056_15820.t7 990.34
R19645 a_8056_15820.n3 a_8056_15820.n2 940.604
R19646 a_8056_15820.n2 a_8056_15820.t5 408.211
R19647 a_8056_15820.n1 a_8056_15820.t6 286.438
R19648 a_8056_15820.n1 a_8056_15820.t4 286.438
R19649 a_8056_15820.t7 a_8056_15820.n1 160.666
R19650 a_8056_15820.n3 a_8056_15820.n0 109.176
R19651 a_8056_15820.n4 a_8056_15820.n3 97.476
R19652 a_8056_15820.n0 a_8056_15820.t3 28.568
R19653 a_8056_15820.n4 a_8056_15820.t2 28.565
R19654 a_8056_15820.t1 a_8056_15820.n4 28.565
R19655 a_8056_15820.n0 a_8056_15820.t0 17.638
R19656 a_11289_6045.n1 a_11289_6045.t6 318.922
R19657 a_11289_6045.n0 a_11289_6045.t7 274.739
R19658 a_11289_6045.n0 a_11289_6045.t5 274.739
R19659 a_11289_6045.n1 a_11289_6045.t4 269.116
R19660 a_11289_6045.t6 a_11289_6045.n0 179.946
R19661 a_11289_6045.n2 a_11289_6045.n1 107.263
R19662 a_11289_6045.n3 a_11289_6045.t1 29.444
R19663 a_11289_6045.n4 a_11289_6045.t0 28.565
R19664 a_11289_6045.t2 a_11289_6045.n4 28.565
R19665 a_11289_6045.n2 a_11289_6045.t3 18.145
R19666 a_11289_6045.n3 a_11289_6045.n2 2.878
R19667 a_11289_6045.n4 a_11289_6045.n3 0.764
R19668 a_31377_6136.t0 a_31377_6136.t1 17.4
R19669 a_19454_10990.t1 a_19454_10990.n0 14.282
R19670 a_19454_10990.n0 a_19454_10990.t2 14.282
R19671 a_19454_10990.n0 a_19454_10990.n1 258.161
R19672 a_19454_10990.n1 a_19454_10990.t3 14.283
R19673 a_19454_10990.n1 a_19454_10990.n7 4.366
R19674 a_19454_10990.n7 a_19454_10990.n5 0.852
R19675 a_19454_10990.n5 a_19454_10990.n6 258.161
R19676 a_19454_10990.n6 a_19454_10990.t5 14.282
R19677 a_19454_10990.n6 a_19454_10990.t6 14.282
R19678 a_19454_10990.n5 a_19454_10990.t4 14.283
R19679 a_19454_10990.n7 a_19454_10990.n4 97.614
R19680 a_19454_10990.n4 a_19454_10990.t8 200.029
R19681 a_19454_10990.t8 a_19454_10990.n3 206.421
R19682 a_19454_10990.n3 a_19454_10990.t9 80.333
R19683 a_19454_10990.n3 a_19454_10990.t10 206.421
R19684 a_19454_10990.n4 a_19454_10990.t11 1527.4
R19685 a_19454_10990.t11 a_19454_10990.n2 657.379
R19686 a_19454_10990.n2 a_19454_10990.t0 8.7
R19687 a_19454_10990.n2 a_19454_10990.t7 8.7
R19688 a_19396_11720.n2 a_19396_11720.t7 990.34
R19689 a_19396_11720.n2 a_19396_11720.t4 408.211
R19690 a_19396_11720.n1 a_19396_11720.t5 286.438
R19691 a_19396_11720.n1 a_19396_11720.t6 286.438
R19692 a_19396_11720.n4 a_19396_11720.n0 185.55
R19693 a_19396_11720.t7 a_19396_11720.n1 160.666
R19694 a_19396_11720.n3 a_19396_11720.n2 70.974
R19695 a_19396_11720.t2 a_19396_11720.n4 28.568
R19696 a_19396_11720.n0 a_19396_11720.t0 28.565
R19697 a_19396_11720.n0 a_19396_11720.t1 28.565
R19698 a_19396_11720.n3 a_19396_11720.t3 21.882
R19699 a_19396_11720.n4 a_19396_11720.n3 1.625
R19700 a_11048_411.t0 a_11048_411.t1 17.4
R19701 a_16545_n2178.n1 a_16545_n2178.t5 990.34
R19702 a_16545_n2178.n1 a_16545_n2178.t7 408.211
R19703 a_16545_n2178.n0 a_16545_n2178.t4 286.438
R19704 a_16545_n2178.n0 a_16545_n2178.t6 286.438
R19705 a_16545_n2178.n4 a_16545_n2178.n3 185.55
R19706 a_16545_n2178.t5 a_16545_n2178.n0 160.666
R19707 a_16545_n2178.n2 a_16545_n2178.n1 46.239
R19708 a_16545_n2178.n3 a_16545_n2178.t1 28.568
R19709 a_16545_n2178.t2 a_16545_n2178.n4 28.565
R19710 a_16545_n2178.n4 a_16545_n2178.t0 28.565
R19711 a_16545_n2178.n2 a_16545_n2178.t3 21.376
R19712 a_16545_n2178.n3 a_16545_n2178.n2 1.637
R19713 a_23071_14428.n2 a_23071_14428.t6 867.497
R19714 a_23071_14428.n2 a_23071_14428.t7 591.811
R19715 a_23071_14428.n1 a_23071_14428.t5 286.438
R19716 a_23071_14428.n1 a_23071_14428.t4 286.438
R19717 a_23071_14428.n4 a_23071_14428.n0 192.754
R19718 a_23071_14428.t6 a_23071_14428.n1 160.666
R19719 a_23071_14428.t0 a_23071_14428.n4 28.568
R19720 a_23071_14428.n0 a_23071_14428.t2 28.565
R19721 a_23071_14428.n0 a_23071_14428.t1 28.565
R19722 a_23071_14428.n3 a_23071_14428.n2 20.232
R19723 a_23071_14428.n3 a_23071_14428.t3 18.713
R19724 a_23071_14428.n4 a_23071_14428.n3 1.312
R19725 a_22598_13724.t0 a_22598_13724.n0 14.283
R19726 a_22598_13724.n0 a_22598_13724.n7 258.161
R19727 a_22598_13724.n7 a_22598_13724.t6 14.282
R19728 a_22598_13724.n7 a_22598_13724.t7 14.282
R19729 a_22598_13724.n0 a_22598_13724.n6 4.366
R19730 a_22598_13724.n6 a_22598_13724.n4 0.852
R19731 a_22598_13724.n4 a_22598_13724.n5 258.161
R19732 a_22598_13724.n5 a_22598_13724.t3 14.282
R19733 a_22598_13724.n5 a_22598_13724.t5 14.282
R19734 a_22598_13724.n4 a_22598_13724.t4 14.283
R19735 a_22598_13724.n6 a_22598_13724.n3 97.614
R19736 a_22598_13724.n3 a_22598_13724.t9 200.029
R19737 a_22598_13724.t9 a_22598_13724.n2 206.421
R19738 a_22598_13724.n2 a_22598_13724.t10 80.333
R19739 a_22598_13724.n2 a_22598_13724.t11 206.421
R19740 a_22598_13724.n3 a_22598_13724.t8 1527.4
R19741 a_22598_13724.t8 a_22598_13724.n1 657.379
R19742 a_22598_13724.n1 a_22598_13724.t1 8.7
R19743 a_22598_13724.n1 a_22598_13724.t2 8.7
R19744 a_23131_14454.n0 a_23131_14454.t8 14.282
R19745 a_23131_14454.t0 a_23131_14454.n0 14.282
R19746 a_23131_14454.n0 a_23131_14454.n9 89.977
R19747 a_23131_14454.n6 a_23131_14454.n7 77.784
R19748 a_23131_14454.n4 a_23131_14454.n6 77.456
R19749 a_23131_14454.n9 a_23131_14454.n4 77.456
R19750 a_23131_14454.n9 a_23131_14454.n2 75.815
R19751 a_23131_14454.n7 a_23131_14454.n8 167.433
R19752 a_23131_14454.n8 a_23131_14454.t5 14.282
R19753 a_23131_14454.n8 a_23131_14454.t4 14.282
R19754 a_23131_14454.n7 a_23131_14454.t6 104.259
R19755 a_23131_14454.n6 a_23131_14454.n5 89.977
R19756 a_23131_14454.n5 a_23131_14454.t3 14.282
R19757 a_23131_14454.n5 a_23131_14454.t2 14.282
R19758 a_23131_14454.n4 a_23131_14454.n3 89.977
R19759 a_23131_14454.n3 a_23131_14454.t1 14.282
R19760 a_23131_14454.n3 a_23131_14454.t7 14.282
R19761 a_23131_14454.n2 a_23131_14454.t9 104.259
R19762 a_23131_14454.n2 a_23131_14454.n1 167.433
R19763 a_23131_14454.n1 a_23131_14454.t10 14.282
R19764 a_23131_14454.n1 a_23131_14454.t11 14.282
R19765 a_23198_1744.n0 a_23198_1744.t2 14.282
R19766 a_23198_1744.t1 a_23198_1744.n0 14.282
R19767 a_23198_1744.n0 a_23198_1744.n1 258.161
R19768 a_23198_1744.n1 a_23198_1744.t3 14.283
R19769 a_23198_1744.n1 a_23198_1744.n5 0.852
R19770 a_23198_1744.n5 a_23198_1744.n6 4.366
R19771 a_23198_1744.n6 a_23198_1744.n7 258.161
R19772 a_23198_1744.n7 a_23198_1744.t4 14.282
R19773 a_23198_1744.n7 a_23198_1744.t5 14.282
R19774 a_23198_1744.n6 a_23198_1744.t6 14.283
R19775 a_23198_1744.n5 a_23198_1744.n4 97.614
R19776 a_23198_1744.n4 a_23198_1744.t9 200.029
R19777 a_23198_1744.t9 a_23198_1744.n3 206.421
R19778 a_23198_1744.n3 a_23198_1744.t11 80.333
R19779 a_23198_1744.n3 a_23198_1744.t8 206.421
R19780 a_23198_1744.n4 a_23198_1744.t10 1527.4
R19781 a_23198_1744.t10 a_23198_1744.n2 657.379
R19782 a_23198_1744.n2 a_23198_1744.t0 8.7
R19783 a_23198_1744.n2 a_23198_1744.t7 8.7
R19784 a_22849_1744.n0 a_22849_1744.n9 167.433
R19785 a_22849_1744.t6 a_22849_1744.n0 14.282
R19786 a_22849_1744.n0 a_22849_1744.t7 14.282
R19787 a_22849_1744.n9 a_22849_1744.n8 75.815
R19788 a_22849_1744.n8 a_22849_1744.n6 77.456
R19789 a_22849_1744.n6 a_22849_1744.n4 77.456
R19790 a_22849_1744.n4 a_22849_1744.n2 77.784
R19791 a_22849_1744.n9 a_22849_1744.t8 104.259
R19792 a_22849_1744.n8 a_22849_1744.n7 89.977
R19793 a_22849_1744.n7 a_22849_1744.t11 14.282
R19794 a_22849_1744.n7 a_22849_1744.t9 14.282
R19795 a_22849_1744.n6 a_22849_1744.n5 89.977
R19796 a_22849_1744.n5 a_22849_1744.t10 14.282
R19797 a_22849_1744.n5 a_22849_1744.t1 14.282
R19798 a_22849_1744.n4 a_22849_1744.n3 89.977
R19799 a_22849_1744.n3 a_22849_1744.t2 14.282
R19800 a_22849_1744.n3 a_22849_1744.t0 14.282
R19801 a_22849_1744.n2 a_22849_1744.t4 104.259
R19802 a_22849_1744.n2 a_22849_1744.n1 167.433
R19803 a_22849_1744.n1 a_22849_1744.t3 14.282
R19804 a_22849_1744.n1 a_22849_1744.t5 14.282
R19805 a_7115_n2148.t9 a_7115_n2148.n0 14.282
R19806 a_7115_n2148.n0 a_7115_n2148.t10 14.282
R19807 a_7115_n2148.n0 a_7115_n2148.n9 89.977
R19808 a_7115_n2148.n9 a_7115_n2148.n7 75.815
R19809 a_7115_n2148.n9 a_7115_n2148.n6 77.456
R19810 a_7115_n2148.n6 a_7115_n2148.n4 77.456
R19811 a_7115_n2148.n4 a_7115_n2148.n2 77.784
R19812 a_7115_n2148.n7 a_7115_n2148.n8 167.433
R19813 a_7115_n2148.n8 a_7115_n2148.t8 14.282
R19814 a_7115_n2148.n8 a_7115_n2148.t7 14.282
R19815 a_7115_n2148.n7 a_7115_n2148.t6 104.259
R19816 a_7115_n2148.n6 a_7115_n2148.n5 89.977
R19817 a_7115_n2148.n5 a_7115_n2148.t11 14.282
R19818 a_7115_n2148.n5 a_7115_n2148.t5 14.282
R19819 a_7115_n2148.n4 a_7115_n2148.n3 89.977
R19820 a_7115_n2148.n3 a_7115_n2148.t4 14.282
R19821 a_7115_n2148.n3 a_7115_n2148.t3 14.282
R19822 a_7115_n2148.n2 a_7115_n2148.t2 104.259
R19823 a_7115_n2148.n2 a_7115_n2148.n1 167.433
R19824 a_7115_n2148.n1 a_7115_n2148.t1 14.282
R19825 a_7115_n2148.n1 a_7115_n2148.t0 14.282
R19826 a_9221_6047.n1 a_9221_6047.t4 318.922
R19827 a_9221_6047.n0 a_9221_6047.t5 274.739
R19828 a_9221_6047.n0 a_9221_6047.t7 274.739
R19829 a_9221_6047.n1 a_9221_6047.t6 269.116
R19830 a_9221_6047.t4 a_9221_6047.n0 179.946
R19831 a_9221_6047.n2 a_9221_6047.n1 107.263
R19832 a_9221_6047.t2 a_9221_6047.n4 29.444
R19833 a_9221_6047.n3 a_9221_6047.t1 28.565
R19834 a_9221_6047.n3 a_9221_6047.t0 28.565
R19835 a_9221_6047.n2 a_9221_6047.t3 18.145
R19836 a_9221_6047.n4 a_9221_6047.n2 2.878
R19837 a_9221_6047.n4 a_9221_6047.n3 0.764
R19838 a_1039_8966.t0 a_1039_8966.n0 14.282
R19839 a_1039_8966.n0 a_1039_8966.t1 14.282
R19840 a_1039_8966.n0 a_1039_8966.n8 122.747
R19841 a_1039_8966.n4 a_1039_8966.n6 74.302
R19842 a_1039_8966.n8 a_1039_8966.n4 50.575
R19843 a_1039_8966.n8 a_1039_8966.n7 157.665
R19844 a_1039_8966.n7 a_1039_8966.t7 8.7
R19845 a_1039_8966.n7 a_1039_8966.t3 8.7
R19846 a_1039_8966.n6 a_1039_8966.n5 90.436
R19847 a_1039_8966.n5 a_1039_8966.t6 14.282
R19848 a_1039_8966.n5 a_1039_8966.t4 14.282
R19849 a_1039_8966.n4 a_1039_8966.n3 90.416
R19850 a_1039_8966.n3 a_1039_8966.t5 14.282
R19851 a_1039_8966.n3 a_1039_8966.t2 14.282
R19852 a_1039_8966.n6 a_1039_8966.n1 2044.64
R19853 a_1039_8966.n1 a_1039_8966.t8 591.811
R19854 a_1039_8966.n1 a_1039_8966.t9 867.497
R19855 a_1039_8966.t9 a_1039_8966.n2 160.666
R19856 a_1039_8966.n2 a_1039_8966.t11 286.438
R19857 a_1039_8966.n2 a_1039_8966.t10 286.438
R19858 a_9761_5354.n0 a_9761_5354.t2 14.282
R19859 a_9761_5354.t0 a_9761_5354.n0 14.282
R19860 a_9761_5354.n0 a_9761_5354.n9 0.999
R19861 a_9761_5354.n6 a_9761_5354.n8 0.2
R19862 a_9761_5354.n9 a_9761_5354.n6 0.575
R19863 a_9761_5354.n9 a_9761_5354.t1 16.058
R19864 a_9761_5354.n8 a_9761_5354.n7 0.999
R19865 a_9761_5354.n7 a_9761_5354.t8 14.282
R19866 a_9761_5354.n7 a_9761_5354.t6 14.282
R19867 a_9761_5354.n8 a_9761_5354.t7 16.058
R19868 a_9761_5354.n6 a_9761_5354.n4 0.227
R19869 a_9761_5354.n4 a_9761_5354.n5 1.511
R19870 a_9761_5354.n5 a_9761_5354.t10 14.282
R19871 a_9761_5354.n5 a_9761_5354.t11 14.282
R19872 a_9761_5354.n4 a_9761_5354.n1 0.669
R19873 a_9761_5354.n1 a_9761_5354.n2 0.001
R19874 a_9761_5354.n1 a_9761_5354.n3 267.767
R19875 a_9761_5354.n3 a_9761_5354.t5 14.282
R19876 a_9761_5354.n3 a_9761_5354.t3 14.282
R19877 a_9761_5354.n2 a_9761_5354.t4 14.282
R19878 a_9761_5354.n2 a_9761_5354.t9 14.282
R19879 a_11133_n2633.n2 a_11133_n2633.t7 867.497
R19880 a_11133_n2633.n2 a_11133_n2633.t5 615.911
R19881 a_11133_n2633.n1 a_11133_n2633.t6 286.438
R19882 a_11133_n2633.n1 a_11133_n2633.t4 286.438
R19883 a_11133_n2633.n4 a_11133_n2633.n0 185.55
R19884 a_11133_n2633.t7 a_11133_n2633.n1 160.666
R19885 a_11133_n2633.t1 a_11133_n2633.n4 28.568
R19886 a_11133_n2633.n0 a_11133_n2633.t3 28.565
R19887 a_11133_n2633.n0 a_11133_n2633.t2 28.565
R19888 a_11133_n2633.n3 a_11133_n2633.n2 22.146
R19889 a_11133_n2633.n3 a_11133_n2633.t0 20.393
R19890 a_11133_n2633.n4 a_11133_n2633.n3 1.835
R19891 a_10259_n2148.n0 a_10259_n2148.n9 167.433
R19892 a_10259_n2148.n0 a_10259_n2148.t2 14.282
R19893 a_10259_n2148.t0 a_10259_n2148.n0 14.282
R19894 a_10259_n2148.n9 a_10259_n2148.n8 75.815
R19895 a_10259_n2148.n8 a_10259_n2148.n6 77.456
R19896 a_10259_n2148.n6 a_10259_n2148.n4 77.456
R19897 a_10259_n2148.n4 a_10259_n2148.n2 77.784
R19898 a_10259_n2148.n9 a_10259_n2148.t1 104.259
R19899 a_10259_n2148.n8 a_10259_n2148.n7 89.977
R19900 a_10259_n2148.n7 a_10259_n2148.t5 14.282
R19901 a_10259_n2148.n7 a_10259_n2148.t4 14.282
R19902 a_10259_n2148.n6 a_10259_n2148.n5 89.977
R19903 a_10259_n2148.n5 a_10259_n2148.t3 14.282
R19904 a_10259_n2148.n5 a_10259_n2148.t11 14.282
R19905 a_10259_n2148.n4 a_10259_n2148.n3 89.977
R19906 a_10259_n2148.n3 a_10259_n2148.t10 14.282
R19907 a_10259_n2148.n3 a_10259_n2148.t9 14.282
R19908 a_10259_n2148.n2 a_10259_n2148.t7 104.259
R19909 a_10259_n2148.n2 a_10259_n2148.n1 167.433
R19910 a_10259_n2148.n1 a_10259_n2148.t6 14.282
R19911 a_10259_n2148.n1 a_10259_n2148.t8 14.282
R19912 a_60766_15769.n0 a_60766_15769.t11 14.282
R19913 a_60766_15769.t9 a_60766_15769.n0 14.282
R19914 a_60766_15769.n0 a_60766_15769.n9 0.999
R19915 a_60766_15769.n9 a_60766_15769.n6 0.2
R19916 a_60766_15769.n6 a_60766_15769.n8 0.575
R19917 a_60766_15769.n8 a_60766_15769.t3 16.058
R19918 a_60766_15769.n8 a_60766_15769.n7 0.999
R19919 a_60766_15769.n7 a_60766_15769.t5 14.282
R19920 a_60766_15769.n7 a_60766_15769.t4 14.282
R19921 a_60766_15769.n9 a_60766_15769.t10 16.058
R19922 a_60766_15769.n6 a_60766_15769.n4 0.227
R19923 a_60766_15769.n4 a_60766_15769.n5 1.511
R19924 a_60766_15769.n5 a_60766_15769.t1 14.282
R19925 a_60766_15769.n5 a_60766_15769.t0 14.282
R19926 a_60766_15769.n4 a_60766_15769.n1 0.669
R19927 a_60766_15769.n1 a_60766_15769.n2 0.001
R19928 a_60766_15769.n1 a_60766_15769.n3 267.767
R19929 a_60766_15769.n3 a_60766_15769.t8 14.282
R19930 a_60766_15769.n3 a_60766_15769.t7 14.282
R19931 a_60766_15769.n2 a_60766_15769.t6 14.282
R19932 a_60766_15769.n2 a_60766_15769.t2 14.282
R19933 a_11947_4620.t0 a_11947_4620.t1 380.209
R19934 a_31375_1763.t0 a_31375_1763.t1 379.845
R19935 a_51337_3364.t0 a_51337_3364.t1 17.4
R19936 a_46233_22680.n2 a_46233_22680.t9 214.335
R19937 a_46233_22680.t7 a_46233_22680.n2 214.335
R19938 a_46233_22680.n3 a_46233_22680.t7 143.851
R19939 a_46233_22680.n3 a_46233_22680.t10 135.658
R19940 a_46233_22680.n2 a_46233_22680.t8 80.333
R19941 a_46233_22680.n4 a_46233_22680.t4 28.565
R19942 a_46233_22680.n4 a_46233_22680.t5 28.565
R19943 a_46233_22680.n0 a_46233_22680.t0 28.565
R19944 a_46233_22680.n0 a_46233_22680.t1 28.565
R19945 a_46233_22680.n7 a_46233_22680.t6 28.565
R19946 a_46233_22680.t2 a_46233_22680.n7 28.565
R19947 a_46233_22680.n1 a_46233_22680.t3 9.714
R19948 a_46233_22680.n1 a_46233_22680.n0 1.003
R19949 a_46233_22680.n6 a_46233_22680.n5 0.833
R19950 a_46233_22680.n5 a_46233_22680.n4 0.653
R19951 a_46233_22680.n7 a_46233_22680.n6 0.653
R19952 a_46233_22680.n6 a_46233_22680.n1 0.341
R19953 a_46233_22680.n5 a_46233_22680.n3 0.032
R19954 a_23316_20259.t0 a_23316_20259.t1 17.4
R19955 a_12808_16408.n0 a_12808_16408.t4 14.282
R19956 a_12808_16408.n0 a_12808_16408.t0 14.282
R19957 a_12808_16408.n1 a_12808_16408.t1 14.282
R19958 a_12808_16408.n1 a_12808_16408.t2 14.282
R19959 a_12808_16408.n3 a_12808_16408.t5 14.282
R19960 a_12808_16408.t3 a_12808_16408.n3 14.282
R19961 a_12808_16408.n3 a_12808_16408.n2 2.538
R19962 a_12808_16408.n2 a_12808_16408.n1 2.375
R19963 a_12808_16408.n2 a_12808_16408.n0 0.001
R19964 a_67370_10757.t0 a_67370_10757.t1 17.4
R19965 a_53304_6816.n1 a_53304_6816.t4 318.922
R19966 a_53304_6816.n0 a_53304_6816.t5 274.739
R19967 a_53304_6816.n0 a_53304_6816.t7 274.739
R19968 a_53304_6816.n1 a_53304_6816.t6 269.116
R19969 a_53304_6816.t4 a_53304_6816.n0 179.946
R19970 a_53304_6816.n2 a_53304_6816.n1 107.263
R19971 a_53304_6816.n3 a_53304_6816.t1 29.444
R19972 a_53304_6816.t2 a_53304_6816.n4 28.565
R19973 a_53304_6816.n4 a_53304_6816.t0 28.565
R19974 a_53304_6816.n2 a_53304_6816.t3 18.145
R19975 a_53304_6816.n3 a_53304_6816.n2 2.878
R19976 a_53304_6816.n4 a_53304_6816.n3 0.764
R19977 a_26279_20719.n2 a_26279_20719.t5 448.381
R19978 a_26279_20719.n1 a_26279_20719.t4 286.438
R19979 a_26279_20719.n1 a_26279_20719.t6 286.438
R19980 a_26279_20719.n0 a_26279_20719.t7 247.69
R19981 a_26279_20719.n4 a_26279_20719.n3 182.117
R19982 a_26279_20719.t5 a_26279_20719.n1 160.666
R19983 a_26279_20719.n3 a_26279_20719.t0 28.568
R19984 a_26279_20719.n4 a_26279_20719.t1 28.565
R19985 a_26279_20719.t2 a_26279_20719.n4 28.565
R19986 a_26279_20719.n0 a_26279_20719.t3 18.127
R19987 a_26279_20719.n2 a_26279_20719.n0 4.036
R19988 a_26279_20719.n3 a_26279_20719.n2 0.937
R19989 a_51699_310.t4 a_51699_310.t6 574.43
R19990 a_51699_310.n1 a_51699_310.t5 285.109
R19991 a_51699_310.n3 a_51699_310.n2 197.217
R19992 a_51699_310.n4 a_51699_310.n0 192.754
R19993 a_51699_310.n1 a_51699_310.t7 160.666
R19994 a_51699_310.n2 a_51699_310.t4 160.666
R19995 a_51699_310.n2 a_51699_310.n1 114.829
R19996 a_51699_310.t2 a_51699_310.n4 28.568
R19997 a_51699_310.n0 a_51699_310.t1 28.565
R19998 a_51699_310.n0 a_51699_310.t0 28.565
R19999 a_51699_310.n3 a_51699_310.t3 18.838
R20000 a_51699_310.n4 a_51699_310.n3 1.129
R20001 a_53307_3873.t7 a_53307_3873.n2 404.877
R20002 a_53307_3873.n1 a_53307_3873.t6 210.902
R20003 a_53307_3873.n3 a_53307_3873.t7 136.943
R20004 a_53307_3873.n2 a_53307_3873.n1 107.801
R20005 a_53307_3873.n1 a_53307_3873.t5 80.333
R20006 a_53307_3873.n2 a_53307_3873.t8 80.333
R20007 a_53307_3873.n0 a_53307_3873.t0 17.4
R20008 a_53307_3873.n0 a_53307_3873.t2 17.4
R20009 a_53307_3873.n4 a_53307_3873.t4 15.032
R20010 a_53307_3873.n5 a_53307_3873.t3 14.282
R20011 a_53307_3873.t1 a_53307_3873.n5 14.282
R20012 a_53307_3873.n5 a_53307_3873.n4 1.65
R20013 a_53307_3873.n3 a_53307_3873.n0 0.672
R20014 a_53307_3873.n4 a_53307_3873.n3 0.665
R20015 a_53425_3873.n1 a_53425_3873.t1 14.282
R20016 a_53425_3873.n1 a_53425_3873.t4 14.282
R20017 a_53425_3873.n0 a_53425_3873.t3 14.282
R20018 a_53425_3873.n0 a_53425_3873.t5 14.282
R20019 a_53425_3873.n3 a_53425_3873.t0 14.282
R20020 a_53425_3873.t2 a_53425_3873.n3 14.282
R20021 a_53425_3873.n2 a_53425_3873.n0 2.546
R20022 a_53425_3873.n3 a_53425_3873.n2 2.367
R20023 a_53425_3873.n2 a_53425_3873.n1 0.001
R20024 a_40101_3874.t8 a_40101_3874.n2 404.877
R20025 a_40101_3874.n1 a_40101_3874.t6 210.902
R20026 a_40101_3874.n3 a_40101_3874.t8 136.943
R20027 a_40101_3874.n2 a_40101_3874.n1 107.801
R20028 a_40101_3874.n1 a_40101_3874.t7 80.333
R20029 a_40101_3874.n2 a_40101_3874.t5 80.333
R20030 a_40101_3874.n0 a_40101_3874.t4 17.4
R20031 a_40101_3874.n0 a_40101_3874.t2 17.4
R20032 a_40101_3874.n4 a_40101_3874.t1 15.032
R20033 a_40101_3874.n5 a_40101_3874.t3 14.282
R20034 a_40101_3874.t0 a_40101_3874.n5 14.282
R20035 a_40101_3874.n5 a_40101_3874.n4 1.65
R20036 a_40101_3874.n3 a_40101_3874.n0 0.672
R20037 a_40101_3874.n4 a_40101_3874.n3 0.665
R20038 a_40365_3291.t5 a_40365_3291.t6 800.071
R20039 a_40365_3291.n3 a_40365_3291.n2 672.951
R20040 a_40365_3291.n1 a_40365_3291.t7 285.109
R20041 a_40365_3291.n2 a_40365_3291.t5 193.602
R20042 a_40365_3291.n1 a_40365_3291.t4 160.666
R20043 a_40365_3291.n2 a_40365_3291.n1 91.507
R20044 a_40365_3291.t2 a_40365_3291.n4 28.57
R20045 a_40365_3291.n0 a_40365_3291.t1 28.565
R20046 a_40365_3291.n0 a_40365_3291.t0 28.565
R20047 a_40365_3291.n4 a_40365_3291.t3 17.638
R20048 a_40365_3291.n3 a_40365_3291.n0 0.69
R20049 a_40365_3291.n4 a_40365_3291.n3 0.6
R20050 a_52465_7535.n2 a_52465_7535.t6 318.922
R20051 a_52465_7535.n1 a_52465_7535.t7 273.935
R20052 a_52465_7535.n1 a_52465_7535.t5 273.935
R20053 a_52465_7535.n2 a_52465_7535.t4 269.116
R20054 a_52465_7535.n4 a_52465_7535.n0 193.227
R20055 a_52465_7535.t6 a_52465_7535.n1 179.142
R20056 a_52465_7535.n3 a_52465_7535.n2 106.999
R20057 a_52465_7535.t2 a_52465_7535.n4 28.568
R20058 a_52465_7535.n0 a_52465_7535.t1 28.565
R20059 a_52465_7535.n0 a_52465_7535.t0 28.565
R20060 a_52465_7535.n3 a_52465_7535.t3 18.149
R20061 a_52465_7535.n4 a_52465_7535.n3 3.726
R20062 a_54358_1734.n1 a_54358_1734.t5 318.922
R20063 a_54358_1734.n0 a_54358_1734.t7 273.935
R20064 a_54358_1734.n0 a_54358_1734.t4 273.935
R20065 a_54358_1734.n1 a_54358_1734.t6 269.116
R20066 a_54358_1734.n4 a_54358_1734.n3 193.227
R20067 a_54358_1734.t5 a_54358_1734.n0 179.142
R20068 a_54358_1734.n2 a_54358_1734.n1 106.999
R20069 a_54358_1734.n3 a_54358_1734.t0 28.568
R20070 a_54358_1734.t2 a_54358_1734.n4 28.565
R20071 a_54358_1734.n4 a_54358_1734.t1 28.565
R20072 a_54358_1734.n2 a_54358_1734.t3 18.149
R20073 a_54358_1734.n3 a_54358_1734.n2 3.726
R20074 a_46219_24330.n0 a_46219_24330.t10 214.335
R20075 a_46219_24330.t8 a_46219_24330.n0 214.335
R20076 a_46219_24330.n1 a_46219_24330.t8 143.851
R20077 a_46219_24330.n1 a_46219_24330.t7 135.658
R20078 a_46219_24330.n0 a_46219_24330.t9 80.333
R20079 a_46219_24330.n2 a_46219_24330.t6 28.565
R20080 a_46219_24330.n2 a_46219_24330.t4 28.565
R20081 a_46219_24330.n4 a_46219_24330.t5 28.565
R20082 a_46219_24330.n4 a_46219_24330.t0 28.565
R20083 a_46219_24330.n7 a_46219_24330.t1 28.565
R20084 a_46219_24330.t2 a_46219_24330.n7 28.565
R20085 a_46219_24330.n6 a_46219_24330.t3 9.714
R20086 a_46219_24330.n7 a_46219_24330.n6 1.003
R20087 a_46219_24330.n5 a_46219_24330.n3 0.833
R20088 a_46219_24330.n3 a_46219_24330.n2 0.653
R20089 a_46219_24330.n5 a_46219_24330.n4 0.653
R20090 a_46219_24330.n6 a_46219_24330.n5 0.341
R20091 a_46219_24330.n3 a_46219_24330.n1 0.032
R20092 a_46809_23893.t6 a_46809_23893.t4 800.071
R20093 a_46809_23893.n2 a_46809_23893.n1 659.097
R20094 a_46809_23893.n0 a_46809_23893.t5 285.109
R20095 a_46809_23893.n1 a_46809_23893.t6 193.602
R20096 a_46809_23893.n4 a_46809_23893.n3 192.754
R20097 a_46809_23893.n0 a_46809_23893.t7 160.666
R20098 a_46809_23893.n1 a_46809_23893.n0 91.507
R20099 a_46809_23893.n3 a_46809_23893.t0 28.568
R20100 a_46809_23893.n4 a_46809_23893.t1 28.565
R20101 a_46809_23893.t2 a_46809_23893.n4 28.565
R20102 a_46809_23893.n2 a_46809_23893.t3 19.061
R20103 a_46809_23893.n3 a_46809_23893.n2 1.005
R20104 a_46356_6910.n0 a_46356_6910.n12 122.999
R20105 a_46356_6910.n0 a_46356_6910.t3 14.282
R20106 a_46356_6910.t1 a_46356_6910.n0 14.282
R20107 a_46356_6910.n12 a_46356_6910.n10 50.575
R20108 a_46356_6910.n10 a_46356_6910.n8 74.302
R20109 a_46356_6910.n12 a_46356_6910.n11 157.665
R20110 a_46356_6910.n11 a_46356_6910.t0 8.7
R20111 a_46356_6910.n11 a_46356_6910.t7 8.7
R20112 a_46356_6910.n10 a_46356_6910.n9 90.416
R20113 a_46356_6910.n9 a_46356_6910.t2 14.282
R20114 a_46356_6910.n9 a_46356_6910.t6 14.282
R20115 a_46356_6910.n8 a_46356_6910.n7 90.436
R20116 a_46356_6910.n7 a_46356_6910.t4 14.282
R20117 a_46356_6910.n7 a_46356_6910.t5 14.282
R20118 a_46356_6910.n8 a_46356_6910.n1 342.688
R20119 a_46356_6910.n1 a_46356_6910.n6 126.566
R20120 a_46356_6910.n6 a_46356_6910.t10 294.653
R20121 a_46356_6910.n6 a_46356_6910.t12 111.663
R20122 a_46356_6910.n1 a_46356_6910.n5 552.333
R20123 a_46356_6910.n5 a_46356_6910.n4 6.615
R20124 a_46356_6910.n4 a_46356_6910.t11 93.989
R20125 a_46356_6910.n5 a_46356_6910.n3 97.816
R20126 a_46356_6910.n3 a_46356_6910.t9 80.333
R20127 a_46356_6910.n3 a_46356_6910.t13 394.151
R20128 a_46356_6910.t13 a_46356_6910.n2 269.523
R20129 a_46356_6910.n2 a_46356_6910.t8 160.666
R20130 a_46356_6910.n2 a_46356_6910.t15 269.523
R20131 a_46356_6910.n4 a_46356_6910.t14 198.043
R20132 a_46238_6910.n3 a_46238_6910.n1 267.767
R20133 a_46238_6910.n7 a_46238_6910.t7 16.058
R20134 a_46238_6910.t2 a_46238_6910.n9 16.058
R20135 a_46238_6910.n2 a_46238_6910.t3 14.282
R20136 a_46238_6910.n2 a_46238_6910.t10 14.282
R20137 a_46238_6910.n1 a_46238_6910.t5 14.282
R20138 a_46238_6910.n1 a_46238_6910.t4 14.282
R20139 a_46238_6910.n4 a_46238_6910.t9 14.282
R20140 a_46238_6910.n4 a_46238_6910.t11 14.282
R20141 a_46238_6910.n0 a_46238_6910.t1 14.282
R20142 a_46238_6910.n0 a_46238_6910.t0 14.282
R20143 a_46238_6910.n6 a_46238_6910.t6 14.282
R20144 a_46238_6910.n6 a_46238_6910.t8 14.282
R20145 a_46238_6910.n5 a_46238_6910.n4 1.511
R20146 a_46238_6910.n9 a_46238_6910.n0 0.999
R20147 a_46238_6910.n7 a_46238_6910.n6 0.999
R20148 a_46238_6910.n5 a_46238_6910.n3 0.669
R20149 a_46238_6910.n9 a_46238_6910.n8 0.575
R20150 a_46238_6910.n8 a_46238_6910.n5 0.227
R20151 a_46238_6910.n8 a_46238_6910.n7 0.2
R20152 a_46238_6910.n3 a_46238_6910.n2 0.001
R20153 a_59322_18605.n0 a_59322_18605.t0 14.282
R20154 a_59322_18605.n0 a_59322_18605.t1 14.282
R20155 a_59322_18605.n1 a_59322_18605.t3 14.282
R20156 a_59322_18605.n1 a_59322_18605.t4 14.282
R20157 a_59322_18605.t2 a_59322_18605.n3 14.282
R20158 a_59322_18605.n3 a_59322_18605.t5 14.282
R20159 a_59322_18605.n2 a_59322_18605.n0 2.546
R20160 a_59322_18605.n2 a_59322_18605.n1 2.367
R20161 a_59322_18605.n3 a_59322_18605.n2 0.001
R20162 a_20290_411.t0 a_20290_411.t1 17.4
R20163 a_20003_20723.n2 a_20003_20723.t5 448.381
R20164 a_20003_20723.n1 a_20003_20723.t4 286.438
R20165 a_20003_20723.n1 a_20003_20723.t7 286.438
R20166 a_20003_20723.n0 a_20003_20723.t6 247.69
R20167 a_20003_20723.n4 a_20003_20723.n3 182.117
R20168 a_20003_20723.t5 a_20003_20723.n1 160.666
R20169 a_20003_20723.n3 a_20003_20723.t0 28.568
R20170 a_20003_20723.n4 a_20003_20723.t1 28.565
R20171 a_20003_20723.t2 a_20003_20723.n4 28.565
R20172 a_20003_20723.n0 a_20003_20723.t3 18.127
R20173 a_20003_20723.n2 a_20003_20723.n0 4.036
R20174 a_20003_20723.n3 a_20003_20723.n2 0.937
R20175 a_71846_4869.t0 a_71846_4869.t1 17.4
R20176 a_22709_16385.n0 a_22709_16385.t8 214.335
R20177 a_22709_16385.t10 a_22709_16385.n0 214.335
R20178 a_22709_16385.n1 a_22709_16385.t10 143.851
R20179 a_22709_16385.n1 a_22709_16385.t7 135.658
R20180 a_22709_16385.n0 a_22709_16385.t9 80.333
R20181 a_22709_16385.n2 a_22709_16385.t3 28.565
R20182 a_22709_16385.n2 a_22709_16385.t4 28.565
R20183 a_22709_16385.n4 a_22709_16385.t5 28.565
R20184 a_22709_16385.n4 a_22709_16385.t0 28.565
R20185 a_22709_16385.n7 a_22709_16385.t1 28.565
R20186 a_22709_16385.t2 a_22709_16385.n7 28.565
R20187 a_22709_16385.n3 a_22709_16385.t6 9.714
R20188 a_22709_16385.n3 a_22709_16385.n2 1.003
R20189 a_22709_16385.n6 a_22709_16385.n5 0.833
R20190 a_22709_16385.n5 a_22709_16385.n4 0.653
R20191 a_22709_16385.n7 a_22709_16385.n6 0.653
R20192 a_22709_16385.n5 a_22709_16385.n3 0.341
R20193 a_22709_16385.n6 a_22709_16385.n1 0.032
R20194 a_64185_771.n5 a_64185_771.n4 465.933
R20195 a_64185_771.t7 a_64185_771.t9 415.315
R20196 a_64185_771.n1 a_64185_771.t13 394.151
R20197 a_64185_771.n4 a_64185_771.t11 294.653
R20198 a_64185_771.n0 a_64185_771.t5 269.523
R20199 a_64185_771.t13 a_64185_771.n0 269.523
R20200 a_64185_771.n7 a_64185_771.t7 220.285
R20201 a_64185_771.n6 a_64185_771.t14 214.335
R20202 a_64185_771.t9 a_64185_771.n6 214.335
R20203 a_64185_771.n2 a_64185_771.t8 198.043
R20204 a_64185_771.n10 a_64185_771.n9 192.754
R20205 a_64185_771.n5 a_64185_771.n3 163.88
R20206 a_64185_771.n0 a_64185_771.t10 160.666
R20207 a_64185_771.n4 a_64185_771.t12 111.663
R20208 a_64185_771.n3 a_64185_771.n1 97.816
R20209 a_64185_771.n2 a_64185_771.t15 93.989
R20210 a_64185_771.n6 a_64185_771.t4 80.333
R20211 a_64185_771.n1 a_64185_771.t6 80.333
R20212 a_64185_771.n7 a_64185_771.n5 61.538
R20213 a_64185_771.n9 a_64185_771.t1 28.568
R20214 a_64185_771.n10 a_64185_771.t0 28.565
R20215 a_64185_771.t2 a_64185_771.n10 28.565
R20216 a_64185_771.n8 a_64185_771.t3 18.824
R20217 a_64185_771.n3 a_64185_771.n2 6.615
R20218 a_64185_771.n8 a_64185_771.n7 4.769
R20219 a_64185_771.n9 a_64185_771.n8 1.105
R20220 Y[4].n1 Y[4].n0 185.55
R20221 Y[4].n1 Y[4].t2 28.568
R20222 Y[4].n0 Y[4].t1 28.565
R20223 Y[4].n0 Y[4].t0 28.565
R20224 Y[4].n2 Y[4].t3 20.393
R20225 Y[4].n2 Y[4].n1 1.829
R20226 Y[4] Y[4].n2 1.121
R20227 a_65224_n537.n1 a_65224_n537.t5 318.922
R20228 a_65224_n537.n0 a_65224_n537.t4 273.935
R20229 a_65224_n537.n0 a_65224_n537.t6 273.935
R20230 a_65224_n537.n1 a_65224_n537.t7 269.116
R20231 a_65224_n537.n4 a_65224_n537.n3 193.227
R20232 a_65224_n537.t5 a_65224_n537.n0 179.142
R20233 a_65224_n537.n2 a_65224_n537.n1 106.999
R20234 a_65224_n537.n3 a_65224_n537.t0 28.568
R20235 a_65224_n537.n4 a_65224_n537.t1 28.565
R20236 a_65224_n537.t2 a_65224_n537.n4 28.565
R20237 a_65224_n537.n2 a_65224_n537.t3 18.149
R20238 a_65224_n537.n3 a_65224_n537.n2 3.726
R20239 a_58986_15769.n0 a_58986_15769.n8 90.436
R20240 a_58986_15769.n0 a_58986_15769.t7 14.282
R20241 a_58986_15769.t5 a_58986_15769.n0 14.282
R20242 a_58986_15769.n8 a_58986_15769.n5 74.302
R20243 a_58986_15769.n5 a_58986_15769.n7 50.575
R20244 a_58986_15769.n7 a_58986_15769.n6 157.665
R20245 a_58986_15769.n6 a_58986_15769.t0 8.7
R20246 a_58986_15769.n6 a_58986_15769.t4 8.7
R20247 a_58986_15769.n5 a_58986_15769.n4 90.416
R20248 a_58986_15769.n4 a_58986_15769.t6 14.282
R20249 a_58986_15769.n4 a_58986_15769.t3 14.282
R20250 a_58986_15769.n7 a_58986_15769.n3 122.746
R20251 a_58986_15769.n3 a_58986_15769.t2 14.282
R20252 a_58986_15769.n3 a_58986_15769.t1 14.282
R20253 a_58986_15769.n8 a_58986_15769.n1 260.998
R20254 a_58986_15769.t9 a_58986_15769.n2 160.666
R20255 a_58986_15769.n1 a_58986_15769.t9 867.393
R20256 a_58986_15769.n2 a_58986_15769.t8 287.241
R20257 a_58986_15769.n2 a_58986_15769.t10 287.241
R20258 a_58986_15769.n1 a_58986_15769.t11 545.094
R20259 a_58986_15037.t0 a_58986_15037.t1 380.209
R20260 a_57736_2352.n0 a_57736_2352.t9 214.335
R20261 a_57736_2352.t8 a_57736_2352.n0 214.335
R20262 a_57736_2352.n1 a_57736_2352.t8 143.851
R20263 a_57736_2352.n1 a_57736_2352.t7 135.658
R20264 a_57736_2352.n0 a_57736_2352.t10 80.333
R20265 a_57736_2352.n2 a_57736_2352.t5 28.565
R20266 a_57736_2352.n2 a_57736_2352.t4 28.565
R20267 a_57736_2352.n4 a_57736_2352.t6 28.565
R20268 a_57736_2352.n4 a_57736_2352.t2 28.565
R20269 a_57736_2352.n7 a_57736_2352.t1 28.565
R20270 a_57736_2352.t3 a_57736_2352.n7 28.565
R20271 a_57736_2352.n6 a_57736_2352.t0 9.714
R20272 a_57736_2352.n7 a_57736_2352.n6 1.003
R20273 a_57736_2352.n5 a_57736_2352.n3 0.833
R20274 a_57736_2352.n3 a_57736_2352.n2 0.653
R20275 a_57736_2352.n5 a_57736_2352.n4 0.653
R20276 a_57736_2352.n6 a_57736_2352.n5 0.341
R20277 a_57736_2352.n3 a_57736_2352.n1 0.032
R20278 a_58326_1915.t5 a_58326_1915.t7 574.43
R20279 a_58326_1915.n0 a_58326_1915.t6 285.109
R20280 a_58326_1915.n2 a_58326_1915.n1 211.136
R20281 a_58326_1915.n4 a_58326_1915.n3 192.754
R20282 a_58326_1915.n0 a_58326_1915.t4 160.666
R20283 a_58326_1915.n1 a_58326_1915.t5 160.666
R20284 a_58326_1915.n1 a_58326_1915.n0 114.829
R20285 a_58326_1915.n3 a_58326_1915.t1 28.568
R20286 a_58326_1915.n4 a_58326_1915.t0 28.565
R20287 a_58326_1915.t2 a_58326_1915.n4 28.565
R20288 a_58326_1915.n2 a_58326_1915.t3 19.084
R20289 a_58326_1915.n3 a_58326_1915.n2 1.051
R20290 a_18243_16385.n0 a_18243_16385.t7 214.335
R20291 a_18243_16385.t10 a_18243_16385.n0 214.335
R20292 a_18243_16385.n1 a_18243_16385.t10 143.851
R20293 a_18243_16385.n1 a_18243_16385.t9 135.658
R20294 a_18243_16385.n0 a_18243_16385.t8 80.333
R20295 a_18243_16385.n2 a_18243_16385.t4 28.565
R20296 a_18243_16385.n2 a_18243_16385.t5 28.565
R20297 a_18243_16385.n4 a_18243_16385.t3 28.565
R20298 a_18243_16385.n4 a_18243_16385.t0 28.565
R20299 a_18243_16385.n7 a_18243_16385.t1 28.565
R20300 a_18243_16385.t2 a_18243_16385.n7 28.565
R20301 a_18243_16385.n3 a_18243_16385.t6 9.714
R20302 a_18243_16385.n3 a_18243_16385.n2 1.003
R20303 a_18243_16385.n6 a_18243_16385.n5 0.833
R20304 a_18243_16385.n5 a_18243_16385.n4 0.653
R20305 a_18243_16385.n7 a_18243_16385.n6 0.653
R20306 a_18243_16385.n5 a_18243_16385.n3 0.341
R20307 a_18243_16385.n6 a_18243_16385.n1 0.032
R20308 a_45055_7783.t4 a_45055_7783.t5 574.43
R20309 a_45055_7783.n0 a_45055_7783.t7 285.109
R20310 a_45055_7783.n2 a_45055_7783.n1 211.136
R20311 a_45055_7783.n4 a_45055_7783.n3 192.754
R20312 a_45055_7783.n0 a_45055_7783.t6 160.666
R20313 a_45055_7783.n1 a_45055_7783.t4 160.666
R20314 a_45055_7783.n1 a_45055_7783.n0 114.829
R20315 a_45055_7783.n3 a_45055_7783.t2 28.568
R20316 a_45055_7783.t0 a_45055_7783.n4 28.565
R20317 a_45055_7783.n4 a_45055_7783.t1 28.565
R20318 a_45055_7783.n2 a_45055_7783.t3 19.084
R20319 a_45055_7783.n3 a_45055_7783.n2 1.051
R20320 a_47918_9746.n1 a_47918_9746.t4 14.282
R20321 a_47918_9746.n1 a_47918_9746.t0 14.282
R20322 a_47918_9746.n0 a_47918_9746.t1 14.282
R20323 a_47918_9746.n0 a_47918_9746.t2 14.282
R20324 a_47918_9746.n3 a_47918_9746.t5 14.282
R20325 a_47918_9746.t3 a_47918_9746.n3 14.282
R20326 a_47918_9746.n2 a_47918_9746.n0 2.546
R20327 a_47918_9746.n3 a_47918_9746.n2 2.367
R20328 a_47918_9746.n2 a_47918_9746.n1 0.001
R20329 a_31375_n2138.t0 a_31375_n2138.t1 17.4
R20330 a_46658_9742.t6 a_46658_9742.n2 404.877
R20331 a_46658_9742.n1 a_46658_9742.t8 210.902
R20332 a_46658_9742.n3 a_46658_9742.t6 136.943
R20333 a_46658_9742.n2 a_46658_9742.n1 107.801
R20334 a_46658_9742.n1 a_46658_9742.t5 80.333
R20335 a_46658_9742.n2 a_46658_9742.t7 80.333
R20336 a_46658_9742.n0 a_46658_9742.t4 17.4
R20337 a_46658_9742.n0 a_46658_9742.t3 17.4
R20338 a_46658_9742.n4 a_46658_9742.t2 15.032
R20339 a_46658_9742.t0 a_46658_9742.n5 14.282
R20340 a_46658_9742.n5 a_46658_9742.t1 14.282
R20341 a_46658_9742.n5 a_46658_9742.n4 1.65
R20342 a_46658_9742.n3 a_46658_9742.n0 0.672
R20343 a_46658_9742.n4 a_46658_9742.n3 0.665
R20344 a_46922_9159.t5 a_46922_9159.t4 800.071
R20345 a_46922_9159.n3 a_46922_9159.n2 672.951
R20346 a_46922_9159.n1 a_46922_9159.t6 285.109
R20347 a_46922_9159.n2 a_46922_9159.t5 193.602
R20348 a_46922_9159.n1 a_46922_9159.t7 160.666
R20349 a_46922_9159.n2 a_46922_9159.n1 91.507
R20350 a_46922_9159.n0 a_46922_9159.t1 28.57
R20351 a_46922_9159.n4 a_46922_9159.t0 28.565
R20352 a_46922_9159.t2 a_46922_9159.n4 28.565
R20353 a_46922_9159.n0 a_46922_9159.t3 17.638
R20354 a_46922_9159.n4 a_46922_9159.n3 0.69
R20355 a_46922_9159.n3 a_46922_9159.n0 0.6
R20356 a_59929_6884.n1 a_59929_6884.t6 318.922
R20357 a_59929_6884.n0 a_59929_6884.t7 274.739
R20358 a_59929_6884.n0 a_59929_6884.t5 274.739
R20359 a_59929_6884.n1 a_59929_6884.t4 269.116
R20360 a_59929_6884.t6 a_59929_6884.n0 179.946
R20361 a_59929_6884.n2 a_59929_6884.n1 107.263
R20362 a_59929_6884.n3 a_59929_6884.t0 29.444
R20363 a_59929_6884.t2 a_59929_6884.n4 28.565
R20364 a_59929_6884.n4 a_59929_6884.t1 28.565
R20365 a_59929_6884.n2 a_59929_6884.t3 18.145
R20366 a_59929_6884.n3 a_59929_6884.n2 2.878
R20367 a_59929_6884.n4 a_59929_6884.n3 0.764
R20368 a_59635_6178.t0 a_59635_6178.t1 380.209
R20369 a_46470_22043.t0 a_46470_22043.t1 17.4
R20370 a_49328_18695.n0 a_49328_18695.t8 214.335
R20371 a_49328_18695.t10 a_49328_18695.n0 214.335
R20372 a_49328_18695.n1 a_49328_18695.t10 143.851
R20373 a_49328_18695.n1 a_49328_18695.t7 135.658
R20374 a_49328_18695.n0 a_49328_18695.t9 80.333
R20375 a_49328_18695.n4 a_49328_18695.t0 28.565
R20376 a_49328_18695.n4 a_49328_18695.t1 28.565
R20377 a_49328_18695.n2 a_49328_18695.t4 28.565
R20378 a_49328_18695.n2 a_49328_18695.t5 28.565
R20379 a_49328_18695.t2 a_49328_18695.n7 28.565
R20380 a_49328_18695.n7 a_49328_18695.t6 28.565
R20381 a_49328_18695.n5 a_49328_18695.t3 9.714
R20382 a_49328_18695.n5 a_49328_18695.n4 1.003
R20383 a_49328_18695.n6 a_49328_18695.n3 0.833
R20384 a_49328_18695.n3 a_49328_18695.n2 0.653
R20385 a_49328_18695.n7 a_49328_18695.n6 0.653
R20386 a_49328_18695.n6 a_49328_18695.n5 0.341
R20387 a_49328_18695.n3 a_49328_18695.n1 0.032
R20388 a_63024_18092.t0 a_63024_18092.t1 17.4
R20389 a_17495_6045.n1 a_17495_6045.t4 318.922
R20390 a_17495_6045.n0 a_17495_6045.t7 274.739
R20391 a_17495_6045.n0 a_17495_6045.t5 274.739
R20392 a_17495_6045.n1 a_17495_6045.t6 269.116
R20393 a_17495_6045.t4 a_17495_6045.n0 179.946
R20394 a_17495_6045.n2 a_17495_6045.n1 107.263
R20395 a_17495_6045.t2 a_17495_6045.n4 29.444
R20396 a_17495_6045.n3 a_17495_6045.t1 28.565
R20397 a_17495_6045.n3 a_17495_6045.t0 28.565
R20398 a_17495_6045.n2 a_17495_6045.t3 18.145
R20399 a_17495_6045.n4 a_17495_6045.n2 2.878
R20400 a_17495_6045.n4 a_17495_6045.n3 0.764
R20401 a_9168_15798.t5 a_9168_15798.n3 406.053
R20402 a_9168_15798.n2 a_9168_15798.t7 188.134
R20403 a_9168_15798.n4 a_9168_15798.t5 136.949
R20404 a_9168_15798.n3 a_9168_15798.n2 107.801
R20405 a_9168_15798.n2 a_9168_15798.t8 80.333
R20406 a_9168_15798.n3 a_9168_15798.t6 80.333
R20407 a_9168_15798.n1 a_9168_15798.t0 17.4
R20408 a_9168_15798.n1 a_9168_15798.t4 17.4
R20409 a_9168_15798.t1 a_9168_15798.n5 15.036
R20410 a_9168_15798.n0 a_9168_15798.t2 14.282
R20411 a_9168_15798.n0 a_9168_15798.t3 14.282
R20412 a_9168_15798.n5 a_9168_15798.n0 1.654
R20413 a_9168_15798.n4 a_9168_15798.n1 0.657
R20414 a_9168_15798.n5 a_9168_15798.n4 0.614
R20415 a_9228_15824.n3 a_9228_15824.n1 1642.26
R20416 a_9228_15824.n1 a_9228_15824.t5 990.34
R20417 a_9228_15824.n1 a_9228_15824.t4 408.211
R20418 a_9228_15824.n0 a_9228_15824.t7 286.438
R20419 a_9228_15824.n0 a_9228_15824.t6 286.438
R20420 a_9228_15824.t5 a_9228_15824.n0 160.666
R20421 a_9228_15824.n3 a_9228_15824.n2 97.131
R20422 a_9228_15824.n4 a_9228_15824.n3 95.622
R20423 a_9228_15824.t2 a_9228_15824.n4 28.568
R20424 a_9228_15824.n2 a_9228_15824.t0 28.565
R20425 a_9228_15824.n2 a_9228_15824.t1 28.565
R20426 a_9228_15824.n4 a_9228_15824.t3 17.641
R20427 a_44465_8220.n4 a_44465_8220.t9 214.335
R20428 a_44465_8220.t8 a_44465_8220.n4 214.335
R20429 a_44465_8220.n5 a_44465_8220.t8 143.851
R20430 a_44465_8220.n5 a_44465_8220.t10 135.658
R20431 a_44465_8220.n4 a_44465_8220.t7 80.333
R20432 a_44465_8220.n0 a_44465_8220.t5 28.565
R20433 a_44465_8220.n0 a_44465_8220.t4 28.565
R20434 a_44465_8220.n2 a_44465_8220.t1 28.565
R20435 a_44465_8220.n2 a_44465_8220.t6 28.565
R20436 a_44465_8220.n7 a_44465_8220.t0 28.565
R20437 a_44465_8220.t2 a_44465_8220.n7 28.565
R20438 a_44465_8220.n1 a_44465_8220.t3 9.714
R20439 a_44465_8220.n1 a_44465_8220.n0 1.003
R20440 a_44465_8220.n6 a_44465_8220.n3 0.833
R20441 a_44465_8220.n3 a_44465_8220.n2 0.653
R20442 a_44465_8220.n7 a_44465_8220.n6 0.653
R20443 a_44465_8220.n3 a_44465_8220.n1 0.341
R20444 a_44465_8220.n6 a_44465_8220.n5 0.032
R20445 a_59517_6910.n0 a_59517_6910.t10 14.282
R20446 a_59517_6910.t9 a_59517_6910.n0 14.282
R20447 a_59517_6910.n0 a_59517_6910.n9 0.999
R20448 a_59517_6910.n9 a_59517_6910.n6 0.575
R20449 a_59517_6910.n6 a_59517_6910.n8 0.2
R20450 a_59517_6910.n8 a_59517_6910.t8 16.058
R20451 a_59517_6910.n8 a_59517_6910.n7 0.999
R20452 a_59517_6910.n7 a_59517_6910.t6 14.282
R20453 a_59517_6910.n7 a_59517_6910.t7 14.282
R20454 a_59517_6910.n9 a_59517_6910.t11 16.058
R20455 a_59517_6910.n6 a_59517_6910.n4 0.227
R20456 a_59517_6910.n4 a_59517_6910.n5 1.511
R20457 a_59517_6910.n5 a_59517_6910.t2 14.282
R20458 a_59517_6910.n5 a_59517_6910.t0 14.282
R20459 a_59517_6910.n4 a_59517_6910.n1 0.669
R20460 a_59517_6910.n1 a_59517_6910.n2 0.001
R20461 a_59517_6910.n1 a_59517_6910.n3 267.767
R20462 a_59517_6910.n3 a_59517_6910.t4 14.282
R20463 a_59517_6910.n3 a_59517_6910.t5 14.282
R20464 a_59517_6910.n2 a_59517_6910.t1 14.282
R20465 a_59517_6910.n2 a_59517_6910.t3 14.282
R20466 a_70455_11391.n2 a_70455_11391.t5 448.381
R20467 a_70455_11391.n1 a_70455_11391.t7 287.241
R20468 a_70455_11391.n1 a_70455_11391.t6 287.241
R20469 a_70455_11391.n0 a_70455_11391.t4 247.733
R20470 a_70455_11391.n4 a_70455_11391.n3 182.117
R20471 a_70455_11391.t5 a_70455_11391.n1 160.666
R20472 a_70455_11391.n3 a_70455_11391.t0 28.568
R20473 a_70455_11391.n4 a_70455_11391.t1 28.565
R20474 a_70455_11391.t2 a_70455_11391.n4 28.565
R20475 a_70455_11391.n0 a_70455_11391.t3 18.127
R20476 a_70455_11391.n2 a_70455_11391.n0 4.036
R20477 a_70455_11391.n3 a_70455_11391.n2 0.937
R20478 a_40621_16458.n1 a_40621_16458.t6 318.922
R20479 a_40621_16458.n0 a_40621_16458.t5 274.739
R20480 a_40621_16458.n0 a_40621_16458.t7 274.739
R20481 a_40621_16458.n1 a_40621_16458.t4 269.116
R20482 a_40621_16458.t6 a_40621_16458.n0 179.946
R20483 a_40621_16458.n2 a_40621_16458.n1 107.263
R20484 a_40621_16458.t2 a_40621_16458.n4 29.444
R20485 a_40621_16458.n3 a_40621_16458.t0 28.565
R20486 a_40621_16458.n3 a_40621_16458.t1 28.565
R20487 a_40621_16458.n2 a_40621_16458.t3 18.145
R20488 a_40621_16458.n4 a_40621_16458.n2 2.878
R20489 a_40621_16458.n4 a_40621_16458.n3 0.764
R20490 a_70513_16782.n2 a_70513_16782.t10 1551.5
R20491 a_70513_16782.t10 a_70513_16782.n0 656.576
R20492 a_70513_16782.n4 a_70513_16782.n3 258.161
R20493 a_70513_16782.n7 a_70513_16782.n6 258.161
R20494 a_70513_16782.n2 a_70513_16782.t11 224.129
R20495 a_70513_16782.n1 a_70513_16782.t9 207.225
R20496 a_70513_16782.t11 a_70513_16782.n1 207.225
R20497 a_70513_16782.n1 a_70513_16782.t8 80.333
R20498 a_70513_16782.n5 a_70513_16782.n2 73.514
R20499 a_70513_16782.n4 a_70513_16782.t4 14.283
R20500 a_70513_16782.n6 a_70513_16782.t1 14.283
R20501 a_70513_16782.n3 a_70513_16782.t5 14.282
R20502 a_70513_16782.n3 a_70513_16782.t3 14.282
R20503 a_70513_16782.t2 a_70513_16782.n7 14.282
R20504 a_70513_16782.n7 a_70513_16782.t0 14.282
R20505 a_70513_16782.n0 a_70513_16782.t7 8.7
R20506 a_70513_16782.n0 a_70513_16782.t6 8.7
R20507 a_70513_16782.n5 a_70513_16782.n4 4.366
R20508 a_70513_16782.n6 a_70513_16782.n5 0.852
R20509 a_20579_1259.n1 a_20579_1259.t6 867.497
R20510 a_20579_1259.n1 a_20579_1259.t7 615.911
R20511 a_20579_1259.n0 a_20579_1259.t5 286.438
R20512 a_20579_1259.n0 a_20579_1259.t4 286.438
R20513 a_20579_1259.n4 a_20579_1259.n3 185.55
R20514 a_20579_1259.t6 a_20579_1259.n0 160.666
R20515 a_20579_1259.n2 a_20579_1259.n1 130.973
R20516 a_20579_1259.n3 a_20579_1259.t0 28.568
R20517 a_20579_1259.n4 a_20579_1259.t1 28.565
R20518 a_20579_1259.t2 a_20579_1259.n4 28.565
R20519 a_20579_1259.n2 a_20579_1259.t3 20.393
R20520 a_20579_1259.n3 a_20579_1259.n2 1.835
R20521 a_44454_746.n4 a_44454_746.t7 214.335
R20522 a_44454_746.t10 a_44454_746.n4 214.335
R20523 a_44454_746.n5 a_44454_746.t10 143.851
R20524 a_44454_746.n5 a_44454_746.t9 135.658
R20525 a_44454_746.n4 a_44454_746.t8 80.333
R20526 a_44454_746.n0 a_44454_746.t3 28.565
R20527 a_44454_746.n0 a_44454_746.t4 28.565
R20528 a_44454_746.n2 a_44454_746.t1 28.565
R20529 a_44454_746.n2 a_44454_746.t5 28.565
R20530 a_44454_746.n7 a_44454_746.t0 28.565
R20531 a_44454_746.t2 a_44454_746.n7 28.565
R20532 a_44454_746.n1 a_44454_746.t6 9.714
R20533 a_44454_746.n1 a_44454_746.n0 1.003
R20534 a_44454_746.n6 a_44454_746.n3 0.833
R20535 a_44454_746.n3 a_44454_746.n2 0.653
R20536 a_44454_746.n7 a_44454_746.n6 0.653
R20537 a_44454_746.n3 a_44454_746.n1 0.341
R20538 a_44454_746.n6 a_44454_746.n5 0.032
R20539 a_1735_10851.n2 a_1735_10851.t6 448.381
R20540 a_1735_10851.n1 a_1735_10851.t5 286.438
R20541 a_1735_10851.n1 a_1735_10851.t4 286.438
R20542 a_1735_10851.n0 a_1735_10851.t7 247.69
R20543 a_1735_10851.n4 a_1735_10851.n3 182.117
R20544 a_1735_10851.t6 a_1735_10851.n1 160.666
R20545 a_1735_10851.n3 a_1735_10851.t0 28.568
R20546 a_1735_10851.n4 a_1735_10851.t1 28.565
R20547 a_1735_10851.t2 a_1735_10851.n4 28.565
R20548 a_1735_10851.n0 a_1735_10851.t3 18.127
R20549 a_1735_10851.n2 a_1735_10851.n0 4.036
R20550 a_1735_10851.n3 a_1735_10851.n2 0.937
R20551 a_13120_11724.n2 a_13120_11724.t4 990.34
R20552 a_13120_11724.n2 a_13120_11724.t7 408.211
R20553 a_13120_11724.n3 a_13120_11724.n2 295.742
R20554 a_13120_11724.n1 a_13120_11724.t5 286.438
R20555 a_13120_11724.n1 a_13120_11724.t6 286.438
R20556 a_13120_11724.n4 a_13120_11724.n0 185.55
R20557 a_13120_11724.t4 a_13120_11724.n1 160.666
R20558 a_13120_11724.t0 a_13120_11724.n4 28.568
R20559 a_13120_11724.n0 a_13120_11724.t3 28.565
R20560 a_13120_11724.n0 a_13120_11724.t1 28.565
R20561 a_13120_11724.n3 a_13120_11724.t2 21.376
R20562 a_13120_11724.n4 a_13120_11724.n3 1.637
R20563 a_59548_23692.t0 a_59548_23692.t1 17.4
R20564 a_37856_8106.n15 a_37856_8106.n14 3522.62
R20565 a_37856_8106.n6 a_37856_8106.n5 501.28
R20566 a_37856_8106.t10 a_37856_8106.t6 437.233
R20567 a_37856_8106.t9 a_37856_8106.t16 415.315
R20568 a_37856_8106.t18 a_37856_8106.n3 313.873
R20569 a_37856_8106.n5 a_37856_8106.t17 294.986
R20570 a_37856_8106.n2 a_37856_8106.t8 272.288
R20571 a_37856_8106.n6 a_37856_8106.t14 236.01
R20572 a_37856_8106.n9 a_37856_8106.t10 216.627
R20573 a_37856_8106.n7 a_37856_8106.t9 216.111
R20574 a_37856_8106.n8 a_37856_8106.t13 214.686
R20575 a_37856_8106.t6 a_37856_8106.n8 214.686
R20576 a_37856_8106.n1 a_37856_8106.t4 214.335
R20577 a_37856_8106.t16 a_37856_8106.n1 214.335
R20578 a_37856_8106.n17 a_37856_8106.n16 192.754
R20579 a_37856_8106.n4 a_37856_8106.t18 190.152
R20580 a_37856_8106.n4 a_37856_8106.t7 190.152
R20581 a_37856_8106.n2 a_37856_8106.t19 160.666
R20582 a_37856_8106.n3 a_37856_8106.t15 160.666
R20583 a_37856_8106.n7 a_37856_8106.n6 148.428
R20584 a_37856_8106.n5 a_37856_8106.t11 110.859
R20585 a_37856_8106.n3 a_37856_8106.n2 96.129
R20586 a_37856_8106.n8 a_37856_8106.t5 80.333
R20587 a_37856_8106.n1 a_37856_8106.t12 80.333
R20588 a_37856_8106.t14 a_37856_8106.n4 80.333
R20589 a_37856_8106.n16 a_37856_8106.t1 28.568
R20590 a_37856_8106.n17 a_37856_8106.t0 28.565
R20591 a_37856_8106.t2 a_37856_8106.n17 28.565
R20592 a_37856_8106.n15 a_37856_8106.t3 18.522
R20593 a_37856_8106.n14 a_37856_8106.n13 5.25
R20594 a_37856_8106.n13 a_37856_8106.n12 3.293
R20595 a_37856_8106.n9 a_37856_8106.n7 2.923
R20596 a_37856_8106.n16 a_37856_8106.n15 1.168
R20597 a_37856_8106.n10 a_37856_8106.n9 0.708
R20598 a_37856_8106.n13 a_37856_8106.n11 0.681
R20599 a_37856_8106.n11 a_37856_8106.n0 0.003
R20600 a_37856_8106.n11 a_37856_8106.n10 0.001
R20601 a_37911_6528.n0 a_37911_6528.t10 214.335
R20602 a_37911_6528.t9 a_37911_6528.n0 214.335
R20603 a_37911_6528.n1 a_37911_6528.t9 143.851
R20604 a_37911_6528.n1 a_37911_6528.t8 135.658
R20605 a_37911_6528.n0 a_37911_6528.t7 80.333
R20606 a_37911_6528.n2 a_37911_6528.t6 28.565
R20607 a_37911_6528.n2 a_37911_6528.t5 28.565
R20608 a_37911_6528.n4 a_37911_6528.t4 28.565
R20609 a_37911_6528.n4 a_37911_6528.t1 28.565
R20610 a_37911_6528.t2 a_37911_6528.n7 28.565
R20611 a_37911_6528.n7 a_37911_6528.t0 28.565
R20612 a_37911_6528.n6 a_37911_6528.t3 9.714
R20613 a_37911_6528.n7 a_37911_6528.n6 1.003
R20614 a_37911_6528.n5 a_37911_6528.n3 0.833
R20615 a_37911_6528.n3 a_37911_6528.n2 0.653
R20616 a_37911_6528.n5 a_37911_6528.n4 0.653
R20617 a_37911_6528.n6 a_37911_6528.n5 0.341
R20618 a_37911_6528.n3 a_37911_6528.n1 0.032
R20619 a_41676_11949.n0 a_41676_11949.t10 214.335
R20620 a_41676_11949.t8 a_41676_11949.n0 214.335
R20621 a_41676_11949.n1 a_41676_11949.t8 143.851
R20622 a_41676_11949.n1 a_41676_11949.t7 135.658
R20623 a_41676_11949.n0 a_41676_11949.t9 80.333
R20624 a_41676_11949.n2 a_41676_11949.t5 28.565
R20625 a_41676_11949.n2 a_41676_11949.t6 28.565
R20626 a_41676_11949.n4 a_41676_11949.t4 28.565
R20627 a_41676_11949.n4 a_41676_11949.t1 28.565
R20628 a_41676_11949.n7 a_41676_11949.t2 28.565
R20629 a_41676_11949.t3 a_41676_11949.n7 28.565
R20630 a_41676_11949.n6 a_41676_11949.t0 9.714
R20631 a_41676_11949.n7 a_41676_11949.n6 1.003
R20632 a_41676_11949.n5 a_41676_11949.n3 0.833
R20633 a_41676_11949.n3 a_41676_11949.n2 0.653
R20634 a_41676_11949.n5 a_41676_11949.n4 0.653
R20635 a_41676_11949.n6 a_41676_11949.n5 0.341
R20636 a_41676_11949.n3 a_41676_11949.n1 0.032
R20637 a_4593_6357.n2 a_4593_6357.t6 990.34
R20638 a_4593_6357.n2 a_4593_6357.t5 408.211
R20639 a_4593_6357.n1 a_4593_6357.t7 286.438
R20640 a_4593_6357.n1 a_4593_6357.t4 286.438
R20641 a_4593_6357.n4 a_4593_6357.n0 197.272
R20642 a_4593_6357.t6 a_4593_6357.n1 160.666
R20643 a_4593_6357.t2 a_4593_6357.n4 28.568
R20644 a_4593_6357.n0 a_4593_6357.t1 28.565
R20645 a_4593_6357.n0 a_4593_6357.t0 28.565
R20646 a_4593_6357.n3 a_4593_6357.n2 19.535
R20647 a_4593_6357.n3 a_4593_6357.t3 18.103
R20648 a_4593_6357.n4 a_4593_6357.n3 0.459
R20649 a_30152_475.n2 a_30152_475.t4 318.119
R20650 a_30152_475.n2 a_30152_475.t7 269.919
R20651 a_30152_475.n1 a_30152_475.t6 267.256
R20652 a_30152_475.n1 a_30152_475.t5 267.256
R20653 a_30152_475.n4 a_30152_475.n0 193.227
R20654 a_30152_475.t4 a_30152_475.n1 160.666
R20655 a_30152_475.n3 a_30152_475.n2 106.999
R20656 a_30152_475.t2 a_30152_475.n4 28.568
R20657 a_30152_475.n0 a_30152_475.t0 28.565
R20658 a_30152_475.n0 a_30152_475.t1 28.565
R20659 a_30152_475.n3 a_30152_475.t3 18.149
R20660 a_30152_475.n4 a_30152_475.n3 3.726
R20661 a_13898_5354.n0 a_13898_5354.t11 14.282
R20662 a_13898_5354.t6 a_13898_5354.n0 14.282
R20663 a_13898_5354.n0 a_13898_5354.n9 0.999
R20664 a_13898_5354.n9 a_13898_5354.n6 0.2
R20665 a_13898_5354.n6 a_13898_5354.n8 0.575
R20666 a_13898_5354.n8 a_13898_5354.t8 16.058
R20667 a_13898_5354.n8 a_13898_5354.n7 0.999
R20668 a_13898_5354.n7 a_13898_5354.t9 14.282
R20669 a_13898_5354.n7 a_13898_5354.t7 14.282
R20670 a_13898_5354.n9 a_13898_5354.t10 16.058
R20671 a_13898_5354.n6 a_13898_5354.n4 0.227
R20672 a_13898_5354.n4 a_13898_5354.n5 1.511
R20673 a_13898_5354.n5 a_13898_5354.t5 14.282
R20674 a_13898_5354.n5 a_13898_5354.t3 14.282
R20675 a_13898_5354.n4 a_13898_5354.n1 0.669
R20676 a_13898_5354.n1 a_13898_5354.n2 0.001
R20677 a_13898_5354.n1 a_13898_5354.n3 267.767
R20678 a_13898_5354.n3 a_13898_5354.t0 14.282
R20679 a_13898_5354.n3 a_13898_5354.t1 14.282
R20680 a_13898_5354.n2 a_13898_5354.t2 14.282
R20681 a_13898_5354.n2 a_13898_5354.t4 14.282
R20682 a_30152_9379.n1 a_30152_9379.t5 318.119
R20683 a_30152_9379.n1 a_30152_9379.t6 269.919
R20684 a_30152_9379.n0 a_30152_9379.t7 267.853
R20685 a_30152_9379.n0 a_30152_9379.t4 267.853
R20686 a_30152_9379.t5 a_30152_9379.n0 160.666
R20687 a_30152_9379.n2 a_30152_9379.n1 107.263
R20688 a_30152_9379.n3 a_30152_9379.t1 29.444
R20689 a_30152_9379.t2 a_30152_9379.n4 28.565
R20690 a_30152_9379.n4 a_30152_9379.t0 28.565
R20691 a_30152_9379.n2 a_30152_9379.t3 18.145
R20692 a_30152_9379.n3 a_30152_9379.n2 2.878
R20693 a_30152_9379.n4 a_30152_9379.n3 0.764
R20694 a_58334_7783.t4 a_58334_7783.t6 574.43
R20695 a_58334_7783.n0 a_58334_7783.t5 285.109
R20696 a_58334_7783.n2 a_58334_7783.n1 211.136
R20697 a_58334_7783.n4 a_58334_7783.n3 192.754
R20698 a_58334_7783.n0 a_58334_7783.t7 160.666
R20699 a_58334_7783.n1 a_58334_7783.t4 160.666
R20700 a_58334_7783.n1 a_58334_7783.n0 114.829
R20701 a_58334_7783.n3 a_58334_7783.t1 28.568
R20702 a_58334_7783.t2 a_58334_7783.n4 28.565
R20703 a_58334_7783.n4 a_58334_7783.t0 28.565
R20704 a_58334_7783.n2 a_58334_7783.t3 19.084
R20705 a_58334_7783.n3 a_58334_7783.n2 1.051
R20706 a_21632_6045.n1 a_21632_6045.t7 318.922
R20707 a_21632_6045.n0 a_21632_6045.t5 274.739
R20708 a_21632_6045.n0 a_21632_6045.t6 274.739
R20709 a_21632_6045.n1 a_21632_6045.t4 269.116
R20710 a_21632_6045.t7 a_21632_6045.n0 179.946
R20711 a_21632_6045.n2 a_21632_6045.n1 107.263
R20712 a_21632_6045.n3 a_21632_6045.t0 29.444
R20713 a_21632_6045.n4 a_21632_6045.t1 28.565
R20714 a_21632_6045.t2 a_21632_6045.n4 28.565
R20715 a_21632_6045.n2 a_21632_6045.t3 18.145
R20716 a_21632_6045.n3 a_21632_6045.n2 2.878
R20717 a_21632_6045.n4 a_21632_6045.n3 0.764
R20718 a_59863_310.t0 a_59863_310.t1 17.4
R20719 a_7995_15753.t5 a_7995_15753.n2 403.87
R20720 a_7995_15753.n1 a_7995_15753.t6 191.682
R20721 a_7995_15753.n3 a_7995_15753.t5 138.556
R20722 a_7995_15753.n2 a_7995_15753.n1 111.349
R20723 a_7995_15753.n1 a_7995_15753.t7 80.333
R20724 a_7995_15753.n2 a_7995_15753.t8 80.333
R20725 a_7995_15753.n0 a_7995_15753.t2 17.4
R20726 a_7995_15753.n0 a_7995_15753.t0 17.4
R20727 a_7995_15753.n4 a_7995_15753.t3 15.036
R20728 a_7995_15753.t1 a_7995_15753.n5 14.282
R20729 a_7995_15753.n5 a_7995_15753.t4 14.282
R20730 a_7995_15753.n5 a_7995_15753.n4 1.654
R20731 a_7995_15753.n3 a_7995_15753.n0 0.664
R20732 a_7995_15753.n4 a_7995_15753.n3 0.614
R20733 a_53571_3290.t4 a_53571_3290.t5 800.071
R20734 a_53571_3290.n3 a_53571_3290.n2 672.951
R20735 a_53571_3290.n1 a_53571_3290.t7 285.109
R20736 a_53571_3290.n2 a_53571_3290.t4 193.602
R20737 a_53571_3290.n1 a_53571_3290.t6 160.666
R20738 a_53571_3290.n2 a_53571_3290.n1 91.507
R20739 a_53571_3290.n0 a_53571_3290.t0 28.57
R20740 a_53571_3290.n4 a_53571_3290.t1 28.565
R20741 a_53571_3290.t2 a_53571_3290.n4 28.565
R20742 a_53571_3290.n0 a_53571_3290.t3 17.638
R20743 a_53571_3290.n4 a_53571_3290.n3 0.69
R20744 a_53571_3290.n3 a_53571_3290.n0 0.6
R20745 a_46823_22243.t5 a_46823_22243.t4 574.43
R20746 a_46823_22243.n0 a_46823_22243.t7 285.109
R20747 a_46823_22243.n2 a_46823_22243.n1 211.136
R20748 a_46823_22243.n4 a_46823_22243.n3 192.754
R20749 a_46823_22243.n0 a_46823_22243.t6 160.666
R20750 a_46823_22243.n1 a_46823_22243.t5 160.666
R20751 a_46823_22243.n1 a_46823_22243.n0 114.829
R20752 a_46823_22243.n3 a_46823_22243.t0 28.568
R20753 a_46823_22243.n4 a_46823_22243.t1 28.565
R20754 a_46823_22243.t2 a_46823_22243.n4 28.565
R20755 a_46823_22243.n2 a_46823_22243.t3 19.084
R20756 a_46823_22243.n3 a_46823_22243.n2 1.051
R20757 a_49568_24206.t5 a_49568_24206.n3 404.877
R20758 a_49568_24206.n2 a_49568_24206.t8 210.902
R20759 a_49568_24206.n4 a_49568_24206.t5 136.943
R20760 a_49568_24206.n3 a_49568_24206.n2 107.801
R20761 a_49568_24206.n2 a_49568_24206.t7 80.333
R20762 a_49568_24206.n3 a_49568_24206.t6 80.333
R20763 a_49568_24206.n1 a_49568_24206.t4 17.4
R20764 a_49568_24206.n1 a_49568_24206.t3 17.4
R20765 a_49568_24206.t2 a_49568_24206.n5 15.032
R20766 a_49568_24206.n0 a_49568_24206.t0 14.282
R20767 a_49568_24206.n0 a_49568_24206.t1 14.282
R20768 a_49568_24206.n5 a_49568_24206.n0 1.65
R20769 a_49568_24206.n4 a_49568_24206.n1 0.672
R20770 a_49568_24206.n5 a_49568_24206.n4 0.665
R20771 a_16378_5326.n1 a_16378_5326.t4 318.922
R20772 a_16378_5326.n0 a_16378_5326.t5 273.935
R20773 a_16378_5326.n0 a_16378_5326.t6 273.935
R20774 a_16378_5326.n1 a_16378_5326.t7 269.116
R20775 a_16378_5326.n4 a_16378_5326.n3 193.227
R20776 a_16378_5326.t4 a_16378_5326.n0 179.142
R20777 a_16378_5326.n2 a_16378_5326.n1 106.999
R20778 a_16378_5326.n3 a_16378_5326.t1 28.568
R20779 a_16378_5326.t2 a_16378_5326.n4 28.565
R20780 a_16378_5326.n4 a_16378_5326.t0 28.565
R20781 a_16378_5326.n2 a_16378_5326.t3 18.149
R20782 a_16378_5326.n3 a_16378_5326.n2 3.726
R20783 a_46456_23693.t0 a_46456_23693.t1 17.4
R20784 a_10115_4622.t0 a_10115_4622.t1 17.4
R20785 a_55139_309.t0 a_55139_309.t1 17.4
R20786 a_53010_6110.t0 a_53010_6110.t1 380.209
R20787 a_41369_9658.n1 a_41369_9658.t2 14.282
R20788 a_41369_9658.n1 a_41369_9658.t5 14.282
R20789 a_41369_9658.n0 a_41369_9658.t4 14.282
R20790 a_41369_9658.n0 a_41369_9658.t3 14.282
R20791 a_41369_9658.t0 a_41369_9658.n3 14.282
R20792 a_41369_9658.n3 a_41369_9658.t1 14.282
R20793 a_41369_9658.n2 a_41369_9658.n0 2.546
R20794 a_41369_9658.n3 a_41369_9658.n2 2.367
R20795 a_41369_9658.n2 a_41369_9658.n1 0.001
R20796 a_22550_8988.n1 a_22550_8988.t7 990.34
R20797 a_22550_8988.n1 a_22550_8988.t4 408.211
R20798 a_22550_8988.n0 a_22550_8988.t6 286.438
R20799 a_22550_8988.n0 a_22550_8988.t5 286.438
R20800 a_22550_8988.n4 a_22550_8988.n3 185.55
R20801 a_22550_8988.t7 a_22550_8988.n0 160.666
R20802 a_22550_8988.n3 a_22550_8988.t1 28.568
R20803 a_22550_8988.n4 a_22550_8988.t0 28.565
R20804 a_22550_8988.t2 a_22550_8988.n4 28.565
R20805 a_22550_8988.n2 a_22550_8988.t3 21.471
R20806 a_22550_8988.n2 a_22550_8988.n1 12.567
R20807 a_22550_8988.n3 a_22550_8988.n2 2.677
R20808 a_13401_n2178.n2 a_13401_n2178.t4 990.34
R20809 a_13401_n2178.n2 a_13401_n2178.t6 408.211
R20810 a_13401_n2178.n1 a_13401_n2178.t7 286.438
R20811 a_13401_n2178.n1 a_13401_n2178.t5 286.438
R20812 a_13401_n2178.n4 a_13401_n2178.n0 185.55
R20813 a_13401_n2178.t4 a_13401_n2178.n1 160.666
R20814 a_13401_n2178.n3 a_13401_n2178.n2 37.035
R20815 a_13401_n2178.t2 a_13401_n2178.n4 28.568
R20816 a_13401_n2178.n0 a_13401_n2178.t0 28.565
R20817 a_13401_n2178.n0 a_13401_n2178.t1 28.565
R20818 a_13401_n2178.n3 a_13401_n2178.t3 21.376
R20819 a_13401_n2178.n4 a_13401_n2178.n3 1.637
R20820 a_13461_n2152.t3 a_13461_n2152.n0 14.282
R20821 a_13461_n2152.n0 a_13461_n2152.t4 14.282
R20822 a_13461_n2152.n0 a_13461_n2152.n9 89.977
R20823 a_13461_n2152.n9 a_13461_n2152.n7 75.815
R20824 a_13461_n2152.n9 a_13461_n2152.n6 77.456
R20825 a_13461_n2152.n6 a_13461_n2152.n4 77.456
R20826 a_13461_n2152.n4 a_13461_n2152.n2 77.784
R20827 a_13461_n2152.n7 a_13461_n2152.n8 167.433
R20828 a_13461_n2152.n8 a_13461_n2152.t0 14.282
R20829 a_13461_n2152.n8 a_13461_n2152.t2 14.282
R20830 a_13461_n2152.n7 a_13461_n2152.t1 104.259
R20831 a_13461_n2152.n6 a_13461_n2152.n5 89.977
R20832 a_13461_n2152.n5 a_13461_n2152.t11 14.282
R20833 a_13461_n2152.n5 a_13461_n2152.t7 14.282
R20834 a_13461_n2152.n4 a_13461_n2152.n3 89.977
R20835 a_13461_n2152.n3 a_13461_n2152.t6 14.282
R20836 a_13461_n2152.n3 a_13461_n2152.t5 14.282
R20837 a_13461_n2152.n2 a_13461_n2152.t10 104.259
R20838 a_13461_n2152.n2 a_13461_n2152.n1 167.433
R20839 a_13461_n2152.n1 a_13461_n2152.t9 14.282
R20840 a_13461_n2152.n1 a_13461_n2152.t8 14.282
R20841 a_26460_20259.t0 a_26460_20259.t1 17.4
R20842 a_45050_6179.t6 a_45050_6179.t7 574.43
R20843 a_45050_6179.n1 a_45050_6179.t4 285.109
R20844 a_45050_6179.n3 a_45050_6179.n2 197.217
R20845 a_45050_6179.n4 a_45050_6179.n0 192.754
R20846 a_45050_6179.n1 a_45050_6179.t5 160.666
R20847 a_45050_6179.n2 a_45050_6179.t6 160.666
R20848 a_45050_6179.n2 a_45050_6179.n1 114.829
R20849 a_45050_6179.t2 a_45050_6179.n4 28.568
R20850 a_45050_6179.n0 a_45050_6179.t1 28.565
R20851 a_45050_6179.n0 a_45050_6179.t0 28.565
R20852 a_45050_6179.n3 a_45050_6179.t3 18.838
R20853 a_45050_6179.n4 a_45050_6179.n3 1.129
R20854 a_46776_9742.n0 a_46776_9742.t4 14.282
R20855 a_46776_9742.n0 a_46776_9742.t3 14.282
R20856 a_46776_9742.n1 a_46776_9742.t2 14.282
R20857 a_46776_9742.n1 a_46776_9742.t1 14.282
R20858 a_46776_9742.t0 a_46776_9742.n3 14.282
R20859 a_46776_9742.n3 a_46776_9742.t5 14.282
R20860 a_46776_9742.n2 a_46776_9742.n0 2.546
R20861 a_46776_9742.n2 a_46776_9742.n1 2.367
R20862 a_46776_9742.n3 a_46776_9742.n2 0.001
R20863 a_13711_14458.n0 a_13711_14458.t7 14.282
R20864 a_13711_14458.t6 a_13711_14458.n0 14.282
R20865 a_13711_14458.n0 a_13711_14458.n9 89.977
R20866 a_13711_14458.n6 a_13711_14458.n7 77.784
R20867 a_13711_14458.n4 a_13711_14458.n6 77.456
R20868 a_13711_14458.n9 a_13711_14458.n4 77.456
R20869 a_13711_14458.n9 a_13711_14458.n2 75.815
R20870 a_13711_14458.n7 a_13711_14458.n8 167.433
R20871 a_13711_14458.n8 a_13711_14458.t9 14.282
R20872 a_13711_14458.n8 a_13711_14458.t10 14.282
R20873 a_13711_14458.n7 a_13711_14458.t11 104.259
R20874 a_13711_14458.n6 a_13711_14458.n5 89.977
R20875 a_13711_14458.n5 a_13711_14458.t5 14.282
R20876 a_13711_14458.n5 a_13711_14458.t4 14.282
R20877 a_13711_14458.n4 a_13711_14458.n3 89.977
R20878 a_13711_14458.n3 a_13711_14458.t3 14.282
R20879 a_13711_14458.n3 a_13711_14458.t8 14.282
R20880 a_13711_14458.n2 a_13711_14458.t0 104.259
R20881 a_13711_14458.n2 a_13711_14458.n1 167.433
R20882 a_13711_14458.n1 a_13711_14458.t2 14.282
R20883 a_13711_14458.n1 a_13711_14458.t1 14.282
R20884 a_13178_13728.t5 a_13178_13728.n0 14.283
R20885 a_13178_13728.n0 a_13178_13728.n5 0.852
R20886 a_13178_13728.n5 a_13178_13728.n6 4.366
R20887 a_13178_13728.n6 a_13178_13728.n7 258.161
R20888 a_13178_13728.n7 a_13178_13728.t4 14.282
R20889 a_13178_13728.n7 a_13178_13728.t3 14.282
R20890 a_13178_13728.n6 a_13178_13728.t2 14.283
R20891 a_13178_13728.n5 a_13178_13728.n4 97.614
R20892 a_13178_13728.n4 a_13178_13728.t9 200.029
R20893 a_13178_13728.t9 a_13178_13728.n3 206.421
R20894 a_13178_13728.n3 a_13178_13728.t10 80.333
R20895 a_13178_13728.n3 a_13178_13728.t11 206.421
R20896 a_13178_13728.n4 a_13178_13728.t8 1527.4
R20897 a_13178_13728.t8 a_13178_13728.n2 657.379
R20898 a_13178_13728.n2 a_13178_13728.t1 8.7
R20899 a_13178_13728.n2 a_13178_13728.t0 8.7
R20900 a_13178_13728.n0 a_13178_13728.n1 258.161
R20901 a_13178_13728.n1 a_13178_13728.t6 14.282
R20902 a_13178_13728.n1 a_13178_13728.t7 14.282
R20903 a_61525_1042.n1 a_61525_1042.t9 989.744
R20904 a_61525_1042.n1 a_61525_1042.t11 408.806
R20905 a_61525_1042.n0 a_61525_1042.t10 287.241
R20906 a_61525_1042.n0 a_61525_1042.t8 287.241
R20907 a_61525_1042.n7 a_61525_1042.n1 224.559
R20908 a_61525_1042.t9 a_61525_1042.n0 160.666
R20909 a_61525_1042.n5 a_61525_1042.n3 157.665
R20910 a_61525_1042.n5 a_61525_1042.n4 122.999
R20911 a_61525_1042.n8 a_61525_1042.n7 90.436
R20912 a_61525_1042.n6 a_61525_1042.n2 90.416
R20913 a_61525_1042.n7 a_61525_1042.n6 74.302
R20914 a_61525_1042.n6 a_61525_1042.n5 50.575
R20915 a_61525_1042.n2 a_61525_1042.t0 14.282
R20916 a_61525_1042.n2 a_61525_1042.t4 14.282
R20917 a_61525_1042.n4 a_61525_1042.t3 14.282
R20918 a_61525_1042.n4 a_61525_1042.t5 14.282
R20919 a_61525_1042.n8 a_61525_1042.t1 14.282
R20920 a_61525_1042.t2 a_61525_1042.n8 14.282
R20921 a_61525_1042.n3 a_61525_1042.t7 8.7
R20922 a_61525_1042.n3 a_61525_1042.t6 8.7
R20923 a_61827_6884.n1 a_61827_6884.t6 318.922
R20924 a_61827_6884.n0 a_61827_6884.t4 274.739
R20925 a_61827_6884.n0 a_61827_6884.t7 274.739
R20926 a_61827_6884.n1 a_61827_6884.t5 269.116
R20927 a_61827_6884.t6 a_61827_6884.n0 179.946
R20928 a_61827_6884.n2 a_61827_6884.n1 105.178
R20929 a_61827_6884.n3 a_61827_6884.t1 29.444
R20930 a_61827_6884.n4 a_61827_6884.t0 28.565
R20931 a_61827_6884.t2 a_61827_6884.n4 28.565
R20932 a_61827_6884.n2 a_61827_6884.t3 18.145
R20933 a_61827_6884.n3 a_61827_6884.n2 2.878
R20934 a_61827_6884.n4 a_61827_6884.n3 0.764
R20935 a_59557_20438.t0 a_59557_20438.t1 17.4
R20936 a_61216_21369.t0 a_61216_21369.n0 14.282
R20937 a_61216_21369.n0 a_61216_21369.t7 14.282
R20938 a_61216_21369.n0 a_61216_21369.n12 90.416
R20939 a_61216_21369.n12 a_61216_21369.n11 50.575
R20940 a_61216_21369.n12 a_61216_21369.n8 74.302
R20941 a_61216_21369.n11 a_61216_21369.n10 157.665
R20942 a_61216_21369.n10 a_61216_21369.t3 8.7
R20943 a_61216_21369.n10 a_61216_21369.t4 8.7
R20944 a_61216_21369.n11 a_61216_21369.n9 122.999
R20945 a_61216_21369.n9 a_61216_21369.t2 14.282
R20946 a_61216_21369.n9 a_61216_21369.t1 14.282
R20947 a_61216_21369.n8 a_61216_21369.n7 90.436
R20948 a_61216_21369.n7 a_61216_21369.t5 14.282
R20949 a_61216_21369.n7 a_61216_21369.t6 14.282
R20950 a_61216_21369.n8 a_61216_21369.n1 342.688
R20951 a_61216_21369.n1 a_61216_21369.n6 126.566
R20952 a_61216_21369.n6 a_61216_21369.t11 294.653
R20953 a_61216_21369.n6 a_61216_21369.t15 111.663
R20954 a_61216_21369.n1 a_61216_21369.n5 552.333
R20955 a_61216_21369.n5 a_61216_21369.n4 6.615
R20956 a_61216_21369.n4 a_61216_21369.t13 93.989
R20957 a_61216_21369.n5 a_61216_21369.n3 97.816
R20958 a_61216_21369.n3 a_61216_21369.t14 80.333
R20959 a_61216_21369.n3 a_61216_21369.t8 394.151
R20960 a_61216_21369.t8 a_61216_21369.n2 269.523
R20961 a_61216_21369.n2 a_61216_21369.t9 160.666
R20962 a_61216_21369.n2 a_61216_21369.t10 269.523
R20963 a_61216_21369.n4 a_61216_21369.t12 198.043
R20964 a_62996_21369.t6 a_62996_21369.n0 14.282
R20965 a_62996_21369.n0 a_62996_21369.t7 14.282
R20966 a_62996_21369.n0 a_62996_21369.n9 0.999
R20967 a_62996_21369.n9 a_62996_21369.n6 0.575
R20968 a_62996_21369.n6 a_62996_21369.n8 0.2
R20969 a_62996_21369.n8 a_62996_21369.t8 16.058
R20970 a_62996_21369.n8 a_62996_21369.n7 0.999
R20971 a_62996_21369.n7 a_62996_21369.t10 14.282
R20972 a_62996_21369.n7 a_62996_21369.t9 14.282
R20973 a_62996_21369.n9 a_62996_21369.t11 16.058
R20974 a_62996_21369.n6 a_62996_21369.n4 0.227
R20975 a_62996_21369.n4 a_62996_21369.n5 1.511
R20976 a_62996_21369.n5 a_62996_21369.t2 14.282
R20977 a_62996_21369.n5 a_62996_21369.t1 14.282
R20978 a_62996_21369.n4 a_62996_21369.n1 0.669
R20979 a_62996_21369.n1 a_62996_21369.n2 0.001
R20980 a_62996_21369.n1 a_62996_21369.n3 267.767
R20981 a_62996_21369.n3 a_62996_21369.t4 14.282
R20982 a_62996_21369.n3 a_62996_21369.t3 14.282
R20983 a_62996_21369.n2 a_62996_21369.t0 14.282
R20984 a_62996_21369.n2 a_62996_21369.t5 14.282
R20985 a_46228_21076.n0 a_46228_21076.t9 214.335
R20986 a_46228_21076.t7 a_46228_21076.n0 214.335
R20987 a_46228_21076.n1 a_46228_21076.t7 143.851
R20988 a_46228_21076.n1 a_46228_21076.t10 135.658
R20989 a_46228_21076.n0 a_46228_21076.t8 80.333
R20990 a_46228_21076.n2 a_46228_21076.t6 28.565
R20991 a_46228_21076.n2 a_46228_21076.t4 28.565
R20992 a_46228_21076.n4 a_46228_21076.t5 28.565
R20993 a_46228_21076.n4 a_46228_21076.t0 28.565
R20994 a_46228_21076.n7 a_46228_21076.t1 28.565
R20995 a_46228_21076.t2 a_46228_21076.n7 28.565
R20996 a_46228_21076.n6 a_46228_21076.t3 9.714
R20997 a_46228_21076.n7 a_46228_21076.n6 1.003
R20998 a_46228_21076.n5 a_46228_21076.n3 0.833
R20999 a_46228_21076.n3 a_46228_21076.n2 0.653
R21000 a_46228_21076.n5 a_46228_21076.n4 0.653
R21001 a_46228_21076.n6 a_46228_21076.n5 0.341
R21002 a_46228_21076.n3 a_46228_21076.n1 0.032
R21003 a_22584_5326.n1 a_22584_5326.t7 318.922
R21004 a_22584_5326.n0 a_22584_5326.t5 273.935
R21005 a_22584_5326.n0 a_22584_5326.t6 273.935
R21006 a_22584_5326.n1 a_22584_5326.t4 269.116
R21007 a_22584_5326.n4 a_22584_5326.n3 193.227
R21008 a_22584_5326.t7 a_22584_5326.n0 179.142
R21009 a_22584_5326.n2 a_22584_5326.n1 106.999
R21010 a_22584_5326.n3 a_22584_5326.t1 28.568
R21011 a_22584_5326.n4 a_22584_5326.t0 28.565
R21012 a_22584_5326.t2 a_22584_5326.n4 28.565
R21013 a_22584_5326.n2 a_22584_5326.t3 18.149
R21014 a_22584_5326.n3 a_22584_5326.n2 3.726
R21015 a_22290_4620.t0 a_22290_4620.t1 380.209
R21016 a_11346_7655.t0 a_11346_7655.t1 17.4
R21017 a_16320_4620.t0 a_16320_4620.t1 17.4
R21018 a_60404_18575.t7 a_60404_18575.t4 800.071
R21019 a_60404_18575.n3 a_60404_18575.n2 659.095
R21020 a_60404_18575.n1 a_60404_18575.t5 285.109
R21021 a_60404_18575.n2 a_60404_18575.t7 193.602
R21022 a_60404_18575.n4 a_60404_18575.n0 192.754
R21023 a_60404_18575.n1 a_60404_18575.t6 160.666
R21024 a_60404_18575.n2 a_60404_18575.n1 91.507
R21025 a_60404_18575.t2 a_60404_18575.n4 28.568
R21026 a_60404_18575.n0 a_60404_18575.t0 28.565
R21027 a_60404_18575.n0 a_60404_18575.t1 28.565
R21028 a_60404_18575.n3 a_60404_18575.t3 19.063
R21029 a_60404_18575.n4 a_60404_18575.n3 1.005
R21030 a_39262_7515.n2 a_39262_7515.t6 318.922
R21031 a_39262_7515.n1 a_39262_7515.t7 273.935
R21032 a_39262_7515.n1 a_39262_7515.t4 273.935
R21033 a_39262_7515.n2 a_39262_7515.t5 269.116
R21034 a_39262_7515.n4 a_39262_7515.n0 193.227
R21035 a_39262_7515.t6 a_39262_7515.n1 179.142
R21036 a_39262_7515.n3 a_39262_7515.n2 106.999
R21037 a_39262_7515.t2 a_39262_7515.n4 28.568
R21038 a_39262_7515.n0 a_39262_7515.t1 28.565
R21039 a_39262_7515.n0 a_39262_7515.t0 28.565
R21040 a_39262_7515.n3 a_39262_7515.t3 18.149
R21041 a_39262_7515.n4 a_39262_7515.n3 3.726
R21042 a_39807_6822.n6 a_39807_6822.n4 552.333
R21043 a_39807_6822.n2 a_39807_6822.t8 394.151
R21044 a_39807_6822.n7 a_39807_6822.n6 342.688
R21045 a_39807_6822.n5 a_39807_6822.t11 294.653
R21046 a_39807_6822.n1 a_39807_6822.t10 269.523
R21047 a_39807_6822.t8 a_39807_6822.n1 269.523
R21048 a_39807_6822.n3 a_39807_6822.t12 198.043
R21049 a_39807_6822.n1 a_39807_6822.t14 160.666
R21050 a_39807_6822.n10 a_39807_6822.n8 157.665
R21051 a_39807_6822.n6 a_39807_6822.n5 126.566
R21052 a_39807_6822.n10 a_39807_6822.n9 122.999
R21053 a_39807_6822.n5 a_39807_6822.t13 111.663
R21054 a_39807_6822.n4 a_39807_6822.n2 97.816
R21055 a_39807_6822.n3 a_39807_6822.t9 93.989
R21056 a_39807_6822.n7 a_39807_6822.n0 90.436
R21057 a_39807_6822.n12 a_39807_6822.n11 90.416
R21058 a_39807_6822.n2 a_39807_6822.t15 80.333
R21059 a_39807_6822.n11 a_39807_6822.n7 74.302
R21060 a_39807_6822.n11 a_39807_6822.n10 50.575
R21061 a_39807_6822.n0 a_39807_6822.t5 14.282
R21062 a_39807_6822.n0 a_39807_6822.t7 14.282
R21063 a_39807_6822.n9 a_39807_6822.t1 14.282
R21064 a_39807_6822.n9 a_39807_6822.t0 14.282
R21065 a_39807_6822.n12 a_39807_6822.t6 14.282
R21066 a_39807_6822.t2 a_39807_6822.n12 14.282
R21067 a_39807_6822.n8 a_39807_6822.t4 8.7
R21068 a_39807_6822.n8 a_39807_6822.t3 8.7
R21069 a_39807_6822.n4 a_39807_6822.n3 6.615
R21070 a_52892_6842.n8 a_52892_6842.n0 267.767
R21071 a_52892_6842.n4 a_52892_6842.t9 16.058
R21072 a_52892_6842.n2 a_52892_6842.t6 16.058
R21073 a_52892_6842.n3 a_52892_6842.t11 14.282
R21074 a_52892_6842.n3 a_52892_6842.t10 14.282
R21075 a_52892_6842.n1 a_52892_6842.t8 14.282
R21076 a_52892_6842.n1 a_52892_6842.t7 14.282
R21077 a_52892_6842.n6 a_52892_6842.t1 14.282
R21078 a_52892_6842.n6 a_52892_6842.t0 14.282
R21079 a_52892_6842.n0 a_52892_6842.t3 14.282
R21080 a_52892_6842.n0 a_52892_6842.t5 14.282
R21081 a_52892_6842.n9 a_52892_6842.t4 14.282
R21082 a_52892_6842.t2 a_52892_6842.n9 14.282
R21083 a_52892_6842.n7 a_52892_6842.n6 1.511
R21084 a_52892_6842.n4 a_52892_6842.n3 0.999
R21085 a_52892_6842.n2 a_52892_6842.n1 0.999
R21086 a_52892_6842.n8 a_52892_6842.n7 0.669
R21087 a_52892_6842.n5 a_52892_6842.n4 0.575
R21088 a_52892_6842.n7 a_52892_6842.n5 0.227
R21089 a_52892_6842.n5 a_52892_6842.n2 0.2
R21090 a_52892_6842.n9 a_52892_6842.n8 0.001
R21091 a_23958_10387.t0 a_23958_10387.t1 17.4
R21092 a_22598_10990.t1 a_22598_10990.n0 14.282
R21093 a_22598_10990.n0 a_22598_10990.t4 14.282
R21094 a_22598_10990.n0 a_22598_10990.n1 258.161
R21095 a_22598_10990.n1 a_22598_10990.t3 14.283
R21096 a_22598_10990.n1 a_22598_10990.n7 4.366
R21097 a_22598_10990.n7 a_22598_10990.n5 0.852
R21098 a_22598_10990.n5 a_22598_10990.n6 258.161
R21099 a_22598_10990.n6 a_22598_10990.t6 14.282
R21100 a_22598_10990.n6 a_22598_10990.t7 14.282
R21101 a_22598_10990.n5 a_22598_10990.t5 14.283
R21102 a_22598_10990.n7 a_22598_10990.n4 97.614
R21103 a_22598_10990.n4 a_22598_10990.t8 200.029
R21104 a_22598_10990.t8 a_22598_10990.n3 206.421
R21105 a_22598_10990.n3 a_22598_10990.t9 80.333
R21106 a_22598_10990.n3 a_22598_10990.t10 206.421
R21107 a_22598_10990.n4 a_22598_10990.t11 1527.4
R21108 a_22598_10990.t11 a_22598_10990.n2 657.379
R21109 a_22598_10990.n2 a_22598_10990.t2 8.7
R21110 a_22598_10990.n2 a_22598_10990.t0 8.7
R21111 a_23131_11720.n0 a_23131_11720.n9 167.433
R21112 a_23131_11720.t9 a_23131_11720.n0 14.282
R21113 a_23131_11720.n0 a_23131_11720.t10 14.282
R21114 a_23131_11720.n9 a_23131_11720.n8 77.784
R21115 a_23131_11720.n8 a_23131_11720.n6 77.456
R21116 a_23131_11720.n6 a_23131_11720.n4 77.456
R21117 a_23131_11720.n4 a_23131_11720.n2 75.815
R21118 a_23131_11720.n9 a_23131_11720.t11 104.259
R21119 a_23131_11720.n8 a_23131_11720.n7 89.977
R21120 a_23131_11720.n7 a_23131_11720.t2 14.282
R21121 a_23131_11720.n7 a_23131_11720.t1 14.282
R21122 a_23131_11720.n6 a_23131_11720.n5 89.977
R21123 a_23131_11720.n5 a_23131_11720.t0 14.282
R21124 a_23131_11720.n5 a_23131_11720.t6 14.282
R21125 a_23131_11720.n4 a_23131_11720.n3 89.977
R21126 a_23131_11720.n3 a_23131_11720.t8 14.282
R21127 a_23131_11720.n3 a_23131_11720.t7 14.282
R21128 a_23131_11720.n2 a_23131_11720.t4 104.259
R21129 a_23131_11720.n2 a_23131_11720.n1 167.433
R21130 a_23131_11720.n1 a_23131_11720.t3 14.282
R21131 a_23131_11720.n1 a_23131_11720.t5 14.282
R21132 a_45041_9433.t4 a_45041_9433.t5 800.071
R21133 a_45041_9433.n2 a_45041_9433.n1 659.097
R21134 a_45041_9433.n0 a_45041_9433.t7 285.109
R21135 a_45041_9433.n1 a_45041_9433.t4 193.602
R21136 a_45041_9433.n4 a_45041_9433.n3 192.754
R21137 a_45041_9433.n0 a_45041_9433.t6 160.666
R21138 a_45041_9433.n1 a_45041_9433.n0 91.507
R21139 a_45041_9433.n3 a_45041_9433.t1 28.568
R21140 a_45041_9433.n4 a_45041_9433.t0 28.565
R21141 a_45041_9433.t2 a_45041_9433.n4 28.565
R21142 a_45041_9433.n2 a_45041_9433.t3 19.061
R21143 a_45041_9433.n3 a_45041_9433.n2 1.005
R21144 a_65649_10704.n0 a_65649_10704.t11 14.282
R21145 a_65649_10704.t3 a_65649_10704.n0 14.282
R21146 a_65649_10704.n0 a_65649_10704.n9 0.999
R21147 a_65649_10704.n6 a_65649_10704.n8 0.575
R21148 a_65649_10704.n9 a_65649_10704.n6 0.2
R21149 a_65649_10704.n9 a_65649_10704.t4 16.058
R21150 a_65649_10704.n8 a_65649_10704.n7 0.999
R21151 a_65649_10704.n7 a_65649_10704.t6 14.282
R21152 a_65649_10704.n7 a_65649_10704.t7 14.282
R21153 a_65649_10704.n8 a_65649_10704.t5 16.058
R21154 a_65649_10704.n6 a_65649_10704.n4 0.227
R21155 a_65649_10704.n4 a_65649_10704.n5 1.511
R21156 a_65649_10704.n5 a_65649_10704.t10 14.282
R21157 a_65649_10704.n5 a_65649_10704.t9 14.282
R21158 a_65649_10704.n4 a_65649_10704.n1 0.669
R21159 a_65649_10704.n1 a_65649_10704.n2 0.001
R21160 a_65649_10704.n1 a_65649_10704.n3 267.767
R21161 a_65649_10704.n3 a_65649_10704.t1 14.282
R21162 a_65649_10704.n3 a_65649_10704.t0 14.282
R21163 a_65649_10704.n2 a_65649_10704.t8 14.282
R21164 a_65649_10704.n2 a_65649_10704.t2 14.282
R21165 a_10844_n3481.t0 a_10844_n3481.t1 17.4
R21166 a_35238_789.t0 a_35238_789.t1 17.4
R21167 a_41905_21347.n1 a_41905_21347.t4 318.922
R21168 a_41905_21347.n0 a_41905_21347.t6 274.739
R21169 a_41905_21347.n0 a_41905_21347.t5 274.739
R21170 a_41905_21347.n1 a_41905_21347.t7 269.116
R21171 a_41905_21347.t4 a_41905_21347.n0 179.946
R21172 a_41905_21347.n2 a_41905_21347.n1 107.263
R21173 a_41905_21347.n3 a_41905_21347.t0 29.444
R21174 a_41905_21347.n4 a_41905_21347.t1 28.565
R21175 a_41905_21347.t2 a_41905_21347.n4 28.565
R21176 a_41905_21347.n2 a_41905_21347.t3 18.145
R21177 a_41905_21347.n3 a_41905_21347.n2 2.878
R21178 a_41905_21347.n4 a_41905_21347.n3 0.764
R21179 a_9928_8988.n2 a_9928_8988.t6 990.34
R21180 a_9928_8988.n2 a_9928_8988.t4 408.211
R21181 a_9928_8988.n1 a_9928_8988.t5 286.438
R21182 a_9928_8988.n1 a_9928_8988.t7 286.438
R21183 a_9928_8988.n4 a_9928_8988.n0 185.55
R21184 a_9928_8988.t6 a_9928_8988.n1 160.666
R21185 a_9928_8988.t2 a_9928_8988.n4 28.568
R21186 a_9928_8988.n0 a_9928_8988.t1 28.565
R21187 a_9928_8988.n0 a_9928_8988.t0 28.565
R21188 a_9928_8988.n3 a_9928_8988.t3 23.433
R21189 a_9928_8988.n3 a_9928_8988.n2 11.507
R21190 a_9928_8988.n4 a_9928_8988.n3 0.002
R21191 a_22322_n2148.n2 a_22322_n2148.t6 448.382
R21192 a_22322_n2148.n1 a_22322_n2148.t4 286.438
R21193 a_22322_n2148.n1 a_22322_n2148.t7 286.438
R21194 a_22322_n2148.n0 a_22322_n2148.t5 247.69
R21195 a_22322_n2148.n4 a_22322_n2148.n3 182.117
R21196 a_22322_n2148.t6 a_22322_n2148.n1 160.666
R21197 a_22322_n2148.n3 a_22322_n2148.t0 28.568
R21198 a_22322_n2148.n4 a_22322_n2148.t1 28.565
R21199 a_22322_n2148.t2 a_22322_n2148.n4 28.565
R21200 a_22322_n2148.n0 a_22322_n2148.t3 18.127
R21201 a_22322_n2148.n2 a_22322_n2148.n0 4.039
R21202 a_22322_n2148.n3 a_22322_n2148.n2 0.937
R21203 a_39254_1735.n2 a_39254_1735.t4 318.922
R21204 a_39254_1735.n1 a_39254_1735.t5 273.935
R21205 a_39254_1735.n1 a_39254_1735.t7 273.935
R21206 a_39254_1735.n2 a_39254_1735.t6 269.116
R21207 a_39254_1735.n4 a_39254_1735.n0 193.227
R21208 a_39254_1735.t4 a_39254_1735.n1 179.142
R21209 a_39254_1735.n3 a_39254_1735.n2 106.999
R21210 a_39254_1735.t2 a_39254_1735.n4 28.568
R21211 a_39254_1735.n0 a_39254_1735.t1 28.565
R21212 a_39254_1735.n0 a_39254_1735.t0 28.565
R21213 a_39254_1735.n3 a_39254_1735.t3 18.149
R21214 a_39254_1735.n4 a_39254_1735.n3 3.726
R21215 a_39717_18601.n1 a_39717_18601.t3 14.282
R21216 a_39717_18601.n1 a_39717_18601.t5 14.282
R21217 a_39717_18601.n0 a_39717_18601.t4 14.282
R21218 a_39717_18601.n0 a_39717_18601.t2 14.282
R21219 a_39717_18601.n3 a_39717_18601.t1 14.282
R21220 a_39717_18601.t0 a_39717_18601.n3 14.282
R21221 a_39717_18601.n2 a_39717_18601.n0 2.546
R21222 a_39717_18601.n3 a_39717_18601.n2 2.367
R21223 a_39717_18601.n2 a_39717_18601.n1 0.001
R21224 a_39582_17945.t6 a_39582_17945.n2 404.877
R21225 a_39582_17945.n1 a_39582_17945.t5 210.902
R21226 a_39582_17945.n3 a_39582_17945.t6 136.949
R21227 a_39582_17945.n2 a_39582_17945.n1 107.801
R21228 a_39582_17945.n1 a_39582_17945.t7 80.333
R21229 a_39582_17945.n2 a_39582_17945.t8 80.333
R21230 a_39582_17945.n0 a_39582_17945.t0 17.4
R21231 a_39582_17945.n0 a_39582_17945.t4 17.4
R21232 a_39582_17945.n4 a_39582_17945.t1 15.032
R21233 a_39582_17945.n5 a_39582_17945.t2 14.282
R21234 a_39582_17945.t3 a_39582_17945.n5 14.282
R21235 a_39582_17945.n5 a_39582_17945.n4 1.65
R21236 a_39582_17945.n3 a_39582_17945.n0 0.657
R21237 a_39582_17945.n4 a_39582_17945.n3 0.614
R21238 a_30154_8749.n2 a_30154_8749.t6 318.119
R21239 a_30154_8749.n2 a_30154_8749.t4 269.919
R21240 a_30154_8749.n1 a_30154_8749.t7 267.256
R21241 a_30154_8749.n1 a_30154_8749.t5 267.256
R21242 a_30154_8749.n4 a_30154_8749.n0 193.227
R21243 a_30154_8749.t6 a_30154_8749.n1 160.666
R21244 a_30154_8749.n3 a_30154_8749.n2 106.999
R21245 a_30154_8749.t2 a_30154_8749.n4 28.568
R21246 a_30154_8749.n0 a_30154_8749.t0 28.565
R21247 a_30154_8749.n0 a_30154_8749.t1 28.565
R21248 a_30154_8749.n3 a_30154_8749.t3 18.149
R21249 a_30154_8749.n4 a_30154_8749.n3 3.726
R21250 a_34985_4186.n4 a_34985_4186.t10 214.335
R21251 a_34985_4186.t9 a_34985_4186.n4 214.335
R21252 a_34985_4186.n5 a_34985_4186.t9 143.851
R21253 a_34985_4186.n5 a_34985_4186.t8 135.658
R21254 a_34985_4186.n4 a_34985_4186.t7 80.333
R21255 a_34985_4186.n0 a_34985_4186.t3 28.565
R21256 a_34985_4186.n0 a_34985_4186.t4 28.565
R21257 a_34985_4186.n2 a_34985_4186.t1 28.565
R21258 a_34985_4186.n2 a_34985_4186.t5 28.565
R21259 a_34985_4186.n7 a_34985_4186.t0 28.565
R21260 a_34985_4186.t2 a_34985_4186.n7 28.565
R21261 a_34985_4186.n1 a_34985_4186.t6 9.714
R21262 a_34985_4186.n1 a_34985_4186.n0 1.003
R21263 a_34985_4186.n6 a_34985_4186.n3 0.833
R21264 a_34985_4186.n3 a_34985_4186.n2 0.653
R21265 a_34985_4186.n7 a_34985_4186.n6 0.653
R21266 a_34985_4186.n3 a_34985_4186.n1 0.341
R21267 a_34985_4186.n6 a_34985_4186.n5 0.032
R21268 a_24652_5324.n1 a_24652_5324.t4 318.922
R21269 a_24652_5324.n0 a_24652_5324.t6 273.935
R21270 a_24652_5324.n0 a_24652_5324.t7 273.935
R21271 a_24652_5324.n1 a_24652_5324.t5 269.116
R21272 a_24652_5324.n4 a_24652_5324.n3 193.227
R21273 a_24652_5324.t4 a_24652_5324.n0 179.142
R21274 a_24652_5324.n2 a_24652_5324.n1 106.999
R21275 a_24652_5324.n3 a_24652_5324.t0 28.568
R21276 a_24652_5324.t2 a_24652_5324.n4 28.565
R21277 a_24652_5324.n4 a_24652_5324.t1 28.565
R21278 a_24652_5324.n2 a_24652_5324.t3 18.149
R21279 a_24652_5324.n3 a_24652_5324.n2 3.726
R21280 a_61452_20637.t0 a_61452_20637.t1 17.4
R21281 a_11155_10847.n2 a_11155_10847.t6 448.381
R21282 a_11155_10847.n1 a_11155_10847.t5 286.438
R21283 a_11155_10847.n1 a_11155_10847.t7 286.438
R21284 a_11155_10847.n0 a_11155_10847.t4 247.69
R21285 a_11155_10847.n4 a_11155_10847.n3 182.117
R21286 a_11155_10847.t6 a_11155_10847.n1 160.666
R21287 a_11155_10847.n3 a_11155_10847.t1 28.568
R21288 a_11155_10847.t2 a_11155_10847.n4 28.565
R21289 a_11155_10847.n4 a_11155_10847.t0 28.565
R21290 a_11155_10847.n0 a_11155_10847.t3 18.127
R21291 a_11155_10847.n2 a_11155_10847.n0 4.036
R21292 a_11155_10847.n3 a_11155_10847.n2 0.937
R21293 a_23777_13581.n3 a_23777_13581.t5 448.381
R21294 a_23777_13581.n2 a_23777_13581.t4 286.438
R21295 a_23777_13581.n2 a_23777_13581.t6 286.438
R21296 a_23777_13581.n1 a_23777_13581.t7 247.69
R21297 a_23777_13581.n4 a_23777_13581.n0 182.117
R21298 a_23777_13581.t5 a_23777_13581.n2 160.666
R21299 a_23777_13581.t2 a_23777_13581.n4 28.568
R21300 a_23777_13581.n0 a_23777_13581.t0 28.565
R21301 a_23777_13581.n0 a_23777_13581.t1 28.565
R21302 a_23777_13581.n1 a_23777_13581.t3 18.127
R21303 a_23777_13581.n3 a_23777_13581.n1 4.036
R21304 a_23777_13581.n4 a_23777_13581.n3 0.937
R21305 a_280_n2152.n3 a_280_n2152.t6 448.382
R21306 a_280_n2152.n2 a_280_n2152.t5 286.438
R21307 a_280_n2152.n2 a_280_n2152.t7 286.438
R21308 a_280_n2152.n1 a_280_n2152.t4 247.69
R21309 a_280_n2152.n4 a_280_n2152.n0 182.117
R21310 a_280_n2152.t6 a_280_n2152.n2 160.666
R21311 a_280_n2152.t2 a_280_n2152.n4 28.568
R21312 a_280_n2152.n0 a_280_n2152.t0 28.565
R21313 a_280_n2152.n0 a_280_n2152.t1 28.565
R21314 a_280_n2152.n1 a_280_n2152.t3 18.127
R21315 a_280_n2152.n3 a_280_n2152.n1 4.039
R21316 a_280_n2152.n4 a_280_n2152.n3 0.937
R21317 a_19705_1744.n0 a_19705_1744.t4 14.282
R21318 a_19705_1744.t3 a_19705_1744.n0 14.282
R21319 a_19705_1744.n0 a_19705_1744.n9 89.977
R21320 a_19705_1744.n9 a_19705_1744.n7 75.815
R21321 a_19705_1744.n9 a_19705_1744.n6 77.456
R21322 a_19705_1744.n6 a_19705_1744.n4 77.456
R21323 a_19705_1744.n4 a_19705_1744.n2 77.784
R21324 a_19705_1744.n7 a_19705_1744.n8 167.433
R21325 a_19705_1744.n8 a_19705_1744.t8 14.282
R21326 a_19705_1744.n8 a_19705_1744.t6 14.282
R21327 a_19705_1744.n7 a_19705_1744.t7 104.259
R21328 a_19705_1744.n6 a_19705_1744.n5 89.977
R21329 a_19705_1744.n5 a_19705_1744.t5 14.282
R21330 a_19705_1744.n5 a_19705_1744.t1 14.282
R21331 a_19705_1744.n4 a_19705_1744.n3 89.977
R21332 a_19705_1744.n3 a_19705_1744.t2 14.282
R21333 a_19705_1744.n3 a_19705_1744.t0 14.282
R21334 a_19705_1744.n2 a_19705_1744.t10 104.259
R21335 a_19705_1744.n2 a_19705_1744.n1 167.433
R21336 a_19705_1744.n1 a_19705_1744.t9 14.282
R21337 a_19705_1744.n1 a_19705_1744.t11 14.282
R21338 a_52753_24325.n0 a_52753_24325.t9 214.335
R21339 a_52753_24325.t7 a_52753_24325.n0 214.335
R21340 a_52753_24325.n1 a_52753_24325.t7 143.851
R21341 a_52753_24325.n1 a_52753_24325.t10 135.658
R21342 a_52753_24325.n0 a_52753_24325.t8 80.333
R21343 a_52753_24325.n2 a_52753_24325.t4 28.565
R21344 a_52753_24325.n2 a_52753_24325.t5 28.565
R21345 a_52753_24325.n4 a_52753_24325.t6 28.565
R21346 a_52753_24325.n4 a_52753_24325.t1 28.565
R21347 a_52753_24325.n7 a_52753_24325.t2 28.565
R21348 a_52753_24325.t3 a_52753_24325.n7 28.565
R21349 a_52753_24325.n6 a_52753_24325.t0 9.714
R21350 a_52753_24325.n7 a_52753_24325.n6 1.003
R21351 a_52753_24325.n5 a_52753_24325.n3 0.833
R21352 a_52753_24325.n3 a_52753_24325.n2 0.653
R21353 a_52753_24325.n5 a_52753_24325.n4 0.653
R21354 a_52753_24325.n6 a_52753_24325.n5 0.341
R21355 a_52753_24325.n3 a_52753_24325.n1 0.032
R21356 a_59937_9742.t6 a_59937_9742.n3 404.877
R21357 a_59937_9742.n2 a_59937_9742.t7 210.902
R21358 a_59937_9742.n4 a_59937_9742.t6 136.943
R21359 a_59937_9742.n3 a_59937_9742.n2 107.801
R21360 a_59937_9742.n2 a_59937_9742.t8 80.333
R21361 a_59937_9742.n3 a_59937_9742.t5 80.333
R21362 a_59937_9742.n1 a_59937_9742.t0 17.4
R21363 a_59937_9742.n1 a_59937_9742.t2 17.4
R21364 a_59937_9742.t1 a_59937_9742.n5 15.032
R21365 a_59937_9742.n0 a_59937_9742.t4 14.282
R21366 a_59937_9742.n0 a_59937_9742.t3 14.282
R21367 a_59937_9742.n5 a_59937_9742.n0 1.65
R21368 a_59937_9742.n4 a_59937_9742.n1 0.672
R21369 a_59937_9742.n5 a_59937_9742.n4 0.665
R21370 a_57731_748.n4 a_57731_748.t8 214.335
R21371 a_57731_748.t9 a_57731_748.n4 214.335
R21372 a_57731_748.n5 a_57731_748.t9 143.851
R21373 a_57731_748.n5 a_57731_748.t10 135.658
R21374 a_57731_748.n4 a_57731_748.t7 80.333
R21375 a_57731_748.n0 a_57731_748.t5 28.565
R21376 a_57731_748.n0 a_57731_748.t3 28.565
R21377 a_57731_748.n2 a_57731_748.t0 28.565
R21378 a_57731_748.n2 a_57731_748.t4 28.565
R21379 a_57731_748.t2 a_57731_748.n7 28.565
R21380 a_57731_748.n7 a_57731_748.t1 28.565
R21381 a_57731_748.n1 a_57731_748.t6 9.714
R21382 a_57731_748.n1 a_57731_748.n0 1.003
R21383 a_57731_748.n6 a_57731_748.n3 0.833
R21384 a_57731_748.n3 a_57731_748.n2 0.653
R21385 a_57731_748.n7 a_57731_748.n6 0.653
R21386 a_57731_748.n3 a_57731_748.n1 0.341
R21387 a_57731_748.n6 a_57731_748.n5 0.032
R21388 a_57968_111.t0 a_57968_111.t1 17.4
R21389 a_39715_21079.n2 a_39715_21079.t7 214.335
R21390 a_39715_21079.t9 a_39715_21079.n2 214.335
R21391 a_39715_21079.n3 a_39715_21079.t9 143.851
R21392 a_39715_21079.n3 a_39715_21079.t8 135.658
R21393 a_39715_21079.n2 a_39715_21079.t10 80.333
R21394 a_39715_21079.n4 a_39715_21079.t0 28.565
R21395 a_39715_21079.n4 a_39715_21079.t1 28.565
R21396 a_39715_21079.n0 a_39715_21079.t4 28.565
R21397 a_39715_21079.n0 a_39715_21079.t5 28.565
R21398 a_39715_21079.t2 a_39715_21079.n7 28.565
R21399 a_39715_21079.n7 a_39715_21079.t3 28.565
R21400 a_39715_21079.n1 a_39715_21079.t6 9.714
R21401 a_39715_21079.n1 a_39715_21079.n0 1.003
R21402 a_39715_21079.n6 a_39715_21079.n5 0.833
R21403 a_39715_21079.n5 a_39715_21079.n4 0.653
R21404 a_39715_21079.n7 a_39715_21079.n6 0.653
R21405 a_39715_21079.n6 a_39715_21079.n1 0.341
R21406 a_39715_21079.n5 a_39715_21079.n3 0.032
R21407 a_39952_20442.t0 a_39952_20442.t1 17.4
R21408 a_61120_15037.t0 a_61120_15037.t1 17.4
R21409 a_6202_20866.t0 a_6202_20866.n0 14.283
R21410 a_6202_20866.n0 a_6202_20866.n7 258.161
R21411 a_6202_20866.n7 a_6202_20866.t2 14.282
R21412 a_6202_20866.n7 a_6202_20866.t1 14.282
R21413 a_6202_20866.n0 a_6202_20866.n6 4.366
R21414 a_6202_20866.n6 a_6202_20866.n4 0.852
R21415 a_6202_20866.n4 a_6202_20866.n5 258.161
R21416 a_6202_20866.n5 a_6202_20866.t5 14.282
R21417 a_6202_20866.n5 a_6202_20866.t7 14.282
R21418 a_6202_20866.n4 a_6202_20866.t6 14.283
R21419 a_6202_20866.n6 a_6202_20866.n3 97.614
R21420 a_6202_20866.n3 a_6202_20866.t10 200.029
R21421 a_6202_20866.t10 a_6202_20866.n2 206.421
R21422 a_6202_20866.n2 a_6202_20866.t11 80.333
R21423 a_6202_20866.n2 a_6202_20866.t8 206.421
R21424 a_6202_20866.n3 a_6202_20866.t9 1527.4
R21425 a_6202_20866.t9 a_6202_20866.n1 657.379
R21426 a_6202_20866.n1 a_6202_20866.t3 8.7
R21427 a_6202_20866.n1 a_6202_20866.t4 8.7
R21428 a_46818_20639.t7 a_46818_20639.t6 574.43
R21429 a_46818_20639.n0 a_46818_20639.t5 285.109
R21430 a_46818_20639.n2 a_46818_20639.n1 197.217
R21431 a_46818_20639.n4 a_46818_20639.n3 192.754
R21432 a_46818_20639.n0 a_46818_20639.t4 160.666
R21433 a_46818_20639.n1 a_46818_20639.t7 160.666
R21434 a_46818_20639.n1 a_46818_20639.n0 114.829
R21435 a_46818_20639.n3 a_46818_20639.t0 28.568
R21436 a_46818_20639.n4 a_46818_20639.t1 28.565
R21437 a_46818_20639.t2 a_46818_20639.n4 28.565
R21438 a_46818_20639.n2 a_46818_20639.t3 18.838
R21439 a_46818_20639.n3 a_46818_20639.n2 1.129
R21440 a_10576_1744.n4 a_10576_1744.t8 1527.4
R21441 a_10576_1744.t8 a_10576_1744.n3 657.379
R21442 a_10576_1744.n1 a_10576_1744.n0 258.161
R21443 a_10576_1744.n7 a_10576_1744.n6 258.161
R21444 a_10576_1744.n2 a_10576_1744.t10 206.421
R21445 a_10576_1744.t9 a_10576_1744.n2 206.421
R21446 a_10576_1744.n4 a_10576_1744.t9 200.029
R21447 a_10576_1744.n5 a_10576_1744.n4 97.614
R21448 a_10576_1744.n2 a_10576_1744.t11 80.333
R21449 a_10576_1744.n6 a_10576_1744.t1 14.283
R21450 a_10576_1744.n1 a_10576_1744.t5 14.283
R21451 a_10576_1744.n0 a_10576_1744.t7 14.282
R21452 a_10576_1744.n0 a_10576_1744.t6 14.282
R21453 a_10576_1744.n7 a_10576_1744.t0 14.282
R21454 a_10576_1744.t2 a_10576_1744.n7 14.282
R21455 a_10576_1744.n3 a_10576_1744.t3 8.7
R21456 a_10576_1744.n3 a_10576_1744.t4 8.7
R21457 a_10576_1744.n6 a_10576_1744.n5 4.366
R21458 a_10576_1744.n5 a_10576_1744.n1 0.852
R21459 a_24157_16385.n0 a_24157_16385.t7 214.335
R21460 a_24157_16385.t9 a_24157_16385.n0 214.335
R21461 a_24157_16385.n1 a_24157_16385.t9 143.851
R21462 a_24157_16385.n1 a_24157_16385.t10 135.658
R21463 a_24157_16385.n0 a_24157_16385.t8 80.333
R21464 a_24157_16385.n2 a_24157_16385.t5 28.565
R21465 a_24157_16385.n2 a_24157_16385.t3 28.565
R21466 a_24157_16385.n4 a_24157_16385.t4 28.565
R21467 a_24157_16385.n4 a_24157_16385.t0 28.565
R21468 a_24157_16385.n7 a_24157_16385.t1 28.565
R21469 a_24157_16385.t2 a_24157_16385.n7 28.565
R21470 a_24157_16385.n3 a_24157_16385.t6 9.714
R21471 a_24157_16385.n3 a_24157_16385.n2 1.003
R21472 a_24157_16385.n6 a_24157_16385.n5 0.833
R21473 a_24157_16385.n5 a_24157_16385.n4 0.653
R21474 a_24157_16385.n7 a_24157_16385.n6 0.653
R21475 a_24157_16385.n5 a_24157_16385.n3 0.341
R21476 a_24157_16385.n6 a_24157_16385.n1 0.032
R21477 a_14303_1255.n1 a_14303_1255.t7 867.497
R21478 a_14303_1255.n1 a_14303_1255.t6 615.911
R21479 a_14303_1255.n0 a_14303_1255.t4 286.438
R21480 a_14303_1255.n0 a_14303_1255.t5 286.438
R21481 a_14303_1255.n4 a_14303_1255.n3 185.55
R21482 a_14303_1255.t7 a_14303_1255.n0 160.666
R21483 a_14303_1255.n2 a_14303_1255.n1 127.305
R21484 a_14303_1255.n3 a_14303_1255.t1 28.568
R21485 a_14303_1255.n4 a_14303_1255.t2 28.565
R21486 a_14303_1255.t0 a_14303_1255.n4 28.565
R21487 a_14303_1255.n2 a_14303_1255.t3 20.393
R21488 a_14303_1255.n3 a_14303_1255.n2 1.832
R21489 a_59090_7603.n1 a_59090_7603.t7 318.922
R21490 a_59090_7603.n0 a_59090_7603.t4 273.935
R21491 a_59090_7603.n0 a_59090_7603.t5 273.935
R21492 a_59090_7603.n1 a_59090_7603.t6 269.116
R21493 a_59090_7603.n4 a_59090_7603.n3 193.227
R21494 a_59090_7603.t7 a_59090_7603.n0 179.142
R21495 a_59090_7603.n2 a_59090_7603.n1 106.999
R21496 a_59090_7603.n3 a_59090_7603.t1 28.568
R21497 a_59090_7603.n4 a_59090_7603.t0 28.565
R21498 a_59090_7603.t2 a_59090_7603.n4 28.565
R21499 a_59090_7603.n2 a_59090_7603.t3 18.149
R21500 a_59090_7603.n3 a_59090_7603.n2 3.726
R21501 a_51704_1914.t4 a_51704_1914.t6 574.43
R21502 a_51704_1914.n0 a_51704_1914.t5 285.109
R21503 a_51704_1914.n2 a_51704_1914.n1 211.136
R21504 a_51704_1914.n4 a_51704_1914.n3 192.754
R21505 a_51704_1914.n0 a_51704_1914.t7 160.666
R21506 a_51704_1914.n1 a_51704_1914.t4 160.666
R21507 a_51704_1914.n1 a_51704_1914.n0 114.829
R21508 a_51704_1914.n3 a_51704_1914.t0 28.568
R21509 a_51704_1914.t2 a_51704_1914.n4 28.565
R21510 a_51704_1914.n4 a_51704_1914.t1 28.565
R21511 a_51704_1914.n2 a_51704_1914.t3 19.084
R21512 a_51704_1914.n3 a_51704_1914.n2 1.051
R21513 a_54449_3877.t8 a_54449_3877.n2 404.877
R21514 a_54449_3877.n1 a_54449_3877.t5 210.902
R21515 a_54449_3877.n3 a_54449_3877.t8 136.943
R21516 a_54449_3877.n2 a_54449_3877.n1 107.801
R21517 a_54449_3877.n1 a_54449_3877.t7 80.333
R21518 a_54449_3877.n2 a_54449_3877.t6 80.333
R21519 a_54449_3877.n0 a_54449_3877.t0 17.4
R21520 a_54449_3877.n0 a_54449_3877.t4 17.4
R21521 a_54449_3877.n4 a_54449_3877.t2 15.032
R21522 a_54449_3877.t1 a_54449_3877.n5 14.282
R21523 a_54449_3877.n5 a_54449_3877.t3 14.282
R21524 a_54449_3877.n5 a_54449_3877.n4 1.65
R21525 a_54449_3877.n3 a_54449_3877.n0 0.672
R21526 a_54449_3877.n4 a_54449_3877.n3 0.665
R21527 a_54567_3877.n0 a_54567_3877.t3 14.282
R21528 a_54567_3877.n0 a_54567_3877.t5 14.282
R21529 a_54567_3877.n1 a_54567_3877.t0 14.282
R21530 a_54567_3877.n1 a_54567_3877.t1 14.282
R21531 a_54567_3877.t2 a_54567_3877.n3 14.282
R21532 a_54567_3877.n3 a_54567_3877.t4 14.282
R21533 a_54567_3877.n2 a_54567_3877.n0 2.546
R21534 a_54567_3877.n2 a_54567_3877.n1 2.367
R21535 a_54567_3877.n3 a_54567_3877.n2 0.001
R21536 a_61079_9746.t8 a_61079_9746.n3 404.877
R21537 a_61079_9746.n2 a_61079_9746.t7 210.902
R21538 a_61079_9746.n4 a_61079_9746.t8 136.943
R21539 a_61079_9746.n3 a_61079_9746.n2 107.801
R21540 a_61079_9746.n2 a_61079_9746.t5 80.333
R21541 a_61079_9746.n3 a_61079_9746.t6 80.333
R21542 a_61079_9746.n1 a_61079_9746.t4 17.4
R21543 a_61079_9746.n1 a_61079_9746.t0 17.4
R21544 a_61079_9746.t3 a_61079_9746.n5 15.032
R21545 a_61079_9746.n0 a_61079_9746.t2 14.282
R21546 a_61079_9746.n0 a_61079_9746.t1 14.282
R21547 a_61079_9746.n5 a_61079_9746.n0 1.65
R21548 a_61079_9746.n4 a_61079_9746.n1 0.672
R21549 a_61079_9746.n5 a_61079_9746.n4 0.665
R21550 a_16046_n2152.n3 a_16046_n2152.t6 448.382
R21551 a_16046_n2152.n2 a_16046_n2152.t5 286.438
R21552 a_16046_n2152.n2 a_16046_n2152.t7 286.438
R21553 a_16046_n2152.n1 a_16046_n2152.t4 247.69
R21554 a_16046_n2152.n4 a_16046_n2152.n0 182.117
R21555 a_16046_n2152.t6 a_16046_n2152.n2 160.666
R21556 a_16046_n2152.t2 a_16046_n2152.n4 28.568
R21557 a_16046_n2152.n0 a_16046_n2152.t0 28.565
R21558 a_16046_n2152.n0 a_16046_n2152.t1 28.565
R21559 a_16046_n2152.n1 a_16046_n2152.t3 18.127
R21560 a_16046_n2152.n3 a_16046_n2152.n1 4.039
R21561 a_16046_n2152.n4 a_16046_n2152.n3 0.937
R21562 a_40219_3874.n0 a_40219_3874.t5 14.282
R21563 a_40219_3874.n0 a_40219_3874.t0 14.282
R21564 a_40219_3874.n1 a_40219_3874.t4 14.282
R21565 a_40219_3874.n1 a_40219_3874.t3 14.282
R21566 a_40219_3874.t2 a_40219_3874.n3 14.282
R21567 a_40219_3874.n3 a_40219_3874.t1 14.282
R21568 a_40219_3874.n3 a_40219_3874.n2 2.546
R21569 a_40219_3874.n2 a_40219_3874.n1 2.367
R21570 a_40219_3874.n2 a_40219_3874.n0 0.001
R21571 a_6735_21596.n2 a_6735_21596.n1 167.433
R21572 a_6735_21596.n6 a_6735_21596.n5 167.433
R21573 a_6735_21596.n2 a_6735_21596.t10 104.259
R21574 a_6735_21596.n6 a_6735_21596.t8 104.259
R21575 a_6735_21596.n3 a_6735_21596.n0 89.977
R21576 a_6735_21596.n7 a_6735_21596.n4 89.977
R21577 a_6735_21596.n9 a_6735_21596.n8 89.977
R21578 a_6735_21596.n7 a_6735_21596.n6 77.784
R21579 a_6735_21596.n8 a_6735_21596.n3 77.456
R21580 a_6735_21596.n8 a_6735_21596.n7 77.456
R21581 a_6735_21596.n3 a_6735_21596.n2 75.815
R21582 a_6735_21596.n1 a_6735_21596.t9 14.282
R21583 a_6735_21596.n1 a_6735_21596.t11 14.282
R21584 a_6735_21596.n0 a_6735_21596.t0 14.282
R21585 a_6735_21596.n0 a_6735_21596.t1 14.282
R21586 a_6735_21596.n4 a_6735_21596.t4 14.282
R21587 a_6735_21596.n4 a_6735_21596.t5 14.282
R21588 a_6735_21596.n5 a_6735_21596.t6 14.282
R21589 a_6735_21596.n5 a_6735_21596.t7 14.282
R21590 a_6735_21596.t2 a_6735_21596.n9 14.282
R21591 a_6735_21596.n9 a_6735_21596.t3 14.282
R21592 a_13358_6047.n1 a_13358_6047.t5 318.922
R21593 a_13358_6047.n0 a_13358_6047.t4 274.739
R21594 a_13358_6047.n0 a_13358_6047.t7 274.739
R21595 a_13358_6047.n1 a_13358_6047.t6 269.116
R21596 a_13358_6047.t5 a_13358_6047.n0 179.946
R21597 a_13358_6047.n2 a_13358_6047.n1 107.263
R21598 a_13358_6047.n3 a_13358_6047.t0 29.444
R21599 a_13358_6047.t2 a_13358_6047.n4 28.565
R21600 a_13358_6047.n4 a_13358_6047.t1 28.565
R21601 a_13358_6047.n2 a_13358_6047.t3 18.145
R21602 a_13358_6047.n3 a_13358_6047.n2 2.878
R21603 a_13358_6047.n4 a_13358_6047.n3 0.764
R21604 a_50316_21344.n1 a_50316_21344.t5 318.922
R21605 a_50316_21344.n0 a_50316_21344.t4 274.739
R21606 a_50316_21344.n0 a_50316_21344.t6 274.739
R21607 a_50316_21344.n1 a_50316_21344.t7 269.116
R21608 a_50316_21344.t5 a_50316_21344.n0 179.946
R21609 a_50316_21344.n2 a_50316_21344.n1 105.178
R21610 a_50316_21344.t2 a_50316_21344.n4 29.444
R21611 a_50316_21344.n3 a_50316_21344.t0 28.565
R21612 a_50316_21344.n3 a_50316_21344.t1 28.565
R21613 a_50316_21344.n2 a_50316_21344.t3 18.145
R21614 a_50316_21344.n4 a_50316_21344.n2 2.878
R21615 a_50316_21344.n4 a_50316_21344.n3 0.764
R21616 a_6524_1744.n2 a_6524_1744.t7 448.382
R21617 a_6524_1744.n1 a_6524_1744.t6 286.438
R21618 a_6524_1744.n1 a_6524_1744.t4 286.438
R21619 a_6524_1744.n0 a_6524_1744.t5 247.69
R21620 a_6524_1744.n4 a_6524_1744.n3 182.117
R21621 a_6524_1744.t7 a_6524_1744.n1 160.666
R21622 a_6524_1744.n3 a_6524_1744.t1 28.568
R21623 a_6524_1744.t2 a_6524_1744.n4 28.565
R21624 a_6524_1744.n4 a_6524_1744.t0 28.565
R21625 a_6524_1744.n0 a_6524_1744.t3 18.127
R21626 a_6524_1744.n2 a_6524_1744.n0 4.039
R21627 a_6524_1744.n3 a_6524_1744.n2 0.937
R21628 a_57981_7583.t0 a_57981_7583.t1 17.4
R21629 a_71846_8013.t0 a_71846_8013.t1 17.4
R21630 a_7365_11720.n0 a_7365_11720.t8 14.282
R21631 a_7365_11720.t6 a_7365_11720.n0 14.282
R21632 a_7365_11720.n0 a_7365_11720.n9 89.977
R21633 a_7365_11720.n6 a_7365_11720.n7 77.784
R21634 a_7365_11720.n4 a_7365_11720.n6 77.456
R21635 a_7365_11720.n9 a_7365_11720.n4 77.456
R21636 a_7365_11720.n9 a_7365_11720.n2 75.815
R21637 a_7365_11720.n7 a_7365_11720.n8 167.433
R21638 a_7365_11720.n8 a_7365_11720.t5 14.282
R21639 a_7365_11720.n8 a_7365_11720.t4 14.282
R21640 a_7365_11720.n7 a_7365_11720.t3 104.259
R21641 a_7365_11720.n6 a_7365_11720.n5 89.977
R21642 a_7365_11720.n5 a_7365_11720.t11 14.282
R21643 a_7365_11720.n5 a_7365_11720.t10 14.282
R21644 a_7365_11720.n4 a_7365_11720.n3 89.977
R21645 a_7365_11720.n3 a_7365_11720.t9 14.282
R21646 a_7365_11720.n3 a_7365_11720.t7 14.282
R21647 a_7365_11720.n2 a_7365_11720.t2 104.259
R21648 a_7365_11720.n2 a_7365_11720.n1 167.433
R21649 a_7365_11720.n1 a_7365_11720.t1 14.282
R21650 a_7365_11720.n1 a_7365_11720.t0 14.282
R21651 a_39720_22683.n0 a_39720_22683.t9 214.335
R21652 a_39720_22683.t7 a_39720_22683.n0 214.335
R21653 a_39720_22683.n1 a_39720_22683.t7 143.851
R21654 a_39720_22683.n1 a_39720_22683.t10 135.658
R21655 a_39720_22683.n0 a_39720_22683.t8 80.333
R21656 a_39720_22683.n2 a_39720_22683.t4 28.565
R21657 a_39720_22683.n2 a_39720_22683.t5 28.565
R21658 a_39720_22683.n4 a_39720_22683.t6 28.565
R21659 a_39720_22683.n4 a_39720_22683.t1 28.565
R21660 a_39720_22683.t2 a_39720_22683.n7 28.565
R21661 a_39720_22683.n7 a_39720_22683.t0 28.565
R21662 a_39720_22683.n6 a_39720_22683.t3 9.714
R21663 a_39720_22683.n7 a_39720_22683.n6 1.003
R21664 a_39720_22683.n5 a_39720_22683.n3 0.833
R21665 a_39720_22683.n3 a_39720_22683.n2 0.653
R21666 a_39720_22683.n5 a_39720_22683.n4 0.653
R21667 a_39720_22683.n6 a_39720_22683.n5 0.341
R21668 a_39720_22683.n3 a_39720_22683.n1 0.032
R21669 a_4889_8119.n3 a_4889_8119.t7 448.381
R21670 a_4889_8119.n2 a_4889_8119.t4 286.438
R21671 a_4889_8119.n2 a_4889_8119.t6 286.438
R21672 a_4889_8119.n1 a_4889_8119.t5 247.69
R21673 a_4889_8119.n4 a_4889_8119.n0 182.117
R21674 a_4889_8119.t7 a_4889_8119.n2 160.666
R21675 a_4889_8119.t2 a_4889_8119.n4 28.568
R21676 a_4889_8119.n0 a_4889_8119.t0 28.565
R21677 a_4889_8119.n0 a_4889_8119.t1 28.565
R21678 a_4889_8119.n1 a_4889_8119.t3 18.127
R21679 a_4889_8119.n3 a_4889_8119.n1 4.036
R21680 a_4889_8119.n4 a_4889_8119.n3 0.937
R21681 a_16573_1740.n0 a_16573_1740.n9 167.433
R21682 a_16573_1740.n0 a_16573_1740.t1 14.282
R21683 a_16573_1740.t0 a_16573_1740.n0 14.282
R21684 a_16573_1740.n9 a_16573_1740.n8 75.815
R21685 a_16573_1740.n8 a_16573_1740.n6 77.456
R21686 a_16573_1740.n6 a_16573_1740.n4 77.456
R21687 a_16573_1740.n4 a_16573_1740.n2 77.784
R21688 a_16573_1740.n9 a_16573_1740.t2 104.259
R21689 a_16573_1740.n8 a_16573_1740.n7 89.977
R21690 a_16573_1740.n7 a_16573_1740.t11 14.282
R21691 a_16573_1740.n7 a_16573_1740.t9 14.282
R21692 a_16573_1740.n6 a_16573_1740.n5 89.977
R21693 a_16573_1740.n5 a_16573_1740.t10 14.282
R21694 a_16573_1740.n5 a_16573_1740.t8 14.282
R21695 a_16573_1740.n4 a_16573_1740.n3 89.977
R21696 a_16573_1740.n3 a_16573_1740.t6 14.282
R21697 a_16573_1740.n3 a_16573_1740.t7 14.282
R21698 a_16573_1740.n2 a_16573_1740.t5 104.259
R21699 a_16573_1740.n2 a_16573_1740.n1 167.433
R21700 a_16573_1740.n1 a_16573_1740.t4 14.282
R21701 a_16573_1740.n1 a_16573_1740.t3 14.282
R21702 a_16922_1740.n2 a_16922_1740.t8 1527.4
R21703 a_16922_1740.t8 a_16922_1740.n1 657.379
R21704 a_16922_1740.n4 a_16922_1740.n3 258.161
R21705 a_16922_1740.n7 a_16922_1740.n6 258.161
R21706 a_16922_1740.n0 a_16922_1740.t11 206.421
R21707 a_16922_1740.t10 a_16922_1740.n0 206.421
R21708 a_16922_1740.n2 a_16922_1740.t10 200.029
R21709 a_16922_1740.n5 a_16922_1740.n2 97.614
R21710 a_16922_1740.n0 a_16922_1740.t9 80.333
R21711 a_16922_1740.n4 a_16922_1740.t6 14.283
R21712 a_16922_1740.n6 a_16922_1740.t0 14.283
R21713 a_16922_1740.n3 a_16922_1740.t5 14.282
R21714 a_16922_1740.n3 a_16922_1740.t7 14.282
R21715 a_16922_1740.n7 a_16922_1740.t1 14.282
R21716 a_16922_1740.t2 a_16922_1740.n7 14.282
R21717 a_16922_1740.n1 a_16922_1740.t4 8.7
R21718 a_16922_1740.n1 a_16922_1740.t3 8.7
R21719 a_16922_1740.n5 a_16922_1740.n4 4.366
R21720 a_16922_1740.n6 a_16922_1740.n5 0.852
R21721 a_59325_22679.n2 a_59325_22679.t7 214.335
R21722 a_59325_22679.t9 a_59325_22679.n2 214.335
R21723 a_59325_22679.n3 a_59325_22679.t9 143.851
R21724 a_59325_22679.n3 a_59325_22679.t8 135.658
R21725 a_59325_22679.n2 a_59325_22679.t10 80.333
R21726 a_59325_22679.n4 a_59325_22679.t0 28.565
R21727 a_59325_22679.n4 a_59325_22679.t1 28.565
R21728 a_59325_22679.n0 a_59325_22679.t5 28.565
R21729 a_59325_22679.n0 a_59325_22679.t6 28.565
R21730 a_59325_22679.t2 a_59325_22679.n7 28.565
R21731 a_59325_22679.n7 a_59325_22679.t4 28.565
R21732 a_59325_22679.n1 a_59325_22679.t3 9.714
R21733 a_59325_22679.n1 a_59325_22679.n0 1.003
R21734 a_59325_22679.n6 a_59325_22679.n5 0.833
R21735 a_59325_22679.n5 a_59325_22679.n4 0.653
R21736 a_59325_22679.n7 a_59325_22679.n6 0.653
R21737 a_59325_22679.n6 a_59325_22679.n1 0.341
R21738 a_59325_22679.n5 a_59325_22679.n3 0.032
R21739 a_4834_7659.t0 a_4834_7659.t1 17.4
R21740 a_40373_9071.t5 a_40373_9071.t6 800.071
R21741 a_40373_9071.n3 a_40373_9071.n2 672.951
R21742 a_40373_9071.n1 a_40373_9071.t7 285.109
R21743 a_40373_9071.n2 a_40373_9071.t5 193.602
R21744 a_40373_9071.n1 a_40373_9071.t4 160.666
R21745 a_40373_9071.n2 a_40373_9071.n1 91.507
R21746 a_40373_9071.t2 a_40373_9071.n4 28.57
R21747 a_40373_9071.n0 a_40373_9071.t1 28.565
R21748 a_40373_9071.n0 a_40373_9071.t0 28.565
R21749 a_40373_9071.n4 a_40373_9071.t3 17.638
R21750 a_40373_9071.n3 a_40373_9071.n0 0.69
R21751 a_40373_9071.n4 a_40373_9071.n3 0.6
R21752 a_66005_5881.t0 a_66005_5881.t1 17.4
R21753 a_13178_10994.t5 a_13178_10994.n0 14.283
R21754 a_13178_10994.n0 a_13178_10994.n5 0.852
R21755 a_13178_10994.n5 a_13178_10994.n6 4.366
R21756 a_13178_10994.n6 a_13178_10994.n7 258.161
R21757 a_13178_10994.n7 a_13178_10994.t1 14.282
R21758 a_13178_10994.n7 a_13178_10994.t0 14.282
R21759 a_13178_10994.n6 a_13178_10994.t2 14.283
R21760 a_13178_10994.n5 a_13178_10994.n4 97.614
R21761 a_13178_10994.n4 a_13178_10994.t8 200.029
R21762 a_13178_10994.t8 a_13178_10994.n3 206.421
R21763 a_13178_10994.n3 a_13178_10994.t9 80.333
R21764 a_13178_10994.n3 a_13178_10994.t11 206.421
R21765 a_13178_10994.n4 a_13178_10994.t10 1527.4
R21766 a_13178_10994.t10 a_13178_10994.n2 657.379
R21767 a_13178_10994.n2 a_13178_10994.t3 8.7
R21768 a_13178_10994.n2 a_13178_10994.t4 8.7
R21769 a_13178_10994.n0 a_13178_10994.n1 258.161
R21770 a_13178_10994.n1 a_13178_10994.t6 14.282
R21771 a_13178_10994.n1 a_13178_10994.t7 14.282
R21772 a_48426_24202.t5 a_48426_24202.n3 404.877
R21773 a_48426_24202.n2 a_48426_24202.t8 210.902
R21774 a_48426_24202.n4 a_48426_24202.t5 136.943
R21775 a_48426_24202.n3 a_48426_24202.n2 107.801
R21776 a_48426_24202.n2 a_48426_24202.t6 80.333
R21777 a_48426_24202.n3 a_48426_24202.t7 80.333
R21778 a_48426_24202.n1 a_48426_24202.t4 17.4
R21779 a_48426_24202.n1 a_48426_24202.t3 17.4
R21780 a_48426_24202.t0 a_48426_24202.n5 15.032
R21781 a_48426_24202.n0 a_48426_24202.t1 14.282
R21782 a_48426_24202.n0 a_48426_24202.t2 14.282
R21783 a_48426_24202.n5 a_48426_24202.n0 1.65
R21784 a_48426_24202.n4 a_48426_24202.n1 0.672
R21785 a_48426_24202.n5 a_48426_24202.n4 0.665
R21786 a_14538_10391.t0 a_14538_10391.t1 17.4
R21787 a_48484_308.t0 a_48484_308.t1 17.4
R21788 a_41573_15739.n1 a_41573_15739.t7 318.922
R21789 a_41573_15739.n0 a_41573_15739.t6 273.935
R21790 a_41573_15739.n0 a_41573_15739.t5 273.935
R21791 a_41573_15739.n1 a_41573_15739.t4 269.116
R21792 a_41573_15739.n4 a_41573_15739.n3 193.227
R21793 a_41573_15739.t7 a_41573_15739.n0 179.142
R21794 a_41573_15739.n2 a_41573_15739.n1 106.999
R21795 a_41573_15739.n3 a_41573_15739.t0 28.568
R21796 a_41573_15739.n4 a_41573_15739.t1 28.565
R21797 a_41573_15739.t2 a_41573_15739.n4 28.565
R21798 a_41573_15739.n2 a_41573_15739.t3 18.149
R21799 a_41573_15739.n3 a_41573_15739.n2 3.726
R21800 a_48265_n1750.n0 a_48265_n1750.t9 214.335
R21801 a_48265_n1750.t8 a_48265_n1750.n0 214.335
R21802 a_48265_n1750.n1 a_48265_n1750.t8 143.85
R21803 a_48265_n1750.n1 a_48265_n1750.t10 135.66
R21804 a_48265_n1750.n0 a_48265_n1750.t7 80.333
R21805 a_48265_n1750.n2 a_48265_n1750.t4 28.565
R21806 a_48265_n1750.n2 a_48265_n1750.t5 28.565
R21807 a_48265_n1750.n4 a_48265_n1750.t6 28.565
R21808 a_48265_n1750.n4 a_48265_n1750.t0 28.565
R21809 a_48265_n1750.n7 a_48265_n1750.t1 28.565
R21810 a_48265_n1750.t2 a_48265_n1750.n7 28.565
R21811 a_48265_n1750.n6 a_48265_n1750.t3 9.714
R21812 a_48265_n1750.n7 a_48265_n1750.n6 1.003
R21813 a_48265_n1750.n5 a_48265_n1750.n3 0.836
R21814 a_48265_n1750.n5 a_48265_n1750.n4 0.653
R21815 a_48265_n1750.n3 a_48265_n1750.n2 0.65
R21816 a_48265_n1750.n6 a_48265_n1750.n5 0.341
R21817 a_48265_n1750.n3 a_48265_n1750.n1 0.032
R21818 a_41243_3878.t5 a_41243_3878.n2 404.877
R21819 a_41243_3878.n1 a_41243_3878.t7 210.902
R21820 a_41243_3878.n3 a_41243_3878.t5 136.943
R21821 a_41243_3878.n2 a_41243_3878.n1 107.801
R21822 a_41243_3878.n1 a_41243_3878.t8 80.333
R21823 a_41243_3878.n2 a_41243_3878.t6 80.333
R21824 a_41243_3878.n0 a_41243_3878.t0 17.4
R21825 a_41243_3878.n0 a_41243_3878.t4 17.4
R21826 a_41243_3878.n4 a_41243_3878.t3 15.032
R21827 a_41243_3878.n5 a_41243_3878.t2 14.282
R21828 a_41243_3878.t1 a_41243_3878.n5 14.282
R21829 a_41243_3878.n5 a_41243_3878.n4 1.65
R21830 a_41243_3878.n3 a_41243_3878.n0 0.672
R21831 a_41243_3878.n4 a_41243_3878.n3 0.665
R21832 a_47357_18567.t7 a_47357_18567.t5 800.071
R21833 a_47357_18567.n3 a_47357_18567.n2 659.095
R21834 a_47357_18567.n1 a_47357_18567.t4 285.109
R21835 a_47357_18567.n2 a_47357_18567.t7 193.602
R21836 a_47357_18567.n4 a_47357_18567.n0 192.754
R21837 a_47357_18567.n1 a_47357_18567.t6 160.666
R21838 a_47357_18567.n2 a_47357_18567.n1 91.507
R21839 a_47357_18567.t2 a_47357_18567.n4 28.568
R21840 a_47357_18567.n0 a_47357_18567.t0 28.565
R21841 a_47357_18567.n0 a_47357_18567.t1 28.565
R21842 a_47357_18567.n3 a_47357_18567.t3 19.063
R21843 a_47357_18567.n4 a_47357_18567.n3 1.005
R21844 a_47417_18593.n1 a_47417_18593.t5 14.282
R21845 a_47417_18593.n1 a_47417_18593.t0 14.282
R21846 a_47417_18593.n0 a_47417_18593.t3 14.282
R21847 a_47417_18593.n0 a_47417_18593.t4 14.282
R21848 a_47417_18593.n3 a_47417_18593.t1 14.282
R21849 a_47417_18593.t2 a_47417_18593.n3 14.282
R21850 a_47417_18593.n2 a_47417_18593.n0 2.546
R21851 a_47417_18593.n3 a_47417_18593.n2 2.367
R21852 a_47417_18593.n2 a_47417_18593.n1 0.001
R21853 a_52809_18602.n0 a_52809_18602.t0 14.282
R21854 a_52809_18602.n0 a_52809_18602.t1 14.282
R21855 a_52809_18602.n1 a_52809_18602.t4 14.282
R21856 a_52809_18602.n1 a_52809_18602.t5 14.282
R21857 a_52809_18602.t2 a_52809_18602.n3 14.282
R21858 a_52809_18602.n3 a_52809_18602.t3 14.282
R21859 a_52809_18602.n2 a_52809_18602.n0 2.546
R21860 a_52809_18602.n2 a_52809_18602.n1 2.367
R21861 a_52809_18602.n3 a_52809_18602.n2 0.001
R21862 a_48225_11948.n2 a_48225_11948.t7 214.335
R21863 a_48225_11948.t9 a_48225_11948.n2 214.335
R21864 a_48225_11948.n3 a_48225_11948.t9 143.851
R21865 a_48225_11948.n3 a_48225_11948.t8 135.658
R21866 a_48225_11948.n2 a_48225_11948.t10 80.333
R21867 a_48225_11948.n4 a_48225_11948.t0 28.565
R21868 a_48225_11948.n4 a_48225_11948.t1 28.565
R21869 a_48225_11948.n0 a_48225_11948.t4 28.565
R21870 a_48225_11948.n0 a_48225_11948.t5 28.565
R21871 a_48225_11948.t2 a_48225_11948.n7 28.565
R21872 a_48225_11948.n7 a_48225_11948.t6 28.565
R21873 a_48225_11948.n1 a_48225_11948.t3 9.714
R21874 a_48225_11948.n1 a_48225_11948.n0 1.003
R21875 a_48225_11948.n6 a_48225_11948.n5 0.833
R21876 a_48225_11948.n5 a_48225_11948.n4 0.653
R21877 a_48225_11948.n7 a_48225_11948.n6 0.653
R21878 a_48225_11948.n6 a_48225_11948.n1 0.341
R21879 a_48225_11948.n5 a_48225_11948.n3 0.032
R21880 a_12672_15792.t6 a_12672_15792.n2 406.221
R21881 a_12672_15792.n1 a_12672_15792.t7 191.682
R21882 a_12672_15792.n3 a_12672_15792.t6 138.556
R21883 a_12672_15792.n2 a_12672_15792.n1 111.349
R21884 a_12672_15792.n1 a_12672_15792.t8 80.333
R21885 a_12672_15792.n2 a_12672_15792.t5 80.333
R21886 a_12672_15792.n0 a_12672_15792.t4 17.4
R21887 a_12672_15792.n0 a_12672_15792.t0 17.4
R21888 a_12672_15792.n4 a_12672_15792.t1 15.036
R21889 a_12672_15792.n5 a_12672_15792.t2 14.282
R21890 a_12672_15792.t3 a_12672_15792.n5 14.282
R21891 a_12672_15792.n5 a_12672_15792.n4 1.654
R21892 a_12672_15792.n3 a_12672_15792.n0 0.664
R21893 a_12672_15792.n4 a_12672_15792.n3 0.614
R21894 a_19396_14454.n2 a_19396_14454.t6 867.497
R21895 a_19396_14454.n2 a_19396_14454.t4 591.811
R21896 a_19396_14454.n1 a_19396_14454.t5 286.438
R21897 a_19396_14454.n1 a_19396_14454.t7 286.438
R21898 a_19396_14454.n4 a_19396_14454.n0 185.55
R21899 a_19396_14454.t6 a_19396_14454.n1 160.666
R21900 a_19396_14454.t2 a_19396_14454.n4 28.568
R21901 a_19396_14454.n0 a_19396_14454.t0 28.565
R21902 a_19396_14454.n0 a_19396_14454.t1 28.565
R21903 a_19396_14454.n3 a_19396_14454.n2 26.014
R21904 a_19396_14454.n3 a_19396_14454.t3 21.376
R21905 a_19396_14454.n4 a_19396_14454.n3 1.637
R21906 a_20578_10387.t0 a_20578_10387.t1 17.4
R21907 a_51704_6111.t7 a_51704_6111.t4 574.43
R21908 a_51704_6111.n0 a_51704_6111.t6 285.109
R21909 a_51704_6111.n2 a_51704_6111.n1 197.217
R21910 a_51704_6111.n4 a_51704_6111.n3 192.754
R21911 a_51704_6111.n0 a_51704_6111.t5 160.666
R21912 a_51704_6111.n1 a_51704_6111.t7 160.666
R21913 a_51704_6111.n1 a_51704_6111.n0 114.829
R21914 a_51704_6111.n3 a_51704_6111.t0 28.568
R21915 a_51704_6111.t2 a_51704_6111.n4 28.565
R21916 a_51704_6111.n4 a_51704_6111.t1 28.565
R21917 a_51704_6111.n2 a_51704_6111.t3 18.838
R21918 a_51704_6111.n3 a_51704_6111.n2 1.129
R21919 a_19987_11720.t0 a_19987_11720.n9 104.259
R21920 a_19987_11720.n6 a_19987_11720.n7 77.784
R21921 a_19987_11720.n4 a_19987_11720.n6 77.456
R21922 a_19987_11720.n2 a_19987_11720.n4 77.456
R21923 a_19987_11720.n9 a_19987_11720.n2 75.815
R21924 a_19987_11720.n7 a_19987_11720.n8 167.433
R21925 a_19987_11720.n8 a_19987_11720.t8 14.282
R21926 a_19987_11720.n8 a_19987_11720.t7 14.282
R21927 a_19987_11720.n7 a_19987_11720.t6 104.259
R21928 a_19987_11720.n6 a_19987_11720.n5 89.977
R21929 a_19987_11720.n5 a_19987_11720.t9 14.282
R21930 a_19987_11720.n5 a_19987_11720.t11 14.282
R21931 a_19987_11720.n4 a_19987_11720.n3 89.977
R21932 a_19987_11720.n3 a_19987_11720.t10 14.282
R21933 a_19987_11720.n3 a_19987_11720.t3 14.282
R21934 a_19987_11720.n2 a_19987_11720.n1 89.977
R21935 a_19987_11720.n1 a_19987_11720.t4 14.282
R21936 a_19987_11720.n1 a_19987_11720.t5 14.282
R21937 a_19987_11720.n9 a_19987_11720.n0 167.433
R21938 a_19987_11720.n0 a_19987_11720.t1 14.282
R21939 a_19987_11720.n0 a_19987_11720.t2 14.282
R21940 a_60884_15037.t0 a_60884_15037.t1 380.209
R21941 a_20558_n3481.t0 a_20558_n3481.t1 17.4
R21942 a_40310_22246.t4 a_40310_22246.t6 574.43
R21943 a_40310_22246.n0 a_40310_22246.t7 285.109
R21944 a_40310_22246.n2 a_40310_22246.n1 211.136
R21945 a_40310_22246.n4 a_40310_22246.n3 192.754
R21946 a_40310_22246.n0 a_40310_22246.t5 160.666
R21947 a_40310_22246.n1 a_40310_22246.t4 160.666
R21948 a_40310_22246.n1 a_40310_22246.n0 114.829
R21949 a_40310_22246.n3 a_40310_22246.t0 28.568
R21950 a_40310_22246.n4 a_40310_22246.t1 28.565
R21951 a_40310_22246.t2 a_40310_22246.n4 28.565
R21952 a_40310_22246.n2 a_40310_22246.t3 19.084
R21953 a_40310_22246.n3 a_40310_22246.n2 1.051
R21954 a_59915_22242.t4 a_59915_22242.t7 574.43
R21955 a_59915_22242.n1 a_59915_22242.t6 285.109
R21956 a_59915_22242.n3 a_59915_22242.n2 211.136
R21957 a_59915_22242.n4 a_59915_22242.n0 192.754
R21958 a_59915_22242.n1 a_59915_22242.t5 160.666
R21959 a_59915_22242.n2 a_59915_22242.t4 160.666
R21960 a_59915_22242.n2 a_59915_22242.n1 114.829
R21961 a_59915_22242.t2 a_59915_22242.n4 28.568
R21962 a_59915_22242.n0 a_59915_22242.t0 28.565
R21963 a_59915_22242.n0 a_59915_22242.t1 28.565
R21964 a_59915_22242.n3 a_59915_22242.t3 19.084
R21965 a_59915_22242.n4 a_59915_22242.n3 1.051
R21966 a_39957_22046.t0 a_39957_22046.t1 17.4
R21967 a_71842_n1407.t0 a_71842_n1407.t1 17.4
R21968 a_71842_1973.t0 a_71842_1973.t1 17.4
R21969 a_7700_n3481.t0 a_7700_n3481.t1 17.4
R21970 a_38140_111.t0 a_38140_111.t1 17.4
R21971 a_59562_22042.t0 a_59562_22042.t1 17.4
R21972 a_56511_18089.t0 a_56511_18089.t1 17.4
R21973 a_17501_13585.n2 a_17501_13585.t6 448.381
R21974 a_17501_13585.n1 a_17501_13585.t5 286.438
R21975 a_17501_13585.n1 a_17501_13585.t4 286.438
R21976 a_17501_13585.n0 a_17501_13585.t7 247.69
R21977 a_17501_13585.n4 a_17501_13585.n3 182.117
R21978 a_17501_13585.t6 a_17501_13585.n1 160.666
R21979 a_17501_13585.n3 a_17501_13585.t0 28.568
R21980 a_17501_13585.n4 a_17501_13585.t1 28.565
R21981 a_17501_13585.t2 a_17501_13585.n4 28.565
R21982 a_17501_13585.n0 a_17501_13585.t3 18.127
R21983 a_17501_13585.n2 a_17501_13585.n0 4.036
R21984 a_17501_13585.n3 a_17501_13585.n2 0.937
R21985 a_16855_14458.t0 a_16855_14458.n0 14.282
R21986 a_16855_14458.n0 a_16855_14458.t1 14.282
R21987 a_16855_14458.n7 a_16855_14458.n8 77.784
R21988 a_16855_14458.n5 a_16855_14458.n7 77.456
R21989 a_16855_14458.n3 a_16855_14458.n5 77.456
R21990 a_16855_14458.n1 a_16855_14458.n3 75.815
R21991 a_16855_14458.n0 a_16855_14458.n1 167.433
R21992 a_16855_14458.n8 a_16855_14458.n9 167.433
R21993 a_16855_14458.n9 a_16855_14458.t6 14.282
R21994 a_16855_14458.n9 a_16855_14458.t8 14.282
R21995 a_16855_14458.n8 a_16855_14458.t7 104.259
R21996 a_16855_14458.n7 a_16855_14458.n6 89.977
R21997 a_16855_14458.n6 a_16855_14458.t5 14.282
R21998 a_16855_14458.n6 a_16855_14458.t4 14.282
R21999 a_16855_14458.n5 a_16855_14458.n4 89.977
R22000 a_16855_14458.n4 a_16855_14458.t3 14.282
R22001 a_16855_14458.n4 a_16855_14458.t10 14.282
R22002 a_16855_14458.n3 a_16855_14458.n2 89.977
R22003 a_16855_14458.n2 a_16855_14458.t9 14.282
R22004 a_16855_14458.n2 a_16855_14458.t11 14.282
R22005 a_16855_14458.n1 a_16855_14458.t2 104.259
R22006 a_16322_13728.t1 a_16322_13728.n0 14.283
R22007 a_16322_13728.n0 a_16322_13728.n5 0.852
R22008 a_16322_13728.n5 a_16322_13728.n6 4.366
R22009 a_16322_13728.n6 a_16322_13728.n7 258.161
R22010 a_16322_13728.n7 a_16322_13728.t5 14.282
R22011 a_16322_13728.n7 a_16322_13728.t4 14.282
R22012 a_16322_13728.n6 a_16322_13728.t6 14.283
R22013 a_16322_13728.n5 a_16322_13728.n4 97.614
R22014 a_16322_13728.n4 a_16322_13728.t8 200.029
R22015 a_16322_13728.t8 a_16322_13728.n3 206.421
R22016 a_16322_13728.n3 a_16322_13728.t9 80.333
R22017 a_16322_13728.n3 a_16322_13728.t10 206.421
R22018 a_16322_13728.n4 a_16322_13728.t11 1527.4
R22019 a_16322_13728.t11 a_16322_13728.n2 657.379
R22020 a_16322_13728.n2 a_16322_13728.t7 8.7
R22021 a_16322_13728.n2 a_16322_13728.t0 8.7
R22022 a_16322_13728.n0 a_16322_13728.n1 258.161
R22023 a_16322_13728.n1 a_16322_13728.t3 14.282
R22024 a_16322_13728.n1 a_16322_13728.t2 14.282
R22025 a_71842_11215.t0 a_71842_11215.t1 17.4
R22026 a_70509_10506.n0 a_70509_10506.t6 14.282
R22027 a_70509_10506.t4 a_70509_10506.n0 14.282
R22028 a_70509_10506.n0 a_70509_10506.n1 258.161
R22029 a_70509_10506.n1 a_70509_10506.t5 14.283
R22030 a_70509_10506.n1 a_70509_10506.n5 0.852
R22031 a_70509_10506.n5 a_70509_10506.n6 4.366
R22032 a_70509_10506.n6 a_70509_10506.n7 258.161
R22033 a_70509_10506.n7 a_70509_10506.t1 14.282
R22034 a_70509_10506.n7 a_70509_10506.t2 14.282
R22035 a_70509_10506.n6 a_70509_10506.t0 14.283
R22036 a_70509_10506.n5 a_70509_10506.n4 73.514
R22037 a_70509_10506.n4 a_70509_10506.t11 1551.5
R22038 a_70509_10506.t11 a_70509_10506.n3 656.576
R22039 a_70509_10506.n3 a_70509_10506.t3 8.7
R22040 a_70509_10506.n3 a_70509_10506.t7 8.7
R22041 a_70509_10506.n4 a_70509_10506.t9 224.129
R22042 a_70509_10506.t9 a_70509_10506.n2 207.225
R22043 a_70509_10506.n2 a_70509_10506.t10 207.225
R22044 a_70509_10506.n2 a_70509_10506.t8 80.333
R22045 a_56556_20633.t0 a_56556_20633.t1 380.209
R22046 a_56556_21365.n0 a_56556_21365.n8 122.999
R22047 a_56556_21365.n0 a_56556_21365.t2 14.282
R22048 a_56556_21365.t1 a_56556_21365.n0 14.282
R22049 a_56556_21365.n8 a_56556_21365.n6 50.575
R22050 a_56556_21365.n6 a_56556_21365.n4 74.302
R22051 a_56556_21365.n8 a_56556_21365.n7 157.665
R22052 a_56556_21365.n7 a_56556_21365.t4 8.7
R22053 a_56556_21365.n7 a_56556_21365.t0 8.7
R22054 a_56556_21365.n6 a_56556_21365.n5 90.416
R22055 a_56556_21365.n5 a_56556_21365.t3 14.282
R22056 a_56556_21365.n5 a_56556_21365.t7 14.282
R22057 a_56556_21365.n4 a_56556_21365.n3 90.436
R22058 a_56556_21365.n3 a_56556_21365.t5 14.282
R22059 a_56556_21365.n3 a_56556_21365.t6 14.282
R22060 a_56556_21365.n4 a_56556_21365.n1 1467.36
R22061 a_56556_21365.t11 a_56556_21365.n2 160.666
R22062 a_56556_21365.n1 a_56556_21365.t11 867.393
R22063 a_56556_21365.n2 a_56556_21365.t9 287.241
R22064 a_56556_21365.n2 a_56556_21365.t8 287.241
R22065 a_56556_21365.n1 a_56556_21365.t10 545.094
R22066 a_60055_9742.n1 a_60055_9742.t1 14.282
R22067 a_60055_9742.n1 a_60055_9742.t5 14.282
R22068 a_60055_9742.n0 a_60055_9742.t4 14.282
R22069 a_60055_9742.n0 a_60055_9742.t3 14.282
R22070 a_60055_9742.n3 a_60055_9742.t0 14.282
R22071 a_60055_9742.t2 a_60055_9742.n3 14.282
R22072 a_60055_9742.n2 a_60055_9742.n0 2.546
R22073 a_60055_9742.n3 a_60055_9742.n2 2.367
R22074 a_60055_9742.n2 a_60055_9742.n1 0.001
R22075 a_16264_14458.n2 a_16264_14458.t5 867.497
R22076 a_16264_14458.n2 a_16264_14458.t6 591.811
R22077 a_16264_14458.n1 a_16264_14458.t7 286.438
R22078 a_16264_14458.n1 a_16264_14458.t4 286.438
R22079 a_16264_14458.n4 a_16264_14458.n0 185.55
R22080 a_16264_14458.t5 a_16264_14458.n1 160.666
R22081 a_16264_14458.t2 a_16264_14458.n4 28.568
R22082 a_16264_14458.n0 a_16264_14458.t0 28.565
R22083 a_16264_14458.n0 a_16264_14458.t1 28.565
R22084 a_16264_14458.n3 a_16264_14458.n2 26.1
R22085 a_16264_14458.n3 a_16264_14458.t3 21.376
R22086 a_16264_14458.n4 a_16264_14458.n3 1.638
R22087 a_22540_11720.n2 a_22540_11720.t5 990.34
R22088 a_22540_11720.n2 a_22540_11720.t7 408.211
R22089 a_22540_11720.n3 a_22540_11720.n2 387.729
R22090 a_22540_11720.n1 a_22540_11720.t4 286.438
R22091 a_22540_11720.n1 a_22540_11720.t6 286.438
R22092 a_22540_11720.n4 a_22540_11720.n0 185.55
R22093 a_22540_11720.t5 a_22540_11720.n1 160.666
R22094 a_22540_11720.t2 a_22540_11720.n4 28.568
R22095 a_22540_11720.n0 a_22540_11720.t0 28.565
R22096 a_22540_11720.n0 a_22540_11720.t1 28.565
R22097 a_22540_11720.n3 a_22540_11720.t3 21.376
R22098 a_22540_11720.n4 a_22540_11720.n3 1.637
R22099 a_14538_13125.t0 a_14538_13125.t1 17.4
R22100 a_61098_21369.n0 a_61098_21369.t11 14.282
R22101 a_61098_21369.t6 a_61098_21369.n0 14.282
R22102 a_61098_21369.n0 a_61098_21369.n9 0.999
R22103 a_61098_21369.n6 a_61098_21369.n8 0.575
R22104 a_61098_21369.n9 a_61098_21369.n6 0.2
R22105 a_61098_21369.n9 a_61098_21369.t7 16.058
R22106 a_61098_21369.n8 a_61098_21369.n7 0.999
R22107 a_61098_21369.n7 a_61098_21369.t1 14.282
R22108 a_61098_21369.n7 a_61098_21369.t0 14.282
R22109 a_61098_21369.n8 a_61098_21369.t2 16.058
R22110 a_61098_21369.n6 a_61098_21369.n4 0.227
R22111 a_61098_21369.n4 a_61098_21369.n5 1.511
R22112 a_61098_21369.n5 a_61098_21369.t5 14.282
R22113 a_61098_21369.n5 a_61098_21369.t4 14.282
R22114 a_61098_21369.n4 a_61098_21369.n1 0.669
R22115 a_61098_21369.n1 a_61098_21369.n2 0.001
R22116 a_61098_21369.n1 a_61098_21369.n3 267.767
R22117 a_61098_21369.n3 a_61098_21369.t8 14.282
R22118 a_61098_21369.n3 a_61098_21369.t10 14.282
R22119 a_61098_21369.n2 a_61098_21369.t3 14.282
R22120 a_61098_21369.n2 a_61098_21369.t9 14.282
R22121 a_19737_n2148.n0 a_19737_n2148.t1 14.282
R22122 a_19737_n2148.t0 a_19737_n2148.n0 14.282
R22123 a_19737_n2148.n7 a_19737_n2148.n8 75.815
R22124 a_19737_n2148.n5 a_19737_n2148.n7 77.456
R22125 a_19737_n2148.n3 a_19737_n2148.n5 77.456
R22126 a_19737_n2148.n1 a_19737_n2148.n3 77.784
R22127 a_19737_n2148.n0 a_19737_n2148.n1 167.433
R22128 a_19737_n2148.n8 a_19737_n2148.n9 167.433
R22129 a_19737_n2148.n9 a_19737_n2148.t6 14.282
R22130 a_19737_n2148.n9 a_19737_n2148.t7 14.282
R22131 a_19737_n2148.n8 a_19737_n2148.t8 104.259
R22132 a_19737_n2148.n7 a_19737_n2148.n6 89.977
R22133 a_19737_n2148.n6 a_19737_n2148.t5 14.282
R22134 a_19737_n2148.n6 a_19737_n2148.t4 14.282
R22135 a_19737_n2148.n5 a_19737_n2148.n4 89.977
R22136 a_19737_n2148.n4 a_19737_n2148.t3 14.282
R22137 a_19737_n2148.n4 a_19737_n2148.t11 14.282
R22138 a_19737_n2148.n3 a_19737_n2148.n2 89.977
R22139 a_19737_n2148.n2 a_19737_n2148.t10 14.282
R22140 a_19737_n2148.n2 a_19737_n2148.t9 14.282
R22141 a_19737_n2148.n1 a_19737_n2148.t2 104.259
R22142 a_8011_10847.n2 a_8011_10847.t6 448.381
R22143 a_8011_10847.n1 a_8011_10847.t5 286.438
R22144 a_8011_10847.n1 a_8011_10847.t7 286.438
R22145 a_8011_10847.n0 a_8011_10847.t4 247.69
R22146 a_8011_10847.n4 a_8011_10847.n3 182.117
R22147 a_8011_10847.t6 a_8011_10847.n1 160.666
R22148 a_8011_10847.n3 a_8011_10847.t1 28.568
R22149 a_8011_10847.t2 a_8011_10847.n4 28.565
R22150 a_8011_10847.n4 a_8011_10847.t0 28.565
R22151 a_8011_10847.n0 a_8011_10847.t3 18.127
R22152 a_8011_10847.n2 a_8011_10847.n0 4.036
R22153 a_8011_10847.n3 a_8011_10847.n2 0.937
R22154 a_59320_21075.n0 a_59320_21075.t7 214.335
R22155 a_59320_21075.t8 a_59320_21075.n0 214.335
R22156 a_59320_21075.n1 a_59320_21075.t8 143.851
R22157 a_59320_21075.n1 a_59320_21075.t10 135.658
R22158 a_59320_21075.n0 a_59320_21075.t9 80.333
R22159 a_59320_21075.n2 a_59320_21075.t4 28.565
R22160 a_59320_21075.n2 a_59320_21075.t5 28.565
R22161 a_59320_21075.n4 a_59320_21075.t6 28.565
R22162 a_59320_21075.n4 a_59320_21075.t0 28.565
R22163 a_59320_21075.n7 a_59320_21075.t1 28.565
R22164 a_59320_21075.t2 a_59320_21075.n7 28.565
R22165 a_59320_21075.n6 a_59320_21075.t3 9.714
R22166 a_59320_21075.n7 a_59320_21075.n6 1.003
R22167 a_59320_21075.n5 a_59320_21075.n3 0.833
R22168 a_59320_21075.n3 a_59320_21075.n2 0.653
R22169 a_59320_21075.n5 a_59320_21075.n4 0.653
R22170 a_59320_21075.n6 a_59320_21075.n5 0.341
R22171 a_59320_21075.n3 a_59320_21075.n1 0.032
R22172 a_63602_n1637.n0 a_63602_n1637.t8 214.335
R22173 a_63602_n1637.t10 a_63602_n1637.n0 214.335
R22174 a_63602_n1637.n1 a_63602_n1637.t10 143.851
R22175 a_63602_n1637.n1 a_63602_n1637.t9 135.658
R22176 a_63602_n1637.n0 a_63602_n1637.t7 80.333
R22177 a_63602_n1637.n2 a_63602_n1637.t4 28.565
R22178 a_63602_n1637.n2 a_63602_n1637.t5 28.565
R22179 a_63602_n1637.n4 a_63602_n1637.t6 28.565
R22180 a_63602_n1637.n4 a_63602_n1637.t0 28.565
R22181 a_63602_n1637.n7 a_63602_n1637.t1 28.565
R22182 a_63602_n1637.t2 a_63602_n1637.n7 28.565
R22183 a_63602_n1637.n6 a_63602_n1637.t3 9.714
R22184 a_63602_n1637.n7 a_63602_n1637.n6 1.003
R22185 a_63602_n1637.n5 a_63602_n1637.n3 0.833
R22186 a_63602_n1637.n3 a_63602_n1637.n2 0.653
R22187 a_63602_n1637.n5 a_63602_n1637.n4 0.653
R22188 a_63602_n1637.n6 a_63602_n1637.n5 0.341
R22189 a_63602_n1637.n3 a_63602_n1637.n1 0.032
R22190 a_20633_13581.n3 a_20633_13581.t5 448.381
R22191 a_20633_13581.n2 a_20633_13581.t4 286.438
R22192 a_20633_13581.n2 a_20633_13581.t7 286.438
R22193 a_20633_13581.n1 a_20633_13581.t6 247.69
R22194 a_20633_13581.n4 a_20633_13581.n0 182.117
R22195 a_20633_13581.t5 a_20633_13581.n2 160.666
R22196 a_20633_13581.t2 a_20633_13581.n4 28.568
R22197 a_20633_13581.n0 a_20633_13581.t0 28.565
R22198 a_20633_13581.n0 a_20633_13581.t1 28.565
R22199 a_20633_13581.n1 a_20633_13581.t3 18.127
R22200 a_20633_13581.n3 a_20633_13581.n1 4.036
R22201 a_20633_13581.n4 a_20633_13581.n3 0.937
R22202 a_58328_16462.n1 a_58328_16462.t4 318.922
R22203 a_58328_16462.n0 a_58328_16462.t6 274.739
R22204 a_58328_16462.n0 a_58328_16462.t5 274.739
R22205 a_58328_16462.n1 a_58328_16462.t7 269.116
R22206 a_58328_16462.t4 a_58328_16462.n0 179.946
R22207 a_58328_16462.n2 a_58328_16462.n1 105.178
R22208 a_58328_16462.n3 a_58328_16462.t0 29.444
R22209 a_58328_16462.n4 a_58328_16462.t1 28.565
R22210 a_58328_16462.t2 a_58328_16462.n4 28.565
R22211 a_58328_16462.n2 a_58328_16462.t3 18.145
R22212 a_58328_16462.n3 a_58328_16462.n2 2.878
R22213 a_58328_16462.n4 a_58328_16462.n3 0.764
R22214 a_17479_n2637.n1 a_17479_n2637.t7 867.497
R22215 a_17479_n2637.n1 a_17479_n2637.t5 615.911
R22216 a_17479_n2637.n0 a_17479_n2637.t6 286.438
R22217 a_17479_n2637.n0 a_17479_n2637.t4 286.438
R22218 a_17479_n2637.n4 a_17479_n2637.n3 185.55
R22219 a_17479_n2637.t7 a_17479_n2637.n0 160.666
R22220 a_17479_n2637.n3 a_17479_n2637.t1 28.568
R22221 a_17479_n2637.t2 a_17479_n2637.n4 28.565
R22222 a_17479_n2637.n4 a_17479_n2637.t0 28.565
R22223 a_17479_n2637.n2 a_17479_n2637.n1 24.086
R22224 a_17479_n2637.n2 a_17479_n2637.t3 20.393
R22225 a_17479_n2637.n3 a_17479_n2637.n2 2.076
R22226 a_41933_310.t0 a_41933_310.t1 17.4
R22227 a_18389_4620.t0 a_18389_4620.t1 17.4
R22228 a_66063_3092.n1 a_66063_3092.t5 318.922
R22229 a_66063_3092.n0 a_66063_3092.t6 274.739
R22230 a_66063_3092.n0 a_66063_3092.t7 274.739
R22231 a_66063_3092.n1 a_66063_3092.t4 269.116
R22232 a_66063_3092.t5 a_66063_3092.n0 179.946
R22233 a_66063_3092.n2 a_66063_3092.n1 107.263
R22234 a_66063_3092.n3 a_66063_3092.t0 29.444
R22235 a_66063_3092.t2 a_66063_3092.n4 28.565
R22236 a_66063_3092.n4 a_66063_3092.t1 28.565
R22237 a_66063_3092.n2 a_66063_3092.t3 18.145
R22238 a_66063_3092.n3 a_66063_3092.n2 2.878
R22239 a_66063_3092.n4 a_66063_3092.n3 0.764
R22240 a_65769_2386.t0 a_65769_2386.t1 380.209
R22241 a_20633_10847.n2 a_20633_10847.t6 448.381
R22242 a_20633_10847.n1 a_20633_10847.t5 286.438
R22243 a_20633_10847.n1 a_20633_10847.t7 286.438
R22244 a_20633_10847.n0 a_20633_10847.t4 247.69
R22245 a_20633_10847.n4 a_20633_10847.n3 182.117
R22246 a_20633_10847.t6 a_20633_10847.n1 160.666
R22247 a_20633_10847.n3 a_20633_10847.t0 28.568
R22248 a_20633_10847.n4 a_20633_10847.t1 28.565
R22249 a_20633_10847.t2 a_20633_10847.n4 28.565
R22250 a_20633_10847.n0 a_20633_10847.t3 18.127
R22251 a_20633_10847.n2 a_20633_10847.n0 4.036
R22252 a_20633_10847.n3 a_20633_10847.n2 0.937
R22253 a_66061_10678.n1 a_66061_10678.t6 318.922
R22254 a_66061_10678.n0 a_66061_10678.t4 274.739
R22255 a_66061_10678.n0 a_66061_10678.t7 274.739
R22256 a_66061_10678.n1 a_66061_10678.t5 269.116
R22257 a_66061_10678.t6 a_66061_10678.n0 179.946
R22258 a_66061_10678.n2 a_66061_10678.n1 107.263
R22259 a_66061_10678.n3 a_66061_10678.t0 29.444
R22260 a_66061_10678.n4 a_66061_10678.t1 28.565
R22261 a_66061_10678.t2 a_66061_10678.n4 28.565
R22262 a_66061_10678.n2 a_66061_10678.t3 18.145
R22263 a_66061_10678.n3 a_66061_10678.n2 2.878
R22264 a_66061_10678.n4 a_66061_10678.n3 0.764
R22265 a_65767_10704.t1 a_65767_10704.n0 14.282
R22266 a_65767_10704.n0 a_65767_10704.t2 14.282
R22267 a_65767_10704.n0 a_65767_10704.n8 122.999
R22268 a_65767_10704.n8 a_65767_10704.n6 50.575
R22269 a_65767_10704.n6 a_65767_10704.n4 74.302
R22270 a_65767_10704.n8 a_65767_10704.n7 157.665
R22271 a_65767_10704.n7 a_65767_10704.t0 8.7
R22272 a_65767_10704.n7 a_65767_10704.t4 8.7
R22273 a_65767_10704.n6 a_65767_10704.n5 90.416
R22274 a_65767_10704.n5 a_65767_10704.t3 14.282
R22275 a_65767_10704.n5 a_65767_10704.t7 14.282
R22276 a_65767_10704.n4 a_65767_10704.n3 90.436
R22277 a_65767_10704.n3 a_65767_10704.t6 14.282
R22278 a_65767_10704.n3 a_65767_10704.t5 14.282
R22279 a_65767_10704.n4 a_65767_10704.n1 1216.25
R22280 a_65767_10704.n1 a_65767_10704.t9 408.806
R22281 a_65767_10704.t10 a_65767_10704.n2 160.666
R22282 a_65767_10704.n1 a_65767_10704.t10 989.744
R22283 a_65767_10704.n2 a_65767_10704.t8 287.241
R22284 a_65767_10704.n2 a_65767_10704.t11 287.241
R22285 a_53299_1015.n1 a_53299_1015.t7 318.922
R22286 a_53299_1015.n0 a_53299_1015.t4 274.739
R22287 a_53299_1015.n0 a_53299_1015.t5 274.739
R22288 a_53299_1015.n1 a_53299_1015.t6 269.116
R22289 a_53299_1015.t7 a_53299_1015.n0 179.946
R22290 a_53299_1015.n2 a_53299_1015.n1 107.263
R22291 a_53299_1015.n3 a_53299_1015.t1 29.444
R22292 a_53299_1015.t2 a_53299_1015.n4 28.565
R22293 a_53299_1015.n4 a_53299_1015.t0 28.565
R22294 a_53299_1015.n2 a_53299_1015.t3 18.145
R22295 a_53299_1015.n3 a_53299_1015.n2 2.878
R22296 a_53299_1015.n4 a_53299_1015.n3 0.764
R22297 a_39943_23696.t0 a_39943_23696.t1 17.4
R22298 a_40305_20642.t5 a_40305_20642.t7 574.43
R22299 a_40305_20642.n1 a_40305_20642.t4 285.109
R22300 a_40305_20642.n3 a_40305_20642.n2 197.217
R22301 a_40305_20642.n4 a_40305_20642.n0 192.754
R22302 a_40305_20642.n1 a_40305_20642.t6 160.666
R22303 a_40305_20642.n2 a_40305_20642.t5 160.666
R22304 a_40305_20642.n2 a_40305_20642.n1 114.829
R22305 a_40305_20642.t2 a_40305_20642.n4 28.568
R22306 a_40305_20642.n0 a_40305_20642.t0 28.565
R22307 a_40305_20642.n0 a_40305_20642.t1 28.565
R22308 a_40305_20642.n3 a_40305_20642.t3 18.838
R22309 a_40305_20642.n4 a_40305_20642.n3 1.129
R22310 a_22540_14454.n2 a_22540_14454.t5 867.497
R22311 a_22540_14454.n2 a_22540_14454.t6 591.811
R22312 a_22540_14454.n1 a_22540_14454.t4 286.438
R22313 a_22540_14454.n1 a_22540_14454.t7 286.438
R22314 a_22540_14454.n4 a_22540_14454.n0 185.55
R22315 a_22540_14454.t5 a_22540_14454.n1 160.666
R22316 a_22540_14454.t2 a_22540_14454.n4 28.568
R22317 a_22540_14454.n0 a_22540_14454.t0 28.565
R22318 a_22540_14454.n0 a_22540_14454.t1 28.565
R22319 a_22540_14454.n3 a_22540_14454.n2 26.067
R22320 a_22540_14454.n3 a_22540_14454.t3 21.376
R22321 a_22540_14454.n4 a_22540_14454.n3 1.637
R22322 a_63769_11165.t0 a_63769_11165.t1 17.4
R22323 a_23958_13121.t0 a_23958_13121.t1 17.4
R22324 a_65222_11397.n2 a_65222_11397.t6 318.922
R22325 a_65222_11397.n1 a_65222_11397.t5 273.935
R22326 a_65222_11397.n1 a_65222_11397.t7 273.935
R22327 a_65222_11397.n2 a_65222_11397.t4 269.116
R22328 a_65222_11397.n4 a_65222_11397.n0 193.227
R22329 a_65222_11397.t6 a_65222_11397.n1 179.142
R22330 a_65222_11397.n3 a_65222_11397.n2 106.999
R22331 a_65222_11397.t2 a_65222_11397.n4 28.568
R22332 a_65222_11397.n0 a_65222_11397.t0 28.565
R22333 a_65222_11397.n0 a_65222_11397.t1 28.565
R22334 a_65222_11397.n3 a_65222_11397.t3 18.149
R22335 a_65222_11397.n4 a_65222_11397.n3 3.726
R22336 a_65767_9972.t0 a_65767_9972.t1 380.209
R22337 a_6556_n2148.n3 a_6556_n2148.t6 448.382
R22338 a_6556_n2148.n2 a_6556_n2148.t5 286.438
R22339 a_6556_n2148.n2 a_6556_n2148.t7 286.438
R22340 a_6556_n2148.n1 a_6556_n2148.t4 247.69
R22341 a_6556_n2148.n4 a_6556_n2148.n0 182.117
R22342 a_6556_n2148.t6 a_6556_n2148.n2 160.666
R22343 a_6556_n2148.t2 a_6556_n2148.n4 28.568
R22344 a_6556_n2148.n0 a_6556_n2148.t0 28.565
R22345 a_6556_n2148.n0 a_6556_n2148.t1 28.565
R22346 a_6556_n2148.n1 a_6556_n2148.t3 18.127
R22347 a_6556_n2148.n3 a_6556_n2148.n1 4.039
R22348 a_6556_n2148.n4 a_6556_n2148.n3 0.937
R22349 a_7936_n3481.t0 a_7936_n3481.t1 17.4
R22350 Cout.n1 Cout.t0 28.57
R22351 Cout.n0 Cout.t1 28.565
R22352 Cout.n0 Cout.t2 28.565
R22353 Cout.n1 Cout.t3 17.638
R22354 Cout Cout.n2 7.386
R22355 Cout.n2 Cout.n0 0.693
R22356 Cout.n2 Cout.n1 0.597
R22357 a_71846_17727.t0 a_71846_17727.t1 17.4
R22358 a_44697_5979.t0 a_44697_5979.t1 17.4
R22359 a_12732_15818.n3 a_12732_15818.n2 3288.61
R22360 a_12732_15818.n2 a_12732_15818.t5 990.34
R22361 a_12732_15818.n2 a_12732_15818.t6 408.211
R22362 a_12732_15818.n1 a_12732_15818.t4 286.438
R22363 a_12732_15818.n1 a_12732_15818.t7 286.438
R22364 a_12732_15818.t5 a_12732_15818.n1 160.666
R22365 a_12732_15818.n3 a_12732_15818.n0 114.449
R22366 a_12732_15818.n4 a_12732_15818.n3 99.011
R22367 a_12732_15818.t2 a_12732_15818.n4 28.568
R22368 a_12732_15818.n0 a_12732_15818.t0 28.565
R22369 a_12732_15818.n0 a_12732_15818.t1 28.565
R22370 a_12732_15818.n4 a_12732_15818.t3 17.641
R22371 a_56792_20633.t0 a_56792_20633.t1 17.4
R22372 a_12902_n2152.n3 a_12902_n2152.t7 448.382
R22373 a_12902_n2152.n2 a_12902_n2152.t6 286.438
R22374 a_12902_n2152.n2 a_12902_n2152.t4 286.438
R22375 a_12902_n2152.n1 a_12902_n2152.t5 247.69
R22376 a_12902_n2152.n4 a_12902_n2152.n0 182.117
R22377 a_12902_n2152.t7 a_12902_n2152.n2 160.666
R22378 a_12902_n2152.t2 a_12902_n2152.n4 28.568
R22379 a_12902_n2152.n0 a_12902_n2152.t0 28.565
R22380 a_12902_n2152.n0 a_12902_n2152.t1 28.565
R22381 a_12902_n2152.n1 a_12902_n2152.t3 18.127
R22382 a_12902_n2152.n3 a_12902_n2152.n1 4.039
R22383 a_12902_n2152.n4 a_12902_n2152.n3 0.937
R22384 a_13810_n2152.n4 a_13810_n2152.t8 1527.4
R22385 a_13810_n2152.t8 a_13810_n2152.n3 657.379
R22386 a_13810_n2152.n1 a_13810_n2152.n0 258.161
R22387 a_13810_n2152.n7 a_13810_n2152.n6 258.161
R22388 a_13810_n2152.n2 a_13810_n2152.t9 206.421
R22389 a_13810_n2152.t11 a_13810_n2152.n2 206.421
R22390 a_13810_n2152.n4 a_13810_n2152.t11 200.029
R22391 a_13810_n2152.n5 a_13810_n2152.n4 97.614
R22392 a_13810_n2152.n2 a_13810_n2152.t10 80.333
R22393 a_13810_n2152.n6 a_13810_n2152.t2 14.283
R22394 a_13810_n2152.n1 a_13810_n2152.t5 14.283
R22395 a_13810_n2152.n0 a_13810_n2152.t6 14.282
R22396 a_13810_n2152.n0 a_13810_n2152.t7 14.282
R22397 a_13810_n2152.t3 a_13810_n2152.n7 14.282
R22398 a_13810_n2152.n7 a_13810_n2152.t1 14.282
R22399 a_13810_n2152.n3 a_13810_n2152.t0 8.7
R22400 a_13810_n2152.n3 a_13810_n2152.t4 8.7
R22401 a_13810_n2152.n6 a_13810_n2152.n5 4.366
R22402 a_13810_n2152.n5 a_13810_n2152.n1 0.852
R22403 a_16605_n2152.t0 a_16605_n2152.n0 14.282
R22404 a_16605_n2152.n0 a_16605_n2152.t2 14.282
R22405 a_16605_n2152.n7 a_16605_n2152.n8 75.815
R22406 a_16605_n2152.n5 a_16605_n2152.n7 77.456
R22407 a_16605_n2152.n3 a_16605_n2152.n5 77.456
R22408 a_16605_n2152.n1 a_16605_n2152.n3 77.784
R22409 a_16605_n2152.n0 a_16605_n2152.n1 167.433
R22410 a_16605_n2152.n8 a_16605_n2152.n9 167.433
R22411 a_16605_n2152.n9 a_16605_n2152.t11 14.282
R22412 a_16605_n2152.n9 a_16605_n2152.t10 14.282
R22413 a_16605_n2152.n8 a_16605_n2152.t9 104.259
R22414 a_16605_n2152.n7 a_16605_n2152.n6 89.977
R22415 a_16605_n2152.n6 a_16605_n2152.t8 14.282
R22416 a_16605_n2152.n6 a_16605_n2152.t7 14.282
R22417 a_16605_n2152.n5 a_16605_n2152.n4 89.977
R22418 a_16605_n2152.n4 a_16605_n2152.t6 14.282
R22419 a_16605_n2152.n4 a_16605_n2152.t4 14.282
R22420 a_16605_n2152.n3 a_16605_n2152.n2 89.977
R22421 a_16605_n2152.n2 a_16605_n2152.t3 14.282
R22422 a_16605_n2152.n2 a_16605_n2152.t5 14.282
R22423 a_16605_n2152.n1 a_16605_n2152.t1 104.259
R22424 a_16954_n2152.n3 a_16954_n2152.t11 1527.4
R22425 a_16954_n2152.t11 a_16954_n2152.n2 657.379
R22426 a_16954_n2152.n5 a_16954_n2152.n4 258.161
R22427 a_16954_n2152.n7 a_16954_n2152.n0 258.161
R22428 a_16954_n2152.n1 a_16954_n2152.t8 206.421
R22429 a_16954_n2152.t10 a_16954_n2152.n1 206.421
R22430 a_16954_n2152.n3 a_16954_n2152.t10 200.029
R22431 a_16954_n2152.n6 a_16954_n2152.n3 97.614
R22432 a_16954_n2152.n1 a_16954_n2152.t9 80.333
R22433 a_16954_n2152.n5 a_16954_n2152.t7 14.283
R22434 a_16954_n2152.t2 a_16954_n2152.n7 14.283
R22435 a_16954_n2152.n4 a_16954_n2152.t5 14.282
R22436 a_16954_n2152.n4 a_16954_n2152.t6 14.282
R22437 a_16954_n2152.n0 a_16954_n2152.t0 14.282
R22438 a_16954_n2152.n0 a_16954_n2152.t1 14.282
R22439 a_16954_n2152.n2 a_16954_n2152.t4 8.7
R22440 a_16954_n2152.n2 a_16954_n2152.t3 8.7
R22441 a_16954_n2152.n6 a_16954_n2152.n5 4.366
R22442 a_16954_n2152.n7 a_16954_n2152.n6 0.852
R22443 a_12870_1740.n2 a_12870_1740.t5 448.382
R22444 a_12870_1740.n1 a_12870_1740.t7 286.438
R22445 a_12870_1740.n1 a_12870_1740.t6 286.438
R22446 a_12870_1740.n0 a_12870_1740.t4 247.69
R22447 a_12870_1740.n4 a_12870_1740.n3 182.117
R22448 a_12870_1740.t5 a_12870_1740.n1 160.666
R22449 a_12870_1740.n3 a_12870_1740.t1 28.568
R22450 a_12870_1740.t2 a_12870_1740.n4 28.565
R22451 a_12870_1740.n4 a_12870_1740.t0 28.565
R22452 a_12870_1740.n0 a_12870_1740.t3 18.127
R22453 a_12870_1740.n2 a_12870_1740.n0 4.039
R22454 a_12870_1740.n3 a_12870_1740.n2 0.937
R22455 a_59871_6178.t0 a_59871_6178.t1 17.4
R22456 a_17190_n3485.t0 a_17190_n3485.t1 17.4
R22457 a_23755_n2633.n1 a_23755_n2633.t5 867.497
R22458 a_23755_n2633.n1 a_23755_n2633.t7 615.911
R22459 a_23755_n2633.n0 a_23755_n2633.t4 286.438
R22460 a_23755_n2633.n0 a_23755_n2633.t6 286.438
R22461 a_23755_n2633.n4 a_23755_n2633.n3 185.55
R22462 a_23755_n2633.t5 a_23755_n2633.n0 160.666
R22463 a_23755_n2633.n3 a_23755_n2633.t1 28.568
R22464 a_23755_n2633.n4 a_23755_n2633.t0 28.565
R22465 a_23755_n2633.t2 a_23755_n2633.n4 28.565
R22466 a_23755_n2633.n2 a_23755_n2633.n1 22.125
R22467 a_23755_n2633.n2 a_23755_n2633.t3 20.393
R22468 a_23755_n2633.n3 a_23755_n2633.n2 1.835
R22469 a_22881_n2148.n0 a_22881_n2148.t1 14.282
R22470 a_22881_n2148.t0 a_22881_n2148.n0 14.282
R22471 a_22881_n2148.n7 a_22881_n2148.n8 75.815
R22472 a_22881_n2148.n5 a_22881_n2148.n7 77.456
R22473 a_22881_n2148.n3 a_22881_n2148.n5 77.456
R22474 a_22881_n2148.n1 a_22881_n2148.n3 77.784
R22475 a_22881_n2148.n0 a_22881_n2148.n1 167.433
R22476 a_22881_n2148.n8 a_22881_n2148.n9 167.433
R22477 a_22881_n2148.n9 a_22881_n2148.t8 14.282
R22478 a_22881_n2148.n9 a_22881_n2148.t4 14.282
R22479 a_22881_n2148.n8 a_22881_n2148.t3 104.259
R22480 a_22881_n2148.n7 a_22881_n2148.n6 89.977
R22481 a_22881_n2148.n6 a_22881_n2148.t11 14.282
R22482 a_22881_n2148.n6 a_22881_n2148.t10 14.282
R22483 a_22881_n2148.n5 a_22881_n2148.n4 89.977
R22484 a_22881_n2148.n4 a_22881_n2148.t9 14.282
R22485 a_22881_n2148.n4 a_22881_n2148.t6 14.282
R22486 a_22881_n2148.n3 a_22881_n2148.n2 89.977
R22487 a_22881_n2148.n2 a_22881_n2148.t5 14.282
R22488 a_22881_n2148.n2 a_22881_n2148.t7 14.282
R22489 a_22881_n2148.n1 a_22881_n2148.t2 104.259
R22490 a_23230_n2148.n2 a_23230_n2148.t9 1527.4
R22491 a_23230_n2148.t9 a_23230_n2148.n1 657.379
R22492 a_23230_n2148.n4 a_23230_n2148.n3 258.161
R22493 a_23230_n2148.n7 a_23230_n2148.n6 258.161
R22494 a_23230_n2148.n0 a_23230_n2148.t8 206.421
R22495 a_23230_n2148.t11 a_23230_n2148.n0 206.421
R22496 a_23230_n2148.n2 a_23230_n2148.t11 200.029
R22497 a_23230_n2148.n5 a_23230_n2148.n2 97.614
R22498 a_23230_n2148.n0 a_23230_n2148.t10 80.333
R22499 a_23230_n2148.n4 a_23230_n2148.t6 14.283
R22500 a_23230_n2148.n6 a_23230_n2148.t0 14.283
R22501 a_23230_n2148.n3 a_23230_n2148.t4 14.282
R22502 a_23230_n2148.n3 a_23230_n2148.t5 14.282
R22503 a_23230_n2148.n7 a_23230_n2148.t1 14.282
R22504 a_23230_n2148.t2 a_23230_n2148.n7 14.282
R22505 a_23230_n2148.n1 a_23230_n2148.t7 8.7
R22506 a_23230_n2148.n1 a_23230_n2148.t3 8.7
R22507 a_23230_n2148.n5 a_23230_n2148.n4 4.366
R22508 a_23230_n2148.n6 a_23230_n2148.n5 0.852
R22509 a_19948_20263.t0 a_19948_20263.t1 17.4
R22510 a_46275_18597.n0 a_46275_18597.t5 14.282
R22511 a_46275_18597.n0 a_46275_18597.t1 14.282
R22512 a_46275_18597.n1 a_46275_18597.t3 14.282
R22513 a_46275_18597.n1 a_46275_18597.t4 14.282
R22514 a_46275_18597.t0 a_46275_18597.n3 14.282
R22515 a_46275_18597.n3 a_46275_18597.t2 14.282
R22516 a_46275_18597.n2 a_46275_18597.n0 2.546
R22517 a_46275_18597.n2 a_46275_18597.n1 2.367
R22518 a_46275_18597.n3 a_46275_18597.n2 0.001
R22519 a_53246_6110.t0 a_53246_6110.t1 17.4
R22520 a_11829_5352.n0 a_11829_5352.t10 14.282
R22521 a_11829_5352.t9 a_11829_5352.n0 14.282
R22522 a_11829_5352.n0 a_11829_5352.n9 0.999
R22523 a_11829_5352.n6 a_11829_5352.n8 0.2
R22524 a_11829_5352.n9 a_11829_5352.n6 0.575
R22525 a_11829_5352.n9 a_11829_5352.t11 16.058
R22526 a_11829_5352.n8 a_11829_5352.n7 0.999
R22527 a_11829_5352.n7 a_11829_5352.t7 14.282
R22528 a_11829_5352.n7 a_11829_5352.t8 14.282
R22529 a_11829_5352.n8 a_11829_5352.t6 16.058
R22530 a_11829_5352.n6 a_11829_5352.n4 0.227
R22531 a_11829_5352.n4 a_11829_5352.n5 1.511
R22532 a_11829_5352.n5 a_11829_5352.t3 14.282
R22533 a_11829_5352.n5 a_11829_5352.t4 14.282
R22534 a_11829_5352.n4 a_11829_5352.n1 0.669
R22535 a_11829_5352.n1 a_11829_5352.n2 0.001
R22536 a_11829_5352.n1 a_11829_5352.n3 267.767
R22537 a_11829_5352.n3 a_11829_5352.t2 14.282
R22538 a_11829_5352.n3 a_11829_5352.t1 14.282
R22539 a_11829_5352.n2 a_11829_5352.t0 14.282
R22540 a_11829_5352.n2 a_11829_5352.t5 14.282
R22541 a_43405_16438.t0 a_43405_16438.t1 17.4
R22542 a_61071_3878.t6 a_61071_3878.n2 404.877
R22543 a_61071_3878.n1 a_61071_3878.t7 210.902
R22544 a_61071_3878.n3 a_61071_3878.t6 136.943
R22545 a_61071_3878.n2 a_61071_3878.n1 107.801
R22546 a_61071_3878.n1 a_61071_3878.t8 80.333
R22547 a_61071_3878.n2 a_61071_3878.t5 80.333
R22548 a_61071_3878.n0 a_61071_3878.t4 17.4
R22549 a_61071_3878.n0 a_61071_3878.t0 17.4
R22550 a_61071_3878.n4 a_61071_3878.t2 15.032
R22551 a_61071_3878.n5 a_61071_3878.t1 14.282
R22552 a_61071_3878.t3 a_61071_3878.n5 14.282
R22553 a_61071_3878.n5 a_61071_3878.n4 1.65
R22554 a_61071_3878.n3 a_61071_3878.n0 0.672
R22555 a_61071_3878.n4 a_61071_3878.n3 0.665
R22556 a_20814_10387.t0 a_20814_10387.t1 17.4
R22557 a_52767_15740.n1 a_52767_15740.t5 318.922
R22558 a_52767_15740.n0 a_52767_15740.t4 273.935
R22559 a_52767_15740.n0 a_52767_15740.t6 273.935
R22560 a_52767_15740.n1 a_52767_15740.t7 269.116
R22561 a_52767_15740.n4 a_52767_15740.n3 193.227
R22562 a_52767_15740.t5 a_52767_15740.n0 179.142
R22563 a_52767_15740.n2 a_52767_15740.n1 106.999
R22564 a_52767_15740.n3 a_52767_15740.t0 28.568
R22565 a_52767_15740.n4 a_52767_15740.t1 28.565
R22566 a_52767_15740.t2 a_52767_15740.n4 28.565
R22567 a_52767_15740.n2 a_52767_15740.t3 18.149
R22568 a_52767_15740.n3 a_52767_15740.n2 3.726
R22569 a_43410_14834.t0 a_43410_14834.t1 17.4
R22570 a_10397_15824.n3 a_10397_15824.n2 2682.61
R22571 a_10397_15824.n2 a_10397_15824.t4 990.34
R22572 a_10397_15824.n2 a_10397_15824.t7 408.211
R22573 a_10397_15824.n1 a_10397_15824.t6 286.438
R22574 a_10397_15824.n1 a_10397_15824.t5 286.438
R22575 a_10397_15824.t4 a_10397_15824.n1 160.666
R22576 a_10397_15824.n4 a_10397_15824.n3 116.875
R22577 a_10397_15824.n3 a_10397_15824.n0 99.45
R22578 a_10397_15824.n0 a_10397_15824.t3 28.568
R22579 a_10397_15824.n4 a_10397_15824.t2 28.565
R22580 a_10397_15824.t1 a_10397_15824.n4 28.565
R22581 a_10397_15824.n0 a_10397_15824.t0 17.64
R22582 a_16322_10994.n4 a_16322_10994.t9 1527.4
R22583 a_16322_10994.t9 a_16322_10994.n3 657.379
R22584 a_16322_10994.n1 a_16322_10994.n0 258.161
R22585 a_16322_10994.n7 a_16322_10994.n6 258.161
R22586 a_16322_10994.n2 a_16322_10994.t8 206.421
R22587 a_16322_10994.t10 a_16322_10994.n2 206.421
R22588 a_16322_10994.n4 a_16322_10994.t10 200.029
R22589 a_16322_10994.n5 a_16322_10994.n4 97.614
R22590 a_16322_10994.n2 a_16322_10994.t11 80.333
R22591 a_16322_10994.n1 a_16322_10994.t5 14.283
R22592 a_16322_10994.n6 a_16322_10994.t1 14.283
R22593 a_16322_10994.n0 a_16322_10994.t7 14.282
R22594 a_16322_10994.n0 a_16322_10994.t6 14.282
R22595 a_16322_10994.n7 a_16322_10994.t2 14.282
R22596 a_16322_10994.t3 a_16322_10994.n7 14.282
R22597 a_16322_10994.n3 a_16322_10994.t4 8.7
R22598 a_16322_10994.n3 a_16322_10994.t0 8.7
R22599 a_16322_10994.n6 a_16322_10994.n5 4.366
R22600 a_16322_10994.n5 a_16322_10994.n1 0.852
R22601 a_16264_11724.n1 a_16264_11724.t5 990.34
R22602 a_16264_11724.n1 a_16264_11724.t4 408.211
R22603 a_16264_11724.n2 a_16264_11724.n1 338.656
R22604 a_16264_11724.n0 a_16264_11724.t6 286.438
R22605 a_16264_11724.n0 a_16264_11724.t7 286.438
R22606 a_16264_11724.n4 a_16264_11724.n3 185.55
R22607 a_16264_11724.t5 a_16264_11724.n0 160.666
R22608 a_16264_11724.n3 a_16264_11724.t1 28.568
R22609 a_16264_11724.t2 a_16264_11724.n4 28.565
R22610 a_16264_11724.n4 a_16264_11724.t0 28.565
R22611 a_16264_11724.n2 a_16264_11724.t3 21.376
R22612 a_16264_11724.n3 a_16264_11724.n2 1.637
R22613 a_16795_14432.n1 a_16795_14432.t7 867.497
R22614 a_16795_14432.n1 a_16795_14432.t6 591.811
R22615 a_16795_14432.n0 a_16795_14432.t4 286.438
R22616 a_16795_14432.n0 a_16795_14432.t5 286.438
R22617 a_16795_14432.n4 a_16795_14432.n3 192.754
R22618 a_16795_14432.t7 a_16795_14432.n0 160.666
R22619 a_16795_14432.n3 a_16795_14432.t3 28.568
R22620 a_16795_14432.n4 a_16795_14432.t2 28.565
R22621 a_16795_14432.t1 a_16795_14432.n4 28.565
R22622 a_16795_14432.n2 a_16795_14432.n1 22.544
R22623 a_16795_14432.n2 a_16795_14432.t0 18.726
R22624 a_16795_14432.n3 a_16795_14432.n2 1.123
R22625 a_14548_7659.t0 a_14548_7659.t1 17.4
R22626 a_7956_10387.t0 a_7956_10387.t1 17.4
R22627 a_47703_1733.n2 a_47703_1733.t7 318.922
R22628 a_47703_1733.n1 a_47703_1733.t4 273.935
R22629 a_47703_1733.n1 a_47703_1733.t5 273.935
R22630 a_47703_1733.n2 a_47703_1733.t6 269.116
R22631 a_47703_1733.n4 a_47703_1733.n0 193.227
R22632 a_47703_1733.t7 a_47703_1733.n1 179.142
R22633 a_47703_1733.n3 a_47703_1733.n2 106.999
R22634 a_47703_1733.t2 a_47703_1733.n4 28.568
R22635 a_47703_1733.n0 a_47703_1733.t1 28.565
R22636 a_47703_1733.n0 a_47703_1733.t0 28.565
R22637 a_47703_1733.n3 a_47703_1733.t3 18.149
R22638 a_47703_1733.n4 a_47703_1733.n3 3.726
R22639 a_41913_11312.t0 a_41913_11312.t1 17.4
R22640 a_10449_14428.n2 a_10449_14428.t5 867.497
R22641 a_10449_14428.n2 a_10449_14428.t7 591.811
R22642 a_10449_14428.n1 a_10449_14428.t4 286.438
R22643 a_10449_14428.n1 a_10449_14428.t6 286.438
R22644 a_10449_14428.n4 a_10449_14428.n0 192.754
R22645 a_10449_14428.t5 a_10449_14428.n1 160.666
R22646 a_10449_14428.t2 a_10449_14428.n4 28.568
R22647 a_10449_14428.n0 a_10449_14428.t0 28.565
R22648 a_10449_14428.n0 a_10449_14428.t1 28.565
R22649 a_10449_14428.n3 a_10449_14428.n2 27.988
R22650 a_10449_14428.n3 a_10449_14428.t3 18.726
R22651 a_10449_14428.n4 a_10449_14428.n3 1.123
R22652 a_38492_9345.t4 a_38492_9345.t6 800.071
R22653 a_38492_9345.n2 a_38492_9345.n1 659.097
R22654 a_38492_9345.n0 a_38492_9345.t5 285.109
R22655 a_38492_9345.n1 a_38492_9345.t4 193.602
R22656 a_38492_9345.n4 a_38492_9345.n3 192.754
R22657 a_38492_9345.n0 a_38492_9345.t7 160.666
R22658 a_38492_9345.n1 a_38492_9345.n0 91.507
R22659 a_38492_9345.n3 a_38492_9345.t1 28.568
R22660 a_38492_9345.n4 a_38492_9345.t0 28.565
R22661 a_38492_9345.t2 a_38492_9345.n4 28.565
R22662 a_38492_9345.n2 a_38492_9345.t3 19.061
R22663 a_38492_9345.n3 a_38492_9345.n2 1.005
R22664 a_19406_8988.n1 a_19406_8988.t6 990.34
R22665 a_19406_8988.n1 a_19406_8988.t4 408.211
R22666 a_19406_8988.n0 a_19406_8988.t5 286.438
R22667 a_19406_8988.n0 a_19406_8988.t7 286.438
R22668 a_19406_8988.n4 a_19406_8988.n3 185.55
R22669 a_19406_8988.t6 a_19406_8988.n0 160.666
R22670 a_19406_8988.n3 a_19406_8988.t1 28.568
R22671 a_19406_8988.n4 a_19406_8988.t0 28.565
R22672 a_19406_8988.t2 a_19406_8988.n4 28.565
R22673 a_19406_8988.n2 a_19406_8988.t3 21.476
R22674 a_19406_8988.n2 a_19406_8988.n1 13.939
R22675 a_19406_8988.n3 a_19406_8988.n2 1.537
R22676 a_4825_1255.n1 a_4825_1255.t7 867.497
R22677 a_4825_1255.n1 a_4825_1255.t4 615.911
R22678 a_4825_1255.n0 a_4825_1255.t5 286.438
R22679 a_4825_1255.n0 a_4825_1255.t6 286.438
R22680 a_4825_1255.n4 a_4825_1255.n3 185.55
R22681 a_4825_1255.t7 a_4825_1255.n0 160.666
R22682 a_4825_1255.n2 a_4825_1255.n1 133.12
R22683 a_4825_1255.t2 a_4825_1255.n4 28.568
R22684 a_4825_1255.n3 a_4825_1255.t0 28.565
R22685 a_4825_1255.n3 a_4825_1255.t1 28.565
R22686 a_4825_1255.n2 a_4825_1255.t3 20.393
R22687 a_4825_1255.n4 a_4825_1255.n2 1.836
R22688 a_4772_407.t0 a_4772_407.t1 17.4
R22689 a_41361_3878.n1 a_41361_3878.t1 14.282
R22690 a_41361_3878.n1 a_41361_3878.t3 14.282
R22691 a_41361_3878.n0 a_41361_3878.t5 14.282
R22692 a_41361_3878.n0 a_41361_3878.t4 14.282
R22693 a_41361_3878.n3 a_41361_3878.t0 14.282
R22694 a_41361_3878.t2 a_41361_3878.n3 14.282
R22695 a_41361_3878.n2 a_41361_3878.n0 2.546
R22696 a_41361_3878.n3 a_41361_3878.n2 2.367
R22697 a_41361_3878.n2 a_41361_3878.n1 0.001
R22698 a_4237_20723.n2 a_4237_20723.t6 448.381
R22699 a_4237_20723.n1 a_4237_20723.t5 286.438
R22700 a_4237_20723.n1 a_4237_20723.t7 286.438
R22701 a_4237_20723.n0 a_4237_20723.t4 247.69
R22702 a_4237_20723.n4 a_4237_20723.n3 182.117
R22703 a_4237_20723.t6 a_4237_20723.n1 160.666
R22704 a_4237_20723.n3 a_4237_20723.t0 28.568
R22705 a_4237_20723.n4 a_4237_20723.t1 28.565
R22706 a_4237_20723.t2 a_4237_20723.n4 28.565
R22707 a_4237_20723.n0 a_4237_20723.t3 18.127
R22708 a_4237_20723.n2 a_4237_20723.n0 4.036
R22709 a_4237_20723.n3 a_4237_20723.n2 0.937
R22710 a_17426_n3485.t0 a_17426_n3485.t1 17.4
R22711 a_1690_7659.t0 a_1690_7659.t1 17.4
R22712 a_20184_20263.t0 a_20184_20263.t1 17.4
R22713 a_51342_9165.t0 a_51342_9165.t1 17.4
R22714 a_39675_15739.n1 a_39675_15739.t7 318.922
R22715 a_39675_15739.n0 a_39675_15739.t6 273.935
R22716 a_39675_15739.n0 a_39675_15739.t4 273.935
R22717 a_39675_15739.n1 a_39675_15739.t5 269.116
R22718 a_39675_15739.n4 a_39675_15739.n3 193.227
R22719 a_39675_15739.t7 a_39675_15739.n0 179.142
R22720 a_39675_15739.n2 a_39675_15739.n1 106.999
R22721 a_39675_15739.n3 a_39675_15739.t2 28.568
R22722 a_39675_15739.n4 a_39675_15739.t1 28.565
R22723 a_39675_15739.t0 a_39675_15739.n4 28.565
R22724 a_39675_15739.n2 a_39675_15739.t3 18.149
R22725 a_39675_15739.n3 a_39675_15739.n2 3.726
R22726 a_13651_14432.n1 a_13651_14432.t5 867.497
R22727 a_13651_14432.n1 a_13651_14432.t7 591.811
R22728 a_13651_14432.n0 a_13651_14432.t4 286.438
R22729 a_13651_14432.n0 a_13651_14432.t6 286.438
R22730 a_13651_14432.n4 a_13651_14432.n3 192.754
R22731 a_13651_14432.t5 a_13651_14432.n0 160.666
R22732 a_13651_14432.n3 a_13651_14432.t1 28.568
R22733 a_13651_14432.t2 a_13651_14432.n4 28.565
R22734 a_13651_14432.n4 a_13651_14432.t0 28.565
R22735 a_13651_14432.n2 a_13651_14432.n1 25.172
R22736 a_13651_14432.n2 a_13651_14432.t3 18.726
R22737 a_13651_14432.n3 a_13651_14432.n2 1.123
R22738 a_15297_16387.n0 a_15297_16387.t7 214.335
R22739 a_15297_16387.t10 a_15297_16387.n0 214.335
R22740 a_15297_16387.n1 a_15297_16387.t10 143.851
R22741 a_15297_16387.n1 a_15297_16387.t8 135.658
R22742 a_15297_16387.n0 a_15297_16387.t9 80.333
R22743 a_15297_16387.n2 a_15297_16387.t3 28.565
R22744 a_15297_16387.n2 a_15297_16387.t4 28.565
R22745 a_15297_16387.n4 a_15297_16387.t5 28.565
R22746 a_15297_16387.n4 a_15297_16387.t1 28.565
R22747 a_15297_16387.t2 a_15297_16387.n7 28.565
R22748 a_15297_16387.n7 a_15297_16387.t0 28.565
R22749 a_15297_16387.n3 a_15297_16387.t6 9.714
R22750 a_15297_16387.n3 a_15297_16387.n2 1.003
R22751 a_15297_16387.n6 a_15297_16387.n5 0.833
R22752 a_15297_16387.n5 a_15297_16387.n4 0.653
R22753 a_15297_16387.n7 a_15297_16387.n6 0.653
R22754 a_15297_16387.n5 a_15297_16387.n3 0.341
R22755 a_15297_16387.n6 a_15297_16387.n1 0.032
R22756 a_54454_9678.t6 a_54454_9678.n2 404.877
R22757 a_54454_9678.n1 a_54454_9678.t8 210.902
R22758 a_54454_9678.n3 a_54454_9678.t6 136.943
R22759 a_54454_9678.n2 a_54454_9678.n1 107.801
R22760 a_54454_9678.n1 a_54454_9678.t5 80.333
R22761 a_54454_9678.n2 a_54454_9678.t7 80.333
R22762 a_54454_9678.n0 a_54454_9678.t0 17.4
R22763 a_54454_9678.n0 a_54454_9678.t4 17.4
R22764 a_54454_9678.n4 a_54454_9678.t2 15.032
R22765 a_54454_9678.n5 a_54454_9678.t1 14.282
R22766 a_54454_9678.t3 a_54454_9678.n5 14.282
R22767 a_54454_9678.n5 a_54454_9678.n4 1.65
R22768 a_54454_9678.n3 a_54454_9678.n0 0.672
R22769 a_54454_9678.n4 a_54454_9678.n3 0.665
R22770 a_31379_12105.t0 a_31379_12105.t1 379.845
R22771 a_3855_6357.n2 a_3855_6357.t4 990.34
R22772 a_3855_6357.n2 a_3855_6357.t5 408.211
R22773 a_3855_6357.n1 a_3855_6357.t6 286.438
R22774 a_3855_6357.n1 a_3855_6357.t7 286.438
R22775 a_3855_6357.n4 a_3855_6357.n0 197.272
R22776 a_3855_6357.t4 a_3855_6357.n1 160.666
R22777 a_3855_6357.t2 a_3855_6357.n4 28.568
R22778 a_3855_6357.n0 a_3855_6357.t0 28.565
R22779 a_3855_6357.n0 a_3855_6357.t1 28.565
R22780 a_3855_6357.n3 a_3855_6357.t3 18.085
R22781 a_3855_6357.n3 a_3855_6357.n2 13.507
R22782 a_3855_6357.n4 a_3855_6357.n3 0.467
R22783 a_41913_24205.t6 a_41913_24205.n2 404.877
R22784 a_41913_24205.n1 a_41913_24205.t8 210.902
R22785 a_41913_24205.n3 a_41913_24205.t6 136.943
R22786 a_41913_24205.n2 a_41913_24205.n1 107.801
R22787 a_41913_24205.n1 a_41913_24205.t7 80.333
R22788 a_41913_24205.n2 a_41913_24205.t5 80.333
R22789 a_41913_24205.n0 a_41913_24205.t4 17.4
R22790 a_41913_24205.n0 a_41913_24205.t0 17.4
R22791 a_41913_24205.n4 a_41913_24205.t2 15.032
R22792 a_41913_24205.n5 a_41913_24205.t3 14.282
R22793 a_41913_24205.t1 a_41913_24205.n5 14.282
R22794 a_41913_24205.n5 a_41913_24205.n4 1.65
R22795 a_41913_24205.n3 a_41913_24205.n0 0.672
R22796 a_41913_24205.n4 a_41913_24205.n3 0.665
R22797 a_7326_20263.t0 a_7326_20263.t1 17.4
R22798 a_19146_1744.n2 a_19146_1744.t4 448.382
R22799 a_19146_1744.n1 a_19146_1744.t6 286.438
R22800 a_19146_1744.n1 a_19146_1744.t7 286.438
R22801 a_19146_1744.n0 a_19146_1744.t5 247.69
R22802 a_19146_1744.n4 a_19146_1744.n3 182.117
R22803 a_19146_1744.t4 a_19146_1744.n1 160.666
R22804 a_19146_1744.n3 a_19146_1744.t1 28.568
R22805 a_19146_1744.n4 a_19146_1744.t0 28.565
R22806 a_19146_1744.t2 a_19146_1744.n4 28.565
R22807 a_19146_1744.n0 a_19146_1744.t3 18.127
R22808 a_19146_1744.n2 a_19146_1744.n0 4.039
R22809 a_19146_1744.n3 a_19146_1744.n2 0.937
R22810 a_31375_1999.t0 a_31375_1999.t1 17.4
R22811 a_41160_7515.n1 a_41160_7515.t7 318.922
R22812 a_41160_7515.n0 a_41160_7515.t4 273.935
R22813 a_41160_7515.n0 a_41160_7515.t5 273.935
R22814 a_41160_7515.n1 a_41160_7515.t6 269.116
R22815 a_41160_7515.n4 a_41160_7515.n3 193.227
R22816 a_41160_7515.t7 a_41160_7515.n0 179.142
R22817 a_41160_7515.n2 a_41160_7515.n1 106.999
R22818 a_41160_7515.n3 a_41160_7515.t1 28.568
R22819 a_41160_7515.n4 a_41160_7515.t0 28.565
R22820 a_41160_7515.t2 a_41160_7515.n4 28.565
R22821 a_41160_7515.n2 a_41160_7515.t3 18.149
R22822 a_41160_7515.n3 a_41160_7515.n2 3.726
R22823 a_56497_16439.t0 a_56497_16439.t1 17.4
R22824 Y[0].n1 Y[0].n0 185.55
R22825 Y[0].n1 Y[0].t0 28.568
R22826 Y[0].n0 Y[0].t1 28.565
R22827 Y[0].n0 Y[0].t2 28.565
R22828 Y[0].n2 Y[0].t3 20.393
R22829 Y[0].n2 Y[0].n1 1.836
R22830 Y[0] Y[0].n2 1.115
R22831 a_14016_4622.t0 a_14016_4622.t1 380.209
R22832 a_10173_5328.n1 a_10173_5328.t4 318.922
R22833 a_10173_5328.n0 a_10173_5328.t6 273.935
R22834 a_10173_5328.n0 a_10173_5328.t5 273.935
R22835 a_10173_5328.n1 a_10173_5328.t7 269.116
R22836 a_10173_5328.n4 a_10173_5328.n3 193.227
R22837 a_10173_5328.t4 a_10173_5328.n0 179.142
R22838 a_10173_5328.n2 a_10173_5328.n1 106.999
R22839 a_10173_5328.n3 a_10173_5328.t1 28.568
R22840 a_10173_5328.n4 a_10173_5328.t0 28.565
R22841 a_10173_5328.t2 a_10173_5328.n4 28.565
R22842 a_10173_5328.n2 a_10173_5328.t3 18.149
R22843 a_10173_5328.n3 a_10173_5328.n2 3.726
R22844 a_10472_16406.n0 a_10472_16406.t4 14.282
R22845 a_10472_16406.n0 a_10472_16406.t0 14.282
R22846 a_10472_16406.n1 a_10472_16406.t1 14.282
R22847 a_10472_16406.n1 a_10472_16406.t2 14.282
R22848 a_10472_16406.n3 a_10472_16406.t5 14.282
R22849 a_10472_16406.t3 a_10472_16406.n3 14.282
R22850 a_10472_16406.n3 a_10472_16406.n2 2.554
R22851 a_10472_16406.n2 a_10472_16406.n1 2.361
R22852 a_10472_16406.n2 a_10472_16406.n0 0.001
R22853 a_48544_24202.n0 a_48544_24202.t4 14.282
R22854 a_48544_24202.n0 a_48544_24202.t1 14.282
R22855 a_48544_24202.n1 a_48544_24202.t5 14.282
R22856 a_48544_24202.n1 a_48544_24202.t3 14.282
R22857 a_48544_24202.t2 a_48544_24202.n3 14.282
R22858 a_48544_24202.n3 a_48544_24202.t0 14.282
R22859 a_48544_24202.n3 a_48544_24202.n2 2.546
R22860 a_48544_24202.n2 a_48544_24202.n1 2.367
R22861 a_48544_24202.n2 a_48544_24202.n0 0.001
R22862 a_35241_6827.t0 a_35241_6827.t1 17.4
R22863 a_48502_n1313.t0 a_48502_n1313.t1 17.4
R22864 a_13120_14458.n2 a_13120_14458.t5 867.497
R22865 a_13120_14458.n2 a_13120_14458.t7 591.811
R22866 a_13120_14458.n1 a_13120_14458.t4 286.438
R22867 a_13120_14458.n1 a_13120_14458.t6 286.438
R22868 a_13120_14458.n4 a_13120_14458.n0 185.55
R22869 a_13120_14458.t5 a_13120_14458.n1 160.666
R22870 a_13120_14458.t2 a_13120_14458.n4 28.568
R22871 a_13120_14458.n0 a_13120_14458.t0 28.565
R22872 a_13120_14458.n0 a_13120_14458.t1 28.565
R22873 a_13120_14458.n3 a_13120_14458.n2 25.767
R22874 a_13120_14458.n3 a_13120_14458.t3 21.376
R22875 a_13120_14458.n4 a_13120_14458.n3 1.64
R22876 a_8130_16410.n1 a_8130_16410.t5 14.282
R22877 a_8130_16410.n1 a_8130_16410.t0 14.282
R22878 a_8130_16410.n0 a_8130_16410.t3 14.282
R22879 a_8130_16410.n0 a_8130_16410.t4 14.282
R22880 a_8130_16410.n3 a_8130_16410.t1 14.282
R22881 a_8130_16410.t2 a_8130_16410.n3 14.282
R22882 a_8130_16410.n2 a_8130_16410.n0 2.538
R22883 a_8130_16410.n3 a_8130_16410.n2 2.375
R22884 a_8130_16410.n2 a_8130_16410.n1 0.001
R22885 a_71846_8249.t0 a_71846_8249.t1 17.4
R22886 a_10199_n2174.n1 a_10199_n2174.t4 990.34
R22887 a_10199_n2174.n1 a_10199_n2174.t6 408.211
R22888 a_10199_n2174.n0 a_10199_n2174.t7 286.438
R22889 a_10199_n2174.n0 a_10199_n2174.t5 286.438
R22890 a_10199_n2174.n4 a_10199_n2174.n3 185.55
R22891 a_10199_n2174.t4 a_10199_n2174.n0 160.666
R22892 a_10199_n2174.n2 a_10199_n2174.n1 35.738
R22893 a_10199_n2174.n3 a_10199_n2174.t1 28.568
R22894 a_10199_n2174.t2 a_10199_n2174.n4 28.565
R22895 a_10199_n2174.n4 a_10199_n2174.t0 28.565
R22896 a_10199_n2174.n2 a_10199_n2174.t3 21.376
R22897 a_10199_n2174.n3 a_10199_n2174.n2 1.637
R22898 a_38131_3365.t0 a_38131_3365.t1 17.4
R22899 a_62778_24205.n0 a_62778_24205.t4 14.282
R22900 a_62778_24205.n0 a_62778_24205.t0 14.282
R22901 a_62778_24205.n1 a_62778_24205.t5 14.282
R22902 a_62778_24205.n1 a_62778_24205.t3 14.282
R22903 a_62778_24205.n3 a_62778_24205.t1 14.282
R22904 a_62778_24205.t2 a_62778_24205.n3 14.282
R22905 a_62778_24205.n3 a_62778_24205.n2 2.546
R22906 a_62778_24205.n2 a_62778_24205.n1 2.367
R22907 a_62778_24205.n2 a_62778_24205.n0 0.001
R22908 a_54960_24197.t5 a_54960_24197.n3 404.877
R22909 a_54960_24197.n2 a_54960_24197.t8 210.902
R22910 a_54960_24197.n4 a_54960_24197.t5 136.943
R22911 a_54960_24197.n3 a_54960_24197.n2 107.801
R22912 a_54960_24197.n2 a_54960_24197.t7 80.333
R22913 a_54960_24197.n3 a_54960_24197.t6 80.333
R22914 a_54960_24197.n1 a_54960_24197.t0 17.4
R22915 a_54960_24197.n1 a_54960_24197.t4 17.4
R22916 a_54960_24197.t1 a_54960_24197.n5 15.032
R22917 a_54960_24197.n0 a_54960_24197.t3 14.282
R22918 a_54960_24197.n0 a_54960_24197.t2 14.282
R22919 a_54960_24197.n5 a_54960_24197.n0 1.65
R22920 a_54960_24197.n4 a_54960_24197.n1 0.672
R22921 a_54960_24197.n5 a_54960_24197.n4 0.665
R22922 a_56438_21365.n2 a_56438_21365.n0 267.767
R22923 a_56438_21365.n6 a_56438_21365.t5 16.058
R22924 a_56438_21365.n4 a_56438_21365.t7 16.058
R22925 a_56438_21365.n5 a_56438_21365.t3 14.282
R22926 a_56438_21365.n5 a_56438_21365.t4 14.282
R22927 a_56438_21365.n3 a_56438_21365.t6 14.282
R22928 a_56438_21365.n3 a_56438_21365.t8 14.282
R22929 a_56438_21365.n1 a_56438_21365.t9 14.282
R22930 a_56438_21365.n1 a_56438_21365.t0 14.282
R22931 a_56438_21365.n0 a_56438_21365.t10 14.282
R22932 a_56438_21365.n0 a_56438_21365.t11 14.282
R22933 a_56438_21365.n9 a_56438_21365.t1 14.282
R22934 a_56438_21365.t2 a_56438_21365.n9 14.282
R22935 a_56438_21365.n9 a_56438_21365.n8 1.511
R22936 a_56438_21365.n6 a_56438_21365.n5 0.999
R22937 a_56438_21365.n4 a_56438_21365.n3 0.999
R22938 a_56438_21365.n8 a_56438_21365.n2 0.669
R22939 a_56438_21365.n7 a_56438_21365.n6 0.575
R22940 a_56438_21365.n8 a_56438_21365.n7 0.227
R22941 a_56438_21365.n7 a_56438_21365.n4 0.2
R22942 a_56438_21365.n2 a_56438_21365.n1 0.001
R22943 a_49977_18084.t0 a_49977_18084.t1 17.4
R22944 a_42031_24205.n0 a_42031_24205.t0 14.282
R22945 a_42031_24205.n0 a_42031_24205.t1 14.282
R22946 a_42031_24205.n1 a_42031_24205.t3 14.282
R22947 a_42031_24205.n1 a_42031_24205.t4 14.282
R22948 a_42031_24205.n3 a_42031_24205.t5 14.282
R22949 a_42031_24205.t2 a_42031_24205.n3 14.282
R22950 a_42031_24205.n2 a_42031_24205.n0 2.546
R22951 a_42031_24205.n2 a_42031_24205.n1 2.367
R22952 a_42031_24205.n3 a_42031_24205.n2 0.001
R22953 Y[7].n1 Y[7].n0 185.55
R22954 Y[7].n1 Y[7].t0 28.568
R22955 Y[7].n0 Y[7].t1 28.565
R22956 Y[7].n0 Y[7].t2 28.565
R22957 Y[7].n2 Y[7].t3 20.393
R22958 Y[7].n2 Y[7].n1 2.161
R22959 Y[7] Y[7].n2 1.127
R22960 a_53352_20634.t4 a_53352_20634.t7 574.43
R22961 a_53352_20634.n0 a_53352_20634.t6 285.109
R22962 a_53352_20634.n2 a_53352_20634.n1 197.217
R22963 a_53352_20634.n4 a_53352_20634.n3 192.754
R22964 a_53352_20634.n0 a_53352_20634.t5 160.666
R22965 a_53352_20634.n1 a_53352_20634.t4 160.666
R22966 a_53352_20634.n1 a_53352_20634.n0 114.829
R22967 a_53352_20634.n3 a_53352_20634.t0 28.568
R22968 a_53352_20634.n4 a_53352_20634.t1 28.565
R22969 a_53352_20634.t2 a_53352_20634.n4 28.565
R22970 a_53352_20634.n2 a_53352_20634.t3 18.838
R22971 a_53352_20634.n3 a_53352_20634.n2 1.129
R22972 a_19677_n2174.n1 a_19677_n2174.t5 990.34
R22973 a_19677_n2174.n1 a_19677_n2174.t6 408.211
R22974 a_19677_n2174.n0 a_19677_n2174.t4 286.438
R22975 a_19677_n2174.n0 a_19677_n2174.t7 286.438
R22976 a_19677_n2174.n4 a_19677_n2174.n3 185.55
R22977 a_19677_n2174.t5 a_19677_n2174.n0 160.666
R22978 a_19677_n2174.n2 a_19677_n2174.n1 48.757
R22979 a_19677_n2174.n3 a_19677_n2174.t0 28.568
R22980 a_19677_n2174.n4 a_19677_n2174.t1 28.565
R22981 a_19677_n2174.t2 a_19677_n2174.n4 28.565
R22982 a_19677_n2174.n2 a_19677_n2174.t3 21.376
R22983 a_19677_n2174.n3 a_19677_n2174.n2 1.637
R22984 a_71842_n1171.t0 a_71842_n1171.t1 17.4
R22985 a_30150_n3032.n1 a_30150_n3032.t5 318.119
R22986 a_30150_n3032.n1 a_30150_n3032.t6 269.919
R22987 a_30150_n3032.n0 a_30150_n3032.t4 267.853
R22988 a_30150_n3032.n0 a_30150_n3032.t7 267.853
R22989 a_30150_n3032.t5 a_30150_n3032.n0 160.666
R22990 a_30150_n3032.n2 a_30150_n3032.n1 107.263
R22991 a_30150_n3032.t2 a_30150_n3032.n4 29.444
R22992 a_30150_n3032.n3 a_30150_n3032.t1 28.565
R22993 a_30150_n3032.n3 a_30150_n3032.t0 28.565
R22994 a_30150_n3032.n2 a_30150_n3032.t3 18.145
R22995 a_30150_n3032.n4 a_30150_n3032.n2 2.878
R22996 a_30150_n3032.n4 a_30150_n3032.n3 0.764
R22997 a_51356_7515.t0 a_51356_7515.t1 17.4
R22998 a_60226_16462.n1 a_60226_16462.t6 318.922
R22999 a_60226_16462.n0 a_60226_16462.t5 274.739
R23000 a_60226_16462.n0 a_60226_16462.t4 274.739
R23001 a_60226_16462.n1 a_60226_16462.t7 269.116
R23002 a_60226_16462.t6 a_60226_16462.n0 179.946
R23003 a_60226_16462.n2 a_60226_16462.n1 107.263
R23004 a_60226_16462.n3 a_60226_16462.t0 29.444
R23005 a_60226_16462.n4 a_60226_16462.t1 28.565
R23006 a_60226_16462.t2 a_60226_16462.n4 28.565
R23007 a_60226_16462.n2 a_60226_16462.t3 18.145
R23008 a_60226_16462.n3 a_60226_16462.n2 2.878
R23009 a_60226_16462.n4 a_60226_16462.n3 0.764
R23010 a_35222_3549.t0 a_35222_3549.t1 17.4
R23011 a_60988_7603.n1 a_60988_7603.t4 318.922
R23012 a_60988_7603.n0 a_60988_7603.t6 273.935
R23013 a_60988_7603.n0 a_60988_7603.t5 273.935
R23014 a_60988_7603.n1 a_60988_7603.t7 269.116
R23015 a_60988_7603.n4 a_60988_7603.n3 193.227
R23016 a_60988_7603.t4 a_60988_7603.n0 179.142
R23017 a_60988_7603.n2 a_60988_7603.n1 106.999
R23018 a_60988_7603.n3 a_60988_7603.t0 28.568
R23019 a_60988_7603.t2 a_60988_7603.n4 28.565
R23020 a_60988_7603.n4 a_60988_7603.t1 28.565
R23021 a_60988_7603.n2 a_60988_7603.t3 18.149
R23022 a_60988_7603.n3 a_60988_7603.n2 3.726
R23023 a_14046_n3485.t0 a_14046_n3485.t1 17.4
R23024 a_21211_16387.n0 a_21211_16387.t7 214.335
R23025 a_21211_16387.t10 a_21211_16387.n0 214.335
R23026 a_21211_16387.n1 a_21211_16387.t10 143.851
R23027 a_21211_16387.n1 a_21211_16387.t8 135.658
R23028 a_21211_16387.n0 a_21211_16387.t9 80.333
R23029 a_21211_16387.n4 a_21211_16387.t4 28.565
R23030 a_21211_16387.n4 a_21211_16387.t5 28.565
R23031 a_21211_16387.n2 a_21211_16387.t0 28.565
R23032 a_21211_16387.n2 a_21211_16387.t1 28.565
R23033 a_21211_16387.n7 a_21211_16387.t3 28.565
R23034 a_21211_16387.t2 a_21211_16387.n7 28.565
R23035 a_21211_16387.n5 a_21211_16387.t6 9.714
R23036 a_21211_16387.n5 a_21211_16387.n4 1.003
R23037 a_21211_16387.n6 a_21211_16387.n3 0.833
R23038 a_21211_16387.n3 a_21211_16387.n2 0.653
R23039 a_21211_16387.n7 a_21211_16387.n6 0.653
R23040 a_21211_16387.n6 a_21211_16387.n5 0.341
R23041 a_21211_16387.n3 a_21211_16387.n1 0.032
R23042 a_4879_13585.n2 a_4879_13585.t6 448.381
R23043 a_4879_13585.n1 a_4879_13585.t5 286.438
R23044 a_4879_13585.n1 a_4879_13585.t7 286.438
R23045 a_4879_13585.n0 a_4879_13585.t4 247.69
R23046 a_4879_13585.n4 a_4879_13585.n3 182.117
R23047 a_4879_13585.t6 a_4879_13585.n1 160.666
R23048 a_4879_13585.n3 a_4879_13585.t1 28.568
R23049 a_4879_13585.t2 a_4879_13585.n4 28.565
R23050 a_4879_13585.n4 a_4879_13585.t0 28.565
R23051 a_4879_13585.n0 a_4879_13585.t3 18.127
R23052 a_4879_13585.n2 a_4879_13585.n0 4.036
R23053 a_4879_13585.n3 a_4879_13585.n2 0.937
R23054 Y[2].n1 Y[2].n0 185.55
R23055 Y[2].n1 Y[2].t0 28.568
R23056 Y[2].n0 Y[2].t1 28.565
R23057 Y[2].n0 Y[2].t2 28.565
R23058 Y[2].n2 Y[2].t3 20.393
R23059 Y[2].n2 Y[2].n1 2.941
R23060 Y[2] Y[2].n2 2.613
R23061 a_9304_16408.n0 a_9304_16408.t0 14.282
R23062 a_9304_16408.n0 a_9304_16408.t3 14.282
R23063 a_9304_16408.n1 a_9304_16408.t4 14.282
R23064 a_9304_16408.n1 a_9304_16408.t5 14.282
R23065 a_9304_16408.n3 a_9304_16408.t1 14.282
R23066 a_9304_16408.t2 a_9304_16408.n3 14.282
R23067 a_9304_16408.n3 a_9304_16408.n2 2.538
R23068 a_9304_16408.n2 a_9304_16408.n1 2.375
R23069 a_9304_16408.n2 a_9304_16408.n0 0.001
R23070 a_55224_23614.t4 a_55224_23614.t7 800.071
R23071 a_55224_23614.n3 a_55224_23614.n2 672.951
R23072 a_55224_23614.n1 a_55224_23614.t6 285.109
R23073 a_55224_23614.n2 a_55224_23614.t4 193.602
R23074 a_55224_23614.n1 a_55224_23614.t5 160.666
R23075 a_55224_23614.n2 a_55224_23614.n1 91.507
R23076 a_55224_23614.t2 a_55224_23614.n4 28.57
R23077 a_55224_23614.n0 a_55224_23614.t0 28.565
R23078 a_55224_23614.n0 a_55224_23614.t1 28.565
R23079 a_55224_23614.n4 a_55224_23614.t3 17.638
R23080 a_55224_23614.n3 a_55224_23614.n0 0.69
R23081 a_55224_23614.n4 a_55224_23614.n3 0.6
R23082 a_10458_20259.t0 a_10458_20259.t1 17.4
R23083 a_12241_5326.n1 a_12241_5326.t4 318.922
R23084 a_12241_5326.n0 a_12241_5326.t6 273.935
R23085 a_12241_5326.n0 a_12241_5326.t7 273.935
R23086 a_12241_5326.n1 a_12241_5326.t5 269.116
R23087 a_12241_5326.n4 a_12241_5326.n3 193.227
R23088 a_12241_5326.t4 a_12241_5326.n0 179.142
R23089 a_12241_5326.n2 a_12241_5326.n1 106.999
R23090 a_12241_5326.n3 a_12241_5326.t0 28.568
R23091 a_12241_5326.t2 a_12241_5326.n4 28.565
R23092 a_12241_5326.n4 a_12241_5326.t1 28.565
R23093 a_12241_5326.n2 a_12241_5326.t3 18.149
R23094 a_12241_5326.n3 a_12241_5326.n2 3.726
R23095 a_38148_5891.t0 a_38148_5891.t1 17.4
R23096 a_61510_21343.n1 a_61510_21343.t6 318.922
R23097 a_61510_21343.n0 a_61510_21343.t5 274.739
R23098 a_61510_21343.n0 a_61510_21343.t7 274.739
R23099 a_61510_21343.n1 a_61510_21343.t4 269.116
R23100 a_61510_21343.t6 a_61510_21343.n0 179.946
R23101 a_61510_21343.n2 a_61510_21343.n1 107.263
R23102 a_61510_21343.n3 a_61510_21343.t0 29.444
R23103 a_61510_21343.n4 a_61510_21343.t1 28.565
R23104 a_61510_21343.t2 a_61510_21343.n4 28.565
R23105 a_61510_21343.n2 a_61510_21343.t3 18.145
R23106 a_61510_21343.n3 a_61510_21343.n2 2.878
R23107 a_61510_21343.n4 a_61510_21343.n3 0.764
R23108 a_4536_407.t0 a_4536_407.t1 17.4
R23109 a_60047_3874.n0 a_60047_3874.t5 14.282
R23110 a_60047_3874.n0 a_60047_3874.t2 14.282
R23111 a_60047_3874.n1 a_60047_3874.t4 14.282
R23112 a_60047_3874.n1 a_60047_3874.t3 14.282
R23113 a_60047_3874.t0 a_60047_3874.n3 14.282
R23114 a_60047_3874.n3 a_60047_3874.t1 14.282
R23115 a_60047_3874.n3 a_60047_3874.n2 2.546
R23116 a_60047_3874.n2 a_60047_3874.n1 2.367
R23117 a_60047_3874.n2 a_60047_3874.n0 0.001
R23118 a_45044_309.t4 a_45044_309.t5 574.43
R23119 a_45044_309.n1 a_45044_309.t6 285.109
R23120 a_45044_309.n3 a_45044_309.n2 197.217
R23121 a_45044_309.n4 a_45044_309.n0 192.754
R23122 a_45044_309.n1 a_45044_309.t7 160.666
R23123 a_45044_309.n2 a_45044_309.t4 160.666
R23124 a_45044_309.n2 a_45044_309.n1 114.829
R23125 a_45044_309.t2 a_45044_309.n4 28.568
R23126 a_45044_309.n0 a_45044_309.t1 28.565
R23127 a_45044_309.n0 a_45044_309.t0 28.565
R23128 a_45044_309.n3 a_45044_309.t3 18.838
R23129 a_45044_309.n4 a_45044_309.n3 1.129
R23130 a_4491_15753.t7 a_4491_15753.n3 406.651
R23131 a_4491_15753.n2 a_4491_15753.t8 207.856
R23132 a_4491_15753.n4 a_4491_15753.t7 136.949
R23133 a_4491_15753.n3 a_4491_15753.n2 111.349
R23134 a_4491_15753.n2 a_4491_15753.t5 80.333
R23135 a_4491_15753.n3 a_4491_15753.t6 80.333
R23136 a_4491_15753.n1 a_4491_15753.t4 17.4
R23137 a_4491_15753.n1 a_4491_15753.t0 17.4
R23138 a_4491_15753.t1 a_4491_15753.n5 15.029
R23139 a_4491_15753.n0 a_4491_15753.t2 14.282
R23140 a_4491_15753.n0 a_4491_15753.t3 14.282
R23141 a_4491_15753.n5 a_4491_15753.n0 1.647
R23142 a_4491_15753.n4 a_4491_15753.n1 0.657
R23143 a_4491_15753.n5 a_4491_15753.n4 0.614
R23144 a_8202_7655.t0 a_8202_7655.t1 17.4
R23145 a_23358_15774.t0 a_23358_15774.t1 17.4
R23146 a_20086_n2148.n2 a_20086_n2148.t11 1527.4
R23147 a_20086_n2148.t11 a_20086_n2148.n1 657.379
R23148 a_20086_n2148.n4 a_20086_n2148.n3 258.161
R23149 a_20086_n2148.n7 a_20086_n2148.n6 258.161
R23150 a_20086_n2148.n0 a_20086_n2148.t8 206.421
R23151 a_20086_n2148.t10 a_20086_n2148.n0 206.421
R23152 a_20086_n2148.n2 a_20086_n2148.t10 200.029
R23153 a_20086_n2148.n5 a_20086_n2148.n2 97.614
R23154 a_20086_n2148.n0 a_20086_n2148.t9 80.333
R23155 a_20086_n2148.n4 a_20086_n2148.t5 14.283
R23156 a_20086_n2148.n6 a_20086_n2148.t0 14.283
R23157 a_20086_n2148.n3 a_20086_n2148.t3 14.282
R23158 a_20086_n2148.n3 a_20086_n2148.t4 14.282
R23159 a_20086_n2148.n7 a_20086_n2148.t1 14.282
R23160 a_20086_n2148.t2 a_20086_n2148.n7 14.282
R23161 a_20086_n2148.n1 a_20086_n2148.t6 8.7
R23162 a_20086_n2148.n1 a_20086_n2148.t7 8.7
R23163 a_20086_n2148.n5 a_20086_n2148.n4 4.366
R23164 a_20086_n2148.n6 a_20086_n2148.n5 0.852
R23165 a_67372_3171.t0 a_67372_3171.t1 17.4
R23166 a_63114_21369.n0 a_63114_21369.n8 122.999
R23167 a_63114_21369.n0 a_63114_21369.t7 14.282
R23168 a_63114_21369.t1 a_63114_21369.n0 14.282
R23169 a_63114_21369.n8 a_63114_21369.n6 50.575
R23170 a_63114_21369.n6 a_63114_21369.n4 74.302
R23171 a_63114_21369.n8 a_63114_21369.n7 157.665
R23172 a_63114_21369.n7 a_63114_21369.t6 8.7
R23173 a_63114_21369.n7 a_63114_21369.t0 8.7
R23174 a_63114_21369.n6 a_63114_21369.n5 90.416
R23175 a_63114_21369.n5 a_63114_21369.t2 14.282
R23176 a_63114_21369.n5 a_63114_21369.t5 14.282
R23177 a_63114_21369.n4 a_63114_21369.n3 90.436
R23178 a_63114_21369.n3 a_63114_21369.t4 14.282
R23179 a_63114_21369.n3 a_63114_21369.t3 14.282
R23180 a_63114_21369.n4 a_63114_21369.n1 449.112
R23181 a_63114_21369.t8 a_63114_21369.n2 160.666
R23182 a_63114_21369.n1 a_63114_21369.t8 867.393
R23183 a_63114_21369.n2 a_63114_21369.t11 287.241
R23184 a_63114_21369.n2 a_63114_21369.t9 287.241
R23185 a_63114_21369.n1 a_63114_21369.t10 545.094
R23186 a_58321_311.t4 a_58321_311.t6 574.43
R23187 a_58321_311.n0 a_58321_311.t5 285.109
R23188 a_58321_311.n2 a_58321_311.n1 197.217
R23189 a_58321_311.n4 a_58321_311.n3 192.754
R23190 a_58321_311.n0 a_58321_311.t7 160.666
R23191 a_58321_311.n1 a_58321_311.t4 160.666
R23192 a_58321_311.n1 a_58321_311.n0 114.829
R23193 a_58321_311.n3 a_58321_311.t1 28.568
R23194 a_58321_311.t2 a_58321_311.n4 28.565
R23195 a_58321_311.n4 a_58321_311.t0 28.565
R23196 a_58321_311.n2 a_58321_311.t3 18.838
R23197 a_58321_311.n3 a_58321_311.n2 1.129
R23198 a_52767_22675.n0 a_52767_22675.t9 214.335
R23199 a_52767_22675.t7 a_52767_22675.n0 214.335
R23200 a_52767_22675.n1 a_52767_22675.t7 143.851
R23201 a_52767_22675.n1 a_52767_22675.t10 135.658
R23202 a_52767_22675.n0 a_52767_22675.t8 80.333
R23203 a_52767_22675.n2 a_52767_22675.t4 28.565
R23204 a_52767_22675.n2 a_52767_22675.t5 28.565
R23205 a_52767_22675.n4 a_52767_22675.t6 28.565
R23206 a_52767_22675.n4 a_52767_22675.t0 28.565
R23207 a_52767_22675.n7 a_52767_22675.t1 28.565
R23208 a_52767_22675.t2 a_52767_22675.n7 28.565
R23209 a_52767_22675.n6 a_52767_22675.t3 9.714
R23210 a_52767_22675.n7 a_52767_22675.n6 1.003
R23211 a_52767_22675.n5 a_52767_22675.n3 0.833
R23212 a_52767_22675.n3 a_52767_22675.n2 0.653
R23213 a_52767_22675.n5 a_52767_22675.n4 0.653
R23214 a_52767_22675.n6 a_52767_22675.n5 0.341
R23215 a_52767_22675.n3 a_52767_22675.n1 0.032
R23216 a_17158_407.t0 a_17158_407.t1 17.4
R23217 a_14250_407.t0 a_14250_407.t1 17.4
R23218 a_38145_1715.t0 a_38145_1715.t1 17.4
R23219 a_50258_20638.t0 a_50258_20638.t1 17.4
R23220 a_5070_7659.t0 a_5070_7659.t1 17.4
R23221 a_61533_6178.t0 a_61533_6178.t1 380.209
R23222 a_20457_4618.t0 a_20457_4618.t1 17.4
R23223 a_10513_20719.n2 a_10513_20719.t6 448.381
R23224 a_10513_20719.n1 a_10513_20719.t5 286.438
R23225 a_10513_20719.n1 a_10513_20719.t7 286.438
R23226 a_10513_20719.n0 a_10513_20719.t4 247.69
R23227 a_10513_20719.n4 a_10513_20719.n3 182.117
R23228 a_10513_20719.t6 a_10513_20719.n1 160.666
R23229 a_10513_20719.n3 a_10513_20719.t0 28.568
R23230 a_10513_20719.n4 a_10513_20719.t1 28.565
R23231 a_10513_20719.t2 a_10513_20719.n4 28.565
R23232 a_10513_20719.n0 a_10513_20719.t3 18.127
R23233 a_10513_20719.n2 a_10513_20719.n0 4.036
R23234 a_10513_20719.n3 a_10513_20719.n2 0.937
R23235 a_48131_15735.n1 a_48131_15735.t5 318.922
R23236 a_48131_15735.n0 a_48131_15735.t4 273.935
R23237 a_48131_15735.n0 a_48131_15735.t6 273.935
R23238 a_48131_15735.n1 a_48131_15735.t7 269.116
R23239 a_48131_15735.n4 a_48131_15735.n3 193.227
R23240 a_48131_15735.t5 a_48131_15735.n0 179.142
R23241 a_48131_15735.n2 a_48131_15735.n1 106.999
R23242 a_48131_15735.n3 a_48131_15735.t0 28.568
R23243 a_48131_15735.n4 a_48131_15735.t1 28.565
R23244 a_48131_15735.t2 a_48131_15735.n4 28.565
R23245 a_48131_15735.n2 a_48131_15735.t3 18.149
R23246 a_48131_15735.n3 a_48131_15735.n2 3.726
R23247 a_1628_407.t0 a_1628_407.t1 17.4
R23248 a_48360_20638.t0 a_48360_20638.t1 17.4
R23249 a_13838_20259.t0 a_13838_20259.t1 17.4
R23250 a_20824_7655.t0 a_20824_7655.t1 17.4
R23251 a_55151_n1325.t0 a_55151_n1325.t1 17.4
R23252 a_71846_20635.t0 a_71846_20635.t1 17.4
R23253 a_10337_15751.t5 a_10337_15751.n2 404.877
R23254 a_10337_15751.n1 a_10337_15751.t6 210.902
R23255 a_10337_15751.n3 a_10337_15751.t5 136.949
R23256 a_10337_15751.n2 a_10337_15751.n1 107.801
R23257 a_10337_15751.n1 a_10337_15751.t7 80.333
R23258 a_10337_15751.n2 a_10337_15751.t8 80.333
R23259 a_10337_15751.n0 a_10337_15751.t1 17.4
R23260 a_10337_15751.n0 a_10337_15751.t0 17.4
R23261 a_10337_15751.n4 a_10337_15751.t2 15.029
R23262 a_10337_15751.n5 a_10337_15751.t3 14.282
R23263 a_10337_15751.t4 a_10337_15751.n5 14.282
R23264 a_10337_15751.n5 a_10337_15751.n4 1.647
R23265 a_10337_15751.n3 a_10337_15751.n0 0.657
R23266 a_10337_15751.n4 a_10337_15751.n3 0.614
R23267 a_54908_6110.t0 a_54908_6110.t1 380.209
R23268 a_11336_10387.t0 a_11336_10387.t1 17.4
R23269 a_57976_5979.t0 a_57976_5979.t1 17.4
R23270 a_4824_10391.t0 a_4824_10391.t1 17.4
R23271 a_17444_15774.t0 a_17444_15774.t1 17.4
R23272 a_55144_6110.t0 a_55144_6110.t1 17.4
R23273 a_39657_18575.t6 a_39657_18575.t7 800.071
R23274 a_39657_18575.n3 a_39657_18575.n2 672.95
R23275 a_39657_18575.n1 a_39657_18575.t4 285.109
R23276 a_39657_18575.n2 a_39657_18575.t6 193.602
R23277 a_39657_18575.n1 a_39657_18575.t5 160.666
R23278 a_39657_18575.n2 a_39657_18575.n1 91.507
R23279 a_39657_18575.n0 a_39657_18575.t0 28.57
R23280 a_39657_18575.n4 a_39657_18575.t1 28.565
R23281 a_39657_18575.t2 a_39657_18575.n4 28.565
R23282 a_39657_18575.n0 a_39657_18575.t3 17.638
R23283 a_39657_18575.n4 a_39657_18575.n3 0.693
R23284 a_39657_18575.n3 a_39657_18575.n0 0.597
R23285 a_4626_16408.n1 a_4626_16408.t5 14.282
R23286 a_4626_16408.n1 a_4626_16408.t0 14.282
R23287 a_4626_16408.n0 a_4626_16408.t3 14.282
R23288 a_4626_16408.n0 a_4626_16408.t4 14.282
R23289 a_4626_16408.n3 a_4626_16408.t1 14.282
R23290 a_4626_16408.t2 a_4626_16408.n3 14.282
R23291 a_4626_16408.n2 a_4626_16408.n0 2.554
R23292 a_4626_16408.n3 a_4626_16408.n2 2.361
R23293 a_4626_16408.n2 a_4626_16408.n1 0.001
R23294 a_47837_15029.t0 a_47837_15029.t1 380.209
R23295 a_10812_411.t0 a_10812_411.t1 17.4
R23296 a_57973_1715.t0 a_57973_1715.t1 17.4
R23297 a_1660_n3485.t0 a_1660_n3485.t1 17.4
R23298 a_38153_7495.t0 a_38153_7495.t1 17.4
R23299 Y[6].n1 Y[6].n0 185.55
R23300 Y[6].n1 Y[6].t1 28.568
R23301 Y[6].n0 Y[6].t2 28.565
R23302 Y[6].n0 Y[6].t0 28.565
R23303 Y[6].n2 Y[6].t3 20.393
R23304 Y[6].n2 Y[6].n1 1.831
R23305 Y[6] Y[6].n2 1.125
R23306 a_4173_14432.n2 a_4173_14432.t7 867.497
R23307 a_4173_14432.n2 a_4173_14432.t4 591.811
R23308 a_4173_14432.n1 a_4173_14432.t6 286.438
R23309 a_4173_14432.n1 a_4173_14432.t5 286.438
R23310 a_4173_14432.n4 a_4173_14432.n0 192.754
R23311 a_4173_14432.t7 a_4173_14432.n1 160.666
R23312 a_4173_14432.n3 a_4173_14432.n2 36.159
R23313 a_4173_14432.t2 a_4173_14432.n4 28.568
R23314 a_4173_14432.n0 a_4173_14432.t0 28.565
R23315 a_4173_14432.n0 a_4173_14432.t1 28.565
R23316 a_4173_14432.n3 a_4173_14432.t3 18.726
R23317 a_4173_14432.n4 a_4173_14432.n3 1.123
R23318 a_4824_13125.t0 a_4824_13125.t1 17.4
R23319 a_11100_13121.t0 a_11100_13121.t1 17.4
R23320 a_24358_4618.t0 a_24358_4618.t1 380.209
R23321 a_22821_n2174.n2 a_22821_n2174.t7 990.34
R23322 a_22821_n2174.n2 a_22821_n2174.t4 408.211
R23323 a_22821_n2174.n1 a_22821_n2174.t5 286.438
R23324 a_22821_n2174.n1 a_22821_n2174.t6 286.438
R23325 a_22821_n2174.n4 a_22821_n2174.n0 185.55
R23326 a_22821_n2174.t7 a_22821_n2174.n1 160.666
R23327 a_22821_n2174.n3 a_22821_n2174.n2 50.538
R23328 a_22821_n2174.t2 a_22821_n2174.n4 28.568
R23329 a_22821_n2174.n0 a_22821_n2174.t0 28.565
R23330 a_22821_n2174.n0 a_22821_n2174.t1 28.565
R23331 a_22821_n2174.n3 a_22821_n2174.t3 21.701
R23332 a_22821_n2174.n4 a_22821_n2174.n3 1.618
R23333 a_40227_9654.n0 a_40227_9654.t5 14.282
R23334 a_40227_9654.n0 a_40227_9654.t4 14.282
R23335 a_40227_9654.n1 a_40227_9654.t1 14.282
R23336 a_40227_9654.n1 a_40227_9654.t0 14.282
R23337 a_40227_9654.t2 a_40227_9654.n3 14.282
R23338 a_40227_9654.n3 a_40227_9654.t3 14.282
R23339 a_40227_9654.n2 a_40227_9654.n0 2.546
R23340 a_40227_9654.n2 a_40227_9654.n1 2.367
R23341 a_40227_9654.n3 a_40227_9654.n2 0.001
R23342 a_14312_7659.t0 a_14312_7659.t1 17.4
R23343 a_41611_20641.t0 a_41611_20641.t1 380.209
R23344 a_51351_1714.t0 a_51351_1714.t1 17.4
R23345 a_43419_18088.t0 a_43419_18088.t1 17.4
R23346 a_66063_n1256.n1 a_66063_n1256.t5 318.922
R23347 a_66063_n1256.n0 a_66063_n1256.t4 274.739
R23348 a_66063_n1256.n0 a_66063_n1256.t7 274.739
R23349 a_66063_n1256.n1 a_66063_n1256.t6 269.116
R23350 a_66063_n1256.t5 a_66063_n1256.n0 179.946
R23351 a_66063_n1256.n2 a_66063_n1256.n1 107.263
R23352 a_66063_n1256.n3 a_66063_n1256.t0 29.444
R23353 a_66063_n1256.t2 a_66063_n1256.n4 28.565
R23354 a_66063_n1256.n4 a_66063_n1256.t1 28.565
R23355 a_66063_n1256.n2 a_66063_n1256.t3 18.145
R23356 a_66063_n1256.n3 a_66063_n1256.n2 2.878
R23357 a_66063_n1256.n4 a_66063_n1256.n3 0.764
R23358 a_39381_15033.t0 a_39381_15033.t1 380.209
R23359 a_62569_22062.n2 a_62569_22062.t6 318.922
R23360 a_62569_22062.n1 a_62569_22062.t5 273.935
R23361 a_62569_22062.n1 a_62569_22062.t7 273.935
R23362 a_62569_22062.n2 a_62569_22062.t4 269.116
R23363 a_62569_22062.n4 a_62569_22062.n0 193.227
R23364 a_62569_22062.t6 a_62569_22062.n1 179.142
R23365 a_62569_22062.n3 a_62569_22062.n2 106.999
R23366 a_62569_22062.t2 a_62569_22062.n4 28.568
R23367 a_62569_22062.n0 a_62569_22062.t0 28.565
R23368 a_62569_22062.n0 a_62569_22062.t1 28.565
R23369 a_62569_22062.n3 a_62569_22062.t3 18.149
R23370 a_62569_22062.n4 a_62569_22062.n3 3.726
R23371 a_41847_20641.t0 a_41847_20641.t1 17.4
R23372 a_61216_20637.t0 a_61216_20637.t1 380.209
R23373 a_14252_4622.t0 a_14252_4622.t1 17.4
R23374 a_39617_15033.t0 a_39617_15033.t1 17.4
R23375 a_20221_4618.t0 a_20221_4618.t1 380.209
R23376 a_12183_4620.t0 a_12183_4620.t1 17.4
R23377 a_41941_6090.t0 a_41941_6090.t1 17.4
R23378 a_31379_8204.t0 a_31379_8204.t1 17.4
R23379 a_31377_3831.t0 a_31377_3831.t1 379.845
R23380 a_7904_411.t0 a_7904_411.t1 17.4
R23381 a_71842_11451.t0 a_71842_11451.t1 17.4
R23382 a_39618_16432.n10 a_39618_16432.n8 552.333
R23383 a_39618_16432.n7 a_39618_16432.t14 394.151
R23384 a_39618_16432.n11 a_39618_16432.n10 342.688
R23385 a_39618_16432.n9 a_39618_16432.t8 294.653
R23386 a_39618_16432.n6 a_39618_16432.t11 269.523
R23387 a_39618_16432.t14 a_39618_16432.n6 269.523
R23388 a_39618_16432.n5 a_39618_16432.t15 198.043
R23389 a_39618_16432.n6 a_39618_16432.t12 160.666
R23390 a_39618_16432.n3 a_39618_16432.n1 157.665
R23391 a_39618_16432.n10 a_39618_16432.n9 126.566
R23392 a_39618_16432.n3 a_39618_16432.n2 122.746
R23393 a_39618_16432.n9 a_39618_16432.t13 111.663
R23394 a_39618_16432.n8 a_39618_16432.n7 97.816
R23395 a_39618_16432.n5 a_39618_16432.t10 93.989
R23396 a_39618_16432.n12 a_39618_16432.n11 90.436
R23397 a_39618_16432.n4 a_39618_16432.n0 90.416
R23398 a_39618_16432.n7 a_39618_16432.t9 80.333
R23399 a_39618_16432.n11 a_39618_16432.n4 74.302
R23400 a_39618_16432.n4 a_39618_16432.n3 50.575
R23401 a_39618_16432.n2 a_39618_16432.t7 14.282
R23402 a_39618_16432.n2 a_39618_16432.t5 14.282
R23403 a_39618_16432.n0 a_39618_16432.t6 14.282
R23404 a_39618_16432.n0 a_39618_16432.t1 14.282
R23405 a_39618_16432.n12 a_39618_16432.t2 14.282
R23406 a_39618_16432.t3 a_39618_16432.n12 14.282
R23407 a_39618_16432.n1 a_39618_16432.t4 8.7
R23408 a_39618_16432.n1 a_39618_16432.t0 8.7
R23409 a_39618_16432.n8 a_39618_16432.n5 6.615
R23410 a_46569_18571.t7 a_46569_18571.t6 574.43
R23411 a_46569_18571.n1 a_46569_18571.t4 285.109
R23412 a_46569_18571.n3 a_46569_18571.n2 211.134
R23413 a_46569_18571.n4 a_46569_18571.n0 192.754
R23414 a_46569_18571.n1 a_46569_18571.t5 160.666
R23415 a_46569_18571.n2 a_46569_18571.t7 160.666
R23416 a_46569_18571.n2 a_46569_18571.n1 114.829
R23417 a_46569_18571.t2 a_46569_18571.n4 28.568
R23418 a_46569_18571.n0 a_46569_18571.t0 28.565
R23419 a_46569_18571.n0 a_46569_18571.t1 28.565
R23420 a_46569_18571.n3 a_46569_18571.t3 19.087
R23421 a_46569_18571.n4 a_46569_18571.n3 1.051
R23422 a_63839_n2274.t0 a_63839_n2274.t1 17.4
R23423 a_44688_9233.t0 a_44688_9233.t1 17.4
R23424 Y[3].n1 Y[3].n0 185.55
R23425 Y[3].n1 Y[3].t0 28.568
R23426 Y[3].n0 Y[3].t1 28.565
R23427 Y[3].n0 Y[3].t2 28.565
R23428 Y[3].n2 Y[3].t3 20.393
R23429 Y[3].n2 Y[3].n1 1.831
R23430 Y[3] Y[3].n2 1.126
R23431 a_26224_20259.t0 a_26224_20259.t1 17.4
R23432 a_31377_10273.t0 a_31377_10273.t1 17.4
R23433 a_41279_15033.t0 a_41279_15033.t1 380.209
R23434 a_40035_310.t0 a_40035_310.t1 17.4
R23435 a_20578_13121.t0 a_20578_13121.t1 17.4
R23436 a_63764_8594.t0 a_63764_8594.t1 17.4
R23437 a_54658_20633.t0 a_54658_20633.t1 380.209
R23438 a_8192_10387.t0 a_8192_10387.t1 17.4
R23439 a_14014_407.t0 a_14014_407.t1 17.4
R23440 a_65769_5881.t0 a_65769_5881.t1 380.209
R23441 a_63764_5561.t0 a_63764_5561.t1 17.4
R23442 a_41515_15033.t0 a_41515_15033.t1 17.4
R23443 a_71842_14359.t0 a_71842_14359.t1 17.4
R23444 a_38139_9145.t0 a_38139_9145.t1 17.4
R23445 a_53241_309.t0 a_53241_309.t1 17.4
R23446 a_1029_14432.n1 a_1029_14432.t5 867.497
R23447 a_1029_14432.n1 a_1029_14432.t7 591.811
R23448 a_1029_14432.n0 a_1029_14432.t4 286.438
R23449 a_1029_14432.n0 a_1029_14432.t6 286.438
R23450 a_1029_14432.n4 a_1029_14432.n3 192.754
R23451 a_1029_14432.t5 a_1029_14432.n0 160.666
R23452 a_1029_14432.n2 a_1029_14432.n1 37.908
R23453 a_1029_14432.n3 a_1029_14432.t1 28.568
R23454 a_1029_14432.t2 a_1029_14432.n4 28.565
R23455 a_1029_14432.n4 a_1029_14432.t0 28.565
R23456 a_1029_14432.n2 a_1029_14432.t3 18.726
R23457 a_1029_14432.n3 a_1029_14432.n2 1.123
R23458 a_54371_15034.t0 a_54371_15034.t1 380.209
R23459 a_71846_20871.t0 a_71846_20871.t1 17.4
R23460 a_66005_2386.t0 a_66005_2386.t1 17.4
R23461 a_20322_n3481.t0 a_20322_n3481.t1 17.4
R23462 a_63835_3641.t0 a_63835_3641.t1 17.4
R23463 a_6962_16408.n1 a_6962_16408.t5 14.282
R23464 a_6962_16408.n1 a_6962_16408.t0 14.282
R23465 a_6962_16408.n0 a_6962_16408.t3 14.282
R23466 a_6962_16408.n0 a_6962_16408.t4 14.282
R23467 a_6962_16408.t2 a_6962_16408.n3 14.282
R23468 a_6962_16408.n3 a_6962_16408.t1 14.282
R23469 a_6962_16408.n2 a_6962_16408.n0 2.554
R23470 a_6962_16408.n3 a_6962_16408.n2 2.361
R23471 a_6962_16408.n2 a_6962_16408.n1 0.001
R23472 a_63832_571.t0 a_63832_571.t1 17.4
R23473 a_54607_15034.t0 a_54607_15034.t1 17.4
R23474 a_20814_13121.t0 a_20814_13121.t1 17.4
R23475 a_60464_18601.n0 a_60464_18601.t0 14.282
R23476 a_60464_18601.n0 a_60464_18601.t1 14.282
R23477 a_60464_18601.n1 a_60464_18601.t4 14.282
R23478 a_60464_18601.n1 a_60464_18601.t5 14.282
R23479 a_60464_18601.t2 a_60464_18601.n3 14.282
R23480 a_60464_18601.n3 a_60464_18601.t3 14.282
R23481 a_60464_18601.n2 a_60464_18601.n0 2.546
R23482 a_60464_18601.n2 a_60464_18601.n1 2.367
R23483 a_60464_18601.n3 a_60464_18601.n2 0.001
R23484 a_23732_7655.t0 a_23732_7655.t1 17.4
R23485 a_23466_n3481.t0 a_23466_n3481.t1 17.4
R23486 a_18153_4620.t0 a_18153_4620.t1 380.209
R23487 a_35249_9412.t0 a_35249_9412.t1 17.4
R23488 a_7956_13121.t0 a_7956_13121.t1 17.4
R23489 a_48490_6178.t0 a_48490_6178.t1 17.4
R23490 a_17446_10391.t0 a_17446_10391.t1 17.4
R23491 a_71846_5105.t0 a_71846_5105.t1 17.4
R23492 a_55116_11332.t0 a_55116_11332.t1 17.4
R23493 a_14282_n3485.t0 a_14282_n3485.t1 17.4
R23494 a_23670_411.t0 a_23670_411.t1 17.4
R23495 a_54894_20633.t0 a_54894_20633.t1 17.4
R23496 a_17446_13125.t0 a_17446_13125.t1 17.4
R23497 a_66005_n1962.t0 a_66005_n1962.t1 17.4
R23498 a_4182_20263.t0 a_4182_20263.t1 17.4
R23499 Y[1].n1 Y[1].n0 185.55
R23500 Y[1].n1 Y[1].t0 28.568
R23501 Y[1].n0 Y[1].t1 28.565
R23502 Y[1].n0 Y[1].t2 28.565
R23503 Y[1].n2 Y[1].t3 20.393
R23504 Y[1].n2 Y[1].n1 1.837
R23505 Y[1] Y[1].n2 1.12
R23506 a_23702_n3481.t0 a_23702_n3481.t1 17.4
R23507 a_39799_310.t0 a_39799_310.t1 380.209
R23508 a_65769_n1962.t0 a_65769_n1962.t1 380.209
R23509 a_53005_309.t0 a_53005_309.t1 380.209
R23510 a_23434_411.t0 a_23434_411.t1 17.4
R23511 a_23722_10387.t0 a_23722_10387.t1 17.4
R23512 a_41705_6090.t0 a_41705_6090.t1 380.209
R23513 a_63015_14838.t0 a_63015_14838.t1 17.4
R23514 a_48462_11311.t0 a_48462_11311.t1 17.4
R23515 a_52473_15034.t0 a_52473_15034.t1 380.209
R23516 a_57967_9233.t0 a_57967_9233.t1 17.4
R23517 a_61525_310.t0 a_61525_310.t1 380.209
R23518 a_40043_6090.t0 a_40043_6090.t1 17.4
R23519 a_48073_15029.t0 a_48073_15029.t1 17.4
R23520 a_51351_5911.t0 a_51351_5911.t1 17.4
R23521 a_48254_6178.t0 a_48254_6178.t1 380.209
R23522 a_7562_20263.t0 a_7562_20263.t1 17.4
R23523 a_5060_10391.t0 a_5060_10391.t1 17.4
R23524 a_9879_4622.t0 a_9879_4622.t1 380.209
R23525 a_31377_5900.t0 a_31377_5900.t1 379.845
R23526 a_20526_411.t0 a_20526_411.t1 17.4
R23527 a_46592_6178.t0 a_46592_6178.t1 17.4
R23528 a_1392_407.t0 a_1392_407.t1 17.4
R23529 a_67372_n1177.t0 a_67372_n1177.t1 17.4
R23530 a_24806_15774.t0 a_24806_15774.t1 17.4
R23531 a_31377_n70.t0 a_31377_n70.t1 17.4
R23532 a_5060_13125.t0 a_5060_13125.t1 17.4
R23533 a_53004_22038.t0 a_53004_22038.t1 17.4
R23534 a_31375_n2374.t0 a_31375_n2374.t1 379.845
R23535 a_11336_13121.t0 a_11336_13121.t1 17.4
R23536 a_10694_20259.t0 a_10694_20259.t1 17.4
R23537 a_1680_10391.t0 a_1680_10391.t1 17.4
R23538 a_23968_7655.t0 a_23968_7655.t1 17.4
R23539 a_18892_15774.t0 a_18892_15774.t1 17.4
R23540 a_71846_17491.t0 a_71846_17491.t1 17.4
R23541 a_46586_308.t0 a_46586_308.t1 17.4
R23542 a_20412_15776.t0 a_20412_15776.t1 17.4
R23543 a_44691_109.t0 a_44691_109.t1 17.4
R23544 a_46465_20439.t0 a_46465_20439.t1 17.4
R23545 a_52990_23688.t0 a_52990_23688.t1 17.4
R23546 a_7668_411.t0 a_7668_411.t1 17.4
R23547 a_61761_310.t0 a_61761_310.t1 17.4
R23548 a_8192_13121.t0 a_8192_13121.t1 17.4
R23549 a_59222_15037.t0 a_59222_15037.t1 17.4
R23550 a_4418_20263.t0 a_4418_20263.t1 17.4
R23551 a_16804_20263.t0 a_16804_20263.t1 17.4
R23552 a_66003_9972.t0 a_66003_9972.t1 17.4
R23553 a_14302_10391.t0 a_14302_10391.t1 17.4
R23554 a_52709_15034.t0 a_52709_15034.t1 17.4
R23555 a_14302_13125.t0 a_14302_13125.t1 17.4
R23556 a_23722_13121.t0 a_23722_13121.t1 17.4
R23557 a_17682_10391.t0 a_17682_10391.t1 17.4
R23558 a_17682_13125.t0 a_17682_13125.t1 17.4
R23559 a_7966_7655.t0 a_7966_7655.t1 17.4
C0 w_42676_18663# A[2] 0.01fF
C1 w_49220_17009# VDD 0.37fF
C2 w_46079_22618# w_46074_21014# 0.02fF
C3 w_49532_24144# A[2] 0.00fF
C4 w_46046_17952# A[3] 0.12fF
C5 w_46074_21014# A[1] 0.20fF
C6 w_39566_22621# VDD 0.37fF
C7 w_39566_22621# Cout 0.00fF
C8 A[1] opcode[0] 10.21fF
C9 VDD A[5] 13.35fF
C10 A[2] A[3] 94.86fF
C11 A[0] A[6] 0.31fF
C12 A[7] opcode[1] 18.01fF
C13 A[1] B[3] 0.11fF
C14 A[2] B[4] 0.09fF
C15 VDD B[1] 6.32fF
C16 A[6] B[7] 0.70fF
C17 A[0] B[2] 0.17fF
C18 w_39561_21017# w_40630_17952# 0.00fF
C19 w_59093_17960# w_60235_17956# 0.03fF
C20 opcode[0] B[6] 1.13fF
C21 A[3] B[5] 54.32fF
C22 VDD Y[0] 0.72fF
C23 B[7] B[2] 0.17fF
C24 B[6] B[3] 0.29fF
C25 B[5] B[4] 44.30fF
C26 A[4] opcode[2] 0.22fF
C27 opcode[1] B[0] 0.14fF
C28 w_55754_17014# A[5] 0.08fF
C29 w_39488_17956# opcode[0] 0.02fF
C30 w_53722_17953# VDD 0.50fF
C31 w_49532_24144# w_47542_22001# 0.01fF
C32 w_52580_17957# A[6] 0.00fF
C33 w_51779_16397# VDD 1.02fF
C34 w_41029_22004# w_39561_21017# 0.00fF
C35 w_59093_17960# A[5] 0.00fF
C36 w_45245_16392# A[6] 0.59fF
C37 w_42676_18663# A[3] 0.09fF
C38 w_59171_22617# VDD 0.37fF
C39 w_46074_21014# w_46046_17952# 0.00fF
C40 w_46074_21014# A[2] 0.01fF
C41 w_39566_22621# A[0] 0.07fF
C42 A[2] opcode[0] 3.00fF
C43 w_40630_17952# VDD 0.54fF
C44 A[0] A[5] 0.31fF
C45 A[1] A[6] 0.32fF
C46 VDD A[7] 11.58fF
C47 A[2] B[3] 0.17fF
C48 A[4] opcode[1] 0.86fF
C49 A[6] B[6] 27.90fF
C50 w_40630_17952# Cout 0.01fF
C51 A[5] B[7] 0.24fF
C52 A[0] B[1] 0.26fF
C53 A[1] B[2] 0.21fF
C54 VDD B[0] 10.21fF
C55 opcode[0] B[5] 1.26fF
C56 A[3] B[4] 2.09fF
C57 w_39552_24271# opcode[0] 0.00fF
C58 B[7] B[1] 0.22fF
C59 B[5] B[3] 0.37fF
C60 B[6] B[2] 0.07fF
C61 w_60634_22000# A[3] 0.60fF
C62 w_43019_24147# VDD 0.67fF
C63 opcode[2] opcode[3] 0.00fF
C64 w_42667_15409# VDD 0.33fF
C65 w_47542_22001# w_46074_21014# 0.00fF
C66 w_62281_18667# A[4] 0.07fF
C67 w_54924_24135# A[2] 0.01fF
C68 w_55768_18664# A[3] 0.08fF
C69 w_41029_22004# VDD 0.93fF
C70 w_52580_17957# w_53722_17953# 0.03fF
C71 w_61482_24139# A[3] 0.01fF
C72 w_42676_18663# opcode[0] 0.00fF
C73 w_47188_17948# VDD 0.50fF
C74 w_52599_24263# w_52613_22613# 0.01fF
C75 w_59157_24267# w_59171_22617# 0.01fF
C76 w_52580_17957# w_51779_16397# 0.01fF
C77 w_38687_16396# A[7] 0.59fF
C78 w_46074_21014# A[3] 0.00fF
C79 w_48390_24140# VDD 0.54fF
C80 A[0] A[7] 0.37fF
C81 A[1] A[5] 0.33fF
C82 A[2] A[6] 0.64fF
C83 A[3] opcode[0] 3.52fF
C84 VDD A[4] 13.33fF
C85 w_55759_15410# VDD 0.33fF
C86 A[5] B[6] 1.56fF
C87 A[6] B[5] 33.06fF
C88 opcode[0] B[4] 1.69fF
C89 A[1] B[1] 16.60fF
C90 VDD opcode[2] 9.23fF
C91 A[2] B[2] 16.18fF
C92 A[3] B[3] 74.47fF
C93 A[7] B[7] 18.59fF
C94 A[0] B[0] 26.81fF
C95 w_54076_21996# w_52608_21009# 0.00fF
C96 B[4] B[3] 48.52fF
C97 B[7] B[0] 9.49fF
C98 B[5] B[2] 0.08fF
C99 B[6] B[1] 0.07fF
C100 w_52599_24263# A[2] 0.06fF
C101 w_62267_17017# w_62272_15413# 0.02fF
C102 w_38687_16396# w_42667_15409# 0.00fF
C103 w_55754_17014# w_55759_15410# 0.02fF
C104 w_49225_15405# A[6] 0.14fF
C105 w_54076_21996# VDD 0.92fF
C106 w_58292_16400# A[5] 0.06fF
C107 w_41029_22004# A[0] 0.60fF
C108 w_49234_18659# VDD 0.36fF
C109 w_56066_24139# w_54076_21996# 0.01fF
C110 w_42676_18663# w_42662_17013# 0.01fF
C111 w_45245_16392# A[7] 0.05fF
C112 w_59166_21013# A[3] 0.20fF
C113 w_46065_24268# VDD 0.40fF
C114 w_60634_22000# w_59166_21013# 0.00fF
C115 w_46074_21014# opcode[0] 0.00fF
C116 w_49220_17009# w_49225_15405# 0.02fF
C117 VDD opcode[1] 26.95fF
C118 A[1] A[7] 0.70fF
C119 A[0] A[4] 0.46fF
C120 A[3] A[6] 1.51fF
C121 A[2] A[5] 0.37fF
C122 w_40630_17952# A[1] 0.01fF
C123 w_39561_21017# VDD 0.34fF
C124 w_39552_24271# w_39566_22621# 0.01fF
C125 A[5] B[5] 43.45fF
C126 A[3] B[2] 19.97fF
C127 opcode[0] B[3] 1.83fF
C128 A[7] B[6] 14.01fF
C129 w_39561_21017# Cout 0.00fF
C130 A[2] B[1] 14.99fF
C131 VDD opcode[3] 8.77fF
C132 A[1] B[0] 16.05fF
C133 A[4] B[7] 0.19fF
C134 A[6] B[4] 3.64fF
C135 B[6] B[0] 0.19fF
C136 B[4] B[2] 0.08fF
C137 B[5] B[1] 0.08fF
C138 w_39488_17956# w_40630_17952# 0.03fF
C139 w_43019_24147# A[1] 0.00fF
C140 opcode[3] Y[7] 0.08fF
C141 w_62281_18667# VDD 0.38fF
C142 w_41029_22004# A[1] 0.07fF
C143 w_62624_24143# VDD 0.67fF
C144 w_41877_24143# w_43019_24147# 0.03fF
C145 w_52608_21009# VDD 0.34fF
C146 w_46046_17952# A[7] 0.00fF
C147 w_48390_24140# A[1] 0.01fF
C148 opcode[0] A[6] 3.62fF
C149 A[2] A[7] 0.41fF
C150 A[1] A[4] 0.43fF
C151 A[0] opcode[1] 0.61fF
C152 A[3] A[5] 1.97fF
C153 VDD Cout 2.64fF
C154 w_39561_21017# A[0] 0.19fF
C155 w_40630_17952# A[2] 0.01fF
C156 w_55754_17014# VDD 0.37fF
C157 A[7] B[5] 0.43fF
C158 A[4] B[6] 1.40fF
C159 VDD Y[7] 0.73fF
C160 A[1] opcode[2] 0.02fF
C161 A[6] B[3] 4.50fF
C162 opcode[0] B[2] 0.93fF
C163 A[5] B[4] 16.86fF
C164 A[2] B[0] 0.35fF
C165 opcode[1] B[7] 0.38fF
C166 A[3] B[1] 0.19fF
C167 B[5] B[0] 0.18fF
C168 B[3] B[2] 44.80fF
C169 B[4] B[1] 0.07fF
C170 opcode[3] Y[6] 0.08fF
C171 w_53722_17953# A[3] 0.10fF
C172 w_56066_24139# VDD 0.67fF
C173 w_58292_16400# A[4] 0.59fF
C174 w_55768_18664# A[5] 0.07fF
C175 w_41029_22004# A[2] 0.00fF
C176 w_59093_17960# VDD 0.66fF
C177 w_46065_24268# w_46079_22618# 0.01fF
C178 w_46046_17952# w_47188_17948# 0.03fF
C179 w_42676_18663# A[7] 0.07fF
C180 w_59171_22617# A[3] 0.08fF
C181 w_46065_24268# A[1] 0.06fF
C182 w_47188_17948# A[2] 0.00fF
C183 w_38687_16396# VDD 1.02fF
C184 w_38687_16396# Cout 0.03fF
C185 w_39566_22621# opcode[0] 0.07fF
C186 VDD A[0] 17.36fF
C187 w_40630_17952# A[3] 0.11fF
C188 A[2] A[4] 1.20fF
C189 A[1] opcode[1] 0.98fF
C190 A[3] A[7] 0.50fF
C191 VDD B[7] 5.36fF
C192 A[0] Cout 0.22fF
C193 w_39561_21017# A[1] 0.03fF
C194 opcode[0] A[5] 3.81fF
C195 w_59157_24267# VDD 0.40fF
C196 A[7] B[4] 0.41fF
C197 A[6] B[2] 0.38fF
C198 A[3] B[0] 0.44fF
C199 A[4] B[5] 1.94fF
C200 VDD Y[6] 0.73fF
C201 opcode[1] B[6] 0.23fF
C202 A[5] B[3] 5.52fF
C203 opcode[0] B[1] 0.85fF
C204 A[2] opcode[2] 0.06fF
C205 B[3] B[1] 0.08fF
C206 B[4] B[0] 0.17fF
C207 w_52608_21009# w_52580_17957# 0.00fF
C208 w_59166_21013# w_60235_17956# 0.00fF
C209 w_39561_21017# w_39488_17956# 0.00fF
C210 opcode[3] Y[5] 0.08fF
C211 w_54076_21996# A[2] 0.60fF
C212 w_52580_17957# VDD 0.63fF
C213 w_49234_18659# A[2] 0.00fF
C214 w_45245_16392# VDD 1.02fF
C215 w_49220_17009# A[6] 0.08fF
C216 w_47188_17948# A[3] 0.10fF
C217 w_46079_22618# VDD 0.37fF
C218 w_48390_24140# w_49532_24144# 0.03fF
C219 VDD A[1] 11.17fF
C220 w_62272_15413# A[4] 0.14fF
C221 w_40630_17952# opcode[0] 0.01fF
C222 A[2] opcode[1] 0.32fF
C223 opcode[0] A[7] 0.81fF
C224 A[6] A[5] 115.99fF
C225 VDD B[6] 10.93fF
C226 A[3] A[4] 90.33fF
C227 A[1] Cout 0.08fF
C228 A[0] B[7] 0.20fF
C229 w_39561_21017# A[2] 0.01fF
C230 A[7] B[3] 0.40fF
C231 opcode[0] B[0] 0.72fF
C232 A[5] B[2] 0.25fF
C233 A[6] B[1] 0.59fF
C234 A[3] opcode[2] 0.08fF
C235 A[4] B[4] 47.59fF
C236 opcode[1] B[5] 0.32fF
C237 VDD Y[5] 0.73fF
C238 w_39488_17956# VDD 0.68fF
C239 B[3] B[0] 0.17fF
C240 B[2] B[1] 38.17fF
C241 w_39488_17956# Cout 0.19fF
C242 w_43019_24147# opcode[0] 0.00fF
C243 opcode[3] Y[4] 0.08fF
C244 w_54076_21996# A[3] 0.05fF
C245 w_41877_24143# VDD 0.54fF
C246 w_58292_16400# VDD 1.02fF
C247 w_52613_22613# w_52608_21009# 0.02fF
C248 w_59171_22617# w_59166_21013# 0.02fF
C249 w_41029_22004# opcode[0] 0.39fF
C250 w_51779_16397# A[6] 0.06fF
C251 w_49234_18659# A[3] 0.08fF
C252 w_52613_22613# VDD 0.37fF
C253 w_52608_21009# A[2] 0.20fF
C254 w_46046_17952# VDD 0.64fF
C255 VDD A[2] 9.88fF
C256 A[0] A[1] 58.38fF
C257 w_39488_17956# w_38687_16396# 0.01fF
C258 w_59093_17960# w_58292_16400# 0.01fF
C259 w_42662_17013# A[7] 0.08fF
C260 VDD B[5] 13.79fF
C261 w_39561_21017# A[3] 0.00fF
C262 opcode[0] A[4] 3.16fF
C263 A[0] B[6] 0.12fF
C264 A[3] opcode[1] 0.51fF
C265 A[6] A[7] 84.34fF
C266 A[2] Cout 0.10fF
C267 A[1] B[7] 0.17fF
C268 w_39552_24271# VDD 0.40fF
C269 A[5] B[1] 0.12fF
C270 A[4] B[3] 16.00fF
C271 VDD Y[4] 0.73fF
C272 B[7] B[6] 46.19fF
C273 opcode[1] B[4] 0.22fF
C274 A[6] B[0] 0.52fF
C275 A[7] B[2] 0.41fF
C276 w_39488_17956# A[0] 0.03fF
C277 w_39552_24271# Cout 0.00fF
C278 B[2] B[0] 0.22fF
C279 w_49225_15405# VDD 0.33fF
C280 opcode[3] Y[3] 0.08fF
C281 w_62267_17017# A[4] 0.08fF
C282 w_53722_17953# A[5] 0.01fF
C283 w_41877_24143# A[0] 0.01fF
C284 w_42662_17013# w_42667_15409# 0.02fF
C285 w_47542_22001# VDD 0.92fF
C286 w_51779_16397# A[5] 0.59fF
C287 w_42676_18663# VDD 0.36fF
C288 w_62624_24143# w_60634_22000# 0.02fF
C289 w_47188_17948# A[6] 0.01fF
C290 w_52608_21009# A[3] 0.00fF
C291 w_46079_22618# A[1] 0.08fF
C292 w_49532_24144# VDD 0.67fF
C293 w_62272_15413# VDD 0.33fF
C294 A[0] A[2] 1.19fF
C295 VDD A[3] 19.28fF
C296 VDD B[4] 10.31fF
C297 w_39561_21017# opcode[0] 0.20fF
C298 A[3] Cout 0.13fF
C299 opcode[0] opcode[1] 38.92fF
C300 A[0] B[5] 0.13fF
C301 A[1] B[6] 0.12fF
C302 A[5] A[7] 1.40fF
C303 A[6] A[4] 5.20fF
C304 A[2] B[7] 0.16fF
C305 w_39552_24271# A[0] 0.06fF
C306 opcode[1] B[3] 0.21fF
C307 B[7] B[5] 0.31fF
C308 A[6] opcode[2] 0.46fF
C309 A[5] B[0] 0.34fF
C310 A[7] B[1] 0.57fF
C311 VDD Y[3] 0.73fF
C312 A[4] B[2] 0.12fF
C313 w_39488_17956# A[1] 0.01fF
C314 w_60634_22000# VDD 0.94fF
C315 w_61482_24139# w_62624_24143# 0.03fF
C316 B[1] B[0] 38.11fF
C317 opcode[3] Y[2] 0.08fF
C318 w_56066_24139# A[3] 0.00fF
C319 w_52580_17957# A[2] 0.02fF
C320 w_55768_18664# VDD 0.36fF
C321 w_60235_17956# A[4] 0.01fF
C322 w_62281_18667# w_62267_17017# 0.01fF
C323 w_46046_17952# w_45245_16392# 0.01fF
C324 w_55768_18664# w_55754_17014# 0.01fF
C325 w_49234_18659# A[6] 0.07fF
C326 w_59093_17960# A[3] 0.02fF
C327 w_61482_24139# VDD 0.54fF
C328 w_45245_16392# w_49225_15405# 0.00fF
C329 w_46046_17952# A[1] 0.02fF
C330 w_46074_21014# VDD 0.34fF
C331 A[1] A[2] 78.96fF
C332 VDD opcode[0] 31.99fF
C333 A[0] A[3] 0.33fF
C334 A[0] B[4] 0.11fF
C335 A[3] B[7] 0.21fF
C336 A[1] B[5] 0.12fF
C337 A[2] B[6] 0.12fF
C338 A[5] A[4] 128.19fF
C339 w_40630_17952# A[7] 0.01fF
C340 A[6] opcode[1] 1.64fF
C341 VDD B[3] 7.87fF
C342 opcode[0] Cout 0.25fF
C343 w_59157_24267# A[3] 0.06fF
C344 w_55759_15410# A[5] 0.14fF
C345 B[7] B[4] 0.24fF
C346 A[5] opcode[2] 0.33fF
C347 A[4] B[1] 0.13fF
C348 opcode[1] B[2] 0.23fF
C349 VDD Y[2] 0.73fF
C350 A[7] B[0] 0.76fF
C351 B[6] B[5] 42.32fF
C352 w_39488_17956# A[2] 0.01fF
C353 w_62267_17017# VDD 0.37fF
C354 opcode[3] Y[1] 0.08fF
C355 w_42667_15409# A[7] 0.14fF
C356 w_49234_18659# w_49220_17009# 0.01fF
C357 w_52580_17957# A[3] 0.12fF
C358 w_47542_22001# A[1] 0.60fF
C359 w_54924_24135# VDD 0.54fF
C360 w_52613_22613# A[2] 0.08fF
C361 w_51779_16397# w_55759_15410# 0.00fF
C362 w_42676_18663# A[1] 0.01fF
C363 w_59166_21013# VDD 0.34fF
C364 w_54924_24135# w_56066_24139# 0.03fF
C365 w_43019_24147# w_41029_22004# 0.01fF
C366 w_46046_17952# A[2] 0.01fF
C367 w_42662_17013# VDD 0.37fF
C368 w_39566_22621# w_39561_21017# 0.02fF
C369 A[0] opcode[0] 6.54fF
C370 VDD A[6] 14.04fF
C371 A[1] A[3] 2.02fF
C372 A[3] B[6] 25.95fF
C373 A[7] A[4] 0.54fF
C374 opcode[0] B[7] 13.72fF
C375 A[0] B[3] 0.14fF
C376 A[1] B[4] 0.11fF
C377 VDD B[2] 5.69fF
C378 A[2] B[5] 0.09fF
C379 A[5] opcode[1] 1.07fF
C380 VDD Y[1] 0.73fF
C381 opcode[1] B[1] 0.21fF
C382 A[7] opcode[2] 0.51fF
C383 B[6] B[4] 27.85fF
C384 A[4] B[0] 0.37fF
C385 B[7] B[3] 0.37fF
C386 w_39488_17956# A[3] 0.12fF
C387 w_52599_24263# VDD 0.40fF
C388 opcode[3] Y[0] 0.01fF
C389 w_59166_21013# w_59093_17960# 0.00fF
C390 w_47542_22001# A[2] 0.06fF
C391 w_58292_16400# w_62272_15413# 0.00fF
C392 w_60235_17956# VDD 0.52fF
.ends

