** sch_path: /home/salih/Desktop/design/xschem/ALU.sch
.subckt ALU A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0]
+ opcode[3] opcode[2] opcode[1] opcode[0] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] VDD VSS flags[0] flags[1]
+ flags[2] flags[3]
*.PININFO A[7:0]:I B[7:0]:I opcode[3:0]:I Y[0:7]:O VDD:B VSS:B flags[0:3]:O
x1 net1 A[7] VDD VSS B[7] xor2
x2 VDD net2 net3 VSS inverter
x3 net3 A[7] VDD VSS Y[7] xor2
x4 flags[2] B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] VSS VDD
+ Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] opcode[0] opcode[1] opcode[2] opcode[3] control_unit
x5 VSS net1 net2 VDD flags[1] and2
x6 Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] VSS VDD flags[3] nor8
.ends

* expanding   symbol:  xor2.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/xor2.sym
** sch_path: /home/salih/Desktop/design/xschem/xor2.sch
.subckt xor2  Y A VDD VSS B
*.PININFO Y:O A:I VDD:B VSS:B B:I
XM7 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Y inv_B net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Y inv_A net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Y A net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y inv_A net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 inv_B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 inv_B B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 inv_B B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 inv_A A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 inv_A A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/salih/Desktop/design/xschem/inverter.sym
** sch_path: /home/salih/Desktop/design/xschem/inverter.sch
.subckt inverter  VDD OUT IN VSS
*.PININFO IN:I VDD:B OUT:O VSS:B
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  control_unit.sym # of pins=7
** sym_path: /home/salih/Desktop/design/xschem/control_unit.sym
** sch_path: /home/salih/Desktop/design/xschem/control_unit.sch
.subckt control_unit  Cout B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] A[0] A[1] A[2] A[3] A[4] A[5]
+ A[6] A[7] VSS VDD Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] opcode[3] opcode[2] opcode[1] opcode[0]
*.PININFO B[0:7]:I A[0:7]:I Y[0:7]:O VDD:B VSS:B opcode[3:0]:I Cout:O
x1 B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] l_u_out[0] l_u_out[1] l_u_out[2] l_u_out[3] l_u_out[4]
+ l_u_out[5] l_u_out[6] l_u_out[7] VDD VSS opcode[0] opcode[1] opcode[2] opcode[3] A[0] A[1] A[2] A[3] A[4] A[5]
+ A[6] A[7] logic_unit
x2 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] s_u_out[0] s_u_out[1] s_u_out[2] s_u_out[3] s_u_out[4]
+ s_u_out[5] s_u_out[6] s_u_out[7] opcode[0] shifter_unit
x3 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] opcode[0]
+ opcode[1] opcode[2] opcode[3] VSS VDD a_u_out[0] a_u_out[1] a_u_out[2] a_u_out[3] a_u_out[4] a_u_out[5]
+ a_u_out[6] a_u_out[7] Cout arithmetic_unit
x4 VSS VDD opcode[2] a_u_out[7] l_u_out[7] net8 2x1_mux
x5 VSS VDD opcode[2] a_u_out[6] l_u_out[6] net7 2x1_mux
x6 VSS VDD opcode[2] a_u_out[5] l_u_out[5] net6 2x1_mux
x7 VSS VDD opcode[2] a_u_out[4] l_u_out[4] net5 2x1_mux
x8 VSS VDD opcode[2] a_u_out[3] l_u_out[3] net4 2x1_mux
x9 VSS VDD opcode[2] a_u_out[2] l_u_out[2] net3 2x1_mux
x10 VSS VDD opcode[2] a_u_out[1] l_u_out[1] net2 2x1_mux
x11 VSS VDD opcode[2] a_u_out[0] l_u_out[0] net1 2x1_mux
x12 VSS VDD opcode[3] net8 s_u_out[7] Y[7] 2x1_mux
x13 VSS VDD opcode[3] net7 s_u_out[6] Y[6] 2x1_mux
x14 VSS VDD opcode[3] net6 s_u_out[5] Y[5] 2x1_mux
x15 VSS VDD opcode[3] net5 s_u_out[4] Y[4] 2x1_mux
x16 VSS VDD opcode[3] net4 s_u_out[3] Y[3] 2x1_mux
x17 VSS VDD opcode[3] net3 s_u_out[2] Y[2] 2x1_mux
x18 VSS VDD opcode[3] net2 s_u_out[1] Y[1] 2x1_mux
x19 VSS VDD opcode[3] net1 s_u_out[0] Y[0] 2x1_mux
.ends


* expanding   symbol:  and2.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/and2.sym
** sch_path: /home/salih/Desktop/design/xschem/and2.sch
.subckt and2  VSS A B VDD OUT
*.PININFO VSS:B A:I B:I VDD:B OUT:O
XM2 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  nor8.sym # of pins=4
** sym_path: /home/salih/Desktop/design/xschem/nor8.sym
** sch_path: /home/salih/Desktop/design/xschem/nor8.sch
.subckt nor8  A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] VSS VDD Y
*.PININFO A[7:0]:I VDD:B VSS:B Y:O
x1 A[0] A[1] VSS VDD net1 or2
x2 A[2] A[3] VSS VDD net2 or2
x3 A[4] A[5] VSS VDD net3 or2
x4 A[6] A[7] VSS VDD net4 or2
x5 net1 net2 VSS VDD net5 or2
x6 net3 net4 VSS VDD net6 or2
x7 net5 net6 VSS VDD net7 or2
x8 VDD Y net7 VSS inverter
.ends


* expanding   symbol:  logic_unit.sym # of pins=6
** sym_path: /home/salih/Desktop/design/xschem/logic_unit.sym
** sch_path: /home/salih/Desktop/design/xschem/logic_unit.sch
.subckt logic_unit  B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
+ VDD VSS opcode[0] opcode[1] opcode[2] opcode[3] A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
*.PININFO B[0:7]:I Y[0:7]:O VDD:B VSS:B opcode[0:3]:I A[0:7]:I
x1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y_or[0] Y_or[1] Y_or[2] Y_or[3] Y_or[4] Y_or[5] Y_or[6]
+ Y_or[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] logic_or
x2 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y_and[0] Y_and[1] Y_and[2] Y_and[3] Y_and[4] Y_and[5]
+ Y_and[6] Y_and[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] logic_and
x3 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y_xor[0] Y_xor[1] Y_xor[2] Y_xor[3] Y_xor[4] Y_xor[5]
+ Y_xor[6] Y_xor[7] VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7] logic_xor
x4 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y_inv[0] Y_inv[1] Y_inv[2] Y_inv[3] Y_inv[4] Y_inv[5]
+ Y_inv[6] Y_inv[7] VSS VDD logic_inverter
x5 VSS VDD opcode[0] Y_and[0] Y_or[0] L1[0] 2x1_mux
x6 VSS VDD opcode[0] Y_and[1] Y_or[1] L1[1] 2x1_mux
x7 VSS VDD opcode[0] Y_and[2] Y_or[2] L1[2] 2x1_mux
x8 VSS VDD opcode[0] Y_and[3] Y_or[3] L1[3] 2x1_mux
x9 VSS VDD opcode[0] Y_and[4] Y_or[4] L1[4] 2x1_mux
x10 VSS VDD opcode[0] Y_and[5] Y_or[5] L1[5] 2x1_mux
x11 VSS VDD opcode[0] Y_and[6] Y_or[6] L1[6] 2x1_mux
x12 VSS VDD opcode[0] Y_and[7] Y_or[7] L1[7] 2x1_mux
x13 VSS VDD opcode[0] Y_xor[0] Y_inv[0] L2[0] 2x1_mux
x14 VSS VDD opcode[0] Y_xor[1] Y_inv[1] L2[1] 2x1_mux
x15 VSS VDD opcode[0] Y_xor[2] Y_inv[2] L2[2] 2x1_mux
x16 VSS VDD opcode[0] Y_xor[3] Y_inv[3] L2[3] 2x1_mux
x17 VSS VDD opcode[0] Y_xor[4] Y_inv[4] L2[4] 2x1_mux
x18 VSS VDD opcode[0] Y_xor[5] Y_inv[5] L2[5] 2x1_mux
x19 VSS VDD opcode[0] Y_xor[6] Y_inv[6] L2[6] 2x1_mux
x20 VSS VDD opcode[0] Y_xor[7] Y_inv[7] L2[7] 2x1_mux
x21 VSS VDD opcode[1] L1[0] L2[0] Y[0] 2x1_mux
x22 VSS VDD opcode[1] L1[1] L2[1] Y[1] 2x1_mux
x23 VSS VDD opcode[1] L1[2] L2[2] Y[2] 2x1_mux
x24 VSS VDD opcode[1] L1[3] L2[3] Y[3] 2x1_mux
x25 VSS VDD opcode[1] L1[4] L2[4] Y[4] 2x1_mux
x26 VSS VDD opcode[1] L1[5] L2[5] Y[5] 2x1_mux
x27 VSS VDD opcode[1] L1[6] L2[6] Y[6] 2x1_mux
x28 VSS VDD opcode[1] L1[7] L2[7] Y[7] 2x1_mux
.ends


* expanding   symbol:  shifter_unit.sym # of pins=3
** sym_path: /home/salih/Desktop/design/xschem/shifter_unit.sym
** sch_path: /home/salih/Desktop/design/xschem/shifter_unit.sch
.subckt shifter_unit  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6]
+ Y[7] dir
*.PININFO A[0:7]:I Y[0:7]:O dir:I
x9 VSS VDD dir A[0] A[0] Y[0] 2x1_mux
x1 VSS VDD dir A[1] A[1] Y[1] 2x1_mux
x2 VSS VDD dir A[2] A[2] Y[2] 2x1_mux
x3 VSS VDD dir A[3] A[3] Y[3] 2x1_mux
x4 VSS VDD dir A[4] A[4] Y[4] 2x1_mux
x5 VSS VDD dir A[5] A[5] Y[5] 2x1_mux
x6 VSS VDD dir A[6] A[6] Y[6] 2x1_mux
x7 VSS VDD dir A[7] A[7] Y[7] 2x1_mux
.ends


* expanding   symbol:  arithmetic_unit.sym # of pins=7
** sym_path: /home/salih/Desktop/design/xschem/arithmetic_unit.sym
** sch_path: /home/salih/Desktop/design/xschem/arithmetic_unit.sch
.subckt arithmetic_unit  A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[7] B[6] B[5] B[4] B[3] B[2] B[1]
+ B[0] opcode[3] opcode[2] opcode[1] opcode[0] VSS VDD Y[7] Y[6] Y[5] Y[4] Y[3] Y[2] Y[1] Y[0] Cout
*.PININFO A[7:0]:I B[7:0]:I opcode[3:0]:I Y[7:0]:O Cout:O VSS:B VDD:B
x1 sub[0] opcode[0] VDD VSS B[0] xor2
x2 sub[1] opcode[0] VDD VSS B[1] xor2
x3 sub[2] opcode[0] VDD VSS B[2] xor2
x4 sub[3] opcode[0] VDD VSS B[3] xor2
x5 sub[4] opcode[0] VDD VSS B[4] xor2
x6 sub[5] opcode[0] VDD VSS B[5] xor2
x7 sub[6] opcode[0] VDD VSS B[6] xor2
x8 sub[7] opcode[0] VDD VSS B[7] xor2
x9 VSS VDD opcode[1] adder[0] multi[0] Y[0] 2x1_mux
x10 VSS VDD opcode[1] adder[1] multi[1] Y[1] 2x1_mux
x11 VSS VDD opcode[1] adder[2] multi[2] Y[2] 2x1_mux
x12 VSS VDD opcode[1] adder[3] multi[3] Y[3] 2x1_mux
x13 VSS VDD opcode[1] adder[4] multi[4] Y[4] 2x1_mux
x14 VSS VDD opcode[1] adder[5] multi[5] Y[5] 2x1_mux
x15 VSS VDD opcode[1] adder[6] multi[6] Y[6] 2x1_mux
x16 VSS VDD opcode[1] adder[7] multi[7] Y[7] 2x1_mux
x17 VSS VDD A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] sub[7] sub[6] sub[5] sub[4] sub[3] sub[2] sub[1]
+ sub[0] opcode[0] adder[7] adder[6] adder[5] adder[4] adder[3] adder[2] adder[1] adder[0] Cout
+ carry_ripple_adder
x18 VSS VDD A[6] A[5] A[4] A[3] B[6] B[5] B[4] B[3] multi[7] multi[6] multi[5] multi[4] multi[3]
+ multi[2] multi[1] multi[0] array_multiplier
.ends


* expanding   symbol:  2x1_mux.sym # of pins=6
** sym_path: /home/salih/Desktop/design/xschem/2x1_mux.sym
** sch_path: /home/salih/Desktop/design/xschem/2x1_mux.sch
.subckt 2x1_mux  VSS VDD S D0 D1 OUT
*.PININFO VSS:B VDD:B S:I D0:I D1:I OUT:O
XM2 net1 S_BAR net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 D1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 D0 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 S_BAR net4 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 D1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net4 S VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 S_BAR S VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 S_BAR S VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 S net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 D0 net4 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  or2.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/or2.sym
** sch_path: /home/salih/Desktop/design/xschem/or2.sch
.subckt or2  A B VSS VDD OUT
*.PININFO A:I B:I VSS:B VDD:B OUT:O
XM3 net1 A net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=6.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  logic_or.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/logic_or.sym
** sch_path: /home/salih/Desktop/design/xschem/logic_or.sch
.subckt logic_or  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
+ VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
*.PININFO A[0:7]:I Y[0:7]:O VSS:B VDD:B B[0:7]:I
x1 A[0] B[0] VSS VDD Y[0] or2
x2 A[1] B[1] VSS VDD Y[1] or2
x3 A[2] B[2] VSS VDD Y[2] or2
x4 A[3] B[3] VSS VDD Y[3] or2
x5 A[4] B[4] VSS VDD Y[4] or2
x6 A[5] B[5] VSS VDD Y[5] or2
x7 A[6] B[6] VSS VDD Y[6] or2
x8 A[7] B[7] VSS VDD Y[7] or2
.ends


* expanding   symbol:  logic_and.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/logic_and.sym
** sch_path: /home/salih/Desktop/design/xschem/logic_and.sch
.subckt logic_and  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
+ VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
*.PININFO A[0:7]:I Y[0:7]:O VSS:B VDD:B B[0:7]:I
x1 VSS A[0] B[0] VDD Y[0] and2
x2 VSS A[1] B[1] VDD Y[1] and2
x3 VSS A[2] B[2] VDD Y[2] and2
x4 VSS A[3] B[3] VDD Y[3] and2
x5 VSS A[4] B[4] VDD Y[4] and2
x6 VSS A[5] B[5] VDD Y[5] and2
x7 VSS A[6] B[6] VDD Y[6] and2
x8 VSS A[7] B[7] VDD Y[7] and2
.ends


* expanding   symbol:  logic_xor.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/logic_xor.sym
** sch_path: /home/salih/Desktop/design/xschem/logic_xor.sch
.subckt logic_xor  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
+ VSS VDD B[0] B[1] B[2] B[3] B[4] B[5] B[6] B[7]
*.PININFO A[0:7]:I Y[0:7]:O VSS:B VDD:B B[0:7]:I
x1 Y[0] A[0] VDD VSS B[0] xor2
x2 Y[1] A[1] VDD VSS B[1] xor2
x3 Y[2] A[2] VDD VSS B[2] xor2
x4 Y[3] A[3] VDD VSS B[3] xor2
x5 Y[4] A[4] VDD VSS B[4] xor2
x6 Y[5] A[5] VDD VSS B[5] xor2
x7 Y[6] A[6] VDD VSS B[6] xor2
x8 Y[7] A[7] VDD VSS B[7] xor2
.ends


* expanding   symbol:  logic_inverter.sym # of pins=4
** sym_path: /home/salih/Desktop/design/xschem/logic_inverter.sym
** sch_path: /home/salih/Desktop/design/xschem/logic_inverter.sch
.subckt logic_inverter  A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6]
+ Y[7] VSS VDD
*.PININFO A[0:7]:I Y[0:7]:O VSS:B VDD:B
x1 VDD Y[0] A[0] VSS inverter
x2 VDD Y[1] A[1] VSS inverter
x3 VDD Y[2] A[2] VSS inverter
x4 VDD Y[3] A[3] VSS inverter
x5 VDD Y[4] A[4] VSS inverter
x6 VDD Y[5] A[5] VSS inverter
x7 VDD Y[6] A[6] VSS inverter
x8 VDD Y[7] A[7] VSS inverter
.ends


* expanding   symbol:  carry_ripple_adder.sym # of pins=7
** sym_path: /home/salih/Desktop/design/xschem/carry_ripple_adder.sym
** sch_path: /home/salih/Desktop/design/xschem/carry_ripple_adder.sch
.subckt carry_ripple_adder  VSS VDD A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4]
+ B[5] B[6] B[7] carry_in Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] carry_out
*.PININFO A[0:7]:I B[0:7]:I carry_in:I VDD:B VSS:B Y[0:7]:O carry_out:O
x1 VDD VSS A[0] B[0] net1 carry_in Y[0] fulladder
x2 VDD VSS A[1] B[1] net2 net1 Y[1] fulladder
x3 VDD VSS A[2] B[2] net3 net2 Y[2] fulladder
x4 VDD VSS A[3] B[3] net4 net3 Y[3] fulladder
x5 VDD VSS A[4] B[4] net5 net4 Y[4] fulladder
x6 VDD VSS A[5] B[5] net6 net5 Y[5] fulladder
x7 VDD VSS A[6] B[6] net7 net6 Y[6] fulladder
x8 VDD VSS A[7] B[7] carry_out net7 Y[7] fulladder
.ends


* expanding   symbol:  array_multiplier.sym # of pins=5
** sym_path: /home/salih/Desktop/design/xschem/array_multiplier.sym
** sch_path: /home/salih/Desktop/design/xschem/array_multiplier.sch
.subckt array_multiplier  VSS VDD A[0] A[1] A[2] A[3] B[0] B[1] B[2] B[3] Y[0] Y[1] Y[2] Y[3] Y[4]
+ Y[5] Y[6] Y[7]
*.PININFO A[0:3]:I B[0:3]:I VDD:B VSS:B Y[0:7]:O
x1 VSS A[1] B[1] VDD net1 and2
x2 VSS A[2] B[0] VDD net2 and2
x3 VSS A[2] B[1] VDD net3 and2
x4 VSS A[3] B[0] VDD net4 and2
x5 VDD VSS net1 net2 net5 net30 net24 fulladder
x6 VDD VSS net3 net4 net10 net5 net7 fulladder
x7 VSS A[1] B[2] VDD net6 and2
x8 VDD VSS net7 net6 net8 net31 net26 fulladder
x9 VSS A[3] B[1] VDD net9 and2
x10 VDD VSS net10 net9 net13 net8 net12 fulladder
x11 VSS A[2] B[2] VDD net11 and2
x12 VDD VSS net12 net11 net15 net32 net20 fulladder
x13 VSS A[3] B[2] VDD net14 and2
x14 VSS A[2] B[3] VDD net17 and2
x15 VSS A[1] B[3] VDD net19 and2
x17 VSS A[0] B[1] VDD net21 and2
x18 VSS A[1] B[0] VDD net22 and2
x19 VSS A[0] B[2] VDD net23 and2
x20 VSS A[0] B[3] VDD net25 and2
x21 VSS A[3] B[3] VDD net28 and2
x22 VDD VSS net16 net17 net29 net18 Y[5] fulladder
x23 VDD VSS net20 Y[4] net19 net18 half_adder
x16 VDD VSS net13 net14 net27 net15 net16 fulladder
x24 VDD VSS net24 Y[2] net23 net31 half_adder
x25 VDD VSS net21 Y[1] net22 net30 half_adder
x26 VSS A[0] B[0] VDD Y[0] and2
x27 VDD VSS net26 Y[3] net25 net32 half_adder
x28 VDD VSS net27 net28 Y[6] net29 Y[7] fulladder
.ends


* expanding   symbol:  fulladder.sym # of pins=7
** sym_path: /home/salih/Desktop/design/xschem/fulladder.sym
** sch_path: /home/salih/Desktop/design/xschem/fulladder.sch
.subckt fulladder  VDD VSS A B carry_out carry_in Y
*.PININFO A:I B:I carry_in:I Y:O carry_out:O VDD:B VSS:B
x1 VSS A B VDD net1 and2
x2 VSS B carry_in VDD net2 and2
x3 VSS A carry_in VDD net3 and2
x4 VDD net1 net3 net2 carry_out VSS or3
x5 VDD A Y B carry_in VSS xor3
.ends


* expanding   symbol:  half_adder.sym # of pins=6
** sym_path: /home/salih/Desktop/design/xschem/half_adder.sym
** sch_path: /home/salih/Desktop/design/xschem/half_adder.sch
.subckt half_adder  VDD VSS A Y B carry_out
*.PININFO A:I B:I Y:O carry_out:O VDD:B VSS:B
x1 Y A VDD VSS B xor2
x2 VSS A B VDD carry_out and2
.ends


* expanding   symbol:  or3.sym # of pins=6
** sym_path: /home/salih/Desktop/design/xschem/or3.sym
** sch_path: /home/salih/Desktop/design/xschem/or3.sch
.subckt or3  VDD A B C OUT VSS
*.PININFO A:I B:I VSS:B VDD:B OUT:O C:I
XM4 net1 A net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 C VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 B net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 C VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xor3.sym # of pins=6
** sym_path: /home/salih/Desktop/design/xschem/xor3.sym
** sch_path: /home/salih/Desktop/design/xschem/xor3.sch
.subckt xor3  VDD A OUT B C VSS
*.PININFO C:I VSS:B A:I B:I OUT:O VDD:B
x1 net1 A VDD VSS B xor2
x2 OUT net1 VDD VSS C xor2
.ends

.end
