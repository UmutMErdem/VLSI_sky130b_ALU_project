* NGSPICE file created from or2_pex.ext - technology: sky130B

.subckt or2 A B VSS VDD OUT
X0 a_612_787.t2 A.t0 a_494_787.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1 VSS.t2 B.t0 a_494_787.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 a_494_787.t1 A.t1 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 VDD.t4 B.t1 a_612_787.t3 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 a_612_787.t1 A.t2 a_494_787.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X5 a_612_787.t4 B.t2 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X6 VDD.t14 B.t3 a_612_787.t5 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 OUT.t2 a_494_787.t5 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8 a_494_787.t0 A.t3 a_612_787.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 VDD.t8 a_494_787.t6 OUT.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10 VDD.t6 a_494_787.t7 OUT.t0 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X11 OUT.t3 a_494_787.t8 VSS.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 A.t0 A.t1 574.43
R1 A.n0 A.t2 285.109
R2 A.n0 A.t3 160.666
R3 A.n1 A.t0 160.666
R4 A A.n1 159.549
R5 A.n1 A.n0 114.829
R6 a_494_787.t8 a_494_787.n2 404.877
R7 a_494_787.n1 a_494_787.t7 210.902
R8 a_494_787.n3 a_494_787.t8 136.943
R9 a_494_787.n2 a_494_787.n1 107.801
R10 a_494_787.n1 a_494_787.t5 80.333
R11 a_494_787.n2 a_494_787.t6 80.333
R12 a_494_787.n0 a_494_787.t4 17.4
R13 a_494_787.n0 a_494_787.t1 17.4
R14 a_494_787.n4 a_494_787.t3 15.032
R15 a_494_787.n5 a_494_787.t2 14.282
R16 a_494_787.t0 a_494_787.n5 14.282
R17 a_494_787.n5 a_494_787.n4 1.65
R18 a_494_787.n3 a_494_787.n0 0.672
R19 a_494_787.n4 a_494_787.n3 0.665
R20 a_612_787.n1 a_612_787.t5 14.282
R21 a_612_787.n1 a_612_787.t1 14.282
R22 a_612_787.n0 a_612_787.t0 14.282
R23 a_612_787.n0 a_612_787.t2 14.282
R24 a_612_787.t3 a_612_787.n3 14.282
R25 a_612_787.n3 a_612_787.t4 14.282
R26 a_612_787.n2 a_612_787.n0 2.546
R27 a_612_787.n3 a_612_787.n2 2.367
R28 a_612_787.n2 a_612_787.n1 0.001
R29 VDD.n1 VDD.n0 602.445
R30 VDD.t9 VDD.t5 406.159
R31 VDD.n0 VDD.t7 404.97
R32 VDD.t13 VDD.t1 143.902
R33 VDD.t1 VDD.t0 143.902
R34 VDD.t0 VDD.t2 143.902
R35 VDD.n5 VDD.t13 137.804
R36 VDD.n6 VDD.t11 60.976
R37 VDD.n2 VDD.n1 29.268
R38 VDD.n9 VDD.t6 28.57
R39 VDD.n8 VDD.t10 28.565
R40 VDD.n8 VDD.t8 28.565
R41 VDD.n10 VDD.t4 14.284
R42 VDD.n11 VDD.t12 14.282
R43 VDD.n11 VDD.t14 14.282
R44 VDD.n3 VDD.t3 13.414
R45 VDD.t11 VDD.n5 6.097
R46 VDD.n4 VDD.n3 5.506
R47 VDD.n10 VDD.n9 2.195
R48 VDD.n9 VDD.n8 1.651
R49 VDD.n12 VDD.n10 1.157
R50 VDD.n12 VDD.n11 1.103
R51 VDD.n13 VDD.n12 0.241
R52 VDD.n13 VDD.n4 0.182
R53 VDD.n0 VDD.t9 0.124
R54 VDD.n4 VDD.n2 0.065
R55 VDD.n14 VDD 0.02
R56 VDD.n14 VDD.n13 0.004
R57 VDD VDD.n14 0.001
R58 VDD.n7 VDD.n6 0.001
R59 VDD.n13 VDD.n7 0.001
R60 B.t3 B.t0 800.071
R61 B B.n1 627.619
R62 B.n0 B.t1 285.109
R63 B.n1 B.t3 193.602
R64 B.n0 B.t2 160.666
R65 B.n1 B.n0 91.507
R66 VSS.n1 VSS.t0 18.459
R67 VSS.n0 VSS.t1 17.4
R68 VSS.n0 VSS.t2 17.4
R69 VSS.n1 VSS.n0 0.533
R70 VSS.n2 VSS.n1 0.17
R71 VSS VSS.n2 0.002
R72 OUT.n0 OUT.t1 28.57
R73 OUT.n1 OUT.t0 28.565
R74 OUT.n1 OUT.t2 28.565
R75 OUT.n0 OUT.t3 17.638
R76 OUT.n2 OUT.n1 0.69
R77 OUT.n2 OUT.n0 0.6
R78 OUT OUT.n2 0.199
R79 OUT OUT.n3 0.043
R80 OUT.n3 OUT 0.041
R81 OUT.n3 OUT 0.022
C0 A VDD 0.13fF
C1 A OUT 0.01fF
C2 B A 0.44fF
C3 OUT VDD 0.85fF
C4 B VDD 0.37fF
C5 B OUT 0.03fF
.ends

