* NGSPICE file created from aritmetic_unit_pex.ext - technology: sky130B

.subckt arithmetic_unit A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7] B[0],B[1],B[2],B[3],B[4],B[5],B[6],B[7] opcode[0],opcode[1] Y[0],Y[1],Y[2],Y[3],Y[4],Y[5],Y[6],Y[7] Cout VSS VDD
X0 VDD.t1424 a_4963_19248.t4 a_8998_20136.t3 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1 a_15556_20132.t6 a_11521_19244.t4 VDD.t2563 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2 a_5917_18826.t2 a_5860_19519.t8 VDD.t2590 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3 VDD.t2570 a_21150_9929.t8 a_31893_6205.t9 VDD.t2569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X4 a_13164_12246.t2 a_12900_12829.t5 VDD.t2613 VDD.t2612 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5 a_17946_9198.t0 a_17356_9635.t7 VSS.t196 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6 a_7735_24460.t2 a_n3111_15192.t8 VDD.t2400 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 a_9415_27296.t2 a_8419_26709.t4 VDD.t2340 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 VDD.t2500 A[3].t0 a_29769_12318.t3 VDD.t2499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X9 a_22462_27288.t5 a_21466_26701.t4 VDD.t2345 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 VDD.t2454 a_30430_6928.t4 a_33377_10390.t2 VDD.t2453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X11 a_31893_1857.t8 a_31466_2550.t4 a_32011_1857.t6 VDD.t2448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X12 VDD.t2523 a_17301_11213.t4 a_17356_9635.t4 VDD.t2522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X13 a_15570_21782.t0 A[6].t0 a_16219_21171.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 a_18991_21663.t3 a_20058_21029.t5 VDD.t2439 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X15 VDD.t2416 a_10641_5411.t4 a_14372_4127.t2 VDD.t2415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 a_14496_9997.t6 a_13951_10690.t4 a_14496_9265.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_8998_20136.t0 a_4963_19248.t5 a_9647_19525.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_12181_18848.t3 a_11523_19541.t4 a_12063_18848.t3 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_12592_4127.t3 a_12886_4101.t4 a_12474_4127.t5 VDD.t2342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 VDD.t2325 a_5899_21662.t4 a_5959_21688.t2 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X21 a_11277_6650.t3 a_10687_7087.t7 VDD.t2320 VDD.t2319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X22 a_13060_23726.t3 a_12470_24163.t7 VDD.t2232 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X23 a_7853_24460.t3 a_7308_25153.t4 a_7735_24460.t11 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X24 a_6966_21028.t3 a_7395_21658.t4 a_7101_21684.t3 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X25 a_4740_5002.t3 a_4150_5439.t7 VDD.t2305 VDD.t2304 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X26 VDD.t2293 a_6041_4129.t8 a_7394_4822.t3 VDD.t2292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X27 a_6552_25333.t0 a_5962_25770.t7 VSS.t393 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X28 VDD.t2370 a_14496_9997.t8 a_17361_11239.t2 VDD.t2369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X29 a_4735_3398.t0 a_4145_3835.t7 VSS.t390 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X30 VSS.t385 a_23918_5413.t4 a_24210_3198.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X31 a_n3111_15192.t4 a_n3604_15973.t4 a_n3804_15135.t2 VDD.t2077 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X32 a_18597_18853.t6 a_18055_19249.t4 VDD.t2080 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X33 a_1246_10551.t4 A[5].t0 VDD.t2124 VDD.t2123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X34 VSS.t360 a_4965_19545.t4 a_5623_18120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X35 a_15097_1774.t3 a_14507_1337.t7 VDD.t2174 VDD.t2173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X36 VDD.t2176 a_7947_9909.t8 a_31891_13791.t5 VDD.t2175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X37 a_14248_24457.t2 A[1].t0 VDD.t2161 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X38 a_33614_1910.t0 a_14490_4127.t8 a_33377_2547.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X39 VDD.t2082 B[5].t0 a_14467_15035.t2 VDD.t2081 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X40 a_10693_12957.t3 a_8508_14599.t4 VDD.t2042 VDD.t2041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X41 a_27000_21662.t3 a_28608_18536.t7 VDD.t1974 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X42 a_7953_1332.t3 B[5].t1 VDD.t2084 VDD.t2083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X43 VDD.t1978 B[4].t0 a_1227_7273.t2 VDD.t1977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X44 a_16074_26710.t0 a_15810_27293.t5 VSS.t338 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X45 VSS.t343 a_36755_23013.t8 Y[0].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X46 a_30359_11881.t3 a_29769_12318.t7 VDD.t2394 VDD.t2393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X47 a_n3115_713.t2 a_n3608_55.t4 a_n3808_656.t2 VDD.t1931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X48 VDD.t1923 a_25465_19523.t8 a_25110_18856.t3 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X49 a_n2381_8987.t0 a_n3606_9768.t4 a_n3113_8987.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X50 VDD.t1752 a_19554_12761.t5 a_19818_12178.t3 VDD.t1751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X51 a_31891_13791.t6 a_31464_14484.t4 a_32009_13791.t5 VDD.t1788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 VDD.t1807 opcode[0].t0 a_5957_24166.t2 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X53 a_36751_13711.t5 a_32011_1857.t8 VDD.t2555 VDD.t2554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X54 a_25759_9997.t8 a_20955_6381.t4 VDD.t1761 VDD.t1760 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X55 VDD.t2442 a_15570_21782.t7 a_13599_21654.t3 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 a_8998_20136.t2 a_4963_19248.t6 VDD.t1423 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 VDD.t2615 a_12900_12829.t6 a_13164_12246.t1 VDD.t2614 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X58 a_17356_5438.t6 a_17296_5412.t4 VDD.t1720 VDD.t1719 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X59 a_5496_4822.t3 a_1833_4076.t4 VDD.t1688 VDD.t1687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X60 VDD.t1658 a_1836_10114.t4 a_4144_12869.t2 VDD.t1657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X61 VDD.t2341 a_8419_26709.t5 a_9415_27296.t1 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X62 a_29769_12318.t2 A[3].t1 VDD.t2502 VDD.t2501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X63 VDD.t2346 a_21466_26701.t5 a_22462_27288.t4 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X64 a_13065_25330.t3 a_12475_25767.t7 VDD.t1644 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X65 a_14490_3395.t0 a_14784_4101.t4 VSS.t296 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X66 VDD.t1609 A[4].t0 a_7953_1332.t4 VDD.t1608 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X67 a_38088_20578.t0 a_16264_24457.t8 VSS.t298 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X68 a_n3606_7699.t0 opcode[0].t1 VSS.t327 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X69 a_14786_27289.t2 a_13051_26980.t4 VDD.t1596 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X70 VDD.t2440 a_20058_21029.t6 a_18991_21663.t2 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X71 a_21145_4128.t7 a_21439_4102.t4 a_21027_4128.t11 VDD.t744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X72 a_28617_21790.t6 a_n3113_6918.t8 VDD.t1401 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X73 a_12063_18848.t8 a_12475_18822.t4 a_12181_18848.t7 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X74 a_36751_16855.t7 opcode[1].t0 VDD.t1477 VDD.t1476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X75 a_16264_24457.t1 a_15719_25150.t4 a_16146_24457.t5 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X76 a_5959_21688.t1 a_5899_21662.t5 VDD.t2326 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X77 VDD.t2233 a_12470_24163.t8 a_13060_23726.t2 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X78 a_n3608_5631.t3 opcode[0].t2 VDD.t1809 VDD.t1808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 a_32305_9674.t0 a_30359_8848.t4 VSS.t266 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X80 a_21032_9929.t7 a_21444_9903.t4 a_21150_9929.t5 VDD.t1380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X81 a_21746_1762.t3 a_21156_1325.t7 VDD.t1471 VDD.t1470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X82 VDD.t558 a_18952_19520.t8 a_18597_18853.t8 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X83 VDD.t2044 a_8508_14599.t5 a_10702_9703.t4 VDD.t2043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X84 VDD.t2126 A[5].t1 a_1246_10551.t3 VDD.t2125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X85 VDD.t2162 A[1].t1 a_14660_24431.t3 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X86 VDD.t2163 A[1].t2 a_14248_24457.t1 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X87 a_29238_24456.t11 a_27458_24456.t8 VDD.t1014 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X88 a_17941_3397.t3 a_17351_3834.t7 VDD.t1030 VDD.t1029 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X89 VSS.t209 a_7939_4129.t8 a_12828_3395.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X90 a_31891_13791.t4 a_7947_9909.t9 VDD.t2178 VDD.t2177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X91 a_28902_27292.t3 a_26157_25329.t4 a_29020_27292.t5 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X92 VDD.t721 a_7749_6382.t4 a_10693_12957.t4 VDD.t720 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X93 VDD.t1975 a_28608_18536.t8 a_27000_21662.t2 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X94 a_n3111_15192.t3 opcode[0].t3 a_n2379_15428.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X95 VDD.t1429 a_4963_19248.t7 a_4965_19545.t3 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X96 VDD.t2396 a_29769_12318.t8 a_30359_11881.t2 VDD.t2395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X97 a_24568_5002.t0 a_23978_5439.t7 VSS.t214 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X98 a_n3808_4793.t5 a_n3608_4192.t4 a_n3115_4850.t2 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X99 a_7611_12745.t4 a_4748_10782.t4 a_7493_12745.t4 VDD.t761 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X100 a_5860_19519.t4 a_6863_19545.t4 a_7403_18852.t11 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X101 a_29356_24456.t6 a_28811_25149.t4 a_29238_24456.t6 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X102 a_38088_23722.t0 a_9751_24460.t8 VSS.t192 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X103 VDD.t854 B[3].t0 a_1243_4513.t6 VDD.t853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X104 a_4734_12432.t0 a_4144_12869.t7 VSS.t304 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X105 a_32009_13791.t4 a_31464_14484.t5 a_31891_13791.t8 VDD.t1790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X106 VDD.t1298 a_21202_27284.t5 a_21466_26701.t0 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X107 a_21027_4128.t6 a_19247_4128.t8 VDD.t869 VDD.t868 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X108 a_7829_9909.t7 a_7402_10602.t4 a_7947_9909.t3 VDD.t764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X109 a_30074_3658.t0 A[4].t1 a_29837_4295.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X110 a_4381_12232.t1 a_1844_12699.t4 a_4144_12869.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X111 VDD.t1422 a_4963_19248.t8 a_8998_20136.t1 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X112 VSS.t271 a_20900_24452.t8 a_22253_25145.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X113 a_25504_21666.t3 a_26571_21032.t5 VDD.t443 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X114 VDD.t2503 A[3].t2 a_27340_24456.t2 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X115 a_15928_27293.t5 a_13065_25330.t4 a_15810_27293.t1 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X116 a_27420_18830.t3 a_n3113_6918.t9 VDD.t1402 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X117 VSS.t177 a_24568_19252.t4 a_24570_19549.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X118 a_4144_12869.t1 a_1836_10114.t5 VDD.t1660 VDD.t1659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X119 a_7402_10602.t0 a_6049_9909.t8 VDD.t1302 VDD.t1301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X120 a_36751_1089.t11 opcode[1].t1 VDD.t1479 VDD.t1478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X121 a_18991_21663.t1 a_20058_21029.t7 VDD.t2441 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X122 VDD.t2180 a_7947_9909.t10 a_33375_14481.t6 VDD.t2179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X123 VDD.t1610 A[4].t2 a_28617_21790.t3 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X124 a_5505_18852.t5 a_5917_18826.t4 a_5623_18852.t6 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X125 a_12181_18848.t6 a_12475_18822.t5 a_12063_18848.t7 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X126 VDD.t1662 a_1836_10114.t6 a_4158_11219.t3 VDD.t1661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X127 a_5824_21032.t4 a_6253_21662.t4 a_5959_21688.t3 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X128 a_6343_9883.t3 a_1844_12699.t5 VDD.t1437 VDD.t1436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X129 a_n3804_10998.t2 a_n3604_10397.t4 a_n3111_11055.t2 VDD.t923 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X130 a_16146_24457.t4 a_15719_25150.t5 a_16264_24457.t2 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X131 a_12517_21684.t5 a_12811_21658.t4 a_12382_21028.t4 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X132 a_13060_23726.t1 a_12470_24163.t9 VDD.t2234 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X133 a_n3113_13124.t4 a_n3606_12466.t4 a_n3806_13067.t5 VDD.t767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X134 VDD.t569 a_n3111_11055.t8 a_20355_25145.t3 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X135 a_10930_12320.t0 a_8508_14599.t6 a_10693_12957.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X136 a_5923_4129.t9 a_1833_4076.t5 VDD.t1690 VDD.t1689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X137 VDD.t2127 A[5].t2 a_22104_21787.t6 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X138 a_1836_10114.t3 a_1246_10551.t7 VDD.t2066 VDD.t2065 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X139 a_14660_24431.t2 A[1].t3 VDD.t2164 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X140 VDD.t1433 a_8998_20136.t7 a_6253_21662.t3 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X141 VDD.t1015 a_27458_24456.t9 a_29238_24456.t10 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X142 a_29837_4295.t4 A[4].t3 VDD.t1612 VDD.t1611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X143 VDD.t1957 a_30359_11881.t4 a_31891_13791.t9 VDD.t1956 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X144 a_29020_27292.t4 a_26157_25329.t5 a_28902_27292.t2 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X145 a_15097_1774.t0 a_14507_1337.t8 VSS.t376 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X146 a_11291_5000.t3 a_10701_5437.t7 VDD.t1292 VDD.t1291 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X147 a_28608_18536.t0 a_24568_19252.t5 VDD.t911 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X148 VSS.t161 a_26468_19549.t4 a_27126_18124.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X149 VDD.t1036 a_7939_4129.t9 a_12886_4101.t0 VDD.t1035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X150 a_4965_19545.t2 a_4963_19248.t9 VDD.t1428 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X151 VDD.t2562 a_11521_19244.t5 a_11523_19541.t3 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X152 a_36755_10391.t5 a_36701_11276.t4 a_36755_10509.t9 VDD.t882 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X153 a_30359_11881.t1 a_29769_12318.t9 VDD.t2398 VDD.t2397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X154 VDD.t2144 a_14490_4127.t9 a_33377_2547.t2 VDD.t2143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X155 a_21145_4128.t0 a_20600_4821.t4 a_21145_3396.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X156 VDD.t680 a_8543_1769.t4 a_12047_4820.t3 VDD.t679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X157 VDD.t2128 A[5].t3 a_20495_18853.t11 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X158 a_n3806_13067.t7 B[1].t0 VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X159 a_28061_4103.t3 a_23918_5413.t5 VDD.t2236 VDD.t2235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X160 a_19134_9929.t2 a_14496_9997.t9 VDD.t2372 VDD.t2371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X161 a_36755_19987.t5 a_36701_20754.t4 a_36755_19869.t5 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X162 VDD.t2262 a_7853_24460.t8 a_9206_25153.t3 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X163 a_23973_3835.t6 a_21145_4128.t8 VDD.t1573 VDD.t1572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X164 a_25869_3397.t0 a_26163_4103.t4 VSS.t250 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X165 VDD.t1283 a_36755_7247.t8 Y[5].t3 VDD.t1282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X166 a_20809_6964.t5 a_19813_6377.t4 VDD.t1118 VDD.t1117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X167 a_8147_24434.t0 A[0].t0 VSS.t218 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X168 VDD.t1341 a_1817_6836.t4 a_5923_4129.t10 VDD.t1340 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X169 VDD.t1155 B[0].t0 a_n3604_14534.t3 VDD.t1154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X170 a_27340_24456.t1 A[3].t3 VDD.t2504 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X171 VDD.t237 a_14932_26706.t4 a_15928_27293.t0 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X172 VDD.t1316 a_21746_1762.t4 a_23978_5439.t6 VDD.t1315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X173 VSS.t318 a_15097_1774.t4 a_17593_4801.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X174 VDD.t689 a_22095_18533.t7 a_20487_21659.t3 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X175 a_24568_19252.t0 a_28902_27292.t5 VSS.t205 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X176 VDD.t1664 a_1836_10114.t7 a_4144_12869.t0 VDD.t1663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X177 VDD.t1304 a_6049_9909.t9 a_7402_10602.t1 VDD.t1303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X178 a_14490_4127.t1 a_13945_4820.t4 a_14372_4127.t3 VDD.t636 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X179 a_19252_9929.t3 a_18707_10622.t4 a_19134_9929.t6 VDD.t1100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X180 a_36697_5000.t3 opcode[1].t2 VDD.t1481 VDD.t1480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X181 a_28069_9971.t3 a_23926_11281.t4 VDD.t1262 VDD.t1261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X182 a_33375_14481.t5 a_7947_9909.t11 VDD.t2182 VDD.t2181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X183 a_28617_21790.t2 A[4].t4 VDD.t1613 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X184 VDD.t1240 a_27775_9997.t8 a_36751_4233.t11 VDD.t1239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X185 a_5959_21688.t4 a_6253_21662.t5 a_5824_21032.t3 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X186 a_16264_24457.t3 a_15719_25150.t6 a_16146_24457.t3 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X187 VDD.t553 a_32011_9700.t8 a_36755_19987.t6 VDD.t552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X188 a_21136_23720.t0 a_n3111_11055.t9 a_20900_24452.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X189 a_22608_26705.t3 a_22344_27288.t5 VDD.t1140 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X190 a_19252_9197.t1 a_19546_9903.t4 VSS.t245 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X191 a_24568_5002.t3 a_23978_5439.t8 VDD.t1059 VDD.t1058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X192 VDD.t1094 A[0].t1 a_5948_27420.t6 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X193 a_12892_9971.t0 a_8508_14599.t7 VSS.t361 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X194 a_32011_5473.t1 a_32305_6179.t4 VSS.t48 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X195 VDD.t1575 a_21145_4128.t9 a_26163_4103.t3 VDD.t1574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X196 a_14496_9997.t5 a_13951_10690.t5 a_14378_9997.t9 VDD.t2353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X197 VDD.t2568 a_21150_9929.t9 a_31893_6205.t8 VDD.t2567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X198 a_26157_25329.t1 a_25567_25766.t7 VDD.t1170 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X199 VDD.t871 a_19247_4128.t9 a_20600_4821.t3 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X200 VSS.t339 a_16074_26710.t4 a_19241_23521.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X201 VDD.t1271 B[7].t0 a_n3608_55.t0 VDD.t1270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X202 a_36755_7365.t7 opcode[1].t3 VDD.t1483 VDD.t1482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X203 a_27878_27288.t5 a_26152_23725.t4 a_27760_27288.t4 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X204 a_20495_18853.t10 A[5].t4 VDD.t2129 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X205 VDD.t2374 a_14496_9997.t10 a_19134_9929.t1 VDD.t2373 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X206 a_n3113_13124.t1 opcode[0].t4 a_n2381_13360.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X207 a_6041_3397.t0 a_6335_4103.t4 VSS.t159 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X208 a_9206_25153.t2 a_7853_24460.t9 VDD.t2263 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X209 a_36755_23131.t3 a_9751_24460.t9 a_36755_23013.t4 VDD.t967 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X210 a_5917_18826.t3 a_5860_19519.t9 VSS.t197 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X211 VDD.t2525 a_17301_11213.t5 a_17356_9635.t5 VDD.t2524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X212 a_15928_27293.t1 a_14932_26706.t5 VDD.t238 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X213 a_17579_6451.t1 a_14306_12250.t4 a_17342_7088.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X214 a_5962_25770.t3 opcode[0].t5 VDD.t1810 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X215 a_36697_17622.t3 opcode[1].t4 VDD.t1485 VDD.t1484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X216 a_36755_7247.t4 a_36701_8132.t4 a_36755_7365.t9 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X217 a_4734_12432.t3 a_4144_12869.t8 VDD.t1648 VDD.t1647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X218 VDD.t81 a_12894_6959.t5 a_13158_6376.t3 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X219 a_19667_6960.t5 a_17941_3397.t4 a_19549_6960.t4 VDD.t1033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X220 VDD.t1264 a_23926_11281.t5 a_28069_9971.t2 VDD.t1263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X221 VDD.t1614 A[4].t5 a_28617_21790.t1 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X222 VDD.t682 a_8543_1769.t5 a_12474_4127.t0 VDD.t681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X223 a_27340_24456.t5 a_27752_24430.t4 a_27458_24456.t3 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X224 a_36701_23898.t3 opcode[1].t5 VDD.t1487 VDD.t1486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X225 a_31893_1857.t0 a_32305_1831.t4 a_32011_1857.t1 VDD.t283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X226 a_26571_21032.t0 a_26646_21662.t4 VSS.t128 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X227 VDD.t610 a_4090_5413.t4 a_4145_3835.t1 VDD.t609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X228 VSS.t127 A[2].t0 a_21136_23720.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X229 a_24576_10870.t0 a_23986_11307.t7 VSS.t96 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X230 VDD.t138 a_1254_13136.t7 a_1844_12699.t0 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X231 a_27321_12833.t3 a_24576_10870.t4 VSS.t251 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X232 a_14154_6963.t5 a_11291_5000.t4 a_14036_6963.t4 VDD.t896 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X233 a_5948_27420.t5 A[0].t2 VDD.t1095 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X234 a_n3606_3562.t3 opcode[0].t6 VDD.t1812 VDD.t1811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X235 a_22798_23720.t1 a_23092_24426.t4 VSS.t220 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X236 a_n3113_6918.t1 a_n3606_6260.t4 a_n3806_6861.t5 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X237 VDD.t645 a_12418_19515.t8 a_12063_18848.t0 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X238 a_12480_9997.t11 a_7749_6382.t5 VDD.t723 VDD.t722 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X239 VSS.t157 a_12382_21028.t5 a_4963_19248.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X240 a_n3115_4850.t3 opcode[0].t7 a_n2383_5086.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X241 VDD.t255 a_17932_6651.t4 a_19667_6960.t0 VDD.t254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X242 a_7939_4129.t4 a_7394_4822.t4 a_7821_4129.t4 VDD.t2285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X243 a_12834_9265.t1 a_7749_6382.t6 a_12598_9997.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X244 VDD.t1171 a_25567_25766.t8 a_26157_25329.t2 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X245 a_n3606_9768.t0 opcode[0].t8 VDD.t1814 VDD.t1813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X246 VDD.t240 a_26143_26979.t4 a_27878_27288.t0 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X247 VDD.t706 B[1].t1 a_n3606_12466.t0 VDD.t705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X248 a_10641_5411.t0 a_33375_14481.t7 VSS.t235 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X249 VDD.t1368 a_n3115_4850.t8 a_20495_18853.t8 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X250 a_n3606_7699.t3 opcode[0].t9 VDD.t1816 VDD.t1815 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X251 a_19134_9929.t0 a_14496_9997.t11 VDD.t2376 VDD.t2375 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X252 VDD.t2238 a_23918_5413.t6 a_27649_4129.t11 VDD.t2237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X253 VDD.t99 a_12598_9997.t8 a_14378_9997.t0 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X254 a_26152_23725.t0 a_25562_24162.t7 VDD.t413 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X255 VSS.t347 a_n3608_55.t5 a_n2383_713.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X256 a_27752_24430.t3 A[3].t4 VDD.t2505 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X257 a_33377_6895.t3 a_21150_9929.t10 VDD.t2566 VDD.t2565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X258 a_6335_4103.t3 a_1817_6836.t5 VDD.t1343 VDD.t1342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X259 a_32009_13791.t3 a_31464_14484.t6 a_31891_13791.t7 VDD.t1789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X260 a_36751_13711.t9 opcode[1].t6 VDD.t1489 VDD.t1488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X261 VSS.t143 a_8543_1769.t6 a_10924_6450.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X262 a_36755_10509.t6 opcode[1].t7 VDD.t1491 VDD.t1490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X263 VDD.t2463 A[6].t1 a_13961_18848.t4 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X264 a_17356_5438.t5 a_17296_5412.t5 VDD.t1722 VDD.t1721 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X265 a_28069_9971.t1 a_23926_11281.t6 VDD.t1266 VDD.t1265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X266 a_1817_6836.t3 a_1227_7273.t7 VDD.t1792 VDD.t1791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X267 VDD.t791 a_10647_11281.t4 a_10702_9703.t5 VDD.t790 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X268 a_27420_18830.t2 a_n3113_6918.t10 VDD.t1403 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X269 VSS.t342 a_27000_21662.t4 a_26571_21032.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X270 a_25465_19523.t3 a_27420_18830.t4 a_27008_18856.t11 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X271 a_36701_23898.t0 opcode[1].t8 VSS.t284 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X272 VDD.t1219 a_36751_971.t8 Y[7].t3 VDD.t1218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X273 VDD.t1345 a_1817_6836.t6 a_4136_7089.t3 VDD.t1344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X274 a_27431_6965.t3 a_24568_5002.t4 a_27313_6965.t3 VDD.t1055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X275 VDD.t1102 a_30427_3858.t4 a_33377_6895.t4 VDD.t1101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X276 VSS.t225 a_n3606_8329.t4 a_n2381_8987.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X277 VDD.t2401 a_n3111_15192.t9 a_5948_27420.t2 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X278 VDD.t2465 A[6].t2 a_1243_4513.t2 VDD.t2464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X279 a_21027_4128.t7 a_19247_4128.t10 VDD.t873 VDD.t872 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X280 VDD.t1616 A[4].t6 a_29769_9285.t3 VDD.t1615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X281 a_25751_4129.t8 a_21746_1762.t5 VDD.t1318 VDD.t1317 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X282 a_10647_11281.t3 a_14036_6963.t5 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X283 a_12063_18848.t1 a_12418_19515.t9 VDD.t646 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X284 a_10701_5437.t3 a_10641_5411.t5 VDD.t2418 VDD.t2417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X285 a_27760_27288.t1 a_26152_23725.t5 VSS.t253 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X286 a_24571_9266.t3 a_23981_9703.t7 VDD.t485 VDD.t484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X287 VDD.t2130 A[5].t5 a_22095_18533.t6 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X288 VDD.t1818 opcode[0].t10 a_n3608_1494.t3 VDD.t1817 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X289 a_26179_12829.t2 a_24571_9266.t4 VSS.t83 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X290 a_26157_25329.t3 a_25567_25766.t9 VDD.t1172 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X291 a_27878_27288.t1 a_26143_26979.t5 VDD.t241 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X292 a_12475_25767.t0 a_9561_26713.t4 VDD.t488 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X293 VDD.t1820 opcode[0].t11 a_n3608_5631.t2 VDD.t1819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X294 VDD.t1666 a_1836_10114.t8 a_5504_10602.t3 VDD.t1665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X295 a_1254_13136.t3 A[4].t7 VDD.t1618 VDD.t1617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X296 VDD.t1938 a_n3115_713.t8 a_7403_18852.t3 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X297 a_16558_24431.t0 a_9561_26713.t5 VSS.t95 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X298 VDD.t660 a_6343_6961.t5 a_6607_6378.t3 VDD.t659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X299 a_n2379_11055.t0 a_n3604_11836.t4 a_n3111_11055.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X300 a_1833_4076.t1 a_1243_4513.t7 VDD.t856 VDD.t855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X301 VDD.t2561 a_11521_19244.t6 a_15561_18528.t6 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X302 a_10696_3833.t6 a_10641_5411.t6 VDD.t2420 VDD.t2419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X303 a_29840_7365.t2 A[3].t5 VDD.t2507 VDD.t2506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X304 a_21032_9929.t1 a_19252_9929.t8 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X305 VDD.t665 a_n3113_13124.t8 a_13821_25150.t3 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X306 a_33614_9753.t0 a_30359_8848.t5 a_33377_10390.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X307 VDD.t1404 a_n3113_6918.t11 a_27420_18830.t1 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X308 a_29837_4295.t6 B[6].t0 VDD.t754 VDD.t753 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X309 a_38088_8192.t1 opcode[1].t9 a_36755_7247.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X310 a_27008_18856.t10 a_27420_18830.t5 a_25465_19523.t4 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X311 VDD.t1980 B[4].t1 a_n3606_6260.t3 VDD.t1979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X312 a_36697_14478.t0 opcode[1].t10 VSS.t285 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X313 a_6049_9909.t5 a_5504_10602.t4 a_5931_9909.t8 VDD.t1012 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X314 a_28608_18536.t3 A[4].t8 a_29257_17925.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X315 a_7603_6965.t5 a_4740_5002.t4 a_7485_6965.t1 VDD.t2290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X316 a_30364_14452.t3 a_29774_14889.t7 VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X317 a_5948_27420.t1 a_n3111_15192.t10 VDD.t2402 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X318 VSS.t313 a_17296_5412.t6 a_21381_3396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X319 a_38084_17682.t1 opcode[1].t11 a_36751_16737.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X320 VDD.t276 a_10696_3833.t7 a_11286_3396.t3 VDD.t275 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X321 VDD.t647 a_12418_19515.t10 a_12063_18848.t2 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X322 a_13012_6959.t5 a_11286_3396.t4 a_12894_6959.t0 VDD.t218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X323 VSS.t54 a_26143_26979.t6 a_27760_27288.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X324 VDD.t1493 opcode[1].t12 a_36697_1856.t3 VDD.t1492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X325 a_17342_7088.t2 a_15097_1774.t5 VDD.t2205 VDD.t2204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X326 a_30011_14252.t1 B[3].t1 a_29774_14889.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X327 a_22095_18533.t5 A[5].t6 VDD.t2131 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X328 VSS.t189 a_24562_12520.t4 a_26179_12829.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X329 a_19594_23721.t0 a_19004_24158.t7 VSS.t229 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X330 VDD.t489 a_9561_26713.t6 a_12475_25767.t1 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X331 VDD.t1982 B[4].t2 a_29840_7365.t6 VDD.t1981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X332 VDD.t912 a_24568_19252.t6 a_28603_20140.t6 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X333 a_12470_24163.t3 A[1].t4 VDD.t2165 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X334 a_14490_4127.t2 a_13945_4820.t5 a_14372_4127.t4 VDD.t880 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X335 a_19549_6960.t1 a_17941_3397.t5 VSS.t208 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X336 a_36751_1089.t6 a_5623_18852.t8 a_36751_971.t4 VDD.t633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X337 a_5504_10602.t2 a_1836_10114.t9 VDD.t1668 VDD.t1667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X338 a_7403_18852.t2 a_n3115_713.t9 VDD.t1939 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X339 a_n3806_13067.t11 a_n3606_13905.t4 a_n3113_13124.t7 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X340 a_27878_27288.t4 a_26152_23725.t6 a_27760_27288.t3 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X341 a_15561_18528.t5 a_11521_19244.t7 VDD.t2560 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X342 a_20849_18121.t1 A[5].t7 VSS.t369 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X343 VSS.t238 a_30427_3858.t5 a_33614_6258.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X344 VDD.t656 a_22104_21787.t7 a_20133_21659.t3 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X345 a_12894_6959.t1 a_11286_3396.t5 a_13012_6959.t4 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X346 VDD.t2193 a_18055_19249.t5 a_22090_20137.t3 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X347 VDD.t402 a_4153_9615.t7 a_4743_9178.t3 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X348 a_19129_4128.t6 a_19541_4102.t4 a_19247_4128.t3 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X349 a_28603_20140.t3 a_24568_19252.t7 a_29252_19529.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X350 VDD.t176 a_19252_9929.t9 a_21032_9929.t2 VDD.t175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X351 a_10687_7087.t3 a_7939_4129.t10 VDD.t1038 VDD.t1037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X352 a_16074_26710.t3 a_15810_27293.t6 VDD.t1757 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X353 VDD.t446 a_22608_26705.t4 a_29650_24430.t3 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X354 VSS.t134 a_9012_21786.t7 a_7041_21658.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X355 VSS.t144 a_8543_1769.t7 a_10938_4800.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X356 VDD.t1933 a_36755_23013.t9 Y[0].t3 VDD.t1932 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X357 a_14373_18822.t0 a_n3113_2781.t8 VSS.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X358 VDD.t1157 B[0].t1 a_n3804_15135.t6 VDD.t1156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X359 VDD.t1495 opcode[1].t13 a_36751_4233.t8 VDD.t1494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X360 a_14507_1337.t3 B[5].t2 VDD.t2086 VDD.t2085 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X361 Y[2].t3 a_36751_16737.t8 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X362 a_5899_21662.t0 a_6966_21028.t5 VDD.t2291 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X363 VSS.t278 a_15556_20132.t7 a_12811_21658.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X364 VDD.t1320 a_21746_1762.t6 a_25324_4822.t3 VDD.t1319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X365 a_36701_11276.t3 opcode[1].t14 VDD.t1497 VDD.t1496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X366 a_4743_9178.t2 a_4153_9615.t8 VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X367 a_20900_24452.t4 a_20355_25145.t4 a_20900_23720.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X368 VSS.t122 a_6607_6378.t4 a_7485_6965.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X369 a_12474_4127.t9 a_12047_4820.t4 a_12592_4127.t4 VDD.t1151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X370 a_28024_26705.t0 a_27760_27288.t5 VSS.t193 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X371 a_12598_9997.t3 a_12053_10690.t4 a_12480_9997.t6 VDD.t600 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X372 a_22680_24452.t8 a_20900_24452.t9 VDD.t1413 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X373 a_26443_12246.t0 a_26179_12829.t5 VSS.t74 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X374 VDD.t1499 opcode[1].t15 a_36701_20754.t3 VDD.t1498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X375 a_12475_25767.t2 a_9561_26713.t7 VDD.t490 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X376 VSS.t305 a_1836_10114.t10 a_5504_10602.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X377 a_5505_18852.t11 a_4963_19248.t10 VDD.t1427 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X378 a_14790_9971.t3 a_10647_11281.t5 VDD.t793 VDD.t792 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X379 a_27767_4129.t7 a_27222_4822.t4 a_27649_4129.t2 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X380 a_19599_25325.t0 a_19009_25762.t7 VSS.t31 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X381 a_15057_14598.t0 a_14467_15035.t7 VSS.t359 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X382 VSS.t216 a_18916_21033.t5 a_11521_19244.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X383 a_9003_18532.t3 A[7].t0 VDD.t206 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X384 VSS.t400 a_11277_6650.t4 a_12894_6959.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X385 a_27230_10690.t3 a_25877_9997.t8 VDD.t221 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X386 a_7829_9909.t8 a_4098_11193.t4 VDD.t981 VDD.t980 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X387 VDD.t1940 a_n3115_713.t10 a_7403_18852.t1 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X388 a_1227_7273.t6 A[5].t8 VDD.t2133 VDD.t2132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X389 a_14704_14398.t1 A[5].t9 a_14467_15035.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X390 a_36755_19987.t7 a_32011_9700.t9 VDD.t555 VDD.t554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X391 a_26171_9971.t3 a_21711_14619.t4 VDD.t400 VDD.t399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X392 a_27760_27288.t2 a_26152_23725.t7 a_27878_27288.t3 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X393 VDD.t970 a_27760_27288.t6 a_28024_26705.t3 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X394 a_20133_21659.t2 a_22104_21787.t8 VDD.t657 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X395 a_25759_9997.t10 a_26171_9971.t4 a_25877_9997.t7 VDD.t974 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X396 a_25228_18856.t7 a_24570_19549.t4 a_25110_18856.t9 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X397 a_n3115_4850.t1 a_n3608_4192.t5 a_n3808_4793.t4 VDD.t1367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X398 a_21032_9929.t3 a_19252_9929.t10 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X399 a_12480_9997.t2 a_12892_9971.t4 a_12598_9997.t2 VDD.t624 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X400 a_10045_24434.t3 opcode[0].t12 VDD.t1821 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X401 a_n3806_2724.t10 B[6].t1 VDD.t756 VDD.t755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X402 VDD.t1758 a_15810_27293.t7 a_16074_26710.t2 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X403 a_29650_24430.t2 a_22608_26705.t5 VDD.t447 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X404 a_27649_4129.t6 a_28061_4103.t4 a_27767_4129.t2 VDD.t1136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X405 VDD.t978 a_9003_18532.t7 a_7395_21658.t3 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X406 VDD.t232 a_25553_27416.t7 a_26143_26979.t1 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X407 a_7735_24460.t1 a_n3111_15192.t11 VDD.t2403 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X408 VSS.t140 a_n3113_13124.t9 a_13821_25150.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X409 VSS.t100 a_13953_21654.t4 a_13524_21024.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X410 a_17598_10602.t1 a_17301_11213.t6 a_17361_11239.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X411 VSS.t78 a_36751_4115.t8 Y[6].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X412 VDD.t2269 a_4145_3835.t8 a_4735_3398.t3 VDD.t2268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X413 a_31893_9700.t5 a_31466_10393.t4 a_32011_9700.t2 VDD.t248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X414 a_17946_9198.t3 a_17356_9635.t8 VDD.t2606 VDD.t2605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X415 a_36755_23013.t5 a_9751_24460.t10 a_36755_23131.t2 VDD.t968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X416 a_14154_6963.t4 a_11291_5000.t5 a_14036_6963.t3 VDD.t897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X417 a_36755_23131.t0 a_30364_14452.t4 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X418 a_1844_12699.t1 a_1254_13136.t8 VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X419 VDD.t1795 a_n3113_8987.t8 a_26913_25149.t3 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X420 VDD.t1823 opcode[0].t13 a_n3806_8930.t5 VDD.t1822 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X421 a_36751_16855.t0 a_22798_24452.t8 a_36751_16737.t0 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X422 a_30359_8848.t0 a_29769_9285.t7 VDD.t1144 VDD.t1143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X423 VSS.t410 a_14496_9997.t12 a_18707_10622.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X424 a_32303_13765.t3 a_30359_11881.t5 VDD.t1959 VDD.t1958 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X425 VDD.t1501 opcode[1].t16 a_36697_17622.t2 VDD.t1500 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X426 a_24554_6652.t0 a_23964_7089.t7 VSS.t34 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X427 VDD.t1825 opcode[0].t14 a_n3806_6861.t2 VDD.t1824 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X428 a_19585_26975.t0 a_18995_27412.t7 VSS.t113 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X429 VDD.t758 B[6].t2 a_21156_1325.t3 VDD.t757 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X430 VDD.t114 a_26171_6961.t5 a_26435_6378.t3 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X431 VDD.t1426 a_4963_19248.t11 a_5505_18852.t10 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X432 a_18715_18853.t6 a_18057_19546.t4 a_18597_18853.t7 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X433 a_23981_9703.t1 a_21711_14619.t5 VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X434 a_18916_21033.t4 a_18991_21663.t4 VSS.t416 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X435 VDD.t564 A[7].t1 a_9003_18532.t2 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X436 VDD.t149 a_25877_9997.t9 a_27230_10690.t2 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X437 VDD.t144 a_4098_11193.t5 a_7829_9909.t0 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X438 a_n2379_15192.t0 a_n3604_15973.t5 a_n3111_15192.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X439 VDD.t45 a_36751_4115.t9 Y[6].t3 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X440 a_17356_5438.t2 a_15097_1774.t6 VDD.t2207 VDD.t2206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X441 a_22680_24452.t11 a_23092_24426.t5 a_22798_24452.t7 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X442 VSS.t324 a_n3113_8987.t9 a_26913_25149.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X443 a_21386_9197.t1 a_19252_9929.t11 a_21150_9929.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X444 VDD.t1619 A[4].t9 a_26468_19549.t3 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X445 a_32305_1831.t3 a_14490_4127.t10 VDD.t2146 VDD.t2145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X446 VSS.t364 B[5].t3 a_14704_14398.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X447 VSS.t119 a_n3111_11055.t10 a_19246_25125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X448 a_n3806_2724.t7 a_n3606_3562.t4 a_n3113_2781.t5 VDD.t1196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X449 a_28024_26705.t2 a_27760_27288.t7 VDD.t971 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X450 VDD.t658 a_22104_21787.t9 a_20133_21659.t1 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X451 a_31893_9700.t11 a_30430_6928.t5 VDD.t2456 VDD.t2455 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X452 a_n2383_713.t1 a_n3608_1494.t4 a_n3115_713.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X453 a_25110_18856.t0 a_25522_18830.t4 a_25228_18856.t0 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X454 VDD.t2134 A[5].t10 a_19955_19546.t3 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X455 a_7821_4129.t0 a_8233_4103.t4 a_7939_4129.t0 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X456 a_7395_21658.t0 a_9003_18532.t8 VDD.t116 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X457 a_17301_11213.t0 a_33377_2547.t7 VSS.t368 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X458 a_19004_24158.t6 a_16074_26710.t5 VDD.t1915 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X459 a_25751_4129.t11 a_21145_4128.t10 VDD.t1577 VDD.t1576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X460 a_32011_6205.t6 a_31466_6898.t4 a_31893_6205.t2 VDD.t215 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X461 a_14036_6963.t1 a_11291_5000.t6 VSS.t173 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X462 VDD.t570 a_n3111_11055.t11 a_19009_25762.t2 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X463 a_8233_4103.t0 a_4090_5413.t5 VSS.t124 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X464 a_26143_26979.t0 a_25553_27416.t8 VDD.t212 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X465 a_13961_18848.t3 A[6].t3 VDD.t2466 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X466 a_10701_5437.t2 a_10641_5411.t7 VDD.t2422 VDD.t2421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X467 a_26706_21688.t2 a_26646_21662.t5 VDD.t622 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X468 VSS.t411 a_14496_9997.t13 a_17598_10602.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X469 a_n2383_949.t0 B[7].t1 VSS.t246 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X470 VDD.t1692 a_1833_4076.t6 a_4136_7089.t6 VDD.t1691 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X471 a_38084_4824.t0 a_12181_18848.t8 VSS.t408 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X472 VDD.t520 a_30434_1013.t4 a_31466_2550.t2 VDD.t519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X473 a_24568_19252.t3 a_28902_27292.t6 VDD.t1020 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X474 VSS.t256 a_21746_1762.t7 a_24201_6452.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X475 VSS.t70 a_4098_11193.t6 a_4390_8978.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X476 a_36751_13593.t6 a_36697_14478.t4 a_36751_13711.t7 VDD.t1168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X477 VDD.t1961 a_30359_11881.t6 a_32303_13765.t2 VDD.t1960 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X478 a_4963_19248.t1 a_12382_21028.t6 VDD.t779 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X479 a_4726_6652.t0 a_4136_7089.t7 VSS.t240 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X480 a_4748_10782.t0 a_4158_11219.t7 VSS.t207 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X481 a_20193_21685.t5 a_20133_21659.t4 VDD.t953 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X482 a_21027_4128.t3 a_17296_5412.t7 VDD.t1724 VDD.t1723 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X483 VSS.t277 a_11521_19244.t8 a_11523_19541.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X484 a_11292_9266.t3 a_10702_9703.t7 VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X485 a_5505_18852.t9 a_4963_19248.t12 VDD.t1425 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X486 VDD.t559 a_18952_19520.t9 a_18597_18853.t9 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X487 a_26171_6961.t0 a_24563_3398.t4 a_26289_6961.t2 VDD.t189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X488 a_36755_10509.t10 a_25228_18856.t8 a_36755_10391.t6 VDD.t979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X489 a_4395_10582.t1 a_4098_11193.t7 a_4158_11219.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X490 a_18597_18853.t2 a_18057_19546.t5 a_18715_18853.t5 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X491 VSS.t112 a_30434_1013.t5 a_31466_2550.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X492 a_8241_9883.t3 a_4098_11193.t8 VDD.t700 VDD.t699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X493 VSS.t0 a_19345_21663.t4 a_18916_21033.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X494 a_30430_6928.t0 a_29840_7365.t7 VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X495 VSS.t319 a_20955_6381.t5 a_25332_10690.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X496 a_27008_18856.t2 A[4].t10 VDD.t1620 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X497 a_26468_19549.t2 A[4].t11 VDD.t1621 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X498 VSS.t195 a_4098_11193.t9 a_8183_9177.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X499 a_27439_12833.t2 a_24576_10870.t5 a_27321_12833.t2 VDD.t1293 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X500 a_38088_11336.t1 opcode[1].t17 a_36755_10391.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X501 VDD.t1827 opcode[0].t15 a_n3804_15135.t9 VDD.t1826 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X502 VDD.t972 a_27760_27288.t8 a_28024_26705.t1 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X503 VSS.t403 a_12592_4127.t8 a_13945_4820.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X504 VDD.t2458 a_30430_6928.t6 a_31893_9700.t10 VDD.t2457 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X505 VDD.t1714 a_19818_12178.t4 a_20814_12765.t5 VDD.t1713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X506 a_7603_6965.t4 a_4740_5002.t5 a_7485_6965.t4 VDD.t2289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X507 a_25228_18856.t4 a_25522_18830.t5 a_25110_18856.t5 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X508 a_36697_5000.t2 opcode[1].t18 VDD.t1503 VDD.t1502 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X509 VDD.t642 a_9012_21786.t8 a_7041_21658.t3 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X510 VSS.t117 a_32011_9700.t10 a_38088_20814.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X511 a_15561_18528.t4 a_11521_19244.t9 VDD.t2564 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X512 a_10944_10670.t1 a_10647_11281.t6 a_10707_11307.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X513 VSS.t29 a_13421_19541.t4 a_14079_18116.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X514 VDD.t1916 a_16074_26710.t6 a_19004_24158.t5 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X515 a_19009_25762.t1 a_n3111_11055.t12 VDD.t571 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X516 VDD.t2166 A[1].t5 a_12461_27417.t3 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X517 a_29844_1450.t6 B[6].t3 VDD.t760 VDD.t759 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X518 VDD.t305 a_26646_21662.t6 a_26706_21688.t1 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X519 a_19672_12761.t5 a_17937_12452.t4 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X520 VDD.t955 a_36755_10391.t8 Y[4].t3 VDD.t954 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X521 VDD.t478 a_30434_1013.t6 a_33377_2547.t4 VDD.t477 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X522 VSS.t434 a_17301_11213.t7 a_17593_8998.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X523 VDD.t1021 a_28902_27292.t7 a_24568_19252.t2 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X524 VSS.t73 a_n3604_10397.t5 a_n2379_11055.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X525 a_20058_21029.t0 a_20487_21659.t4 a_20193_21685.t2 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X526 a_6343_6961.t0 a_4735_3398.t4 a_6461_6961.t2 VDD.t2259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X527 VDD.t2591 a_5860_19519.t10 a_5505_18852.t8 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X528 VSS.t306 a_1836_10114.t11 a_4395_10582.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X529 a_18715_18853.t4 a_18057_19546.t6 a_18597_18853.t0 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X530 VDD.t1322 a_21746_1762.t8 a_23978_5439.t5 VDD.t1321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X531 a_25522_18830.t0 a_25465_19523.t9 VSS.t341 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X532 a_12900_12829.t4 a_11292_9266.t4 a_13018_12829.t3 VDD.t984 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X533 Y[4].t2 a_36755_10391.t9 VDD.t957 VDD.t956 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X534 a_19129_4128.t5 a_19541_4102.t5 a_19247_4128.t0 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X535 VDD.t1622 A[4].t12 a_27008_18856.t1 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X536 a_28608_18536.t1 a_24568_19252.t8 VDD.t913 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X537 VDD.t1623 A[4].t13 a_26468_19549.t1 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X538 VDD.t347 a_20691_6964.t5 a_20955_6381.t3 VDD.t346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X539 a_10933_3196.t0 a_7939_4129.t11 a_10696_3833.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X540 VDD.t716 a_30434_1013.t7 a_31893_1857.t4 VDD.t715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X541 VDD.t169 a_26443_12246.t4 a_27439_12833.t5 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X542 a_17301_11213.t1 a_33377_2547.t8 VDD.t2118 VDD.t2117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X543 VSS.t171 a_25869_4129.t8 a_27222_4822.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X544 a_27657_9997.t2 a_27230_10690.t4 a_27775_9997.t7 VDD.t1001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X545 a_19252_9929.t5 a_19546_9903.t5 a_19134_9929.t7 VDD.t1267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X546 a_4743_9178.t0 a_4153_9615.t9 VSS.t33 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X547 a_14490_4127.t5 a_14784_4101.t5 a_14372_4127.t6 VDD.t1599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X548 a_31893_9700.t9 a_30430_6928.t7 VDD.t2460 VDD.t2459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X549 a_20814_12765.t4 a_19818_12178.t5 VDD.t1716 VDD.t1715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X550 a_n3806_6861.t8 B[4].t3 VDD.t1984 VDD.t1983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X551 VSS.t116 B[6].t4 a_21358_14419.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X552 a_22798_24452.t3 a_22253_25145.t4 a_22680_24452.t3 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X553 a_36755_7365.t3 a_18715_18853.t8 a_36755_7247.t0 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X554 a_9012_21786.t3 a_n3115_713.t11 VDD.t1941 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X555 a_36701_23898.t2 opcode[1].t19 VDD.t1505 VDD.t1504 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X556 a_27420_18830.t0 a_n3113_6918.t12 VSS.t268 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X557 a_6461_6961.t5 a_4726_6652.t4 VDD.t990 VDD.t989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X558 a_17356_9635.t0 a_15057_14598.t4 VDD.t261 VDD.t260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X559 a_19594_23721.t3 a_19004_24158.t8 VDD.t963 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X560 a_14315_18116.t0 A[6].t4 VSS.t424 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X561 a_14372_4127.t9 a_12592_4127.t9 VDD.t2329 VDD.t2328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X562 VDD.t496 a_23972_12957.t7 a_24562_12520.t3 VDD.t495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X563 a_22090_20137.t2 a_18055_19249.t6 VDD.t2194 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X564 a_12461_27417.t2 A[1].t6 VDD.t2167 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X565 a_12474_4127.t4 a_12886_4101.t5 a_12592_4127.t2 VDD.t2343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X566 a_n3113_2781.t0 a_n3606_2123.t4 a_n3806_2724.t0 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X567 a_1464_6636.t1 A[5].t11 a_1227_7273.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X568 a_26706_21688.t0 a_26646_21662.t7 VDD.t306 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X569 a_14372_4127.t7 a_14784_4101.t6 a_14490_4127.t6 VDD.t1600 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X570 a_31893_1857.t9 a_14490_4127.t11 VDD.t2148 VDD.t2147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X571 a_17937_12452.t3 a_17347_12889.t7 VSS.t105 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X572 VDD.t2209 a_15097_1774.t7 a_19129_4128.t2 VDD.t2208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X573 a_8233_4103.t3 a_4090_5413.t6 VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X574 VDD.t38 a_14366_24457.t8 a_16146_24457.t1 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X575 a_n3113_6918.t2 a_n3606_6260.t5 a_n3806_6861.t4 VDD.t309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X576 a_17584_12252.t1 a_15057_14598.t5 a_17347_12889.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X577 a_20782_24452.t2 a_n3111_11055.t13 VDD.t572 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X578 a_32011_1857.t5 a_31466_2550.t5 a_31893_1857.t7 VDD.t2447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X579 a_4145_3835.t4 a_1817_6836.t7 VDD.t1347 VDD.t1346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X580 VSS.t212 a_n3608_4192.t6 a_n2383_4850.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X581 VDD.t1439 a_1844_12699.t6 a_5931_9909.t11 VDD.t1438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X582 VDD.t1694 a_1833_4076.t7 a_4150_5439.t4 VDD.t1693 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X583 VSS.t241 a_23926_11281.t7 a_28011_9265.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X584 a_n3804_10998.t8 B[2].t0 VDD.t512 VDD.t511 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X585 a_17347_12889.t2 a_14496_9997.t14 VDD.t2378 VDD.t2377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X586 a_21466_26701.t1 a_21202_27284.t6 VSS.t252 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X587 a_25869_4129.t3 a_25324_4822.t4 a_25751_4129.t5 VDD.t904 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X588 VDD.t1226 a_23926_11281.t8 a_23986_11307.t6 VDD.t1225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X589 a_13018_12829.t2 a_11292_9266.t5 a_12900_12829.t2 VDD.t380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X590 VDD.t1829 opcode[0].t16 a_n3806_13067.t3 VDD.t1828 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X591 VDD.t1414 a_20900_24452.t10 a_22680_24452.t7 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X592 VDD.t2467 A[6].t5 a_15570_21782.t3 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X593 a_27008_18856.t0 A[4].t14 VDD.t1624 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X594 a_n3806_6861.t11 a_n3606_7699.t4 a_n3113_6918.t6 VDD.t1602 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X595 a_16205_19521.t0 a_n3113_2781.t9 VSS.t35 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X596 a_27439_12833.t4 a_26443_12246.t5 VDD.t171 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X597 a_29356_23724.t0 a_29650_24430.t4 VSS.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X598 VDD.t1384 a_30359_8848.t6 a_31893_9700.t2 VDD.t1383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X599 a_12382_21028.t0 a_12457_21658.t4 VSS.t13 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X600 a_27649_4129.t5 a_28061_4103.t5 a_27767_4129.t1 VDD.t1137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X601 a_6199_25133.t0 opcode[0].t17 a_5962_25770.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X602 VDD.t1718 a_19818_12178.t6 a_20814_12765.t3 VDD.t1717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X603 a_1227_7273.t5 A[5].t12 VDD.t2136 VDD.t2135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X604 a_25877_9997.t0 a_25332_10690.t4 a_25877_9265.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X605 VDD.t133 a_36751_16737.t9 Y[2].t2 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X606 a_19541_4102.t3 a_14306_12250.t5 VDD.t823 VDD.t822 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X607 a_10707_11307.t2 a_7749_6382.t7 VDD.t725 VDD.t724 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X608 a_9633_24460.t8 a_9206_25153.t4 a_9751_24460.t3 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X609 a_22680_24452.t4 a_22253_25145.t5 a_22798_24452.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X610 a_18952_19520.t5 a_19955_19546.t4 a_20495_18853.t4 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X611 VDD.t2088 B[5].t4 a_n3608_4192.t3 VDD.t2087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X612 VDD.t1942 a_n3115_713.t12 a_9012_21786.t2 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X613 a_36755_19987.t11 opcode[1].t20 VDD.t1507 VDD.t1506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X614 a_14490_4127.t3 a_13945_4820.t6 a_14490_3395.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X615 a_14366_23725.t1 a_14660_24431.t4 VSS.t202 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X616 a_27649_4129.t7 a_25869_4129.t9 VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X617 VDD.t2090 B[5].t5 a_n3808_4793.t2 VDD.t2089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X618 a_n3604_11836.t3 opcode[0].t18 VDD.t1831 VDD.t1830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X619 VDD.t964 a_19004_24158.t9 a_19594_23721.t2 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X620 a_12418_19515.t0 a_n3113_2781.t10 a_14315_18116.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X621 a_24562_12520.t0 a_23972_12957.t8 VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X622 VDD.t1324 a_21746_1762.t9 a_23964_7089.t2 VDD.t1323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X623 a_14154_6963.t2 a_13158_6376.t4 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X624 VDD.t1833 opcode[0].t19 a_n3606_13905.t3 VDD.t1832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X625 a_36751_4115.t5 a_36697_5000.t4 a_36751_4233.t5 VDD.t1139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X626 a_36701_20754.t2 opcode[1].t21 VDD.t1509 VDD.t1508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X627 a_36751_13593.t3 a_36697_14478.t5 a_38084_14302.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X628 VDD.t666 a_n3113_13124.t10 a_12461_27417.t6 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X629 VDD.t2184 a_7947_9909.t12 a_31464_14484.t3 VDD.t2183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X630 a_5962_25770.t5 opcode[0].t20 VDD.t1834 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X631 a_32247_1125.t1 a_30434_1013.t8 a_32011_1857.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X632 a_19483_3396.t0 a_15097_1774.t8 a_19247_4128.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X633 a_26113_9265.t1 a_20955_6381.t6 a_25877_9997.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X634 VSS.t115 a_24554_6652.t4 a_26171_6961.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X635 VDD.t2404 a_n3111_15192.t12 a_7735_24460.t0 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X636 a_16146_24457.t0 a_14366_24457.t9 VDD.t37 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X637 a_21027_4128.t0 a_20600_4821.t5 a_21145_4128.t1 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X638 a_31893_9700.t8 a_32305_9674.t4 a_32011_9700.t4 VDD.t948 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X639 VSS.t412 a_14496_9997.t15 a_17584_12252.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X640 a_14160_12833.t5 a_11297_10870.t4 a_14042_12833.t3 VDD.t531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X641 VSS.t145 B[1].t2 a_n3606_12466.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X642 a_11283_12520.t0 a_10693_12957.t7 VSS.t357 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X643 a_11291_5000.t0 a_10701_5437.t8 VSS.t80 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X644 a_4098_11193.t0 a_33377_10390.t7 VSS.t421 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X645 a_33377_10390.t1 a_30430_6928.t8 VDD.t2462 VDD.t2461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X646 VDD.t386 a_21711_14619.t6 a_23972_12957.t3 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X647 a_25869_4129.t6 a_26163_4103.t5 a_25751_4129.t3 VDD.t1288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X648 a_6538_26983.t0 a_5948_27420.t7 VSS.t132 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X649 a_36755_23131.t11 opcode[1].t22 VDD.t1511 VDD.t1510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X650 VDD.t2380 a_14496_9997.t16 a_17347_12889.t1 VDD.t2379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X651 a_23986_11307.t5 a_23926_11281.t9 VDD.t1228 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X652 a_6185_26783.t1 A[0].t3 a_5948_27420.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X653 VDD.t1405 a_n3113_6918.t13 a_27008_18856.t8 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X654 a_15556_20132.t3 a_11521_19244.t10 a_16205_19521.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X655 VDD.t1726 a_17296_5412.t8 a_17351_3834.t4 VDD.t1725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X656 a_7947_9909.t4 a_7402_10602.t5 a_7829_9909.t6 VDD.t765 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X657 a_10693_12957.t5 a_7749_6382.t8 VDD.t727 VDD.t726 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X658 a_7821_4129.t8 a_8233_4103.t5 a_7939_4129.t6 VDD.t521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X659 a_31893_9700.t1 a_30359_8848.t7 VDD.t1386 VDD.t1385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X660 VDD.t1230 a_23926_11281.t10 a_23981_9703.t6 VDD.t1229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X661 a_n3604_11836.t0 opcode[0].t21 VSS.t328 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X662 VSS.t180 a_12811_21658.t5 a_12382_21028.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X663 VSS.t414 a_n3111_15192.t13 a_6199_25133.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X664 a_5859_18120.t1 a_4963_19248.t13 VSS.t274 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X665 a_n3115_4850.t7 a_n3608_5631.t4 a_n3808_4793.t11 VDD.t946 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X666 a_9751_24460.t4 a_9206_25153.t5 a_9633_24460.t7 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X667 a_n3806_2724.t3 opcode[0].t22 VDD.t1836 VDD.t1835 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X668 VDD.t729 a_7749_6382.t9 a_10707_11307.t1 VDD.t728 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X669 a_14467_15035.t1 B[5].t6 VDD.t2092 VDD.t2091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X670 VDD.t1369 a_n3115_4850.t9 a_20495_18853.t7 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X671 a_22798_24452.t1 a_22253_25145.t6 a_22680_24452.t5 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X672 a_20495_18853.t3 a_19955_19546.t5 a_18952_19520.t4 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X673 a_27767_4129.t4 a_27222_4822.t5 a_27767_3397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X674 VDD.t2572 a_21150_9929.t11 a_32305_6179.t3 VDD.t2571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X675 a_24571_9266.t0 a_23981_9703.t8 VSS.t71 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X676 a_7821_4129.t11 a_6041_4129.t9 VDD.t2295 VDD.t2294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X677 a_14079_18116.t0 a_14373_18822.t4 a_12418_19515.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X678 a_n3608_5631.t1 opcode[0].t23 VDD.t1838 VDD.t1837 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X679 VDD.t340 a_26179_12829.t6 a_26443_12246.t3 VDD.t339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X680 a_5860_19519.t7 a_n3115_713.t13 a_7757_18120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X681 a_27431_6965.t0 a_26435_6378.t4 VDD.t286 VDD.t285 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X682 VDD.t1696 a_1833_4076.t8 a_4136_7089.t5 VDD.t1695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X683 VSS.t125 a_4090_5413.t7 a_4382_3198.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X684 VDD.t1211 a_30427_3858.t6 a_31466_6898.t3 VDD.t1210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X685 a_19818_12178.t2 a_19554_12761.t6 VDD.t1754 VDD.t1753 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X686 a_12461_27417.t5 a_n3113_13124.t11 VDD.t667 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X687 a_5957_24166.t1 opcode[0].t24 VDD.t1839 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X688 a_31464_14484.t2 a_7947_9909.t13 VDD.t2186 VDD.t2185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X689 VDD.t2405 a_n3111_15192.t14 a_5962_25770.t2 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X690 VDD.t526 a_21711_14619.t7 a_25759_9997.t5 VDD.t525 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X691 a_13599_21654.t2 a_15570_21782.t8 VDD.t2443 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X692 a_18702_4821.t3 a_15097_1774.t9 VDD.t2211 VDD.t2210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X693 a_32011_6205.t2 a_32305_6179.t5 a_31893_6205.t3 VDD.t229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X694 VDD.t1040 a_7939_4129.t12 a_10696_3833.t3 VDD.t1039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X695 VDD.t1684 a_17356_5438.t7 a_17946_5001.t3 VDD.t1683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X696 VSS.t365 B[5].t7 a_n3608_4192.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X697 VSS.t200 a_4726_6652.t5 a_6343_6961.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X698 a_20809_6964.t1 a_17946_5001.t4 a_20691_6964.t1 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X699 a_11292_9266.t2 a_10702_9703.t8 VDD.t1051 VDD.t1050 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X700 VDD.t2509 A[3].t6 a_29844_1450.t2 VDD.t2508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X701 Y[6].t2 a_36751_4115.t10 VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X702 a_19813_6377.t0 a_19549_6960.t5 VDD.t1081 VDD.t1080 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X703 a_32305_6179.t2 a_21150_9929.t12 VDD.t2580 VDD.t2579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X704 VDD.t2297 a_6041_4129.t10 a_7821_4129.t10 VDD.t2296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X705 VDD.t1441 a_1844_12699.t7 a_6343_9883.t2 VDD.t1440 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X706 a_9297_27296.t1 a_6552_25333.t4 VSS.t392 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X707 a_6041_4129.t0 a_6335_4103.t5 a_5923_4129.t1 VDD.t787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X708 a_23918_5413.t0 a_33377_6895.t7 VDD.t1093 VDD.t1092 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X709 VSS.t130 a_36755_19869.t8 Y[1].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X710 VDD.t225 B[2].t1 a_n3604_10397.t0 VDD.t224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X711 a_7493_12745.t1 a_4748_10782.t5 VSS.t153 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X712 a_17937_12452.t2 a_17347_12889.t8 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X713 VDD.t549 B[6].t5 a_21121_15056.t6 VDD.t548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X714 a_27458_24456.t0 a_26913_25149.t4 a_27458_23724.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X715 a_14784_4101.t3 a_10641_5411.t8 VDD.t2424 VDD.t2423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X716 VDD.t1763 a_20955_6381.t7 a_23986_11307.t2 VDD.t1762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X717 a_1833_4076.t2 a_1243_4513.t8 VDD.t858 VDD.t857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X718 a_7918_15036.t6 B[4].t4 VDD.t1986 VDD.t1985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X719 a_n3113_8987.t5 a_n3606_8329.t5 a_n3806_8930.t2 VDD.t1134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X720 VDD.t2068 a_1246_10551.t8 a_1836_10114.t2 VDD.t2067 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X721 VSS.t415 a_n3111_15192.t15 a_6185_26783.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X722 a_6253_21662.t2 a_8998_20136.t8 VDD.t1432 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X723 a_27008_18856.t7 a_n3113_6918.t14 VDD.t1406 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X724 a_6049_9909.t6 a_5504_10602.t5 a_6049_9177.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X725 VDD.t731 a_7749_6382.t10 a_10693_12957.t6 VDD.t730 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X726 a_18995_27412.t2 a_n3111_11055.t14 VDD.t573 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X727 VDD.t684 a_8543_1769.t8 a_10701_5437.t4 VDD.t683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X728 a_13961_18848.t6 a_14373_18822.t5 a_12418_19515.t2 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X729 a_13945_4820.t3 a_12592_4127.t10 VDD.t2331 VDD.t2330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X730 a_30430_6928.t1 a_29840_7365.t8 VDD.t398 VDD.t397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X731 a_23926_11281.t0 a_27313_6965.t5 VSS.t223 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X732 a_19051_21689.t5 a_18991_21663.t5 VDD.t2413 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X733 VDD.t2137 A[5].t13 a_22095_18533.t4 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X734 a_n3606_9768.t1 opcode[0].t25 VDD.t1841 VDD.t1840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X735 a_11297_10870.t3 a_10707_11307.t7 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X736 VDD.t2094 B[5].t8 a_14467_15035.t0 VDD.t2093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X737 VDD.t157 a_19585_26975.t4 a_21320_27284.t5 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X738 Y[1].t3 a_36755_19869.t9 VDD.t628 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X739 a_26443_12246.t2 a_26179_12829.t7 VDD.t342 VDD.t341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X740 a_7521_18120.t1 a_7815_18826.t4 a_5860_19519.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X741 VDD.t1843 opcode[0].t26 a_n3808_656.t9 VDD.t1842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X742 a_7493_12745.t3 a_4748_10782.t6 a_7611_12745.t3 VDD.t762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X743 a_7403_18852.t10 a_6863_19545.t5 a_5860_19519.t5 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X744 VDD.t1756 a_19554_12761.t7 a_19818_12178.t1 VDD.t1755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X745 VDD.t668 a_n3113_13124.t12 a_12461_27417.t4 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X746 VDD.t1844 opcode[0].t27 a_5957_24166.t0 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X747 a_36751_13711.t10 opcode[1].t23 VDD.t1513 VDD.t1512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X748 a_5962_25770.t1 a_n3111_15192.t16 VDD.t2406 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X749 a_25759_9997.t3 a_21711_14619.t8 VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X750 a_6049_9177.t0 a_6343_9883.t4 VSS.t206 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X751 a_4153_9615.t5 a_1844_12699.t8 VDD.t1443 VDD.t1442 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X752 VSS.t307 a_1836_10114.t12 a_4381_12232.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X753 VDD.t444 a_26571_21032.t6 a_25504_21666.t2 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X754 a_32009_13791.t6 a_31464_14484.t7 a_32009_13059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X755 a_36697_14478.t3 opcode[1].t24 VDD.t1515 VDD.t1514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X756 a_8175_3397.t1 a_6041_4129.t11 a_7939_4129.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X757 a_n2381_7154.t1 B[4].t5 VSS.t352 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X758 a_16558_24431.t3 a_9561_26713.t8 VDD.t885 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X759 a_27222_4822.t1 a_25869_4129.t10 VDD.t599 VDD.t598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X760 Y[0].t2 a_36755_23013.t10 VDD.t1935 VDD.t1934 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X761 a_32011_6205.t3 a_31466_6898.t5 a_32011_5473.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X762 a_21393_1762.t0 B[6].t6 a_21156_1325.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X763 VDD.t582 a_6607_6378.t5 a_7603_6965.t2 VDD.t581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X764 VSS.t404 a_8419_26709.t6 a_9297_27296.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X765 a_n3804_15135.t7 B[0].t2 VDD.t1159 VDD.t1158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X766 a_25110_18856.t6 a_24568_19252.t9 VDD.t914 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X767 a_17296_5412.t2 a_20696_12765.t5 VSS.t79 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X768 VDD.t2468 A[6].t6 a_13421_19541.t3 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X769 VSS.t222 a_19813_6377.t5 a_20691_6964.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X770 a_21121_15056.t5 B[6].t7 VDD.t551 VDD.t550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X771 a_23092_24426.t3 a_16074_26710.t7 VDD.t1917 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X772 a_27694_23724.t1 a_n3113_8987.t10 a_27458_24456.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X773 VDD.t1517 opcode[1].t25 a_36701_11276.t2 VDD.t1516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X774 a_1836_10114.t1 a_1246_10551.t9 VDD.t2070 VDD.t2069 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X775 VDD.t1431 a_8998_20136.t9 a_6253_21662.t1 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X776 a_19252_9929.t4 a_18707_10622.t5 a_19252_9197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X777 VSS.t149 a_7749_6382.t11 a_10930_12320.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X778 a_6041_4129.t3 a_5496_4822.t4 a_6041_3397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X779 VDD.t2313 a_11277_6650.t5 a_13012_6959.t2 VDD.t2312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X780 a_32305_9674.t3 a_30359_8848.t8 VDD.t1388 VDD.t1387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X781 VDD.t925 a_4098_11193.t10 a_4153_9615.t1 VDD.t924 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X782 a_11283_12520.t3 a_10693_12957.t8 VDD.t2020 VDD.t2019 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X783 VDD.t574 a_n3111_11055.t15 a_18995_27412.t1 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X784 VDD.t2510 A[3].t7 a_25553_27416.t3 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X785 a_8155_27292.t2 a_6547_23729.t4 VSS.t42 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X786 a_21746_1762.t0 a_21156_1325.t8 VSS.t283 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X787 a_9415_27296.t3 a_6552_25333.t5 a_9297_27296.t4 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X788 a_29238_24456.t9 a_27458_24456.t10 VDD.t1016 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X789 VDD.t379 a_10707_11307.t8 a_11297_10870.t2 VDD.t378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X790 a_13018_12829.t1 a_11292_9266.t6 a_12900_12829.t3 VDD.t983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X791 a_31891_13791.t10 a_30359_11881.t7 VDD.t1963 VDD.t1962 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X792 VDD.t9 a_20691_6964.t6 a_20955_6381.t0 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X793 a_14373_18822.t3 a_n3113_2781.t11 VDD.t567 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X794 a_18715_18853.t3 a_18952_19520.t10 a_18951_18121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X795 a_n3604_15973.t0 opcode[0].t28 VDD.t1846 VDD.t1845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X796 a_21320_27284.t4 a_19585_26975.t5 VDD.t41 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X797 a_31893_6205.t11 a_30427_3858.t7 VDD.t1213 VDD.t1212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X798 a_27775_9997.t5 a_28069_9971.t4 a_27657_9997.t11 VDD.t1186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X799 VDD.t419 a_10647_11281.t7 a_14378_9997.t4 VDD.t418 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X800 VDD.t1430 a_4963_19248.t14 a_4965_19545.t1 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X801 a_13659_21680.t5 a_13599_21654.t4 VDD.t1653 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X802 VDD.t825 a_14306_12250.t6 a_19129_4128.t11 VDD.t824 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X803 VSS.t399 a_6966_21028.t6 a_5899_21662.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X804 a_14507_1337.t2 A[6].t7 VDD.t2470 VDD.t2469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X805 a_7611_12745.t2 a_4748_10782.t7 a_7493_12745.t2 VDD.t763 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X806 a_5860_19519.t6 a_6863_19545.t6 a_7403_18852.t9 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X807 a_21444_9903.t3 a_17301_11213.t8 VDD.t2527 VDD.t2526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X808 VDD.t1326 a_21746_1762.t10 a_25324_4822.t2 VDD.t1325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X809 VDD.t2407 a_n3111_15192.t17 a_5962_25770.t0 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X810 VDD.t998 a_21711_14619.t9 a_25759_9997.t11 VDD.t997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X811 a_14372_4127.t10 a_12592_4127.t11 VDD.t2333 VDD.t2332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X812 a_17356_9635.t2 a_15057_14598.t6 VDD.t354 VDD.t353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X813 VDD.t1744 a_32009_13791.t8 a_36751_16855.t4 VDD.t1743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X814 a_1246_10551.t6 B[3].t2 VDD.t1469 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X815 a_18055_19249.t0 a_25429_21036.t5 VDD.t14 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X816 a_14248_24457.t3 a_n3113_13124.t13 VDD.t669 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X817 VDD.t2322 a_10687_7087.t8 a_11277_6650.t2 VDD.t2321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X818 VSS.t437 a_30430_6928.t9 a_31466_10393.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X819 a_32245_13059.t1 a_7947_9909.t14 a_32009_13791.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X820 a_12886_4101.t1 a_7939_4129.t13 VSS.t210 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X821 a_8147_24434.t3 A[0].t4 VDD.t1096 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X822 VDD.t799 B[3].t3 a_n3606_8329.t3 VDD.t798 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X823 a_10641_5411.t1 a_33375_14481.t8 VDD.t1181 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X824 a_4748_10782.t1 a_4158_11219.t8 VDD.t1024 VDD.t1023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X825 VDD.t1988 B[4].t6 a_n3606_6260.t2 VDD.t1987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X826 VDD.t2382 a_14496_9997.t17 a_18707_10622.t3 VDD.t2381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X827 VDD.t2472 A[6].t8 a_14507_1337.t1 VDD.t2471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X828 VDD.t1990 B[4].t7 a_n3806_6861.t7 VDD.t1989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X829 a_13421_19541.t2 A[6].t9 VDD.t2473 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X830 a_5824_21032.t2 a_6253_21662.t6 a_5959_21688.t5 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X831 a_22753_21176.t0 a_n3115_4850.t10 VSS.t262 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X832 VDD.t124 B[6].t8 a_21121_15056.t4 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X833 VDD.t1918 a_16074_26710.t8 a_23092_24426.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X834 a_16146_24457.t9 a_16558_24431.t4 a_16264_24457.t5 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X835 VSS.t429 A[3].t8 a_27694_23724.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X836 a_4145_3835.t5 a_1817_6836.t8 VDD.t1349 VDD.t1348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X837 a_32247_8968.t1 a_30430_6928.t10 a_32011_9700.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X838 a_1227_7273.t1 B[4].t8 VDD.t1992 VDD.t1991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X839 a_36755_23131.t1 a_9751_24460.t11 a_36755_23013.t6 VDD.t969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X840 a_36751_1089.t0 a_36697_1856.t4 a_36751_971.t0 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X841 a_8998_20136.t4 a_n3115_713.t14 VDD.t1943 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X842 a_23092_24426.t0 a_16074_26710.t9 VSS.t340 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X843 VDD.t901 a_30364_14452.t5 a_36755_23131.t7 VDD.t900 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X844 VSS.t85 a_10647_11281.t8 a_14732_9265.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X845 VSS.t425 A[6].t10 a_1480_3876.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X846 a_25759_9997.t9 a_26171_9971.t5 a_25877_9997.t6 VDD.t973 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X847 a_n3804_10998.t9 a_n3604_11836.t5 a_n3111_11055.t5 VDD.t608 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X848 a_19585_26975.t3 a_18995_27412.t8 VDD.t48 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X849 a_12480_9997.t1 a_12892_9971.t5 a_12598_9997.t1 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X850 VSS.t43 a_6538_26983.t4 a_8155_27292.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X851 a_20900_24452.t5 a_20355_25145.t5 a_20782_24452.t11 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X852 a_9297_27296.t3 a_6552_25333.t6 a_9415_27296.t4 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X853 a_n3806_2724.t11 a_n3606_2123.t5 a_n3113_2781.t7 VDD.t1004 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X854 a_23986_11307.t4 a_23926_11281.t11 VDD.t1232 VDD.t1231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X855 a_11297_10870.t1 a_10707_11307.t9 VDD.t435 VDD.t434 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X856 VDD.t1965 a_30359_11881.t8 a_31891_13791.t11 VDD.t1964 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X857 a_n3608_1494.t0 opcode[0].t29 VSS.t329 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X858 VDD.t884 a_6538_26983.t5 a_8273_27292.t2 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X859 a_18715_18121.t0 a_19009_18827.t4 a_18715_18853.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X860 VDD.t1351 a_1817_6836.t9 a_6335_4103.t2 VDD.t1350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X861 a_17296_5412.t0 a_20696_12765.t6 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X862 VDD.t375 a_19585_26975.t6 a_21320_27284.t3 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X863 a_4158_11219.t0 a_4098_11193.t11 VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X864 a_19247_3396.t0 a_19541_4102.t6 VSS.t9 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X865 a_n3804_15135.t3 a_n3604_14534.t4 a_n3111_15192.t0 VDD.t942 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X866 a_15097_1774.t2 a_14507_1337.t9 VDD.t2229 VDD.t2228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X867 a_25877_9265.t0 a_26171_9971.t6 VSS.t77 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X868 a_36751_1089.t7 a_5623_18852.t9 a_36751_971.t3 VDD.t634 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X869 a_36697_1856.t2 opcode[1].t26 VDD.t1519 VDD.t1518 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X870 VDD.t1698 a_1833_4076.t9 a_5496_4822.t2 VDD.t1697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X871 VDD.t523 a_27585_12250.t4 a_36751_1089.t5 VDD.t522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X872 a_7953_1332.t5 A[4].t15 VDD.t1626 VDD.t1625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X873 VDD.t1794 a_1227_7273.t8 a_1817_6836.t2 VDD.t1793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X874 a_21027_4128.t10 a_21439_4102.t5 a_21145_4128.t6 VDD.t745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X875 VDD.t460 a_25429_21036.t6 a_18055_19249.t1 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X876 VDD.t371 a_23964_7089.t8 a_24554_6652.t3 VDD.t370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X877 VDD.t670 a_n3113_13124.t14 a_14248_24457.t4 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X878 a_29769_9285.t6 B[3].t4 VDD.t1359 VDD.t1358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X879 a_26163_4103.t0 a_21145_4128.t11 VSS.t293 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X880 a_8508_14599.t1 a_7918_15036.t7 VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X881 VDD.t239 a_14932_26706.t6 a_15928_27293.t2 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X882 a_13060_23726.t0 a_12470_24163.t10 VSS.t384 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X883 a_32011_1125.t0 a_32305_1831.t5 VSS.t62 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X884 a_21150_9929.t2 a_20605_10622.t4 a_21032_9929.t4 VDD.t207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X885 a_n3806_13067.t2 opcode[0].t30 VDD.t1848 VDD.t1847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X886 VDD.t2583 a_11521_19244.t11 a_15556_20132.t5 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X887 VDD.t1183 a_33375_14481.t9 a_10641_5411.t2 VDD.t1182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X888 VDD.t2096 B[5].t9 a_29769_12318.t4 VDD.t2095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X889 a_10702_9703.t3 a_8508_14599.t8 VDD.t2046 VDD.t2045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X890 a_18707_10622.t2 a_14496_9997.t18 VDD.t2384 VDD.t2383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X891 a_12828_3395.t1 a_8543_1769.t9 a_12592_4127.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X892 VDD.t1328 a_21746_1762.t11 a_25751_4129.t7 VDD.t1327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X893 VSS.t26 B[6].t9 a_n3606_2123.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X894 a_16264_24457.t6 a_16558_24431.t5 a_16146_24457.t10 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X895 a_27458_23724.t1 a_27752_24430.t5 VSS.t232 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X896 a_n3608_4192.t2 B[5].t10 VDD.t2098 VDD.t2097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X897 a_36751_13711.t0 a_29356_24456.t8 a_36751_13593.t2 VDD.t844 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X898 VDD.t1944 a_n3115_713.t15 a_8998_20136.t5 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X899 a_36751_4233.t2 a_12181_18848.t9 a_36751_4115.t2 VDD.t2347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X900 a_n3808_4793.t1 B[5].t11 VDD.t2100 VDD.t2099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X901 a_23972_12957.t2 a_21711_14619.t10 VDD.t384 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X902 a_7101_21684.t2 a_7395_21658.t5 a_6966_21028.t2 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X903 VDD.t213 a_18995_27412.t9 a_19585_26975.t2 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X904 a_7735_24460.t9 a_7308_25153.t5 a_7853_24460.t2 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X905 a_1844_12699.t2 a_1254_13136.t9 VDD.t211 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X906 a_21032_9929.t6 a_21444_9903.t5 a_21150_9929.t6 VDD.t1381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X907 a_4144_12869.t4 a_1844_12699.t9 VDD.t1445 VDD.t1444 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X908 a_38084_14538.t0 opcode[1].t27 a_36751_13593.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X909 a_32303_13765.t1 a_30359_11881.t9 VDD.t1967 VDD.t1966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X910 a_9415_27296.t5 a_6552_25333.t7 a_9297_27296.t2 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X911 a_26152_23725.t1 a_25562_24162.t8 VSS.t84 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X912 a_n3808_656.t6 B[7].t2 VDD.t1273 VDD.t1272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X913 a_7918_15036.t5 B[4].t9 VDD.t1994 VDD.t1993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X914 VDD.t2318 a_15556_20132.t8 a_12811_21658.t3 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X915 VDD.t1234 a_23926_11281.t12 a_23981_9703.t5 VDD.t1233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X916 VDD.t1850 opcode[0].t31 a_n3808_4793.t8 VDD.t1849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X917 a_12517_21684.t0 a_12457_21658.t5 VDD.t235 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X918 VSS.t72 a_5824_21032.t5 Cout.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X919 a_1833_4076.t3 a_1243_4513.t9 VSS.t168 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X920 a_27767_3397.t0 a_28061_4103.t6 VSS.t226 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X921 a_20495_18853.t6 a_n3115_4850.t11 VDD.t1370 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X922 a_9652_17921.t1 a_4963_19248.t15 VSS.t273 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X923 VDD.t1221 a_4136_7089.t8 a_4726_6652.t3 VDD.t1220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X924 a_18055_19249.t2 a_25429_21036.t7 VDD.t524 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X925 a_14378_9997.t10 a_12598_9997.t9 VDD.t1246 VDD.t1245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X926 VDD.t414 a_25562_24162.t9 a_26152_23725.t2 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X927 VDD.t1924 a_25465_19523.t10 a_25522_18830.t3 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X928 a_36755_23013.t0 a_36701_23898.t4 a_36755_23131.t4 VDD.t620 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X929 VSS.t426 A[6].t11 a_14744_1774.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X930 a_n3808_656.t3 a_n3608_1494.t5 a_n3115_713.t4 VDD.t782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X931 a_7829_9909.t1 a_8241_9883.t4 a_7947_9909.t0 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X932 a_36751_16855.t9 a_36697_17622.t4 a_36751_16737.t5 VDD.t1222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X933 a_29769_12318.t5 B[5].t12 VDD.t2102 VDD.t2101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X934 a_14366_24457.t3 a_13821_25150.t4 a_14248_24457.t6 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X935 VSS.t137 a_22104_21787.t10 a_20133_21659.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X936 a_19541_4102.t0 a_14306_12250.t7 VSS.t164 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X937 VDD.t1851 opcode[0].t32 a_9633_24460.t2 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X938 VDD.t365 a_29844_1450.t7 a_30434_1013.t3 VDD.t364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X939 VDD.t539 a_24554_6652.t5 a_26289_6961.t5 VDD.t538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X940 VSS.t430 A[3].t9 a_30081_813.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X941 a_13961_18848.t2 A[6].t12 VDD.t2474 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X942 VDD.t388 a_10701_5437.t9 a_11291_5000.t2 VDD.t387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X943 VSS.t150 a_7749_6382.t12 a_12053_10690.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X944 a_16146_24457.t11 a_16558_24431.t6 a_16264_24457.t7 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X945 a_12707_23526.t0 A[1].t7 a_12470_24163.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X946 VDD.t1597 a_13051_26980.t5 a_14786_27289.t1 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X947 a_12886_4101.t2 a_7939_4129.t14 VDD.t1042 VDD.t1041 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X948 a_4726_6652.t2 a_4136_7089.t9 VDD.t1200 VDD.t1199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X949 Y[3].t3 a_36751_13593.t8 VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X950 a_27340_24456.t8 a_n3113_8987.t11 VDD.t1796 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X951 a_33377_2547.t1 a_14490_4127.t12 VDD.t2150 VDD.t2149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X952 a_6966_21028.t1 a_7395_21658.t6 a_7101_21684.t1 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X953 a_36701_8132.t3 opcode[1].t28 VDD.t1521 VDD.t1520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X954 VSS.t38 a_19252_9929.t12 a_20605_10622.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X955 VSS.t86 a_10647_11281.t9 a_10939_9066.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X956 a_9633_24460.t11 a_10045_24434.t4 a_9751_24460.t1 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X957 VDD.t13 a_27767_4129.t8 a_36755_7365.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X958 VDD.t1853 opcode[0].t33 a_n3806_8930.t4 VDD.t1852 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X959 VDD.t2240 a_23918_5413.t7 a_28061_4103.t2 VDD.t2239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X960 VSS.t102 a_27585_12250.t5 a_38084_1916.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X961 VDD.t1996 B[4].t10 a_7918_15036.t4 VDD.t1995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X962 VSS.t294 a_21145_4128.t12 a_26105_3397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X963 VDD.t1120 a_19813_6377.t6 a_20809_6964.t4 VDD.t1119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X964 a_12811_21658.t2 a_15556_20132.t9 VDD.t2607 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X965 a_5923_4129.t8 a_1833_4076.t10 VDD.t1700 VDD.t1699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X966 VDD.t827 a_14306_12250.t8 a_17342_7088.t6 VDD.t826 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X967 a_30359_8848.t1 a_29769_9285.t8 VSS.t228 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X968 a_5623_18852.t2 a_4965_19545.t5 a_5505_18852.t2 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X969 a_27657_9997.t5 a_25877_9997.t10 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X970 a_27458_24456.t2 a_26913_25149.t5 a_27340_24456.t4 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X971 VDD.t959 a_36755_10391.t10 Y[4].t1 VDD.t958 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X972 a_32305_9674.t2 a_30359_8848.t9 VDD.t1390 VDD.t1389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X973 VDD.t614 a_12457_21658.t6 a_12517_21684.t2 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X974 a_26157_25329.t0 a_25567_25766.t10 VSS.t219 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X975 a_5824_21032.t0 a_5899_21662.t6 VSS.t402 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X976 a_17593_4801.t1 a_17296_5412.t9 a_17356_5438.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X977 a_19247_4128.t6 a_18702_4821.t4 a_19129_4128.t8 VDD.t544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X978 a_n3604_15973.t1 opcode[0].t34 VSS.t330 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X979 VSS.t120 a_n3111_11055.t16 a_20355_25145.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X980 a_29238_24456.t7 a_28811_25149.t5 a_29356_24456.t5 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X981 VDD.t994 a_30434_1013.t9 a_33377_2547.t6 VDD.t993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X982 a_31891_13791.t2 a_32303_13765.t4 a_32009_13791.t2 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X983 a_21466_26701.t2 a_21202_27284.t7 VDD.t1299 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X984 a_26152_23725.t3 a_25562_24162.t10 VDD.t415 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X985 a_25522_18830.t2 a_25465_19523.t11 VDD.t1925 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X986 VDD.t421 a_10647_11281.t10 a_14378_9997.t5 VDD.t420 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X987 VDD.t686 a_8543_1769.t10 a_12047_4820.t2 VDD.t685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X988 VDD.t1415 a_20900_24452.t11 a_22253_25145.t3 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X989 a_12475_18822.t3 a_12418_19515.t11 VSS.t135 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X990 a_23973_3835.t2 a_23918_5413.t8 VDD.t2242 VDD.t2241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X991 a_14248_24457.t10 a_13821_25150.t5 a_14366_24457.t2 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X992 VSS.t389 a_7853_24460.t10 a_9206_25153.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X993 VSS.t37 a_15057_14598.t7 a_19488_9197.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X994 a_9633_24460.t1 opcode[0].t35 VDD.t1854 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X995 VDD.t1061 a_23978_5439.t9 a_24568_5002.t2 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X996 VSS.t107 a_21150_9929.t13 a_32247_5473.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X997 VSS.t172 a_9561_26713.t9 a_12707_23526.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X998 a_21439_4102.t3 a_17296_5412.t10 VDD.t1728 VDD.t1727 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X999 a_26163_4103.t2 a_21145_4128.t13 VDD.t1579 VDD.t1578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1000 a_12063_18848.t6 a_12475_18822.t6 a_12181_18848.t5 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1001 a_4748_10782.t2 a_4158_11219.t9 VDD.t1026 VDD.t1025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1002 a_n3804_10998.t3 B[2].t2 VDD.t243 VDD.t242 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1003 VDD.t1628 A[4].t16 a_29837_4295.t3 VDD.t1627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1004 VDD.t257 a_17932_6651.t5 a_19667_6960.t1 VDD.t256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1005 a_n3804_15135.t1 a_n3604_15973.t6 a_n3111_15192.t6 VDD.t2078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1006 a_14378_9997.t8 a_13951_10690.t6 a_14496_9997.t4 VDD.t2352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1007 VDD.t1797 a_n3113_8987.t12 a_27340_24456.t7 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1008 a_9751_24460.t0 a_10045_24434.t5 a_9633_24460.t10 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1009 VSS.t255 a_24570_19549.t5 a_25228_18124.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1010 a_n3113_2781.t1 opcode[0].t36 a_n2381_3017.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1011 VDD.t180 a_19252_9929.t13 a_20605_10622.t3 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1012 VDD.t2408 a_n3111_15192.t18 a_5948_27420.t0 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1013 VSS.t259 a_1817_6836.t10 a_6277_3397.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1014 a_26143_26979.t2 a_25553_27416.t9 VSS.t174 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1015 VDD.t2602 a_15556_20132.t10 a_12811_21658.t1 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1016 VDD.t0 a_28024_26705.t4 a_29020_27292.t0 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1017 VDD.t2595 a_5860_19519.t11 a_5505_18852.t7 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1018 a_5505_18852.t1 a_4965_19545.t6 a_5623_18852.t1 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1019 a_n3808_656.t1 a_n3608_55.t6 a_n3115_713.t1 VDD.t1950 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1020 a_36755_10509.t11 a_25228_18856.t9 a_36755_10391.t7 VDD.t982 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1021 VDD.t952 a_25877_9997.t11 a_27657_9997.t4 VDD.t951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1022 a_17356_9635.t6 a_17301_11213.t9 VDD.t2529 VDD.t2528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1023 a_14372_4127.t1 a_10641_5411.t9 VDD.t2426 VDD.t2425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1024 VDD.t1392 a_30359_8848.t10 a_32305_9674.t1 VDD.t1391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1025 a_12517_21684.t1 a_12457_21658.t7 VDD.t613 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1026 VDD.t2557 a_32011_1857.t9 a_36751_13711.t4 VDD.t2556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1027 a_27362_18124.t0 A[4].t17 VSS.t300 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1028 VDD.t1730 a_17296_5412.t11 a_21439_4102.t2 VDD.t1729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1029 VDD.t312 a_32011_6205.t8 a_36755_10509.t2 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1030 VDD.t2409 a_n3111_15192.t19 a_7308_25153.t3 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1031 a_21444_9903.t0 a_17301_11213.t10 VSS.t435 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1032 VDD.t1856 opcode[0].t37 a_n3804_15135.t10 VDD.t1855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1033 a_29356_24456.t4 a_28811_25149.t6 a_29238_24456.t8 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1034 a_32009_13791.t1 a_32303_13765.t5 a_31891_13791.t1 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1035 VDD.t1300 a_21202_27284.t8 a_21466_26701.t3 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1036 VSS.t156 a_28617_21790.t7 a_26646_21662.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1037 VDD.t829 a_14306_12250.t9 a_19129_4128.t10 VDD.t828 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1038 a_14378_9997.t3 a_10647_11281.t11 VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1039 a_28603_20140.t5 a_24568_19252.t10 VDD.t915 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1040 a_8233_4103.t2 a_4090_5413.t8 VDD.t1065 VDD.t1064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1041 VDD.t2168 A[1].t8 a_12470_24163.t5 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1042 a_20613_18121.t1 a_20907_18827.t4 a_18952_19520.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1043 VDD.t875 a_19247_4128.t11 a_20600_4821.t2 VDD.t874 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1044 VDD.t1670 a_1836_10114.t13 a_5504_10602.t1 VDD.t1669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1045 a_36755_19869.t6 a_36701_20754.t5 a_38088_20578.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1046 a_4145_3835.t2 a_4090_5413.t9 VDD.t1067 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1047 VDD.t2586 a_11521_19244.t12 a_11523_19541.t2 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1048 VDD.t2428 a_10641_5411.t10 a_14372_4127.t0 VDD.t2427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1049 VDD.t2475 A[6].t13 a_15561_18528.t3 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1050 VDD.t1523 opcode[1].t29 a_36751_16855.t6 VDD.t1522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1051 a_14366_24457.t1 a_13821_25150.t6 a_14248_24457.t11 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1052 a_20487_21659.t2 a_22095_18533.t8 VDD.t690 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1053 VDD.t2307 a_4150_5439.t8 a_4740_5002.t2 VDD.t2306 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1054 VSS.t104 A[7].t2 a_6863_19545.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1055 a_30430_6928.t2 a_29840_7365.t9 VSS.t82 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1056 VDD.t1028 a_4158_11219.t10 a_4748_10782.t3 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1057 VDD.t2188 a_7947_9909.t15 a_33375_14481.t4 VDD.t2187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1058 a_30427_3858.t0 a_29837_4295.t7 VSS.t169 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1059 a_19667_6960.t4 a_17941_3397.t6 a_19549_6960.t3 VDD.t1034 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1060 a_27340_24456.t6 a_n3113_8987.t13 VDD.t1798 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1061 a_9633_24460.t9 a_10045_24434.t6 a_9751_24460.t2 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1062 VDD.t1044 a_7939_4129.t15 a_12474_4127.t6 VDD.t1043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1063 a_12598_9997.t4 a_12053_10690.t5 a_12598_9265.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1064 a_32011_8968.t1 a_32305_9674.t5 VSS.t184 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1065 a_8241_9883.t0 a_4098_11193.t12 VSS.t66 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1066 a_19541_4102.t2 a_14306_12250.t10 VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1067 a_8190_1769.t0 B[5].t13 a_7953_1332.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1068 a_31893_1857.t1 a_32305_1831.t6 a_32011_1857.t2 VDD.t284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1069 VSS.t279 a_8998_20136.t10 a_6253_21662.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1070 a_20605_10622.t2 a_19252_9929.t14 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1071 a_6538_26983.t3 a_5948_27420.t8 VDD.t639 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1072 a_32011_9700.t1 a_31466_10393.t5 a_31893_9700.t4 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1073 a_4740_5002.t1 a_4150_5439.t9 VDD.t2309 VDD.t2308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1074 a_29020_27292.t1 a_28024_26705.t5 VDD.t1 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1075 a_36755_23013.t1 a_36701_23898.t5 a_38088_23722.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1076 a_25465_19523.t7 a_n3113_6918.t15 a_27362_18124.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1077 VDD.t1919 a_16074_26710.t10 a_22680_24452.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1078 a_10924_6450.t0 a_7939_4129.t16 a_10687_7087.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1079 a_7308_25153.t2 a_n3111_15192.t20 VDD.t2410 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1080 a_25465_19523.t0 a_26468_19549.t5 a_27008_18856.t5 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1081 VDD.t671 a_n3113_13124.t15 a_12475_25767.t3 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1082 a_8543_1769.t0 a_7953_1332.t7 VSS.t356 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1083 a_12474_4127.t7 a_7939_4129.t17 VDD.t1046 VDD.t1045 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1084 a_29238_24456.t0 a_29650_24430.t5 a_29356_24456.t0 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1085 VDD.t776 a_28617_21790.t8 a_26646_21662.t3 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1086 VDD.t1732 a_17296_5412.t12 a_17356_5438.t4 VDD.t1731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1087 VDD.t197 a_10647_11281.t12 a_14790_9971.t2 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1088 VDD.t2512 A[3].t10 a_29774_14889.t2 VDD.t2511 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1089 a_10702_9703.t2 a_8508_14599.t9 VDD.t2048 VDD.t2047 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1090 VDD.t916 a_24568_19252.t11 a_28603_20140.t4 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1091 a_12470_24163.t6 A[1].t9 VDD.t2169 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1092 a_8543_1769.t3 a_7953_1332.t8 VDD.t2014 VDD.t2013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1093 VDD.t2264 a_7853_24460.t11 a_9206_25153.t1 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1094 VDD.t2244 a_23918_5413.t9 a_27649_4129.t10 VDD.t2243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1095 VDD.t1525 opcode[1].t30 a_36751_1089.t10 VDD.t1524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1096 a_36755_7365.t4 a_18715_18853.t9 a_36755_7247.t1 VDD.t508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1097 a_12063_18848.t11 a_11521_19244.t13 VDD.t2587 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1098 VDD.t529 a_21711_14619.t11 a_26171_9971.t2 VDD.t528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1099 a_11297_10870.t0 a_10707_11307.t10 VSS.t8 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1100 a_15561_18528.t2 A[6].t14 VDD.t2476 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1101 a_4136_7089.t2 a_1817_6836.t11 VDD.t1353 VDD.t1352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1102 a_14248_24457.t7 a_14660_24431.t5 a_14366_24457.t6 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1103 a_33377_6895.t2 a_21150_9929.t14 VDD.t2578 VDD.t2577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1104 a_n3111_11055.t1 a_n3604_10397.t6 a_n3804_10998.t1 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1105 VDD.t691 a_22095_18533.t9 a_20487_21659.t1 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1106 VSS.t431 A[3].t11 a_30077_6728.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1107 VDD.t1650 a_4144_12869.t9 a_4734_12432.t2 VDD.t1649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1108 a_12457_21658.t3 a_13524_21024.t5 VDD.t534 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1109 a_1243_4513.t5 B[3].t5 VDD.t1465 VDD.t1464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1110 a_29769_9285.t2 A[4].t18 VDD.t1630 VDD.t1629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1111 VDD.t91 a_14036_6963.t6 a_10647_11281.t2 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1112 VDD.t330 a_23981_9703.t9 a_24571_9266.t2 VDD.t329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1113 a_n3111_15192.t1 a_n3604_14534.t5 a_n3804_15135.t4 VDD.t943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1114 a_n3113_8987.t6 a_n3606_8329.t6 a_n3806_8930.t1 VDD.t1135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1115 a_20900_23720.t0 a_21194_24426.t4 VSS.t101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1116 a_9661_21175.t0 a_n3115_713.t16 VSS.t344 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1117 a_11292_9266.t0 a_10702_9703.t9 VSS.t211 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1118 a_36755_10509.t8 a_36701_11276.t5 a_36755_10391.t4 VDD.t883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1119 VSS.t21 a_26443_12246.t6 a_27321_12833.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1120 a_12712_25130.t1 a_9561_26713.t10 a_12475_25767.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1121 VDD.t202 a_28024_26705.t6 a_29020_27292.t2 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1122 VDD.t708 B[1].t3 a_n3806_13067.t8 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1123 a_22680_24452.t1 a_16074_26710.t11 VDD.t1920 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1124 a_36755_19869.t4 a_36701_20754.t6 a_36755_19987.t4 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1125 a_27008_18856.t4 a_26468_19549.t6 a_25465_19523.t1 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1126 VDD.t2478 A[6].t15 a_1243_4513.t1 VDD.t2477 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1127 VDD.t733 a_7749_6382.t13 a_12480_9997.t10 VDD.t732 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1128 a_12475_25767.t4 a_n3113_13124.t16 VDD.t672 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1129 a_17941_3397.t2 a_17351_3834.t8 VDD.t1032 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1130 a_7829_9909.t2 a_8241_9883.t5 a_7947_9909.t1 VDD.t307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1131 VDD.t317 a_9297_27296.t5 a_9561_26713.t1 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1132 VDD.t2514 A[3].t12 a_29840_7365.t1 VDD.t2513 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1133 a_26646_21662.t2 a_28617_21790.t9 VDD.t777 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1134 a_14790_9971.t1 a_10647_11281.t13 VDD.t199 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1135 VDD.t1361 a_7493_12745.t5 a_4090_5413.t3 VDD.t1360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1136 a_29774_14889.t1 A[3].t13 VDD.t2516 VDD.t2515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1137 VDD.t886 a_9561_26713.t11 a_12470_24163.t1 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1138 VSS.t382 a_15097_1774.t10 a_18702_4821.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1139 VDD.t406 a_15057_14598.t8 a_19134_9929.t4 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1140 VDD.t1069 a_4090_5413.t10 a_7821_4129.t7 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1141 a_5931_9909.t7 a_5504_10602.t6 a_6049_9909.t7 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1142 VDD.t2588 a_11521_19244.t14 a_12063_18848.t10 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1143 VSS.t30 a_9003_18532.t9 a_7395_21658.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1144 a_26171_9971.t1 a_21711_14619.t12 VDD.t217 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1145 a_36751_4233.t10 a_27775_9997.t9 VDD.t1242 VDD.t1241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1146 a_22104_21787.t2 a_n3115_4850.t12 VDD.t1371 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1147 VSS.t239 a_36751_971.t9 Y[7].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1148 a_25522_18830.t1 a_25465_19523.t12 VDD.t1926 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1149 a_36755_19869.t2 a_16264_24457.t9 a_36755_19987.t2 VDD.t1605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1150 VSS.t151 a_7749_6382.t14 a_10944_10670.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1151 VDD.t359 a_13524_21024.t6 a_12457_21658.t2 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1152 VDD.t1124 a_27313_6965.t6 a_23926_11281.t1 VDD.t1123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1153 a_11286_3396.t2 a_10696_3833.t8 VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1154 VDD.t1122 a_19813_6377.t7 a_20809_6964.t3 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1155 VDD.t1527 opcode[1].t31 a_36697_14478.t2 VDD.t1526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1156 a_13051_26980.t2 a_12461_27417.t7 VSS.t55 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1157 a_27752_24430.t2 A[3].t14 VDD.t2517 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1158 VDD.t975 a_9003_18532.t10 a_7395_21658.t2 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1159 a_27313_6965.t2 a_24568_5002.t5 VSS.t213 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1160 VDD.t2213 a_15097_1774.t11 a_17342_7088.t1 VDD.t2212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1161 a_n3113_6918.t0 opcode[0].t38 a_n2381_7154.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1162 VDD.t2547 a_30430_6928.t11 a_31466_10393.t3 VDD.t2546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1163 a_25567_25766.t6 a_22608_26705.t6 VDD.t448 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1164 a_30427_3858.t3 a_29837_4295.t8 VDD.t865 VDD.t864 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1165 a_6049_9909.t2 a_6343_9883.t5 a_5931_9909.t5 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1166 VSS.t370 A[5].t14 a_1483_9914.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1167 a_27585_12250.t0 a_27321_12833.t5 VSS.t139 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1168 VSS.t141 a_n3113_13124.t17 a_12712_25130.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1169 a_14372_4127.t5 a_13945_4820.t7 a_14490_4127.t4 VDD.t881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1170 a_28069_9971.t0 a_23926_11281.t13 VSS.t242 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1171 a_n3608_55.t1 B[7].t3 VDD.t1275 VDD.t1274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1172 a_36755_23131.t10 opcode[1].t32 VDD.t1529 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1173 VDD.t1531 opcode[1].t33 a_36755_7365.t6 VDD.t1530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1174 VDD.t1921 a_16074_26710.t12 a_22680_24452.t0 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1175 VSS.t88 a_26571_21032.t7 a_25504_21666.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1176 a_n2381_13124.t0 a_n3606_13905.t5 a_n3113_13124.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1177 a_5923_4129.t11 a_1817_6836.t12 VDD.t1355 VDD.t1354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1178 a_12480_9997.t9 a_7749_6382.t15 VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1179 a_8155_14399.t1 B[4].t11 a_7918_15036.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1180 a_36751_16737.t4 a_36697_17622.t5 a_36751_16855.t10 VDD.t1223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1181 a_33614_6258.t0 a_21150_9929.t15 a_33377_6895.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1182 a_4153_9615.t4 a_1844_12699.t10 VDD.t1447 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1183 a_19247_4128.t2 a_18702_4821.t5 a_19129_4128.t3 VDD.t167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1184 VDD.t778 a_28617_21790.t10 a_26646_21662.t1 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1185 a_14660_24431.t0 A[1].t10 VSS.t374 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1186 a_17932_6651.t3 a_17342_7088.t7 VDD.t593 VDD.t592 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1187 VDD.t1104 a_7939_4129.t18 a_10687_7087.t5 VDD.t1103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1188 a_12470_24163.t2 a_9561_26713.t12 VDD.t887 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1189 a_n3115_4850.t0 a_n3608_4192.t7 a_n3808_4793.t3 VDD.t1054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1190 a_36755_7365.t10 a_36701_8132.t5 a_36755_7247.t5 VDD.t1087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1191 a_19134_9929.t3 a_15057_14598.t9 VDD.t272 VDD.t271 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1192 a_36755_19987.t1 a_16264_24457.t10 a_36755_19869.t1 VDD.t1606 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1193 a_10938_4800.t0 a_10641_5411.t11 a_10701_5437.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1194 a_19134_9929.t10 a_18707_10622.t6 a_19252_9929.t2 VDD.t1296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1195 a_26163_4103.t1 a_21145_4128.t14 VDD.t1581 VDD.t1580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1196 VDD.t1632 A[4].t19 a_1254_13136.t2 VDD.t1631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1197 VDD.t374 a_8155_27292.t5 a_8419_26709.t1 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1198 a_19813_6377.t1 a_19549_6960.t6 VSS.t215 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1199 VSS.t309 a_1833_4076.t11 a_4373_6452.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1200 VDD.t1372 a_n3115_4850.t13 a_22104_21787.t1 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1201 a_12457_21658.t1 a_13524_21024.t7 VDD.t129 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1202 a_25110_18856.t4 a_25522_18830.t6 a_25228_18856.t2 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1203 a_24563_3398.t3 a_23973_3835.t7 VDD.t889 VDD.t888 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1204 a_n3113_13124.t3 a_n3606_12466.t5 a_n3806_13067.t4 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1205 a_36751_16855.t3 a_32009_13791.t9 VDD.t1746 VDD.t1745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1206 a_38084_1680.t1 a_5623_18852.t10 VSS.t131 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1207 a_9003_18532.t6 a_4963_19248.t16 VDD.t1420 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1208 a_12592_4127.t5 a_12047_4820.t5 a_12474_4127.t10 VDD.t1152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1209 a_7485_6965.t2 a_4740_5002.t6 VSS.t395 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1210 a_26571_21032.t4 a_27000_21662.t5 a_26706_21688.t5 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1211 a_31466_10393.t2 a_30430_6928.t12 VDD.t2549 VDD.t2548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1212 VDD.t575 a_n3111_11055.t17 a_19009_25762.t0 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1213 VDD.t449 a_22608_26705.t7 a_25567_25766.t5 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1214 a_27752_24430.t0 A[3].t15 VSS.t432 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1215 VDD.t1858 opcode[0].t39 a_n3606_3562.t2 VDD.t1857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1216 a_13158_6376.t2 a_12894_6959.t6 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1217 a_25562_24162.t3 A[3].t16 VDD.t2518 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1218 a_27649_4129.t1 a_27222_4822.t6 a_27767_4129.t6 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1219 a_n2383_4850.t1 a_n3608_5631.t5 a_n3115_4850.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1220 VDD.t576 a_n3111_11055.t18 a_20782_24452.t1 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1221 a_12894_6959.t2 a_11286_3396.t6 VSS.t59 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1222 VDD.t1248 a_12598_9997.t10 a_13951_10690.t1 VDD.t1247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1223 VDD.t607 B[2].t3 a_n3604_10397.t3 VDD.t606 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1224 a_14507_1337.t4 B[5].t14 VDD.t2104 VDD.t2103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1225 VDD.t1860 opcode[0].t40 a_n3606_7699.t2 VDD.t1859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1226 a_n3606_12466.t2 B[1].t4 VDD.t710 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1227 a_30006_11681.t0 A[3].t17 a_29769_12318.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1228 a_28011_9265.t0 a_25877_9997.t12 a_27775_9997.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1229 a_14496_9265.t0 a_14790_9971.t4 VSS.t133 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1230 a_28617_21790.t5 a_n3113_6918.t16 VDD.t1407 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1231 a_5505_18852.t6 a_5860_19519.t12 VDD.t2594 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1232 a_12598_9997.t5 a_12053_10690.t6 a_12480_9997.t7 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1233 a_17951_10802.t3 a_17361_11239.t7 VDD.t2277 VDD.t2276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1234 VSS.t423 a_n3111_15192.t21 a_7308_25153.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1235 a_14373_18822.t2 a_n3113_2781.t12 VDD.t568 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1236 VDD.t56 a_14366_24457.t10 a_15719_25150.t0 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1237 a_25804_25129.t1 a_22608_26705.t8 a_25567_25766.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1238 a_9751_24460.t5 a_9206_25153.t6 a_9751_23728.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1239 VSS.t397 a_6041_4129.t12 a_7394_4822.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1240 a_1254_13136.t1 A[4].t20 VDD.t1634 VDD.t1633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1241 a_8419_26709.t3 a_8155_27292.t6 VDD.t506 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1242 a_22104_21787.t0 a_n3115_4850.t14 VDD.t1373 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1243 a_30081_813.t1 B[6].t10 a_29844_1450.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1244 a_18952_19520.t7 a_n3115_4850.t15 a_20849_18121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1245 VDD.t1285 a_36755_7247.t9 Y[5].t2 VDD.t1284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1246 VDD.t2599 a_17356_9635.t9 a_17946_9198.t2 VDD.t2598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1247 Y[7].t2 a_36751_971.t10 VDD.t1258 VDD.t1257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1248 a_23964_7089.t6 a_21145_4128.t15 VDD.t1583 VDD.t1582 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1249 a_n3115_713.t0 a_n3608_55.t7 a_n3808_656.t0 VDD.t1951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1250 a_14036_6963.t2 a_11291_5000.t7 a_14154_6963.t3 VDD.t898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1251 VDD.t1421 a_4963_19248.t17 a_9003_18532.t5 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1252 VDD.t1306 a_6049_9909.t10 a_7829_9909.t9 VDD.t1305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1253 a_n2381_9223.t1 B[3].t6 VSS.t167 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1254 a_19599_25325.t3 a_19009_25762.t8 VDD.t345 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1255 VSS.t257 a_21746_1762.t12 a_24215_4802.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1256 VDD.t2551 a_30430_6928.t13 a_31466_10393.t1 VDD.t2550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1257 a_25567_25766.t4 a_22608_26705.t9 VDD.t450 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1258 a_26435_6378.t2 a_26171_6961.t6 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1259 VDD.t2519 A[3].t18 a_25562_24162.t2 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1260 a_20782_24452.t0 a_n3111_11055.t19 VDD.t577 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1261 a_n3608_1494.t2 opcode[0].t41 VDD.t1862 VDD.t1861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1262 a_13951_10690.t2 a_12598_9997.t11 VDD.t1250 VDD.t1249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1263 a_21150_9929.t4 a_20605_10622.t5 a_21150_9197.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1264 a_8543_1769.t2 a_7953_1332.t9 VDD.t2016 VDD.t2015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1265 a_12892_9971.t3 a_8508_14599.t10 VDD.t2050 VDD.t2049 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1266 a_25332_10690.t3 a_20955_6381.t8 VDD.t1765 VDD.t1764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1267 a_5931_9909.t10 a_1844_12699.t11 VDD.t1449 VDD.t1448 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1268 a_7853_24460.t1 a_7308_25153.t6 a_7735_24460.t10 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1269 a_19345_21663.t3 a_22090_20137.t7 VDD.t862 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1270 a_20900_24452.t6 a_20355_25145.t6 a_20782_24452.t10 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1271 a_27313_6965.t0 a_24568_5002.t6 a_27431_6965.t2 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1272 a_21150_9929.t0 a_20605_10622.t6 a_21032_9929.t0 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1273 a_33377_6895.t6 a_30427_3858.t8 VDD.t1215 VDD.t1214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1274 a_38088_7956.t0 a_18715_18853.t10 VSS.t99 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1275 a_30359_8848.t2 a_29769_9285.t9 VDD.t1146 VDD.t1145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1276 VDD.t2279 a_17361_11239.t8 a_17951_10802.t2 VDD.t2278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1277 a_25790_26779.t0 A[3].t19 a_25553_27416.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1278 VDD.t322 a_27321_12833.t6 a_27585_12250.t3 VDD.t321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1279 a_7939_4129.t3 a_7394_4822.t5 a_7821_4129.t3 VDD.t2286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1280 VDD.t2139 A[5].t15 a_21156_1325.t6 VDD.t2138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1281 a_12598_9265.t0 a_12892_9971.t6 VSS.t129 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1282 a_15719_25150.t3 a_14366_24457.t11 VDD.t537 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1283 VSS.t325 a_n3113_8987.t14 a_25804_25129.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1284 a_31893_6205.t6 a_31466_6898.t6 a_32011_6205.t5 VDD.t502 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1285 VDD.t93 a_14036_6963.t7 a_10647_11281.t1 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1286 VDD.t95 a_26443_12246.t7 a_27439_12833.t3 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1287 a_9987_23728.t1 a_7853_24460.t12 a_9751_24460.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1288 VDD.t2430 a_10641_5411.t12 a_10701_5437.t1 VDD.t2429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1289 VSS.t1 a_27767_4129.t9 a_38088_8192.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1290 a_21150_9197.t0 a_21444_9903.t6 VSS.t265 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1291 VSS.t182 a_n3604_14534.t6 a_n2379_15192.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1292 a_14042_12833.t2 a_11297_10870.t5 VSS.t28 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1293 a_17941_3397.t0 a_17351_3834.t9 VSS.t221 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1294 a_4136_7089.t1 a_1817_6836.t13 VDD.t1357 VDD.t1356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1295 VDD.t2531 a_17301_11213.t11 a_21032_9929.t10 VDD.t2530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1296 VDD.t1863 opcode[0].t42 a_10045_24434.t2 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1297 a_38088_23958.t0 opcode[1].t34 a_36755_23013.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1298 a_9003_18532.t4 a_4963_19248.t18 VDD.t1419 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1299 a_5923_4129.t6 a_5496_4822.t5 a_6041_4129.t4 VDD.t1654 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1300 a_7829_9909.t10 a_6049_9909.t11 VDD.t1308 VDD.t1307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1301 a_19554_12761.t3 a_17946_9198.t4 VSS.t433 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1302 a_26297_12829.t2 a_24562_12520.t5 VDD.t893 VDD.t892 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1303 a_19594_23721.t1 a_19004_24158.t10 VDD.t252 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1304 VSS.t310 a_1833_4076.t12 a_4387_4802.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1305 VDD.t34 a_19009_25762.t9 a_19599_25325.t2 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1306 a_31466_2550.t0 a_30434_1013.t10 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1307 VDD.t1799 a_n3113_8987.t15 a_25567_25766.t2 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1308 VSS.t316 a_32009_13791.t10 a_38084_17682.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1309 a_6607_6378.t2 a_6343_6961.t6 VDD.t662 VDD.t661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1310 VDD.t201 a_10647_11281.t14 a_10702_9703.t0 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1311 a_29844_1450.t5 B[6].t11 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1312 a_26289_6961.t1 a_24563_3398.t5 a_26171_6961.t3 VDD.t542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1313 VDD.t1097 A[0].t5 a_7735_24460.t3 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1314 VDD.t785 a_28603_20140.t7 a_25858_21666.t3 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1315 a_10647_11281.t0 a_14036_6963.t8 VSS.t20 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1316 VDD.t615 A[2].t1 a_20782_24452.t8 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1317 VDD.t1252 a_12598_9997.t12 a_13951_10690.t3 VDD.t1251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1318 a_4098_11193.t3 a_33377_10390.t8 VDD.t2450 VDD.t2449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1319 a_25564_21692.t2 a_25504_21666.t4 VDD.t440 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1320 a_8183_9177.t1 a_6049_9909.t12 a_7947_9909.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1321 a_29650_24430.t1 a_22608_26705.t10 VDD.t464 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1322 VDD.t122 a_36751_13593.t9 Y[3].t2 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1323 a_28902_27292.t4 a_26157_25329.t6 VSS.t188 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1324 a_36751_1089.t9 opcode[1].t35 VDD.t1533 VDD.t1532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1325 VDD.t2052 a_8508_14599.t11 a_12892_9971.t2 VDD.t2051 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1326 a_14042_12833.t4 a_11297_10870.t6 a_14160_12833.t4 VDD.t161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1327 VDD.t166 a_17347_12889.t9 a_17937_12452.t0 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1328 VDD.t616 A[2].t2 a_19004_24158.t3 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1329 a_36755_7365.t0 a_27767_4129.t10 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1330 VDD.t1767 a_20955_6381.t9 a_25332_10690.t2 VDD.t1766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1331 VDD.t1451 a_1844_12699.t12 a_5931_9909.t9 VDD.t1450 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1332 a_23972_12957.t1 a_21711_14619.t13 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1333 a_7735_24460.t6 a_8147_24434.t4 a_7853_24460.t5 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1334 VDD.t863 a_22090_20137.t8 a_19345_21663.t2 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1335 a_n3804_10998.t10 a_n3604_11836.t6 a_n3111_11055.t6 VDD.t820 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1336 VDD.t1800 a_n3113_8987.t16 a_25553_27416.t6 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1337 a_20782_24452.t3 a_21194_24426.t5 a_20900_24452.t0 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1338 a_17951_10802.t1 a_17361_11239.t9 VDD.t2281 VDD.t2280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1339 VDD.t917 a_24568_19252.t12 a_24570_19549.t3 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1340 a_n3113_13124.t6 a_n3606_13905.t6 a_n3806_13067.t10 VDD.t1090 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1341 VDD.t664 a_6343_6961.t7 a_6607_6378.t1 VDD.t663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1342 a_5623_18120.t1 a_5917_18826.t5 a_5623_18852.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1343 VDD.t251 a_24554_6652.t6 a_26289_6961.t4 VDD.t250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1344 a_15057_14598.t3 a_14467_15035.t8 VDD.t2072 VDD.t2071 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1345 a_22798_24452.t6 a_23092_24426.t6 a_22680_24452.t10 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1346 VDD.t1394 a_30359_8848.t11 a_31893_9700.t0 VDD.t1393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1347 VSS.t314 a_17296_5412.t13 a_17588_3197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1348 VSS.t420 a_20058_21029.t8 a_18991_21663.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1349 a_18952_19520.t6 a_19955_19546.t6 a_20495_18853.t5 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1350 a_7939_4129.t5 a_7394_4822.t6 a_7939_3397.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1351 VSS.t243 a_23926_11281.t14 a_24218_9066.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1352 VDD.t1535 opcode[1].t36 a_36755_10509.t5 VDD.t1534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1353 a_10045_24434.t1 opcode[0].t43 VDD.t1864 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1354 a_36751_4233.t7 opcode[1].t37 VDD.t1537 VDD.t1536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1355 a_17593_8998.t0 a_15057_14598.t10 a_17356_9635.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1356 VSS.t5 a_17937_12452.t5 a_19554_12761.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1357 VDD.t895 a_24562_12520.t6 a_26297_12829.t1 VDD.t894 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1358 a_19599_25325.t1 a_19009_25762.t10 VDD.t63 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1359 VSS.t249 a_36755_7247.t10 Y[5].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1360 VDD.t1017 a_27458_24456.t11 a_28811_25149.t3 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1361 VDD.t2190 a_7947_9909.t16 a_31464_14484.t1 VDD.t2189 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1362 a_7735_24460.t4 A[0].t6 VDD.t1098 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1363 a_23978_5439.t3 a_23918_5413.t10 VDD.t2246 VDD.t2245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1364 a_13012_6959.t3 a_11286_3396.t7 a_12894_6959.t3 VDD.t273 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1365 a_25858_21666.t2 a_28603_20140.t8 VDD.t786 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1366 VSS.t109 a_n3606_2123.t6 a_n2381_2781.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1367 a_19247_4128.t7 a_19541_4102.t7 a_19129_4128.t4 VDD.t1203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1368 a_30427_3858.t2 a_29837_4295.t9 VDD.t867 VDD.t866 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1369 VDD.t2452 a_33377_10390.t9 a_4098_11193.t2 VDD.t2451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1370 VDD.t441 a_25504_21666.t5 a_25564_21692.t1 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1371 a_31893_1857.t3 a_30434_1013.t11 VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1372 a_4740_5002.t0 a_4150_5439.t10 VSS.t398 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1373 a_14160_12833.t3 a_11297_10870.t7 a_14042_12833.t1 VDD.t507 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1374 VDD.t279 a_15561_18528.t7 a_13953_21654.t3 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1375 a_6343_9883.t1 a_1844_12699.t13 VDD.t1453 VDD.t1452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1376 a_17937_12452.t1 a_17347_12889.t10 VDD.t227 VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1377 a_19004_24158.t2 A[2].t3 VDD.t617 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1378 a_29650_24430.t0 a_22608_26705.t11 VSS.t90 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1379 a_27775_9997.t2 a_27230_10690.t5 a_27657_9997.t1 VDD.t527 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1380 a_19134_9929.t8 a_19546_9903.t6 a_19252_9929.t6 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1381 VDD.t2559 a_32011_1857.t10 a_36751_13711.t3 VDD.t2558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1382 VDD.t1769 a_20955_6381.t10 a_23972_12957.t6 VDD.t1768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1383 a_7853_24460.t6 a_8147_24434.t5 a_7735_24460.t7 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1384 a_22090_20137.t6 a_n3115_4850.t16 VDD.t1374 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1385 VDD.t780 a_12382_21028.t7 a_4963_19248.t2 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1386 a_24570_19549.t2 a_24568_19252.t13 VDD.t918 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1387 VSS.t36 a_6615_12158.t4 a_7493_12745.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1388 VDD.t557 a_32011_9700.t11 a_36755_19987.t8 VDD.t556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1389 a_23986_11307.t1 a_20955_6381.t11 VDD.t1771 VDD.t1770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1390 VDD.t1408 a_n3113_6918.t17 a_27008_18856.t6 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1391 VDD.t103 a_4726_6652.t6 a_6461_6961.t4 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1392 a_24563_3398.t2 a_23973_3835.t8 VDD.t891 VDD.t890 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1393 VDD.t423 B[6].t12 a_n3606_2123.t3 VDD.t422 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1394 a_19546_9903.t0 a_15057_14598.t11 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1395 a_19672_12761.t2 a_17946_9198.t5 a_19554_12761.t4 VDD.t2520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1396 VDD.t2074 a_14467_15035.t9 a_15057_14598.t2 VDD.t2073 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1397 a_10687_7087.t0 a_8543_1769.t11 VDD.t688 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1398 VDD.t425 B[6].t13 a_n3806_2724.t9 VDD.t424 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1399 a_7749_6382.t1 a_7485_6965.t5 VSS.t162 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1400 a_12592_4127.t6 a_12047_4820.t6 a_12474_4127.t11 VDD.t1153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1401 a_6351_12741.t1 a_4743_9178.t4 VSS.t183 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1402 a_20058_21029.t4 a_20133_21659.t5 VSS.t185 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1403 VSS.t406 a_11523_19541.t5 a_12181_18116.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1404 VDD.t2152 a_14490_4127.t13 a_31893_1857.t10 VDD.t2151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1405 a_17301_11213.t2 a_33377_2547.t9 VDD.t2120 VDD.t2119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1406 VSS.t379 a_18055_19249.t7 a_18057_19546.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1407 a_19129_4128.t1 a_15097_1774.t12 VDD.t2215 VDD.t2214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1408 VDD.t2533 a_17301_11213.t12 a_21444_9903.t2 VDD.t2532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1409 a_17347_12889.t6 a_15057_14598.t12 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1410 a_36751_16855.t8 a_22798_24452.t9 a_36751_16737.t7 VDD.t1010 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1411 VDD.t1277 B[7].t4 a_n3608_55.t2 VDD.t1276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1412 a_n3808_656.t4 a_n3608_1494.t6 a_n3115_713.t5 VDD.t783 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1413 VDD.t1255 a_n3113_2781.t13 a_15570_21782.t6 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1414 a_28811_25149.t2 a_27458_24456.t12 VDD.t1018 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1415 a_36697_5000.t0 opcode[1].t38 VSS.t286 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1416 a_36751_16855.t5 opcode[1].t39 VDD.t1539 VDD.t1538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1417 a_4150_5439.t2 a_4090_5413.t11 VDD.t1071 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1418 a_38084_17446.t1 a_22798_24452.t10 VSS.t198 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1419 VDD.t1099 A[0].t7 a_7735_24460.t5 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1420 VDD.t264 a_17937_12452.t6 a_19672_12761.t4 VDD.t263 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1421 a_36755_23131.t5 a_36701_23898.t6 a_36755_23013.t2 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1422 a_36697_17622.t1 opcode[1].t40 VDD.t1541 VDD.t1540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1423 a_n3806_6861.t1 opcode[0].t44 VDD.t1866 VDD.t1865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1424 a_36755_7247.t6 a_36701_8132.t6 a_36755_7365.t11 VDD.t1088 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1425 a_4098_11193.t1 a_33377_10390.t10 VDD.t2275 VDD.t2274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1426 a_25564_21692.t0 a_25504_21666.t6 VDD.t442 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1427 a_12900_12829.t0 a_11292_9266.t7 VSS.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1428 VDD.t2609 a_13164_12246.t4 a_14160_12833.t2 VDD.t2608 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1429 a_27767_4129.t0 a_28061_4103.t7 a_27649_4129.t4 VDD.t1138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1430 a_23972_12957.t5 a_20955_6381.t12 VDD.t1773 VDD.t1772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1431 a_7735_24460.t8 a_8147_24434.t6 a_7853_24460.t7 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1432 VDD.t1375 a_n3115_4850.t17 a_22090_20137.t5 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1433 VDD.t471 a_12418_19515.t12 a_12475_18822.t0 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1434 a_20193_21685.t1 a_20487_21659.t5 a_20058_21029.t1 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1435 VDD.t919 a_24568_19252.t14 a_25110_18856.t7 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1436 VDD.t920 a_24568_19252.t15 a_24570_19549.t1 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1437 a_4090_5413.t0 a_7493_12745.t6 VSS.t261 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1438 a_n3113_2781.t4 a_n3606_3562.t5 a_n3806_2724.t6 VDD.t1197 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1439 a_16264_24457.t4 a_15719_25150.t7 a_16264_23725.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1440 a_36751_971.t1 a_36697_1856.t5 a_38084_1680.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1441 VDD.t1702 a_1833_4076.t13 a_4150_5439.t5 VDD.t1701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1442 a_7394_4822.t2 a_6041_4129.t13 VDD.t2299 VDD.t2298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1443 a_19554_12761.t1 a_17946_9198.t6 a_19672_12761.t1 VDD.t2521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1444 a_15057_14598.t1 a_14467_15035.t10 VDD.t2076 VDD.t2075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1445 a_23964_7089.t1 a_21746_1762.t13 VDD.t1330 VDD.t1329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1446 VDD.t2022 a_10693_12957.t9 a_11283_12520.t2 VDD.t2021 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1447 VDD.t1635 A[4].t21 a_28608_18536.t4 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1448 VDD.t31 a_13158_6376.t5 a_14154_6963.t1 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1449 a_25553_27416.t2 A[3].t20 VDD.t2354 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1450 a_24210_3198.t1 a_21145_4128.t16 a_23973_3835.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1451 a_n3606_3562.t1 opcode[0].t45 VDD.t1868 VDD.t1867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1452 a_32011_1857.t4 a_31466_2550.t6 a_32011_1125.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1453 VDD.t324 a_27321_12833.t7 a_27585_12250.t2 VDD.t323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1454 VSS.t152 a_4734_12432.t4 a_6351_12741.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1455 a_19247_4128.t4 a_18702_4821.t6 a_19247_3396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1456 a_7815_18826.t3 a_n3115_713.t17 VDD.t1945 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1457 VDD.t1256 a_n3113_2781.t14 a_14373_18822.t1 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1458 a_12417_18116.t1 a_11521_19244.t15 VSS.t276 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1459 a_7611_12745.t5 a_6615_12158.t5 VDD.t1007 VDD.t1006 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1460 a_26171_6961.t2 a_24563_3398.t6 VSS.t114 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1461 a_21444_9903.t1 a_17301_11213.t13 VDD.t2535 VDD.t2534 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1462 a_22744_17922.t0 a_18055_19249.t8 VSS.t380 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1463 VDD.t2106 B[5].t15 a_7953_1332.t2 VDD.t2105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1464 a_15570_21782.t4 a_n3113_2781.t15 VDD.t818 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1465 VSS.t417 a_10641_5411.t13 a_14726_3395.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1466 VDD.t737 a_7749_6382.t16 a_12053_10690.t3 VDD.t736 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1467 a_12418_19515.t5 a_13421_19541.t5 a_13961_18848.t9 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1468 a_25751_4129.t1 a_26163_4103.t6 a_25869_4129.t5 VDD.t1289 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1469 VSS.t247 B[7].t5 a_n3608_55.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1470 a_36751_4115.t6 a_36697_5000.t5 a_38084_4824.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1471 a_7829_9909.t11 a_6049_9909.t13 VDD.t1310 VDD.t1309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1472 a_4734_12432.t1 a_4144_12869.t10 VDD.t1652 VDD.t1651 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1473 a_36751_13711.t8 a_36697_14478.t6 a_36751_13593.t5 VDD.t1169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1474 VDD.t2386 a_14496_9997.t19 a_18707_10622.t1 VDD.t2385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1475 VSS.t75 a_11283_12520.t4 a_12900_12829.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1476 a_17351_3834.t5 a_14306_12250.t11 VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1477 a_14160_12833.t1 a_13164_12246.t5 VDD.t2604 VDD.t2603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1478 a_23981_9703.t0 a_21711_14619.t14 VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1479 VDD.t2141 A[5].t16 a_21156_1325.t5 VDD.t2140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1480 a_22090_20137.t4 a_n3115_4850.t18 VDD.t1376 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1481 a_20058_21029.t2 a_20487_21659.t6 a_20193_21685.t0 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1482 a_25110_18856.t8 a_24568_19252.t16 VDD.t921 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1483 a_6469_12741.t2 a_4743_9178.t5 a_6351_12741.t0 VDD.t945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1484 a_31893_9700.t7 a_32305_9674.t6 a_32011_9700.t5 VDD.t949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1485 a_36755_10391.t3 a_36701_11276.t6 a_36755_10509.t7 VDD.t1047 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1486 a_21711_14619.t0 a_21121_15056.t7 VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1487 a_7853_24460.t4 a_7308_25153.t7 a_7853_23728.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1488 a_23092_24426.t1 a_16074_26710.t13 VDD.t1922 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1489 a_32305_6179.t1 a_21150_9929.t16 VDD.t2576 VDD.t2575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1490 a_16500_23725.t0 a_14366_24457.t12 a_16264_24457.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1491 VSS.t63 a_32011_6205.t9 a_38088_11336.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1492 VDD.t1000 a_11283_12520.t5 a_13018_12829.t5 VDD.t999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1493 VDD.t1009 a_26435_6378.t5 a_27431_6965.t5 VDD.t1008 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1494 a_4136_7089.t4 a_1833_4076.t14 VDD.t1704 VDD.t1703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1495 a_11283_12520.t1 a_10693_12957.t10 VDD.t2024 VDD.t2023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1496 a_28608_18536.t5 A[4].t22 VDD.t1636 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1497 a_4382_3198.t1 a_1817_6836.t14 a_4145_3835.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1498 a_8419_26709.t2 a_8155_27292.t7 VSS.t81 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1499 VDD.t1801 a_n3113_8987.t17 a_25553_27416.t5 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1500 a_20782_24452.t9 a_20355_25145.t7 a_20900_24452.t7 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1501 a_1243_4513.t4 B[3].t7 VDD.t852 VDD.t851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1502 a_27585_12250.t1 a_27321_12833.t8 VDD.t326 VDD.t325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1503 a_6615_12158.t0 a_6351_12741.t5 VSS.t50 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1504 VDD.t1946 a_n3115_713.t18 a_7815_18826.t2 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1505 a_12181_18848.t0 a_12418_19515.t13 a_12417_18116.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1506 a_10696_3833.t2 a_7939_4129.t19 VDD.t1106 VDD.t1105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1507 VDD.t1734 a_17296_5412.t14 a_17351_3834.t3 VDD.t1733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1508 a_31893_6205.t4 a_32305_6179.t6 a_32011_6205.t1 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1509 a_17946_5001.t2 a_17356_5438.t8 VDD.t1686 VDD.t1685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1510 a_23918_5413.t1 a_33377_6895.t8 VSS.t217 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1511 VDD.t996 a_20696_12765.t7 a_17296_5412.t3 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1512 VDD.t53 a_6615_12158.t6 a_7611_12745.t0 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1513 a_7403_18852.t0 a_7815_18826.t5 a_5860_19519.t0 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1514 VDD.t1053 a_10702_9703.t10 a_11292_9266.t1 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1515 a_4090_5413.t2 a_7493_12745.t7 VDD.t1363 VDD.t1362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1516 a_29844_1450.t1 A[3].t21 VDD.t2356 VDD.t2355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1517 a_32305_6179.t0 a_21150_9929.t17 VSS.t106 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1518 a_21202_27284.t1 a_19594_23721.t4 VSS.t60 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1519 VDD.t1083 a_19549_6960.t7 a_19813_6377.t2 VDD.t1082 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1520 a_9012_21786.t1 a_n3115_713.t19 VDD.t1947 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1521 a_36751_4233.t0 a_12181_18848.t10 a_36751_4115.t1 VDD.t2348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1522 VDD.t1244 a_27775_9997.t10 a_36751_4233.t9 VDD.t1243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1523 a_7947_9177.t1 a_8241_9883.t6 VSS.t23 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1524 a_5923_4129.t2 a_6335_4103.t6 a_6041_4129.t1 VDD.t788 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1525 VDD.t1165 a_33377_6895.t9 a_23918_5413.t2 VDD.t1164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1526 a_13961_18848.t8 a_13421_19541.t6 a_12418_19515.t4 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1527 a_18597_18853.t5 a_18055_19249.t9 VDD.t2195 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1528 a_14248_24457.t5 a_n3113_13124.t18 VDD.t673 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1529 VDD.t2432 a_10641_5411.t14 a_14784_4101.t2 VDD.t2431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1530 a_6335_4103.t0 a_1817_6836.t15 VSS.t260 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1531 VDD.t771 a_1243_4513.t10 a_1833_4076.t0 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1532 VDD.t1217 a_30427_3858.t9 a_31466_6898.t2 VDD.t1216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1533 a_n2379_11291.t1 B[2].t4 VSS.t67 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1534 a_10641_5411.t3 a_33375_14481.t10 VDD.t1185 VDD.t1184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1535 VDD.t2434 a_10641_5411.t15 a_10696_3833.t5 VDD.t2433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1536 VDD.t2597 a_13164_12246.t6 a_14160_12833.t0 VDD.t2596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1537 a_10701_5437.t5 a_8543_1769.t12 VDD.t929 VDD.t928 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1538 VDD.t2335 a_12592_4127.t12 a_13945_4820.t2 VDD.t2334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1539 VDD.t638 a_29840_7365.t10 a_30430_6928.t3 VDD.t637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1540 a_20809_6964.t0 a_17946_5001.t5 a_20691_6964.t0 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1541 a_n3606_13905.t0 opcode[0].t46 VSS.t331 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1542 VDD.t692 a_9561_26713.t13 a_16146_24457.t6 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1543 VDD.t1927 a_25465_19523.t13 a_25110_18856.t2 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1544 VDD.t2553 a_30430_6928.t14 a_33377_10390.t0 VDD.t2552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1545 a_6351_12741.t3 a_4743_9178.t6 a_6469_12741.t1 VDD.t438 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1546 a_n2379_15428.t1 B[0].t3 VSS.t231 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1547 VDD.t1073 a_4090_5413.t12 a_7821_4129.t6 VDD.t1072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1548 VDD.t338 a_21121_15056.t8 a_21711_14619.t1 VDD.t337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1549 VSS.t332 opcode[0].t47 a_9987_23728.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1550 a_22344_27288.t0 a_19599_25325.t4 VSS.t49 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1551 a_1817_6836.t0 a_1227_7273.t9 VSS.t323 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1552 a_8998_20136.t6 a_n3115_713.t20 VDD.t1948 w_8904_20100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1553 a_13018_12829.t0 a_11283_12520.t6 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1554 a_19004_24158.t1 A[2].t4 VDD.t618 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1555 VDD.t2611 a_12900_12829.t7 a_13164_12246.t0 VDD.t2610 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1556 a_19585_26975.t1 a_18995_27412.t10 VDD.t50 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1557 a_25553_27416.t4 a_n3113_8987.t18 VDD.t1802 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1558 VDD.t926 a_18916_21033.t6 a_11521_19244.t1 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1559 a_36701_20754.t0 opcode[1].t41 VSS.t287 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1560 VDD.t1637 A[4].t23 a_28608_18536.t6 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1561 a_23973_3835.t5 a_21145_4128.t17 VDD.t1585 VDD.t1584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1562 VDD.t1543 opcode[1].t42 a_36701_23898.t1 VDD.t1542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1563 VSS.t190 a_36755_10391.t11 Y[4].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1564 a_13659_21680.t2 a_13953_21654.t5 a_13524_21024.t3 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1565 a_12181_18116.t1 a_12475_18822.t7 a_12181_18848.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1566 VSS.t280 a_1844_12699.t14 a_6285_9177.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1567 a_5623_18852.t7 a_5860_19519.t13 a_5859_18120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1568 a_9647_19525.t1 a_n3115_713.t21 VSS.t345 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1569 a_21121_15056.t3 A[6].t16 VDD.t2480 VDD.t2479 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1570 VDD.t427 B[6].t14 a_29844_1450.t4 VDD.t426 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1571 VDD.t147 A[7].t3 a_9012_21786.t0 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1572 a_7603_6965.t1 a_6607_6378.t6 VDD.t584 VDD.t583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1573 VDD.t619 A[2].t5 a_18995_27412.t6 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1574 a_12418_19515.t6 a_13421_19541.t7 a_13961_18848.t10 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1575 a_14790_9971.t0 a_10647_11281.t15 VSS.t39 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1576 a_20691_6964.t2 a_17946_5001.t6 VSS.t108 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1577 a_17361_11239.t6 a_17301_11213.t14 VDD.t2537 VDD.t2536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1578 a_n3806_6861.t3 a_n3606_6260.t6 a_n3113_6918.t3 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1579 a_9751_24460.t6 a_9206_25153.t7 a_9633_24460.t6 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1580 VDD.t1587 a_21145_4128.t18 a_23973_3835.t4 VDD.t1586 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1581 VDD.t2444 a_15570_21782.t9 a_13599_21654.t1 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1582 VSS.t371 A[5].t17 a_19955_19546.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1583 a_n3608_5631.t0 opcode[0].t48 VSS.t333 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1584 a_8273_27292.t5 a_6547_23729.t5 a_8155_27292.t4 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1585 a_21320_27284.t2 a_19594_23721.t5 a_21202_27284.t3 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1586 a_13012_6959.t1 a_11277_6650.t6 VDD.t2315 VDD.t2314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1587 a_4153_9615.t0 a_4098_11193.t13 VDD.t462 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1588 VDD.t1870 opcode[0].t49 a_n3804_10998.t6 VDD.t1869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1589 VDD.t2108 B[5].t16 a_29769_12318.t6 VDD.t2107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1590 a_17932_6651.t2 a_17342_7088.t8 VDD.t595 VDD.t594 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1591 a_16146_24457.t7 a_9561_26713.t14 VDD.t693 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1592 a_7939_3397.t1 a_8233_4103.t6 VSS.t32 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1593 a_25110_18856.t1 a_25465_19523.t14 VDD.t1928 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1594 a_n3113_6918.t5 a_n3606_7699.t5 a_n3806_6861.t10 VDD.t1603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1595 a_6469_12741.t0 a_4743_9178.t7 a_6351_12741.t2 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1596 a_9751_23728.t1 a_10045_24434.t7 VSS.t51 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1597 VSS.t407 a_21466_26701.t6 a_22344_27288.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1598 VDD.t1175 a_30427_3858.t10 a_31893_6205.t10 VDD.t1174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1599 a_27657_9997.t10 a_28069_9971.t5 a_27775_9997.t6 VDD.t1187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1600 a_36755_10509.t4 opcode[1].t43 VDD.t1545 VDD.t1544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1601 VSS.t25 a_22090_20137.t9 a_19345_21663.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1602 VDD.t2154 a_14490_4127.t14 a_31893_1857.t11 VDD.t2153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1603 VSS.t377 a_7947_9909.t17 a_31464_14484.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1604 VDD.t2482 A[6].t17 a_7918_15036.t2 VDD.t2481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1605 a_11521_19244.t0 a_18916_21033.t7 VDD.t483 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1606 a_36755_19869.t3 a_36701_20754.t7 a_36755_19987.t3 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1607 VDD.t2337 a_12592_4127.t13 a_14372_4127.t11 VDD.t2336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1608 VDD.t860 a_15057_14598.t13 a_17356_9635.t3 VDD.t859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1609 a_12480_9997.t5 a_8508_14599.t12 VDD.t2054 VDD.t2053 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1610 VDD.t1872 opcode[0].t50 a_n3604_11836.t2 VDD.t1871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1611 VSS.t353 B[4].t12 a_n3606_6260.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1612 a_11277_6650.t1 a_10687_7087.t9 VDD.t2324 VDD.t2323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1613 VDD.t1409 a_n3113_6918.t18 a_28617_21790.t4 w_28523_21754# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1614 VSS.t258 a_21746_1762.t14 a_25324_4822.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1615 a_25759_9997.t2 a_25332_10690.t5 a_25877_9997.t3 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1616 a_22462_27288.t2 a_19599_25325.t5 a_22344_27288.t3 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1617 VDD.t1803 a_n3113_8987.t19 a_26913_25149.t2 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1618 VSS.t191 a_6253_21662.t7 a_5824_21032.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1619 VDD.t344 a_26179_12829.t8 a_26443_12246.t1 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1620 VDD.t1547 opcode[1].t44 a_36697_5000.t1 VDD.t1546 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1621 a_31893_6205.t7 a_21150_9929.t18 VDD.t2574 VDD.t2573 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1622 a_18995_27412.t5 A[2].t6 VDD.t70 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1623 a_13961_18848.t7 a_14373_18822.t6 a_12418_19515.t3 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1624 a_6547_23729.t3 a_5957_24166.t7 VDD.t1784 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1625 a_12474_4127.t1 a_8543_1769.t13 VDD.t931 VDD.t930 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1626 VDD.t453 a_1817_6836.t16 a_4145_3835.t0 VDD.t452 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1627 a_32011_9700.t0 a_31466_10393.t6 a_32011_8968.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1628 VDD.t394 a_6351_12741.t6 a_6615_12158.t3 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1629 VSS.t282 B[3].t8 a_30006_8648.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1630 a_15570_21782.t5 a_n3113_2781.t16 VDD.t819 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1631 a_32011_1857.t7 a_31466_2550.t7 a_31893_1857.t6 VDD.t2446 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1632 a_8155_27292.t3 a_6547_23729.t6 a_8273_27292.t4 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1633 a_22253_25145.t2 a_20900_24452.t12 VDD.t1416 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1634 a_25504_21666.t1 a_26571_21032.t8 VDD.t445 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1635 a_n3606_2123.t2 B[6].t15 VDD.t429 VDD.t428 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1636 a_14732_9265.t1 a_12598_9997.t13 a_14496_9997.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1637 a_12474_4127.t3 a_12886_4101.t6 a_12592_4127.t1 VDD.t2344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1638 a_25877_9997.t2 a_25332_10690.t6 a_25759_9997.t1 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1639 VDD.t1873 opcode[0].t51 a_9633_24460.t0 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1640 VDD.t694 a_9561_26713.t15 a_16558_24431.t2 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1641 a_21194_24426.t3 A[2].t7 VDD.t71 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1642 a_20814_12765.t1 a_17951_10802.t4 a_20696_12765.t1 VDD.t509 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1643 VDD.t695 a_9561_26713.t16 a_16146_24457.t8 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1644 VDD.t748 a_4734_12432.t5 a_6469_12741.t5 VDD.t747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1645 a_6335_4103.t1 a_1817_6836.t17 VDD.t455 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1646 a_9561_26713.t3 a_9297_27296.t6 VSS.t98 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1647 a_13065_25330.t0 a_12475_25767.t8 VSS.t303 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1648 VDD.t2231 a_14507_1337.t10 a_15097_1774.t1 VDD.t2230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1649 a_n3806_8930.t8 B[3].t9 VDD.t1467 VDD.t1466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1650 VSS.t186 a_30434_1013.t12 a_33614_1910.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1651 a_n3808_4793.t10 a_n3608_5631.t6 a_n3115_4850.t6 VDD.t947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1652 a_7918_15036.t1 A[6].t18 VDD.t2484 VDD.t2483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1653 a_12475_18822.t1 a_12418_19515.t14 VDD.t472 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1654 VDD.t1875 opcode[0].t52 a_n3806_2724.t2 VDD.t1874 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1655 VDD.t1639 A[4].t24 a_7953_1332.t6 VDD.t1638 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1656 a_1817_6836.t1 a_1227_7273.t10 VDD.t1930 VDD.t1929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1657 VDD.t2056 a_8508_14599.t13 a_12480_9997.t4 VDD.t2055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1658 a_24554_6652.t2 a_23964_7089.t9 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1659 VDD.t465 a_22608_26705.t12 a_29238_24456.t3 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1660 a_5623_18852.t0 a_4965_19545.t7 a_5505_18852.t0 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1661 VDD.t1461 B[3].t10 a_29769_9285.t5 VDD.t1460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1662 a_22344_27288.t2 a_19599_25325.t6 a_22462_27288.t1 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1663 a_25751_4129.t2 a_26163_4103.t7 a_25869_4129.t4 VDD.t1290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1664 a_21032_9929.t11 a_20605_10622.t7 a_21150_9929.t3 VDD.t510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1665 VSS.t372 a_14490_4127.t15 a_32247_1125.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1666 a_36755_7365.t5 opcode[1].t45 VDD.t1549 VDD.t1548 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1667 VSS.t301 A[4].t25 a_26468_19549.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1668 a_1844_12699.t3 a_1254_13136.t10 VSS.t44 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1669 a_7101_21684.t5 a_7041_21658.t4 VDD.t244 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1670 VDD.t1682 a_13599_21654.t5 a_13659_21680.t4 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1671 a_6966_21028.t4 a_7041_21658.t5 VSS.t46 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1672 a_7403_18852.t4 a_7815_18826.t6 a_5860_19519.t2 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1673 a_12418_19515.t1 a_14373_18822.t7 a_13961_18848.t5 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1674 VSS.t148 a_22095_18533.t10 a_20487_21659.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1675 a_25751_4129.t6 a_21746_1762.t15 VDD.t1332 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1676 VDD.t518 a_6615_12158.t7 a_7611_12745.t1 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1677 VDD.t533 a_36751_4115.t11 Y[6].t1 VDD.t532 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1678 a_8241_9883.t2 a_4098_11193.t14 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1679 a_1491_12499.t0 A[4].t26 a_1254_13136.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1680 a_31891_13791.t0 a_32303_13765.t6 a_32009_13791.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1681 VDD.t1785 a_5957_24166.t8 a_6547_23729.t2 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1682 a_16210_17917.t1 a_11521_19244.t16 VSS.t275 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1683 a_6552_25333.t3 a_5962_25770.t8 VDD.t2282 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1684 a_27649_4129.t0 a_25869_4129.t11 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1685 VDD.t1706 a_1833_4076.t15 a_5496_4822.t1 VDD.t1705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1686 VDD.t1463 B[3].t11 a_1246_10551.t5 VDD.t1462 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1687 VDD.t1417 a_20900_24452.t13 a_22253_25145.t1 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1688 a_21027_4128.t9 a_21439_4102.t6 a_21145_4128.t5 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1689 VSS.t349 a_30359_11881.t10 a_32245_13059.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1690 a_11523_19541.t1 a_11521_19244.t17 VDD.t2584 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1691 VDD.t650 A[0].t8 a_8147_24434.t2 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1692 a_16558_24431.t1 a_9561_26713.t17 VDD.t696 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1693 VDD.t72 A[2].t8 a_21194_24426.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1694 a_20696_12765.t0 a_17951_10802.t5 a_20814_12765.t0 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1695 a_21150_9929.t7 a_21444_9903.t7 a_21032_9929.t5 VDD.t1382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1696 a_n3806_8930.t11 a_n3606_9768.t5 a_n3113_8987.t1 VDD.t1787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1697 a_10707_11307.t6 a_10647_11281.t16 VDD.t1189 VDD.t1188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1698 a_21194_24426.t0 A[2].t9 VSS.t17 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1699 a_6469_12741.t4 a_4734_12432.t6 VDD.t750 VDD.t749 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1700 a_20495_18853.t9 A[5].t18 VDD.t2142 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1701 VDD.t1473 a_21156_1325.t9 a_21746_1762.t2 VDD.t1472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1702 VDD.t2485 A[6].t19 a_13421_19541.t1 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1703 a_22104_21787.t3 A[5].t19 a_22753_21176.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1704 a_n2383_5086.t0 B[5].t17 VSS.t366 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1705 VDD.t1877 opcode[0].t53 a_n3606_9768.t2 VDD.t1876 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1706 VDD.t630 a_36755_19869.t10 Y[1].t2 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1707 VDD.t184 a_19252_9929.t15 a_20605_10622.t1 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1708 a_1836_10114.t0 a_1246_10551.t10 VSS.t363 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1709 a_29238_24456.t4 a_22608_26705.t13 VDD.t466 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1710 a_6049_9909.t0 a_5504_10602.t7 a_5931_9909.t6 VDD.t352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1711 VDD.t674 a_n3113_13124.t19 a_12475_25767.t5 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1712 VDD.t877 a_19247_4128.t12 a_21027_4128.t8 VDD.t876 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1713 a_7947_9909.t5 a_7402_10602.t6 a_7829_9909.t5 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1714 VDD.t1551 opcode[1].t46 a_36751_13711.t11 VDD.t1550 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1715 a_27126_18124.t1 a_27420_18830.t6 a_25465_19523.t5 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1716 VSS.t64 B[6].t16 a_30074_3658.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1717 a_12181_18848.t2 a_11523_19541.t6 a_12063_18848.t4 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1718 a_21746_1762.t1 a_21156_1325.t10 VDD.t1475 VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1719 VDD.t1003 a_4098_11193.t15 a_4158_11219.t6 VDD.t1002 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1720 a_13659_21680.t3 a_13599_21654.t6 VDD.t1681 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1721 a_25869_4129.t0 a_25324_4822.t5 a_25869_3397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1722 VSS.t394 a_7395_21658.t7 a_6966_21028.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1723 a_5860_19519.t3 a_7815_18826.t7 a_7403_18852.t5 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1724 a_11291_5000.t1 a_10701_5437.t10 VDD.t390 VDD.t389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1725 a_29356_24456.t1 a_29650_24430.t6 a_29238_24456.t1 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1726 a_6547_23729.t1 a_5957_24166.t9 VDD.t1786 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1727 VDD.t2339 a_12592_4127.t14 a_13945_4820.t1 VDD.t2338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1728 VDD.t1937 a_36755_23013.t11 Y[0].t1 VDD.t1936 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1729 a_n3606_13905.t2 opcode[0].t54 VDD.t1879 VDD.t1878 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1730 a_11286_3396.t0 a_10696_3833.t9 VSS.t61 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1731 a_1246_10551.t0 B[3].t12 VDD.t801 VDD.t800 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1732 a_38088_11100.t0 a_25228_18856.t10 VSS.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1733 a_33612_13844.t0 a_30359_11881.t11 a_33375_14481.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1734 a_10939_9066.t0 a_8508_14599.t14 a_10702_9703.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1735 a_32009_13059.t1 a_32303_13765.t7 VSS.t56 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1736 a_10693_12957.t2 a_8508_14599.t15 VDD.t2058 VDD.t2057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1737 a_8147_24434.t1 A[0].t9 VDD.t651 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1738 a_14366_24457.t5 a_14660_24431.t6 a_14248_24457.t8 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1739 a_21194_24426.t1 A[2].t10 VDD.t73 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1740 a_36701_11276.t1 opcode[1].t47 VDD.t1553 VDD.t1552 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1741 a_20814_12765.t2 a_17951_10802.t6 a_20696_12765.t2 VDD.t899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1742 a_22095_18533.t2 a_18055_19249.t10 VDD.t2196 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1743 VDD.t1804 a_n3113_8987.t20 a_25567_25766.t1 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1744 VDD.t1191 a_10647_11281.t17 a_10707_11307.t5 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1745 a_26105_3397.t0 a_21746_1762.t16 a_25869_4129.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1746 a_n3606_3562.t0 opcode[0].t55 VSS.t334 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1747 VDD.t1708 a_1833_4076.t16 a_5923_4129.t7 VDD.t1707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1748 VDD.t291 B[6].t17 a_29837_4295.t5 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1749 a_n3608_1494.t1 opcode[0].t56 VDD.t1881 VDD.t1880 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1750 a_12698_26780.t0 A[1].t11 a_12461_27417.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1751 a_5957_24166.t3 A[0].t10 VDD.t652 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1752 a_12886_4101.t3 a_7939_4129.t20 VDD.t1108 VDD.t1107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1753 a_9012_21786.t4 A[7].t4 a_9661_21175.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1754 a_33377_2547.t0 a_14490_4127.t16 VDD.t2156 VDD.t2155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1755 a_7815_18826.t0 a_n3115_713.t22 VSS.t346 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1756 VDD.t1455 a_1844_12699.t15 a_4144_12869.t5 VDD.t1454 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1757 VDD.t467 a_22608_26705.t14 a_29238_24456.t5 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1758 a_21381_3396.t0 a_19247_4128.t13 a_21145_4128.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1759 VSS.t351 a_28608_18536.t9 a_27000_21662.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1760 a_13065_25330.t2 a_12475_25767.t9 VDD.t1645 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1761 a_12047_4820.t1 a_8543_1769.t14 VDD.t933 VDD.t932 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1762 a_n3111_11055.t3 opcode[0].t57 a_n2379_11291.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1763 a_11521_19244.t2 a_18916_21033.t8 VDD.t1089 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1764 VSS.t409 A[3].t22 a_30011_14252.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1765 a_4158_11219.t4 a_4098_11193.t16 VDD.t367 VDD.t366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1766 a_33375_14481.t3 a_30359_11881.t12 VDD.t1969 VDD.t1968 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1767 a_18597_18853.t11 a_19009_18827.t5 a_18715_18853.t7 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1768 VDD.t2248 a_23918_5413.t11 a_23973_3835.t1 VDD.t2247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1769 VDD.t717 a_9561_26713.t18 a_12470_24163.t0 w_12316_24101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1770 a_19488_9197.t0 a_14496_9997.t20 a_19252_9929.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1771 a_13524_21024.t1 a_13953_21654.t6 a_13659_21680.t1 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1772 a_n3806_2724.t8 B[6].t18 VDD.t293 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1773 a_24568_5002.t1 a_23978_5439.t10 VDD.t1063 VDD.t1062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1774 VDD.t475 a_25869_4129.t12 a_27222_4822.t0 VDD.t474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1775 a_29840_7365.t5 B[4].t13 VDD.t1998 VDD.t1997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1776 a_29238_24456.t2 a_29650_24430.t7 a_29356_24456.t2 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1777 a_25799_23525.t0 A[3].t23 a_25562_24162.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1778 VDD.t649 a_26143_26979.t7 a_27878_27288.t2 w_27724_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1779 a_9003_18532.t0 A[7].t5 a_9652_17921.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1780 a_24563_3398.t0 a_23973_3835.t9 VSS.t47 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1781 a_17932_6651.t0 a_17342_7088.t9 VSS.t123 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1782 a_36755_7247.t7 a_36701_8132.t7 a_38088_7956.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1783 a_n3606_6260.t1 B[4].t14 VDD.t2000 VDD.t1999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1784 VDD.t2026 A[5].t20 a_1246_10551.t2 VDD.t2025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1785 a_19667_6960.t2 a_17932_6651.t6 VDD.t259 VDD.t258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1786 a_29837_4295.t2 A[4].t27 VDD.t1641 VDD.t1640 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1787 a_14496_9997.t3 a_13951_10690.t7 a_14378_9997.t7 VDD.t2351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1788 VSS.t378 a_7947_9909.t18 a_33612_13844.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1789 a_36751_16737.t1 a_22798_24452.t11 a_36751_16855.t1 VDD.t253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1790 VSS.t348 a_16074_26710.t14 a_23034_23720.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1791 VDD.t2060 a_8508_14599.t16 a_10693_12957.t1 VDD.t2059 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1792 a_18995_27412.t4 A[2].t11 VDD.t74 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1793 VSS.t254 a_6049_9909.t14 a_7402_10602.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1794 a_14248_24457.t9 a_14660_24431.t7 a_14366_24457.t4 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1795 VDD.t2197 a_18055_19249.t11 a_22095_18533.t1 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1796 VDD.t300 a_6351_12741.t7 a_6615_12158.t1 VDD.t299 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1797 a_6277_3397.t1 a_1833_4076.t17 a_6041_4129.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1798 a_10707_11307.t4 a_10647_11281.t18 VDD.t1193 VDD.t1192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1799 VDD.t795 a_7485_6965.t6 a_7749_6382.t2 VDD.t794 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1800 a_36751_16737.t2 a_36697_17622.t6 a_38084_17446.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1801 a_4743_9178.t1 a_4153_9615.t10 VDD.t678 VDD.t677 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1802 VDD.t150 a_n3113_2781.t17 a_13961_18848.t0 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1803 a_15810_27293.t2 a_13065_25330.t5 VSS.t299 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1804 VDD.t468 a_22608_26705.t15 a_25562_24162.t6 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1805 a_14378_9997.t11 a_12598_9997.t14 VDD.t1254 VDD.t1253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1806 a_36697_1856.t1 opcode[1].t48 VDD.t1555 VDD.t1554 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1807 VSS.t175 a_30364_14452.t6 a_38088_23958.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1808 a_n3113_2781.t2 a_n3606_2123.t7 a_n3806_2724.t4 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1809 VSS.t142 a_n3113_13124.t20 a_12698_26780.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1810 a_27657_9997.t9 a_28069_9971.t6 a_27775_9997.t4 VDD.t1131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1811 a_25759_9997.t7 a_20955_6381.t13 VDD.t1775 VDD.t1774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1812 a_14378_9997.t6 a_14790_9971.t5 a_14496_9997.t2 VDD.t641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1813 a_19129_4128.t9 a_14306_12250.t12 VDD.t835 VDD.t834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1814 a_36751_971.t2 a_5623_18852.t11 a_36751_1089.t8 VDD.t635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1815 a_4144_12869.t6 a_1844_12699.t16 VDD.t1457 VDD.t1456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1816 a_20600_4821.t1 a_19247_4128.t14 VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1817 a_25324_4822.t1 a_21746_1762.t17 VDD.t1334 VDD.t1333 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1818 VDD.t1646 a_12475_25767.t10 a_13065_25330.t1 w_12321_25705# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1819 a_n3806_2724.t5 a_n3606_3562.t6 a_n3113_2781.t6 VDD.t1198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1820 a_36751_1089.t4 a_27585_12250.t6 VDD.t498 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1821 a_7749_6382.t3 a_7485_6965.t7 VDD.t797 VDD.t796 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1822 a_19009_18827.t3 a_18952_19520.t11 VDD.t560 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1823 VDD.t1598 a_13051_26980.t6 a_14786_27289.t0 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1824 VDD.t1075 a_4090_5413.t13 a_4145_3835.t3 VDD.t1074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1825 VDD.t1672 a_1836_10114.t14 a_4158_11219.t2 VDD.t1671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1826 VDD.t1971 a_30359_11881.t13 a_33375_14481.t2 VDD.t1970 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1827 a_27340_24456.t3 a_26913_25149.t6 a_27458_24456.t1 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1828 a_18715_18853.t2 a_19009_18827.t6 a_18597_18853.t3 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1829 a_4150_5439.t3 a_4090_5413.t14 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1830 VDD.t2062 a_8508_14599.t17 a_12480_9997.t3 VDD.t2061 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1831 a_25877_9997.t4 a_26171_9971.t7 a_25759_9997.t4 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1832 VDD.t1883 opcode[0].t58 a_n3806_13067.t1 VDD.t1882 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1833 VDD.t578 a_n3111_11055.t20 a_20355_25145.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1834 VSS.t91 a_22608_26705.t16 a_25799_23525.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1835 a_5959_21688.t0 a_5899_21662.t7 VDD.t2327 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1836 VSS.t383 a_15097_1774.t13 a_17579_6451.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1837 a_n3806_6861.t9 a_n3606_7699.t6 a_n3113_6918.t4 VDD.t1604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1838 a_24223_10670.t1 a_23926_11281.t15 a_23986_11307.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1839 VDD.t605 a_15057_14598.t14 a_19134_9929.t5 VDD.t604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1840 a_14660_24431.t1 A[1].t12 VDD.t2170 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1841 a_19549_6960.t2 a_17941_3397.t7 a_19667_6960.t3 VDD.t1339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1842 a_12474_4127.t2 a_8543_1769.t15 VDD.t935 VDD.t934 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1843 a_n3804_15135.t8 B[0].t4 VDD.t1161 VDD.t1160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1844 VSS.t267 a_30359_8848.t12 a_32247_8968.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1845 a_36751_4233.t6 opcode[1].t49 VDD.t1557 VDD.t1556 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1846 VDD.t135 a_36751_16737.t10 Y[2].t1 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1847 a_22095_18533.t0 a_18055_19249.t12 VDD.t2198 w_22001_18497# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1848 a_32011_1857.t3 a_32305_1831.t7 a_31893_1857.t5 VDD.t966 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1849 VDD.t2110 B[5].t18 a_n3608_4192.t1 VDD.t2109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1850 a_6615_12158.t2 a_6351_12741.t8 VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1851 a_36751_4115.t0 a_12181_18848.t11 a_36751_4233.t1 VDD.t2349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1852 a_4735_3398.t2 a_4145_3835.t9 VDD.t2271 VDD.t2270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1853 a_36755_19987.t10 opcode[1].t50 VDD.t1559 VDD.t1558 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1854 a_13961_18848.t1 a_n3113_2781.t18 VDD.t151 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1855 VSS.t52 a_14932_26706.t7 a_15810_27293.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1856 a_36751_13593.t4 a_36697_14478.t7 a_36751_13711.t6 VDD.t1091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1857 VDD.t1410 a_n3113_6918.t19 a_28603_20140.t2 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1858 a_24554_6652.t1 a_23964_7089.t10 VDD.t437 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1859 VSS.t439 a_32011_1857.t11 a_38084_14538.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1860 a_26706_21688.t4 a_27000_21662.t6 a_26571_21032.t1 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1861 a_36751_4115.t4 a_36697_5000.t6 a_36751_4233.t3 VDD.t1132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1862 a_36701_20754.t1 opcode[1].t51 VDD.t1561 VDD.t1560 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1863 VDD.t1885 opcode[0].t59 a_n3808_656.t10 VDD.t1884 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1864 VDD.t803 B[3].t13 a_29769_9285.t4 VDD.t802 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1865 VDD.t1777 a_20955_6381.t14 a_25759_9997.t6 VDD.t1776 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1866 a_21156_1325.t1 B[6].t19 VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1867 a_25464_18124.t1 a_24568_19252.t17 VSS.t178 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1868 a_7821_4129.t2 a_7394_4822.t7 a_7939_4129.t2 VDD.t2287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1869 VSS.t362 a_8508_14599.t18 a_12834_9265.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1870 a_14668_27289.t4 a_13060_23726.t4 VSS.t396 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1871 VDD.t1312 a_6049_9909.t15 a_7402_10602.t3 VDD.t1311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1872 a_15928_27293.t4 a_13065_25330.t6 a_15810_27293.t3 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1873 a_15556_20132.t2 a_n3113_2781.t19 VDD.t1208 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1874 VDD.t561 a_18952_19520.t12 a_19009_18827.t2 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1875 a_8089_23728.t0 a_n3111_15192.t22 a_7853_24460.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1876 a_27649_4129.t9 a_23918_5413.t12 VDD.t2250 VDD.t2249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1877 a_4158_11219.t1 a_1836_10114.t15 VDD.t1674 VDD.t1673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1878 a_33375_14481.t1 a_30359_11881.t14 VDD.t1973 VDD.t1972 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1879 a_27458_24456.t5 a_26913_25149.t7 a_27340_24456.t9 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1880 a_18597_18853.t1 a_19009_18827.t7 a_18715_18853.t0 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1881 a_12382_21028.t3 a_12811_21658.t6 a_12517_21684.t4 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1882 a_30006_8648.t0 A[4].t28 a_29769_9285.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1883 VDD.t2582 a_21150_9929.t19 a_33377_6895.t1 VDD.t2581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1884 VDD.t1887 opcode[0].t60 a_n3604_15973.t2 VDD.t1886 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1885 a_29257_17925.t1 a_24568_19252.t18 VSS.t179 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1886 a_30077_6728.t1 B[4].t15 a_29840_7365.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1887 VDD.t164 a_14366_24457.t13 a_15719_25150.t1 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1888 a_20355_25145.t1 a_n3111_11055.t21 VDD.t579 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1889 VSS.t320 a_20955_6381.t15 a_24223_10670.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1890 a_17351_3834.t6 a_14306_12250.t13 VDD.t837 VDD.t836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1891 VDD.t805 B[3].t14 a_n3606_8329.t2 VDD.t804 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1892 a_32011_6205.t4 a_31466_6898.t7 a_31893_6205.t0 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1893 VSS.t272 a_4963_19248.t19 a_4965_19545.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1894 VDD.t2217 a_15097_1774.t14 a_17356_5438.t1 VDD.t2216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1895 a_24571_9266.t1 a_23981_9703.t10 VDD.t332 VDD.t331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1896 VDD.t807 B[3].t15 a_n3806_8930.t7 VDD.t806 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1897 VDD.t2002 B[4].t16 a_1254_13136.t6 VDD.t2001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1898 VDD.t247 a_8155_27292.t8 a_8419_26709.t0 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1899 VDD.t1209 a_n3113_2781.t20 a_13961_18848.t11 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1900 VSS.t89 a_25877_9997.t13 a_27230_10690.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1901 VDD.t903 a_30364_14452.t7 a_36755_23131.t8 VDD.t902 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1902 a_6041_4129.t5 a_5496_4822.t6 a_5923_4129.t5 VDD.t1655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1903 a_28603_20140.t1 a_n3113_6918.t20 VDD.t1411 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1904 a_n3806_8930.t3 opcode[0].t61 VDD.t1889 VDD.t1888 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1905 a_26571_21032.t2 a_27000_21662.t7 a_26706_21688.t3 w_26477_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1906 a_n3806_6861.t6 B[4].t17 VDD.t2004 VDD.t2003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1907 a_25429_21036.t3 a_25858_21666.t4 a_25564_21692.t5 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1908 a_1243_4513.t0 A[6].t20 VDD.t2487 VDD.t2486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1909 VDD.t1736 a_17296_5412.t15 a_21027_4128.t2 VDD.t1735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1910 VDD.t1116 a_17351_3834.t10 a_17941_3397.t1 VDD.t1115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1911 a_12592_3395.t1 a_12886_4101.t7 VSS.t405 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1912 a_29769_9285.t1 A[4].t29 VDD.t1643 VDD.t1642 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1913 a_7947_9909.t2 a_8241_9883.t7 a_7829_9909.t3 VDD.t327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1914 VDD.t1589 a_21145_4128.t19 a_25751_4129.t10 VDD.t1588 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1915 a_29840_7365.t4 B[4].t18 VDD.t2006 VDD.t2005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1916 a_36751_971.t5 a_36697_1856.t6 a_36751_1089.t2 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1917 VDD.t965 A[7].t6 a_6863_19545.t2 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1918 a_25228_18856.t1 a_25465_19523.t15 a_25464_18124.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1919 a_25562_24162.t1 A[3].t24 VDD.t2357 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1920 VSS.t295 a_13051_26980.t7 a_14668_27289.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1921 a_30434_1013.t0 a_29844_1450.t8 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1922 VDD.t640 a_5948_27420.t9 a_6538_26983.t2 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1923 a_25228_18856.t6 a_24570_19549.t6 a_25110_18856.t10 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1924 a_29252_19529.t0 a_n3113_6918.t21 VSS.t269 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1925 a_15810_27293.t4 a_13065_25330.t7 a_15928_27293.t3 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1926 a_19009_18827.t1 a_18952_19520.t13 VDD.t562 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1927 a_7821_4129.t5 a_4090_5413.t15 VDD.t1079 VDD.t1078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1928 a_30364_14452.t0 a_29774_14889.t8 VSS.t236 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1929 VDD.t1759 a_15810_27293.t8 a_16074_26710.t1 w_15774_27231# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1930 VSS.t136 A[0].t11 a_8089_23728.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1931 a_25429_21036.t0 a_25504_21666.t7 VSS.t87 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1932 a_27340_24456.t10 a_27752_24430.t6 a_27458_24456.t6 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1933 a_n3115_713.t7 opcode[0].t62 a_n2383_949.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1934 a_24201_6452.t1 a_21145_4128.t20 a_23964_7089.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1935 a_4390_8978.t1 a_1844_12699.t17 a_4153_9615.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1936 VDD.t2445 a_n3111_15192.t23 a_7308_25153.t1 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1937 VDD.t2310 a_6966_21028.t7 a_5899_21662.t2 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1938 a_n3113_8987.t2 a_n3606_9768.t6 a_n3806_8930.t10 VDD.t1750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1939 VSS.t326 a_n3113_8987.t21 a_25790_26779.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1940 a_14786_27289.t3 a_13060_23726.t5 a_14668_27289.t3 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1941 VDD.t1141 a_22344_27288.t6 a_22608_26705.t2 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1942 VDD.t2436 a_10641_5411.t16 a_10696_3833.t4 VDD.t2435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1943 VDD.t2359 A[3].t25 a_29840_7365.t0 VDD.t2358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1944 VDD.t2412 a_18991_21663.t6 a_19051_21689.t4 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1945 VDD.t1163 B[0].t5 a_n3604_14534.t2 VDD.t1162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1946 a_17342_7088.t5 a_14306_12250.t14 VDD.t839 VDD.t838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1947 a_1254_13136.t5 B[4].t19 VDD.t2008 VDD.t2007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1948 VSS.t438 a_30430_6928.t15 a_33614_9753.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1949 VDD.t17 B[6].t20 a_29837_4295.t0 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1950 VDD.t2488 A[6].t21 a_15561_18528.t1 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1951 a_1483_9914.t0 B[3].t16 a_1246_10551.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1952 a_5931_9909.t4 a_6343_9883.t6 a_6049_9909.t3 VDD.t432 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1953 VSS.t19 a_13164_12246.t7 a_14042_12833.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1954 VSS.t14 a_18057_19546.t7 a_18715_18121.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1955 a_7485_6965.t3 a_4740_5002.t7 a_7603_6965.t3 VDD.t2288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1956 a_19241_23521.t0 A[2].t12 a_19004_24158.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1957 a_22798_24452.t0 a_22253_25145.t7 a_22798_23720.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1958 a_21032_9929.t9 a_17301_11213.t15 VDD.t2539 VDD.t2538 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1959 a_13051_26980.t1 a_12461_27417.t8 VDD.t205 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1960 a_n2381_2781.t1 a_n3606_3562.t7 a_n3113_2781.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1961 a_33377_2547.t5 a_30434_1013.t13 VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1962 a_36697_1856.t0 opcode[1].t52 VSS.t288 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1963 VDD.t541 a_25877_9997.t14 a_27230_10690.t1 VDD.t540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1964 VDD.t516 a_4098_11193.t17 a_7829_9909.t4 VDD.t515 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1965 a_21145_3396.t1 a_21439_4102.t7 VSS.t292 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1966 a_29774_14889.t6 B[3].t17 VDD.t809 VDD.t808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1967 a_25567_25766.t0 a_n3113_8987.t22 VDD.t1805 w_25413_25704# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1968 a_11286_3396.t1 a_10696_3833.t10 VDD.t698 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1969 a_n3808_656.t7 B[7].t6 VDD.t1279 VDD.t1278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1970 a_n3804_10998.t5 opcode[0].t63 VDD.t1891 VDD.t1890 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1971 a_7403_18852.t8 A[7].t7 VDD.t962 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1972 a_19129_4128.t7 a_18702_4821.t7 a_19247_4128.t5 VDD.t535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1973 a_36755_10391.t0 a_25228_18856.t11 a_36755_10509.t0 VDD.t262 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1974 a_25228_18124.t0 a_25522_18830.t7 a_25228_18856.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1975 VDD.t2219 a_15097_1774.t15 a_17342_7088.t0 VDD.t2218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1976 a_10687_7087.t6 a_7939_4129.t21 VDD.t1110 VDD.t1109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1977 VDD.t469 a_22608_26705.t17 a_25562_24162.t5 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1978 VDD.t1893 opcode[0].t64 a_n3808_4793.t7 VDD.t1892 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1979 a_36755_10509.t1 a_32011_6205.t10 VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1980 a_14932_26706.t2 a_14668_27289.t5 VSS.t97 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1981 a_20782_24452.t7 A[2].t13 VDD.t75 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1982 a_38084_5060.t0 opcode[1].t53 a_36751_4115.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1983 a_6538_26983.t1 a_5948_27420.t10 VDD.t648 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1984 a_25110_18856.t11 a_24570_19549.t7 a_25228_18856.t5 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1985 a_30359_11881.t0 a_29769_12318.t10 VSS.t413 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1986 VSS.t45 a_25858_21666.t5 a_25429_21036.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1987 a_7853_23728.t0 a_8147_24434.t7 VSS.t237 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1988 a_36755_10391.t2 a_36701_11276.t7 a_38088_11100.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1989 a_n3804_15135.t11 opcode[0].t65 VDD.t1895 VDD.t1894 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1990 VSS.t40 a_28024_26705.t7 a_28902_27292.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1991 a_27458_24456.t7 a_27752_24430.t7 a_27340_24456.t11 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1992 a_12892_9971.t1 a_8508_14599.t19 VDD.t2064 VDD.t2063 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1993 a_8508_14599.t3 a_7918_15036.t8 VSS.t187 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1994 a_4373_6452.t0 a_1817_6836.t18 a_4136_7089.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1995 a_14372_4127.t8 a_14784_4101.t7 a_14490_4127.t7 VDD.t1601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1996 VSS.t57 a_17932_6651.t7 a_19549_6960.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1997 VDD.t1952 a_16074_26710.t15 a_19009_25762.t6 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1998 a_25465_19523.t2 a_26468_19549.t7 a_27008_18856.t3 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X1999 a_9561_26713.t2 a_9297_27296.t7 VDD.t320 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2000 VDD.t2252 a_23918_5413.t13 a_23973_3835.t0 VDD.t2251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2001 a_6461_6961.t1 a_4735_3398.t5 a_6343_6961.t3 VDD.t2260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2002 a_38088_20814.t1 opcode[1].t54 a_36755_19869.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2003 a_14668_27289.t2 a_13060_23726.t6 a_14786_27289.t5 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2004 VSS.t154 a_n3606_12466.t6 a_n2381_13124.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2005 VDD.t2361 A[3].t26 a_29774_14889.t0 VDD.t2360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2006 VDD.t1011 a_14668_27289.t6 a_14932_26706.t3 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2007 a_19051_21689.t3 a_18991_21663.t7 VDD.t2411 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2008 a_20907_18827.t3 a_n3115_4850.t19 VDD.t1377 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2009 VDD.t937 a_8543_1769.t16 a_10687_7087.t1 VDD.t936 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2010 a_26913_25149.t1 a_n3113_8987.t23 VDD.t1806 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2011 VDD.t2010 B[4].t20 a_1254_13136.t4 VDD.t2009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2012 a_22680_24452.t9 a_23092_24426.t7 a_22798_24452.t5 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2013 a_18952_19520.t1 a_20907_18827.t5 a_20495_18853.t1 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2014 a_12063_18848.t9 a_11521_19244.t18 VDD.t2589 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2015 a_5948_27420.t4 A[0].t12 VDD.t653 w_5794_27358# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2016 a_14306_12250.t2 a_14042_12833.t5 VSS.t65 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2017 a_18951_18121.t0 a_18055_19249.t13 VSS.t381 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2018 a_27767_4129.t5 a_27222_4822.t7 a_27649_4129.t3 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2019 a_23034_23720.t1 a_20900_24452.t14 a_22798_24452.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2020 VDD.t2112 B[5].t19 a_14507_1337.t5 VDD.t2111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2021 VDD.t2541 a_17301_11213.t16 a_21032_9929.t8 VDD.t2540 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2022 VDD.t543 a_12461_27417.t9 a_13051_26980.t3 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2023 VDD.t1019 a_27458_24456.t13 a_28811_25149.t1 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2024 a_19818_12178.t0 a_19554_12761.t8 VSS.t317 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2025 VDD.t811 B[3].t18 a_29774_14889.t5 VDD.t810 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2026 VDD.t2199 a_18055_19249.t14 a_18057_19546.t3 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2027 VDD.t19 B[6].t21 a_n3606_2123.t1 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2028 VDD.t2362 A[3].t27 a_27752_24430.t1 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2029 a_19246_25125.t1 a_16074_26710.t16 a_19009_25762.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2030 a_27775_9997.t1 a_27230_10690.t6 a_27775_9265.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2031 a_27439_12833.t1 a_24576_10870.t6 a_27321_12833.t4 VDD.t1294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2032 VDD.t719 A[7].t8 a_7403_18852.t7 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2033 a_17946_5001.t0 a_17356_5438.t9 VSS.t308 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2034 a_21439_4102.t1 a_17296_5412.t16 VDD.t1738 VDD.t1737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2035 a_23964_7089.t5 a_21145_4128.t21 VDD.t1591 VDD.t1590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2036 a_25562_24162.t4 a_22608_26705.t18 VDD.t470 w_25408_24100# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2037 a_12480_9997.t8 a_12053_10690.t7 a_12598_9997.t6 VDD.t773 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2038 VDD.t1173 a_28603_20140.t9 a_25858_21666.t1 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2039 VDD.t718 A[2].t14 a_20782_24452.t6 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2040 a_24209_12320.t0 a_21711_14619.t15 a_23972_12957.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2041 a_n3111_11055.t0 a_n3604_10397.t7 a_n3804_10998.t0 VDD.t908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2042 VSS.t367 B[5].t20 a_30006_11681.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2043 a_13953_21654.t2 a_15561_18528.t8 VDD.t280 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2044 VDD.t1953 a_16074_26710.t17 a_19004_24158.t4 w_18850_24096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2045 a_19009_25762.t5 a_16074_26710.t18 VDD.t1954 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2046 a_4963_19248.t3 a_12382_21028.t8 VDD.t781 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2047 a_27008_18856.t9 a_27420_18830.t7 a_25465_19523.t6 w_24534_19487# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2048 VDD.t2028 A[5].t21 a_1227_7273.t4 VDD.t2027 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2049 VSS.t427 A[6].t22 a_8155_14399.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2050 VDD.t58 a_14306_12250.t15 a_19541_4102.t1 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2051 a_17946_9198.t1 a_17356_9635.t10 VDD.t2601 VDD.t2600 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2052 VSS.t302 A[4].t30 a_8190_1769.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2053 a_7953_1332.t1 B[5].t21 VDD.t2114 VDD.t2113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2054 a_36755_7247.t3 a_18715_18853.t11 a_36755_7365.t8 VDD.t1005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2055 a_14786_27289.t4 a_13060_23726.t7 a_14668_27289.t1 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2056 VSS.t194 a_36751_13593.t10 Y[3].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2057 VDD.t1593 a_21145_4128.t22 a_23964_7089.t4 VDD.t1592 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2058 a_30364_14452.t2 a_29774_14889.t9 VDD.t1205 VDD.t1204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2059 a_14932_26706.t1 a_14668_27289.t7 VDD.t188 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2060 a_18916_21033.t2 a_19345_21663.t5 a_19051_21689.t2 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2061 VDD.t1378 a_n3115_4850.t20 a_20907_18827.t2 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2062 a_19546_9903.t3 a_15057_14598.t15 VSS.t204 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2063 a_24215_4802.t0 a_23918_5413.t14 a_23978_5439.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2064 a_20495_18853.t2 a_20907_18827.t6 a_18952_19520.t3 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2065 VDD.t1022 a_28902_27292.t8 a_24568_19252.t1 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2066 VDD.t362 a_26171_6961.t7 a_26435_6378.t1 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2067 a_5931_9909.t2 a_1836_10114.t16 VDD.t1676 VDD.t1675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2068 a_n3804_15135.t0 a_n3604_15973.t7 a_n3111_15192.t7 VDD.t2079 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2069 VDD.t1112 a_7939_4129.t22 a_12474_4127.t8 VDD.t1111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2070 a_13051_26980.t0 a_12461_27417.t10 VDD.t187 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2071 a_19232_26775.t1 A[2].t15 a_18995_27412.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2072 VDD.t302 a_27585_12250.t7 a_36751_1089.t1 VDD.t301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2073 a_29774_14889.t4 B[3].t19 VDD.t813 VDD.t812 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2074 a_18057_19546.t2 a_18055_19249.t15 VDD.t2200 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2075 a_21145_4128.t2 a_20600_4821.t6 a_21027_4128.t4 VDD.t847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2076 VDD.t2018 a_7953_1332.t10 a_8543_1769.t1 VDD.t2017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2077 a_32011_9700.t3 a_31466_10393.t7 a_31893_9700.t3 VDD.t530 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2078 a_27321_12833.t1 a_24576_10870.t7 a_27439_12833.t0 VDD.t287 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2079 VSS.t428 A[6].t23 a_13421_19541.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2080 a_29266_21179.t1 a_n3113_6918.t22 VSS.t270 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2081 a_7403_18852.t6 A[7].t9 VDD.t643 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2082 VDD.t459 B[2].t5 a_n3804_10998.t7 VDD.t458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2083 a_13164_12246.t3 a_12900_12829.t8 VSS.t41 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2084 VSS.t126 a_36751_16737.t11 Y[2].t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2085 a_28603_20140.t0 a_n3113_6918.t23 VDD.t1412 w_28509_20104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2086 VDD.t1148 a_29769_9285.t10 a_30359_8848.t3 VDD.t1147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2087 a_n3806_13067.t9 B[1].t5 VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2088 a_6343_9883.t0 a_1844_12699.t18 VSS.t281 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2089 VSS.t321 a_20955_6381.t16 a_24209_12320.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2090 a_25429_21036.t4 a_25858_21666.t6 a_25564_21692.t4 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2091 a_21156_1325.t0 B[6].t22 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2092 VDD.t281 a_15561_18528.t9 a_13953_21654.t1 w_15467_18492# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2093 a_26297_12829.t5 a_24571_9266.t5 a_26179_12829.t3 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2094 Cout.t3 a_5824_21032.t6 VDD.t333 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2095 VDD.t2221 a_15097_1774.t16 a_17356_5438.t0 VDD.t2220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2096 a_12475_18822.t2 a_12418_19515.t15 VDD.t473 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2097 VSS.t436 a_17301_11213.t17 a_21386_9197.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2098 VDD.t2158 a_14490_4127.t17 a_32305_1831.t2 VDD.t2157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2099 a_36751_13711.t1 a_29356_24456.t9 a_36751_13593.t1 VDD.t845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2100 VDD.t675 a_n3113_13124.t21 a_13821_25150.t2 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2101 VDD.t1563 opcode[1].t55 a_36755_19987.t9 VDD.t1562 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2102 VSS.t163 B[3].t20 a_n3606_8329.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2103 VDD.t1207 a_29774_14889.t10 a_30364_14452.t1 VDD.t1206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2104 VDD.t49 a_14668_27289.t8 a_14932_26706.t0 w_14632_27227# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2105 a_n3808_4793.t0 B[5].t22 VDD.t2116 VDD.t2115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2106 VSS.t68 a_n3606_6260.t7 a_n2381_6918.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2107 a_19051_21689.t1 a_19345_21663.t6 a_18916_21033.t3 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2108 a_36755_19987.t0 a_16264_24457.t11 a_36755_19869.t0 VDD.t1607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2109 a_20907_18827.t1 a_n3115_4850.t21 VDD.t1379 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2110 a_4387_4802.t0 a_4090_5413.t16 a_4150_5439.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2111 a_n3606_13905.t1 opcode[0].t66 VDD.t1897 VDD.t1896 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2112 a_36751_4233.t4 a_36697_5000.t7 a_36751_4115.t3 VDD.t1133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2113 VDD.t377 a_30434_1013.t14 a_31466_2550.t1 VDD.t376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2114 a_19672_12761.t0 a_17946_9198.t7 a_19554_12761.t2 VDD.t2350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2115 a_38084_14302.t0 a_29356_24456.t10 VSS.t166 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2116 a_22739_19526.t1 a_n3115_4850.t22 VSS.t263 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2117 a_7939_4129.t1 a_8233_4103.t7 a_7821_4129.t1 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2118 a_10702_9703.t6 a_10647_11281.t19 VDD.t1195 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2119 VDD.t2029 A[5].t22 a_22104_21787.t5 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2120 VDD.t1678 a_1836_10114.t17 a_5931_9909.t1 VDD.t1677 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2121 a_36697_14478.t1 opcode[1].t56 VDD.t1565 VDD.t1564 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2122 VDD.t1595 a_21145_4128.t23 a_25751_4129.t9 VDD.t1594 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2123 VSS.t11 a_13158_6376.t6 a_14036_6963.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2124 a_n3604_11836.t1 opcode[0].t67 VDD.t1899 VDD.t1898 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2125 a_n2381_6918.t1 a_n3606_7699.t7 a_n3113_6918.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2126 a_29020_27292.t3 a_26157_25329.t7 a_28902_27292.t1 w_28866_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2127 a_32305_1831.t1 a_14490_4127.t18 VDD.t2160 VDD.t2159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2128 VSS.t121 a_n3111_11055.t22 a_19232_26775.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2129 VDD.t939 a_8543_1769.t17 a_10701_5437.t6 VDD.t938 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2130 a_7947_9909.t6 a_7402_10602.t7 a_7947_9177.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2131 VDD.t2489 A[6].t24 a_15570_21782.t2 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2132 VDD.t2201 a_18055_19249.t16 a_18057_19546.t1 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2133 a_12053_10690.t2 a_7749_6382.t17 VDD.t739 VDD.t738 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2134 a_n3604_15973.t3 opcode[0].t68 VDD.t1901 VDD.t1900 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2135 a_28617_21790.t0 A[4].t31 a_29266_21179.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2136 VDD.t1567 opcode[1].t57 a_36755_23131.t9 VDD.t1566 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2137 VSS.t22 a_19955_19546.t7 a_20613_18121.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2138 VDD.t2223 a_15097_1774.t17 a_18702_4821.t2 VDD.t2222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2139 VDD.t1740 a_17296_5412.t17 a_21027_4128.t1 VDD.t1739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2140 a_6343_6961.t2 a_4735_3398.t6 VSS.t388 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2141 a_21358_14419.t0 A[6].t25 a_21121_15056.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2142 a_25564_21692.t3 a_25858_21666.t7 a_25429_21036.t2 w_25335_21047# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2143 a_23926_11281.t2 a_27313_6965.t7 VDD.t1126 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2144 a_19009_18827.t0 a_18952_19520.t14 VSS.t118 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2145 a_26289_6961.t0 a_24563_3398.t7 a_26171_6961.t1 VDD.t536 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2146 a_26179_12829.t1 a_24571_9266.t6 a_26297_12829.t4 VDD.t602 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2147 a_21711_14619.t3 a_21121_15056.t9 VDD.t907 VDD.t906 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2148 a_23978_5439.t2 a_23918_5413.t15 VDD.t2254 VDD.t2253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2149 VDD.t2202 a_18055_19249.t17 a_22090_20137.t1 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2150 a_n3808_4793.t9 a_n3608_5631.t7 a_n3115_4850.t5 VDD.t1313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2151 VSS.t201 a_26435_6378.t6 a_27313_6965.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2152 VSS.t422 a_15570_21782.t10 a_13599_21654.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2153 VDD.t1903 opcode[0].t69 a_n3806_2724.t1 VDD.t1902 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2154 a_17588_3197.t1 a_14306_12250.t16 a_17351_3834.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2155 a_13821_25150.t1 a_n3113_13124.t22 VDD.t676 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2156 a_24218_9066.t0 a_21711_14619.t16 a_23981_9703.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2157 VSS.t110 a_25429_21036.t8 a_18055_19249.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2158 VSS.t147 a_9561_26713.t19 a_16500_23725.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2159 a_36701_8132.t2 opcode[1].t58 VDD.t1569 VDD.t1568 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2160 a_5931_9909.t3 a_6343_9883.t7 a_6049_9909.t4 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2161 a_18916_21033.t0 a_19345_21663.t7 a_19051_21689.t0 w_18822_21044# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2162 VSS.t12 a_13524_21024.t8 a_12457_21658.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2163 VDD.t586 a_6607_6378.t7 a_7603_6965.t0 VDD.t585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2164 VDD.t192 a_17937_12452.t7 a_19672_12761.t3 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2165 a_22090_20137.t0 a_18055_19249.t18 a_22739_19526.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2166 VDD.t1150 a_27313_6965.t8 a_23926_11281.t3 VDD.t1149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2167 a_n3806_13067.t6 a_n3606_12466.t7 a_n3113_13124.t2 VDD.t769 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2168 VDD.t1748 a_32009_13791.t11 a_36751_16855.t2 VDD.t1747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2169 a_5899_21662.t3 a_6966_21028.t8 VDD.t2311 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2170 a_22104_21787.t4 A[5].t23 VDD.t2030 w_22010_21751# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2171 VDD.t457 a_1817_6836.t19 a_5923_4129.t0 VDD.t456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2172 VDD.t2256 a_23918_5413.t16 a_23978_5439.t1 VDD.t2255 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2173 a_5931_9909.t0 a_1836_10114.t18 VDD.t1680 VDD.t1679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2174 a_7815_18826.t1 a_n3115_713.t23 VDD.t1949 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2175 VDD.t1435 a_29837_4295.t10 a_30427_3858.t1 VDD.t1434 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2176 VSS.t24 a_19585_26975.t7 a_21202_27284.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2177 a_9633_24460.t5 a_7853_24460.t13 VDD.t2265 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2178 VSS.t230 a_15561_18528.t10 a_13953_21654.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2179 a_22680_24452.t6 a_20900_24452.t15 VDD.t1418 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2180 a_15570_21782.t1 A[6].t26 VDD.t2490 w_15476_21746# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2181 VDD.t909 A[7].t10 a_9003_18532.t1 w_8909_18496# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2182 a_19252_9929.t1 a_18707_10622.t7 a_19134_9929.t11 VDD.t1297 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2183 VDD.t741 a_7749_6382.t18 a_12053_10690.t1 VDD.t740 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2184 a_n3604_10397.t1 B[2].t6 VDD.t487 VDD.t486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2185 VDD.t714 B[1].t6 a_n3606_12466.t3 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2186 a_n3606_7699.t1 opcode[0].t70 VDD.t1905 VDD.t1904 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2187 a_n3806_8930.t0 a_n3606_8329.t7 a_n3113_8987.t0 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2188 VDD.t1459 a_1844_12699.t19 a_4153_9615.t3 VDD.t1458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2189 a_10045_24434.t0 opcode[0].t71 VSS.t335 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2190 a_36701_8132.t0 opcode[1].t59 VSS.t289 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2191 VDD.t223 a_23973_3835.t10 a_24563_3398.t1 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2192 a_6461_6961.t0 a_4735_3398.t7 a_6343_6961.t1 VDD.t2261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2193 VSS.t181 a_8543_1769.t18 a_12047_4820.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2194 a_23978_5439.t4 a_21746_1762.t18 VDD.t1336 VDD.t1335 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2195 a_32305_1831.t0 a_14490_4127.t19 VSS.t373 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2196 VDD.t961 a_25869_4129.t13 a_27222_4822.t3 VDD.t960 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2197 a_26297_12829.t3 a_24571_9266.t7 a_26179_12829.t0 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2198 VDD.t2031 A[5].t24 a_19955_19546.t2 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2199 VSS.t160 a_6863_19545.t7 a_7521_18120.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2200 a_26171_9971.t0 a_21711_14619.t17 VSS.t10 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2201 a_20955_6381.t1 a_20691_6964.t7 VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2202 VDD.t632 a_36755_19869.t11 Y[1].t1 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2203 VSS.t418 a_10641_5411.t17 a_10933_3196.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2204 a_31893_1857.t2 a_30434_1013.t15 VDD.t404 VDD.t403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2205 VDD.t2122 a_33377_2547.t10 a_17301_11213.t3 VDD.t2121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2206 a_27775_9997.t3 a_27230_10690.t7 a_27657_9997.t0 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2207 a_19134_9929.t9 a_19546_9903.t7 a_19252_9929.t7 VDD.t1269 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2208 a_26143_26979.t3 a_25553_27416.t10 VDD.t927 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2209 a_20900_24452.t1 a_21194_24426.t6 a_20782_24452.t4 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2210 a_16264_23725.t1 a_16558_24431.t7 VSS.t158 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2211 a_14784_4101.t0 a_10641_5411.t18 VSS.t419 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2212 a_14496_9997.t0 a_14790_9971.t6 a_14378_9997.t1 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2213 a_36697_17622.t0 opcode[1].t60 VSS.t290 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2214 a_13524_21024.t4 a_13599_21654.t7 VSS.t297 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2215 a_n3808_656.t11 opcode[0].t72 VDD.t1907 VDD.t1906 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2216 VDD.t514 a_11283_12520.t7 a_13018_12829.t4 VDD.t513 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2217 Y[5].t1 a_36755_7247.t11 VDD.t1287 VDD.t1286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2218 a_19009_25762.t4 a_16074_26710.t19 VDD.t1955 w_18855_25700# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2219 VDD.t356 a_7485_6965.t8 a_7749_6382.t0 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2220 VDD.t1260 a_36751_971.t11 Y[7].t1 VDD.t1259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2221 a_27657_9997.t3 a_25877_9997.t15 VDD.t266 VDD.t265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2222 VDD.t1909 opcode[0].t73 a_n3804_10998.t4 VDD.t1908 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2223 VDD.t841 a_4090_5413.t17 a_4150_5439.t1 VDD.t840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2224 VDD.t986 a_4726_6652.t7 a_6461_6961.t3 VDD.t985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2225 VDD.t1779 a_20955_6381.t17 a_25332_10690.t1 VDD.t1778 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2226 a_13524_21024.t0 a_13953_21654.t7 a_13659_21680.t0 w_13430_21035# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2227 VDD.t118 a_22090_20137.t10 a_19345_21663.t1 w_21996_20101# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2228 a_n3113_8987.t7 opcode[0].t74 a_n2381_9223.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2229 a_20193_21685.t4 a_20133_21659.t6 VDD.t86 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2230 VDD.t349 a_32011_6205.t11 a_36755_10509.t3 VDD.t348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2231 VSS.t244 a_27775_9997.t11 a_38084_5060.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2232 a_11277_6650.t0 a_10687_7087.t10 VSS.t401 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2233 VDD.t2492 A[6].t27 a_21121_15056.t2 VDD.t2491 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2234 VDD.t2266 a_7853_24460.t14 a_9633_24460.t4 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2235 a_20495_18853.t0 a_20907_18827.t7 a_18952_19520.t0 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2236 VSS.t354 B[4].t21 a_1464_6636.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2237 VDD.t85 a_12894_6959.t7 a_13158_6376.t1 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2238 a_9012_21786.t6 A[7].t11 VDD.t910 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2239 a_14378_9997.t2 a_14790_9971.t7 a_14496_9997.t1 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2240 a_19129_4128.t0 a_15097_1774.t18 VDD.t2225 VDD.t2224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2241 VDD.t2494 A[6].t28 a_14507_1337.t0 VDD.t2493 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2242 a_13158_6376.t0 a_12894_6959.t8 VSS.t18 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2243 VDD.t843 a_4090_5413.t18 a_8233_4103.t1 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2244 VSS.t111 B[2].t7 a_n3604_10397.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2245 VDD.t2543 a_17301_11213.t18 a_17361_11239.t5 VDD.t2542 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2246 a_24562_12520.t2 a_23972_12957.t9 VSS.t93 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2247 VSS.t170 a_19247_4128.t15 a_20600_4821.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2248 a_27775_9265.t1 a_28069_9971.t7 VSS.t224 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2249 a_21202_27284.t4 a_19594_23721.t6 a_21320_27284.t1 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2250 a_4150_5439.t6 a_1833_4076.t18 VDD.t1710 VDD.t1709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2251 VDD.t2301 a_6041_4129.t14 a_7394_4822.t1 VDD.t2300 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2252 VDD.t1338 a_21746_1762.t19 a_23964_7089.t0 VDD.t1337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2253 VDD.t51 a_9297_27296.t8 a_9561_26713.t0 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2254 VDD.t65 a_24562_12520.t7 a_26297_12829.t0 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2255 a_19955_19546.t1 A[5].t25 VDD.t2032 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2256 a_25751_4129.t4 a_25324_4822.t6 a_25869_4129.t2 VDD.t430 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2257 VDD.t76 a_9012_21786.t9 a_7041_21658.t2 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2258 a_7757_18120.t1 A[7].t12 VSS.t94 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2259 a_n3606_9768.t3 opcode[0].t75 VSS.t336 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2260 a_17951_10802.t0 a_17361_11239.t10 VSS.t391 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2261 a_28061_4103.t0 a_23918_5413.t17 VSS.t386 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2262 a_22608_26705.t0 a_22344_27288.t7 VSS.t227 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2263 a_20782_24452.t5 a_21194_24426.t7 a_20900_24452.t2 w_20318_25083# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2264 VSS.t234 a_30427_3858.t11 a_31466_6898.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2265 VDD.t2012 B[4].t22 a_1227_7273.t0 VDD.t2011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2266 VDD.t1781 a_20955_6381.t18 a_23986_11307.t0 VDD.t1780 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2267 Cout.t2 a_5824_21032.t7 VDD.t334 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2268 VDD.t587 a_n3113_2781.t21 a_15556_20132.t0 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2269 a_4735_3398.t1 a_4145_3835.t10 VDD.t2273 VDD.t2272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2270 a_14726_3395.t0 a_12592_4127.t15 a_14490_4127.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2271 a_1480_3876.t1 B[3].t21 a_1243_4513.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2272 VDD.t1236 a_23926_11281.t16 a_27657_9997.t8 VDD.t1235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2273 VDD.t97 a_15057_14598.t16 a_19546_9903.t1 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2274 a_12598_9997.t0 a_12892_9971.t7 a_12480_9997.t0 VDD.t626 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2275 a_6547_23729.t0 a_5957_24166.t10 VSS.t322 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2276 VDD.t566 a_25869_4129.t14 a_27649_4129.t8 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2277 a_25869_4129.t1 a_25324_4822.t7 a_25751_4129.t0 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2278 VDD.t33 a_13158_6376.t7 a_14154_6963.t0 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2279 VDD.t87 a_20133_21659.t7 a_20193_21685.t3 w_19964_21040# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2280 VSS.t311 a_1833_4076.t19 a_5496_4822.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2281 a_20696_12765.t4 a_17951_10802.t7 VSS.t199 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2282 a_6194_23529.t1 A[0].t13 a_5957_24166.t4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2283 a_33377_10390.t4 a_30359_8848.t13 VDD.t1396 VDD.t1395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2284 VSS.t176 a_20487_21659.t7 a_20058_21029.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2285 a_n3606_8329.t1 B[3].t22 VDD.t815 VDD.t814 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2286 a_21121_15056.t1 A[6].t29 VDD.t2496 VDD.t2495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2287 a_9633_24460.t3 a_7853_24460.t15 VDD.t2267 w_7271_25091# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2288 VSS.t103 a_14366_24457.t14 a_15719_25150.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2289 VDD.t644 A[7].t13 a_9012_21786.t5 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2290 a_18597_18853.t10 a_18952_19520.t15 VDD.t563 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2291 VDD.t60 a_14306_12250.t17 a_17351_3834.t1 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2292 VSS.t15 a_14306_12250.t18 a_19483_3396.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2293 VDD.t417 a_15057_14598.t17 a_17347_12889.t5 VDD.t416 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2294 VSS.t53 a_21711_14619.t18 a_26113_9265.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2295 VDD.t369 a_21711_14619.t19 a_23981_9703.t3 VDD.t368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2296 a_21156_1325.t4 A[5].t26 VDD.t2034 VDD.t2033 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2297 a_26435_6378.t0 a_26171_6961.t8 VSS.t16 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2298 VDD.t580 a_n3111_11055.t23 a_18995_27412.t0 w_18841_27350# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2299 a_17361_11239.t4 a_17301_11213.t19 VDD.t2545 VDD.t2544 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2300 a_29356_24456.t3 a_28811_25149.t7 a_29356_23724.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2301 a_21145_4128.t3 a_20600_4821.t7 a_21027_4128.t5 VDD.t848 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2302 a_32011_9700.t6 a_32305_9674.t7 a_31893_9700.t6 VDD.t950 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2303 a_36751_971.t6 a_36697_1856.t7 a_36751_1089.t3 VDD.t412 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2304 a_8273_27292.t3 a_6547_23729.t7 a_8155_27292.t1 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2305 VDD.t5 a_27767_4129.t11 a_36755_7365.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2306 a_21320_27284.t0 a_19594_23721.t7 a_21202_27284.t2 w_21166_27222# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2307 a_n3111_11055.t7 a_n3604_11836.t7 a_n3804_10998.t11 VDD.t821 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2308 a_27431_6965.t1 a_24568_5002.t7 a_27313_6965.t1 VDD.t1057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2309 a_14467_15035.t6 A[5].t27 VDD.t2036 VDD.t2035 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2310 VDD.t1177 a_30427_3858.t12 a_33377_6895.t5 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2311 VSS.t233 a_28603_20140.t10 a_25858_21666.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2312 a_n3806_13067.t0 a_n3606_13905.t7 a_n3113_13124.t0 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2313 a_7041_21658.t1 a_9012_21786.t10 VDD.t77 w_8918_21750# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2314 a_14366_24457.t0 a_13821_25150.t7 a_14366_23725.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2315 VDD.t304 a_14042_12833.t6 a_14306_12250.t1 VDD.t303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2316 VSS.t203 a_27458_24456.t14 a_28811_25149.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2317 a_17351_3834.t2 a_17296_5412.t18 VDD.t1742 VDD.t1741 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2318 a_12592_4127.t7 a_12047_4820.t7 a_12592_3395.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2319 VDD.t1783 a_20955_6381.t19 a_23972_12957.t4 VDD.t1782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2320 a_23981_9703.t4 a_23926_11281.t17 VDD.t1238 VDD.t1237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2321 a_12461_27417.t1 A[1].t13 VDD.t2171 w_12307_27355# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2322 a_6863_19545.t0 A[7].t14 VDD.t451 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2323 VDD.t2364 A[3].t28 a_29844_1450.t0 VDD.t2363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2324 a_n3111_15192.t2 a_n3604_14534.t7 a_n3804_15135.t5 VDD.t944 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2325 a_24576_10870.t3 a_23986_11307.t8 VDD.t492 VDD.t491 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2326 VDD.t2498 A[6].t30 a_7918_15036.t0 VDD.t2497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2327 VDD.t335 a_5824_21032.t8 Cout.t1 w_5730_21043# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2328 a_20907_18827.t0 a_n3115_4850.t23 VSS.t264 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2329 a_15556_20132.t1 a_n3113_2781.t22 VDD.t588 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2330 a_5917_18826.t1 a_5860_19519.t14 VDD.t2593 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2331 a_21439_4102.t0 a_17296_5412.t19 VSS.t315 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2332 a_28003_3397.t0 a_25869_4129.t15 a_27767_4129.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2333 a_5623_18852.t5 a_5917_18826.t6 a_5505_18852.t4 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2334 a_27657_9997.t7 a_23926_11281.t18 VDD.t1128 VDD.t1127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2335 a_19546_9903.t2 a_15057_14598.t18 VDD.t358 VDD.t357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2336 a_23918_5413.t3 a_33377_6895.t10 VDD.t1167 VDD.t1166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2337 a_12382_21028.t2 a_12811_21658.t7 a_12517_21684.t3 w_12288_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2338 a_6041_4129.t6 a_5496_4822.t7 a_5923_4129.t4 VDD.t1656 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2339 VSS.t58 a_12598_9997.t15 a_13951_10690.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2340 a_4726_6652.t1 a_4136_7089.t10 VDD.t1202 VDD.t1201 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2341 VDD.t850 a_26435_6378.t7 a_27431_6965.t4 VDD.t849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2342 a_14784_4101.t1 a_10641_5411.t19 VDD.t2438 VDD.t2437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2343 a_n3806_8930.t9 a_n3606_9768.t7 a_n3113_8987.t3 VDD.t1749 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2344 a_14744_1774.t0 B[5].t23 a_14507_1337.t6 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2345 VSS.t312 a_19818_12178.t7 a_20696_12765.t3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2346 VSS.t337 opcode[0].t76 a_6194_23529.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2347 a_31466_6898.t1 a_30427_3858.t13 VDD.t1179 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2348 VDD.t1398 a_30359_8848.t14 a_33377_10390.t5 VDD.t1397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2349 a_22462_27288.t0 a_19599_25325.t7 a_22344_27288.t1 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2350 a_22095_18533.t3 A[5].t28 a_22744_17922.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2351 a_10696_3833.t1 a_7939_4129.t23 VDD.t1114 VDD.t1113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2352 VDD.t2227 a_15097_1774.t19 a_18702_4821.t1 VDD.t2226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2353 a_31893_6205.t5 a_32305_6179.t7 a_32011_6205.t0 VDD.t231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2354 a_17946_5001.t1 a_17356_5438.t10 VDD.t1712 VDD.t1711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2355 a_17347_12889.t4 a_15057_14598.t19 VDD.t186 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2356 a_n3604_14534.t1 B[0].t6 VDD.t775 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2357 a_n2381_3017.t1 B[6].t23 VSS.t2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2358 a_6607_6378.t0 a_6343_6961.t8 VSS.t138 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2359 a_20691_6964.t3 a_17946_5001.t7 a_20809_6964.t2 VDD.t905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2360 a_32303_13765.t0 a_30359_11881.t15 VSS.t350 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2361 VDD.t214 a_7041_21658.t6 a_7101_21684.t4 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2362 a_30434_1013.t2 a_29844_1450.t9 VDD.t314 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2363 VDD.t922 a_24568_19252.t19 a_28608_18536.t2 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2364 VDD.t1085 a_19549_6960.t8 a_19813_6377.t3 VDD.t1084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2365 a_25553_27416.t1 A[3].t29 VDD.t2365 w_25399_27354# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2366 VSS.t387 a_23918_5413.t18 a_28003_3397.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2367 VDD.t992 a_4098_11193.t18 a_8241_9883.t1 VDD.t991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2368 VDD.t2388 a_14496_9997.t21 a_17361_11239.t1 VDD.t2387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2369 VSS.t355 B[4].t23 a_1491_12499.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2370 a_29592_23724.t1 a_27458_24456.t15 a_29356_24456.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2371 a_15561_18528.t0 A[6].t31 a_16210_17917.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2372 a_7821_4129.t9 a_6041_4129.t15 VDD.t2303 VDD.t2302 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2373 a_36751_13593.t0 a_29356_24456.t11 a_36751_13711.t2 VDD.t846 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2374 VDD.t2283 a_5962_25770.t9 a_6552_25333.t2 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2375 a_21711_14619.t2 a_21121_15056.t10 VSS.t76 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2376 VDD.t282 a_6538_26983.t6 a_8273_27292.t1 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2377 a_30434_1013.t1 a_29844_1450.t10 VSS.t27 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2378 a_5923_4129.t3 a_6335_4103.t7 a_6041_4129.t2 VDD.t789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2379 VDD.t2038 A[5].t29 a_14467_15035.t5 VDD.t2037 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2380 a_14602_23725.t1 a_n3113_13124.t23 a_14366_24457.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2381 VDD.t1281 B[7].t7 a_n3808_656.t8 VDD.t1280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2382 a_14306_12250.t0 a_14042_12833.t7 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2383 a_26289_6961.t3 a_24554_6652.t7 VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2384 VDD.t2366 A[3].t30 a_27340_24456.t0 w_26876_25087# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2385 a_6285_9177.t0 a_1836_10114.t19 a_6049_9909.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2386 a_24562_12520.t1 a_23972_12957.t10 VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2387 VDD.t752 a_4734_12432.t7 a_6469_12741.t3 VDD.t751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2388 a_n3808_4793.t6 opcode[0].t77 VDD.t1911 VDD.t1910 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2389 a_17342_7088.t4 a_14306_12250.t19 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2390 VDD.t654 A[0].t14 a_5957_24166.t5 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2391 VDD.t1314 A[7].t15 a_6863_19545.t3 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2392 VDD.t494 a_23986_11307.t9 a_24576_10870.t2 VDD.t493 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2393 a_8508_14599.t2 a_7918_15036.t9 VDD.t351 VDD.t350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2394 VDD.t2585 a_11521_19244.t19 a_15556_20132.t4 w_15462_20096# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2395 VDD.t2592 a_5860_19519.t15 a_5917_18826.t0 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2396 a_5505_18852.t3 a_5917_18826.t7 a_5623_18852.t4 w_4929_19483# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2397 VDD.t1130 a_23926_11281.t19 a_27657_9997.t6 VDD.t1129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2398 a_28061_4103.t1 a_23918_5413.t19 VDD.t2258 VDD.t2257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2399 a_16146_24457.t2 a_14366_24457.t15 VDD.t360 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2400 a_n3115_713.t6 a_n3608_1494.t7 a_n3808_656.t5 VDD.t784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2401 VDD.t2399 a_8419_26709.t7 a_9415_27296.t0 w_9261_27234# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2402 a_29769_12318.t1 A[3].t31 VDD.t2368 VDD.t2367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2403 VDD.t2414 a_21466_26701.t7 a_22462_27288.t3 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2404 a_33377_10390.t6 a_30359_8848.t15 VDD.t1400 VDD.t1399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2405 a_n2381_13360.t1 B[1].t7 VSS.t146 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2406 a_36751_16737.t3 a_36697_17622.t7 a_36751_16855.t11 VDD.t1224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2407 VDD.t1142 a_22344_27288.t8 a_22608_26705.t1 w_22308_27226# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2408 a_16219_21171.t1 a_n3113_2781.t23 VSS.t248 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2409 a_12063_18848.t5 a_11523_19541.t7 a_12181_18848.t1 w_11487_19479# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2410 VDD.t2317 a_11277_6650.t7 a_13012_6959.t0 VDD.t2316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2411 VDD.t977 a_4098_11193.t19 a_4153_9615.t6 VDD.t976 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2412 VDD.t1365 a_7493_12745.t8 a_4090_5413.t1 VDD.t1364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2413 VDD.t2390 a_14496_9997.t22 a_17347_12889.t0 VDD.t2389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2414 VDD.t597 a_17342_7088.t10 a_17932_6651.t1 VDD.t596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2415 a_36701_11276.t0 opcode[1].t61 VSS.t291 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2416 a_7101_21684.t0 a_7041_21658.t7 VDD.t24 w_6872_21039# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2417 VSS.t155 B[0].t7 a_n3604_14534.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2418 a_36755_23013.t3 a_36701_23898.t7 a_36755_23131.t6 VDD.t861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2419 VSS.t165 a_4090_5413.t19 a_8175_3397.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2420 VDD.t1913 opcode[0].t78 a_n3806_6861.t0 VDD.t1912 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2421 a_17361_11239.t0 a_14496_9997.t23 VDD.t2392 VDD.t2391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2422 VSS.t92 a_22608_26705.t19 a_29592_23724.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2423 a_6552_25333.t1 a_5962_25770.t10 VDD.t2284 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2424 a_32247_5473.t1 a_30427_3858.t14 a_32011_6205.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2425 VDD.t2203 a_18055_19249.t19 a_18597_18853.t4 w_18021_19484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2426 VSS.t358 A[5].t30 a_21393_1762.t1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2427 a_31893_6205.t1 a_30427_3858.t15 VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2428 VDD.t988 a_36751_13593.t11 Y[3].t1 VDD.t987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2429 a_8273_27292.t0 a_6538_26983.t7 VDD.t190 w_8119_27230# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2430 VDD.t111 a_20696_12765.t8 a_17296_5412.t1 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2431 VDD.t1571 opcode[1].t62 a_36701_8132.t1 VDD.t1570 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2432 a_31891_13791.t3 a_7947_9909.t19 VDD.t2192 VDD.t2191 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2433 VDD.t2172 A[1].t14 a_14248_24457.t0 w_13784_25088# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2434 VDD.t743 a_7749_6382.t19 a_10707_11307.t0 VDD.t742 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2435 a_14467_15035.t4 A[5].t31 VDD.t2040 VDD.t2039 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2436 a_20955_6381.t2 a_20691_6964.t8 VSS.t69 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2437 VDD.t1976 a_28608_18536.t10 a_27000_21662.t1 w_28514_18500# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2438 a_n3806_8930.t6 B[3].t23 VDD.t817 VDD.t816 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2439 VSS.t375 A[1].t15 a_14602_23725.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2440 a_38084_1916.t1 opcode[1].t63 a_36751_971.t7 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2441 VDD.t480 a_14042_12833.t8 a_14306_12250.t3 VDD.t479 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2442 VDD.t941 a_8543_1769.t19 a_10687_7087.t2 VDD.t940 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2443 a_5957_24166.t6 A[0].t15 VDD.t655 w_5803_24104# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2444 a_25877_9997.t1 a_25332_10690.t7 a_25759_9997.t0 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X2445 VDD.t1914 opcode[0].t79 a_5962_25770.t6 w_5808_25708# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2446 a_24576_10870.t1 a_23986_11307.t10 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2447 VDD.t47 a_7918_15036.t10 a_8508_14599.t0 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
R0 a_4963_19248.n6 a_4963_19248.n5 501.28
R1 a_4963_19248.t5 a_4963_19248.t4 437.233
R2 a_4963_19248.t15 a_4963_19248.t18 415.315
R3 a_4963_19248.t14 a_4963_19248.n3 313.873
R4 a_4963_19248.n5 a_4963_19248.t13 294.986
R5 a_4963_19248.n2 a_4963_19248.t12 272.288
R6 a_4963_19248.n6 a_4963_19248.t9 236.009
R7 a_4963_19248.n9 a_4963_19248.t5 216.627
R8 a_4963_19248.n7 a_4963_19248.t15 216.111
R9 a_4963_19248.n8 a_4963_19248.t8 214.686
R10 a_4963_19248.t4 a_4963_19248.n8 214.686
R11 a_4963_19248.n1 a_4963_19248.t16 214.335
R12 a_4963_19248.t18 a_4963_19248.n1 214.335
R13 a_4963_19248.n4 a_4963_19248.t7 190.152
R14 a_4963_19248.n4 a_4963_19248.t14 190.152
R15 a_4963_19248.n2 a_4963_19248.t11 160.666
R16 a_4963_19248.n3 a_4963_19248.t10 160.666
R17 a_4963_19248.n7 a_4963_19248.n6 148.428
R18 a_4963_19248.n5 a_4963_19248.t19 110.859
R19 a_4963_19248.n3 a_4963_19248.n2 96.129
R20 a_4963_19248.n8 a_4963_19248.t6 80.333
R21 a_4963_19248.n1 a_4963_19248.t17 80.333
R22 a_4963_19248.t9 a_4963_19248.n4 80.333
R23 a_4963_19248.n0 a_4963_19248.t3 28.57
R24 a_4963_19248.n11 a_4963_19248.t2 28.565
R25 a_4963_19248.t1 a_4963_19248.n11 28.565
R26 a_4963_19248.n0 a_4963_19248.t0 17.638
R27 a_4963_19248.n10 a_4963_19248.n9 5.638
R28 a_4963_19248.n9 a_4963_19248.n7 2.923
R29 a_4963_19248.n11 a_4963_19248.n10 0.693
R30 a_4963_19248.n10 a_4963_19248.n0 0.597
R31 a_8998_20136.n0 a_8998_20136.t7 214.335
R32 a_8998_20136.t9 a_8998_20136.n0 214.335
R33 a_8998_20136.n1 a_8998_20136.t9 143.851
R34 a_8998_20136.n1 a_8998_20136.t10 135.658
R35 a_8998_20136.n0 a_8998_20136.t8 80.333
R36 a_8998_20136.n2 a_8998_20136.t5 28.565
R37 a_8998_20136.n2 a_8998_20136.t4 28.565
R38 a_8998_20136.n4 a_8998_20136.t3 28.565
R39 a_8998_20136.n4 a_8998_20136.t6 28.565
R40 a_8998_20136.t1 a_8998_20136.n7 28.565
R41 a_8998_20136.n7 a_8998_20136.t2 28.565
R42 a_8998_20136.n6 a_8998_20136.t0 9.714
R43 a_8998_20136.n7 a_8998_20136.n6 1.003
R44 a_8998_20136.n5 a_8998_20136.n3 0.833
R45 a_8998_20136.n3 a_8998_20136.n2 0.653
R46 a_8998_20136.n5 a_8998_20136.n4 0.653
R47 a_8998_20136.n6 a_8998_20136.n5 0.341
R48 a_8998_20136.n3 a_8998_20136.n1 0.032
R49 VDD.t2347 VDD.t532 95474.9
R50 VDD.t508 VDD.t1282 95474.9
R51 VDD.t982 VDD.t958 95474.9
R52 VDD.t845 VDD.t121 95474.9
R53 VDD.t1010 VDD.t132 95474.9
R54 VDD.t1606 VDD.t629 95474.9
R55 VDD.t967 VDD.t1936 95474.9
R56 VDD.t634 VDD.t1259 95474.9
R57 VDD.t1436 VDD.t1450 2079.61
R58 VDD.t2049 VDD.t2055 2079.61
R59 VDD.t54 VDD.t604 2079.61
R60 VDD.t399 VDD.t997 2079.61
R61 VDD.t1578 VDD.t1594 2079.61
R62 VDD.t830 VDD.t828 2079.61
R63 VDD.t1041 VDD.t1111 2079.61
R64 VDD.t454 VDD.t456 2079.61
R65 VDD.n1064 VDD.n1063 1412.62
R66 VDD.n726 VDD.n725 1412.62
R67 VDD.n869 VDD.n868 1412.59
R68 VDD.n503 VDD.n491 1408.41
R69 VDD.n555 VDD.n554 1404.25
R70 VDD.n937 VDD.n936 1239.11
R71 VDD.n638 VDD.n637 1235.85
R72 VDD.n1000 VDD.n999 1235.85
R73 VDD.n971 VDD.n970 1033.17
R74 VDD.n618 VDD.n612 1033.13
R75 VDD.n737 VDD.n731 1033.13
R76 VDD.n694 VDD.n693 1033.13
R77 VDD.n469 VDD.n468 1033.13
R78 VDD.n760 VDD.n754 1033.12
R79 VDD.n902 VDD.n901 1029.24
R80 VDD.n603 VDD.n599 1029.22
R81 VDD.n1038 VDD.n1037 1029.21
R82 VDD.n1172 VDD.n1171 1029.21
R83 VDD.n841 VDD.n840 1025.33
R84 VDD.n456 VDD.n452 1025.3
R85 VDD.t1311 VDD.t1452 999.845
R86 VDD.t1247 VDD.t2063 999.845
R87 VDD.t179 VDD.t357 999.845
R88 VDD.t540 VDD.t216 999.845
R89 VDD.t960 VDD.t1580 999.845
R90 VDD.t870 VDD.t822 999.845
R91 VDD.t2334 VDD.t1107 999.845
R92 VDD.t2300 VDD.t1342 999.845
R93 VDD.n979 VDD.n973 880.922
R94 VDD.n1031 VDD.n1030 874.899
R95 VDD.n681 VDD.n675 874.857
R96 VDD.n526 VDD.n522 874.804
R97 VDD.n1196 VDD.n1195 871.829
R98 VDD.n1695 VDD.n1694 871.827
R99 VDD.n642 VDD.n641 871.827
R100 VDD.n1107 VDD.n1101 871.811
R101 VDD.n849 VDD.n843 871.81
R102 VDD.n914 VDD.n909 871.809
R103 VDD.n1142 VDD.n1141 871.808
R104 VDD.n535 VDD.n534 871.808
R105 VDD.n1147 VDD.n1146 809.201
R106 VDD.n656 VDD.n655 805.926
R107 VDD.n1710 VDD.n1709 805.926
R108 VDD.n768 VDD.n767 805.925
R109 VDD.n1210 VDD.n1209 802.65
R110 VDD.n1178 VDD.n1177 687.118
R111 VDD.n1116 VDD.n1114 687.068
R112 VDD.n743 VDD.n741 684.693
R113 VDD.n1254 VDD.n1253 600.209
R114 VDD.n1391 VDD.n1390 600.209
R115 VDD.n1240 VDD.n1239 600.207
R116 VDD.n399 VDD.n398 600.207
R117 VDD.t1278 VDD.t1276 541.402
R118 VDD.t755 VDD.t18 541.402
R119 VDD.t2115 VDD.t2109 541.402
R120 VDD.t1983 VDD.t1979 541.402
R121 VDD.t1466 VDD.t798 541.402
R122 VDD.t242 VDD.t224 541.402
R123 VDD.t703 VDD.t713 541.402
R124 VDD.t1160 VDD.t1154 541.402
R125 VDD.n1094 VDD.n1093 491.958
R126 VDD.n1702 VDD.t1362 479.013
R127 VDD.n665 VDD.t68 479.01
R128 VDD.n748 VDD.t25 479.007
R129 VDD.n1128 VDD.t796 479.006
R130 VDD.n1159 VDD.t88 479.006
R131 VDD.n1188 VDD.t162 479.006
R132 VDD.n773 VDD.t325 424.731
R133 VDD.t143 VDD.t127 422.41
R134 VDD.t418 VDD.t792 422.41
R135 VDD.t2540 VDD.t2526 422.41
R136 VDD.t1129 VDD.t1261 422.41
R137 VDD.t2243 VDD.t2257 422.41
R138 VDD.t1739 VDD.t1727 422.41
R139 VDD.t2427 VDD.t2437 422.41
R140 VDD.t1068 VDD.t611 422.41
R141 VDD.n1217 VDD.t1125 422.371
R142 VDD.t2149 VDD.t2159 394.32
R143 VDD.t2565 VDD.t2579 394.32
R144 VDD.t1395 VDD.t1387 394.32
R145 VDD.t1968 VDD.t1966 394.32
R146 VDD.t1243 VDD.t1502 382.217
R147 VDD.t4 VDD.t1568 382.217
R148 VDD.t348 VDD.t1496 382.217
R149 VDD.t2556 VDD.t1514 382.217
R150 VDD.t1747 VDD.t1484 382.217
R151 VDD.t556 VDD.t1560 382.217
R152 VDD.t900 VDD.t1504 382.217
R153 VDD.t301 VDD.t1554 382.217
R154 VDD.t2153 VDD.t2145 352.102
R155 VDD.t2567 VDD.t2575 352.102
R156 VDD.t1393 VDD.t1389 352.102
R157 VDD.t1964 VDD.t1958 352.102
R158 VDD.t1649 VDD.t1651 345.987
R159 VDD.t1647 VDD.t1649 345.987
R160 VDD.t1663 VDD.t1647 345.987
R161 VDD.t1659 VDD.t1663 345.987
R162 VDD.t1657 VDD.t1456 345.987
R163 VDD.t1456 VDD.t1454 345.987
R164 VDD.t1454 VDD.t1444 345.987
R165 VDD.t1817 VDD.t1861 345.987
R166 VDD.t1880 VDD.t1817 345.987
R167 VDD.t1276 VDD.t1274 345.987
R168 VDD.t1274 VDD.t1270 345.987
R169 VDD.t1857 VDD.t1867 345.987
R170 VDD.t1811 VDD.t1857 345.987
R171 VDD.t18 VDD.t428 345.987
R172 VDD.t428 VDD.t422 345.987
R173 VDD.t1819 VDD.t1837 345.987
R174 VDD.t1808 VDD.t1819 345.987
R175 VDD.t2109 VDD.t2097 345.987
R176 VDD.t2097 VDD.t2087 345.987
R177 VDD.t1859 VDD.t1904 345.987
R178 VDD.t1815 VDD.t1859 345.987
R179 VDD.t1979 VDD.t1999 345.987
R180 VDD.t1999 VDD.t1987 345.987
R181 VDD.t1876 VDD.t1813 345.987
R182 VDD.t1840 VDD.t1876 345.987
R183 VDD.t798 VDD.t814 345.987
R184 VDD.t814 VDD.t804 345.987
R185 VDD.t1871 VDD.t1898 345.987
R186 VDD.t1830 VDD.t1871 345.987
R187 VDD.t224 VDD.t486 345.987
R188 VDD.t486 VDD.t606 345.987
R189 VDD.t1832 VDD.t1878 345.987
R190 VDD.t1896 VDD.t1832 345.987
R191 VDD.t713 VDD.t709 345.987
R192 VDD.t709 VDD.t705 345.987
R193 VDD.t1886 VDD.t1900 345.987
R194 VDD.t1845 VDD.t1886 345.987
R195 VDD.t1154 VDD.t774 345.987
R196 VDD.t774 VDD.t1162 345.987
R197 VDD.t1220 VDD.t1199 345.987
R198 VDD.t1201 VDD.t1220 345.987
R199 VDD.t1695 VDD.t1201 345.987
R200 VDD.t1703 VDD.t1695 345.987
R201 VDD.t1691 VDD.t1356 345.987
R202 VDD.t1356 VDD.t1344 345.987
R203 VDD.t1344 VDD.t1352 345.987
R204 VDD.t2321 VDD.t2319 345.987
R205 VDD.t2323 VDD.t2321 345.987
R206 VDD.t940 VDD.t2323 345.987
R207 VDD.t687 VDD.t940 345.987
R208 VDD.t936 VDD.t1037 345.987
R209 VDD.t1037 VDD.t1103 345.987
R210 VDD.t1103 VDD.t1109 345.987
R211 VDD.t596 VDD.t594 345.987
R212 VDD.t592 VDD.t596 345.987
R213 VDD.t2218 VDD.t592 345.987
R214 VDD.t2204 VDD.t2218 345.987
R215 VDD.t2212 VDD.t838 345.987
R216 VDD.t838 VDD.t826 345.987
R217 VDD.t826 VDD.t61 345.987
R218 VDD.t370 VDD.t436 345.987
R219 VDD.t318 VDD.t370 345.987
R220 VDD.t1323 VDD.t318 345.987
R221 VDD.t1329 VDD.t1323 345.987
R222 VDD.t1337 VDD.t1582 345.987
R223 VDD.t1582 VDD.t1592 345.987
R224 VDD.t1592 VDD.t1590 345.987
R225 VDD.t2017 VDD.t2015 345.987
R226 VDD.t2013 VDD.t2017 345.987
R227 VDD.t1608 VDD.t2013 345.987
R228 VDD.t1625 VDD.t1608 345.987
R229 VDD.t1638 VDD.t2083 345.987
R230 VDD.t2083 VDD.t2105 345.987
R231 VDD.t2105 VDD.t2113 345.987
R232 VDD.t495 VDD.t245 345.987
R233 VDD.t372 VDD.t495 345.987
R234 VDD.t1782 VDD.t372 345.987
R235 VDD.t1772 VDD.t1782 345.987
R236 VDD.t1768 VDD.t381 345.987
R237 VDD.t381 VDD.t385 345.987
R238 VDD.t385 VDD.t383 345.987
R239 VDD.t165 VDD.t226 345.987
R240 VDD.t481 VDD.t165 345.987
R241 VDD.t2379 VDD.t481 345.987
R242 VDD.t2377 VDD.t2379 345.987
R243 VDD.t2389 VDD.t185 345.987
R244 VDD.t185 VDD.t416 345.987
R245 VDD.t416 VDD.t22 345.987
R246 VDD.t2021 VDD.t2023 345.987
R247 VDD.t2019 VDD.t2021 345.987
R248 VDD.t730 VDD.t2019 345.987
R249 VDD.t726 VDD.t730 345.987
R250 VDD.t720 VDD.t2041 345.987
R251 VDD.t2041 VDD.t2059 345.987
R252 VDD.t2059 VDD.t2057 345.987
R253 VDD.t1303 VDD.t1301 345.987
R254 VDD.t1301 VDD.t1311 345.987
R255 VDD.t1452 VDD.t1440 345.987
R256 VDD.t1440 VDD.t1436 345.987
R257 VDD.t991 VDD.t699 345.987
R258 VDD.t127 VDD.t991 345.987
R259 VDD.t1027 VDD.t1023 345.987
R260 VDD.t1025 VDD.t1027 345.987
R261 VDD.t1661 VDD.t1025 345.987
R262 VDD.t1673 VDD.t1661 345.987
R263 VDD.t1671 VDD.t366 345.987
R264 VDD.t366 VDD.t1002 345.987
R265 VDD.t1002 VDD.t296 345.987
R266 VDD.t401 VDD.t145 345.987
R267 VDD.t677 VDD.t401 345.987
R268 VDD.t924 VDD.t677 345.987
R269 VDD.t461 VDD.t924 345.987
R270 VDD.t976 VDD.t1442 345.987
R271 VDD.t1442 VDD.t1458 345.987
R272 VDD.t1458 VDD.t1446 345.987
R273 VDD.t1251 VDD.t1249 345.987
R274 VDD.t1249 VDD.t1247 345.987
R275 VDD.t2063 VDD.t2051 345.987
R276 VDD.t2051 VDD.t2049 345.987
R277 VDD.t196 VDD.t198 345.987
R278 VDD.t792 VDD.t196 345.987
R279 VDD.t378 VDD.t434 345.987
R280 VDD.t158 VDD.t378 345.987
R281 VDD.t728 VDD.t158 345.987
R282 VDD.t724 VDD.t728 345.987
R283 VDD.t742 VDD.t1192 345.987
R284 VDD.t1192 VDD.t1190 345.987
R285 VDD.t1190 VDD.t1188 345.987
R286 VDD.t1052 VDD.t1050 345.987
R287 VDD.t1048 VDD.t1052 345.987
R288 VDD.t200 VDD.t1048 345.987
R289 VDD.t1194 VDD.t200 345.987
R290 VDD.t790 VDD.t2047 345.987
R291 VDD.t2047 VDD.t2043 345.987
R292 VDD.t2043 VDD.t2045 345.987
R293 VDD.t183 VDD.t181 345.987
R294 VDD.t181 VDD.t179 345.987
R295 VDD.t357 VDD.t96 345.987
R296 VDD.t96 VDD.t54 345.987
R297 VDD.t2532 VDD.t2534 345.987
R298 VDD.t2526 VDD.t2532 345.987
R299 VDD.t2278 VDD.t2280 345.987
R300 VDD.t2276 VDD.t2278 345.987
R301 VDD.t2369 VDD.t2276 345.987
R302 VDD.t2391 VDD.t2369 345.987
R303 VDD.t2387 VDD.t2544 345.987
R304 VDD.t2544 VDD.t2542 345.987
R305 VDD.t2542 VDD.t2536 345.987
R306 VDD.t2598 VDD.t2605 345.987
R307 VDD.t2600 VDD.t2598 345.987
R308 VDD.t2524 VDD.t2600 345.987
R309 VDD.t2528 VDD.t2524 345.987
R310 VDD.t2522 VDD.t353 345.987
R311 VDD.t353 VDD.t859 345.987
R312 VDD.t859 VDD.t260 345.987
R313 VDD.t1546 VDD.t1480 345.987
R314 VDD.t1502 VDD.t1546 345.987
R315 VDD.t532 VDD.t409 345.987
R316 VDD.t409 VDD.t44 345.987
R317 VDD.t1570 VDD.t1520 345.987
R318 VDD.t1568 VDD.t1570 345.987
R319 VDD.t1282 VDD.t1286 345.987
R320 VDD.t1286 VDD.t1284 345.987
R321 VDD.t1516 VDD.t1552 345.987
R322 VDD.t1496 VDD.t1516 345.987
R323 VDD.t958 VDD.t956 345.987
R324 VDD.t956 VDD.t954 345.987
R325 VDD.t1526 VDD.t1564 345.987
R326 VDD.t1514 VDD.t1526 345.987
R327 VDD.t121 VDD.t139 345.987
R328 VDD.t139 VDD.t987 345.987
R329 VDD.t1500 VDD.t1540 345.987
R330 VDD.t1484 VDD.t1500 345.987
R331 VDD.t132 VDD.t130 345.987
R332 VDD.t130 VDD.t134 345.987
R333 VDD.t1498 VDD.t1508 345.987
R334 VDD.t1560 VDD.t1498 345.987
R335 VDD.t629 VDD.t627 345.987
R336 VDD.t627 VDD.t631 345.987
R337 VDD.t1542 VDD.t1486 345.987
R338 VDD.t1504 VDD.t1542 345.987
R339 VDD.t1936 VDD.t1934 345.987
R340 VDD.t1934 VDD.t1932 345.987
R341 VDD.t1492 VDD.t1518 345.987
R342 VDD.t1554 VDD.t1492 345.987
R343 VDD.t1259 VDD.t1257 345.987
R344 VDD.t1257 VDD.t1218 345.987
R345 VDD.t148 VDD.t220 345.987
R346 VDD.t220 VDD.t540 345.987
R347 VDD.t216 VDD.t528 345.987
R348 VDD.t528 VDD.t399 345.987
R349 VDD.t1263 VDD.t1265 345.987
R350 VDD.t1261 VDD.t1263 345.987
R351 VDD.t493 VDD.t6 345.987
R352 VDD.t491 VDD.t493 345.987
R353 VDD.t1780 VDD.t491 345.987
R354 VDD.t1770 VDD.t1780 345.987
R355 VDD.t1762 VDD.t1227 345.987
R356 VDD.t1227 VDD.t1225 345.987
R357 VDD.t1225 VDD.t1231 345.987
R358 VDD.t329 VDD.t484 345.987
R359 VDD.t331 VDD.t329 345.987
R360 VDD.t1233 VDD.t331 345.987
R361 VDD.t1237 VDD.t1233 345.987
R362 VDD.t1229 VDD.t153 345.987
R363 VDD.t153 VDD.t368 345.987
R364 VDD.t368 VDD.t233 345.987
R365 VDD.t474 VDD.t598 345.987
R366 VDD.t598 VDD.t960 345.987
R367 VDD.t1580 VDD.t1574 345.987
R368 VDD.t1574 VDD.t1578 345.987
R369 VDD.t2239 VDD.t2235 345.987
R370 VDD.t2257 VDD.t2239 345.987
R371 VDD.t1060 VDD.t1058 345.987
R372 VDD.t1062 VDD.t1060 345.987
R373 VDD.t1315 VDD.t1062 345.987
R374 VDD.t1335 VDD.t1315 345.987
R375 VDD.t1321 VDD.t2245 345.987
R376 VDD.t2245 VDD.t2255 345.987
R377 VDD.t2255 VDD.t2253 345.987
R378 VDD.t222 VDD.t890 345.987
R379 VDD.t888 VDD.t222 345.987
R380 VDD.t2251 VDD.t888 345.987
R381 VDD.t2241 VDD.t2251 345.987
R382 VDD.t2247 VDD.t1572 345.987
R383 VDD.t1572 VDD.t1586 345.987
R384 VDD.t1586 VDD.t1584 345.987
R385 VDD.t874 VDD.t878 345.987
R386 VDD.t878 VDD.t870 345.987
R387 VDD.t822 VDD.t57 345.987
R388 VDD.t57 VDD.t830 345.987
R389 VDD.t1729 VDD.t1737 345.987
R390 VDD.t1727 VDD.t1729 345.987
R391 VDD.t1683 VDD.t1711 345.987
R392 VDD.t1685 VDD.t1683 345.987
R393 VDD.t2220 VDD.t1685 345.987
R394 VDD.t2206 VDD.t2220 345.987
R395 VDD.t2216 VDD.t1721 345.987
R396 VDD.t1721 VDD.t1731 345.987
R397 VDD.t1731 VDD.t1719 345.987
R398 VDD.t1115 VDD.t1031 345.987
R399 VDD.t1029 VDD.t1115 345.987
R400 VDD.t1733 VDD.t1029 345.987
R401 VDD.t1741 VDD.t1733 345.987
R402 VDD.t1725 VDD.t832 345.987
R403 VDD.t832 VDD.t59 345.987
R404 VDD.t59 VDD.t836 345.987
R405 VDD.t2338 VDD.t2330 345.987
R406 VDD.t2330 VDD.t2334 345.987
R407 VDD.t1107 VDD.t1035 345.987
R408 VDD.t1035 VDD.t1041 345.987
R409 VDD.t2431 VDD.t2423 345.987
R410 VDD.t2437 VDD.t2431 345.987
R411 VDD.t387 VDD.t1291 345.987
R412 VDD.t389 VDD.t387 345.987
R413 VDD.t683 VDD.t389 345.987
R414 VDD.t928 VDD.t683 345.987
R415 VDD.t938 VDD.t2421 345.987
R416 VDD.t2421 VDD.t2429 345.987
R417 VDD.t2429 VDD.t2417 345.987
R418 VDD.t275 VDD.t697 345.987
R419 VDD.t277 VDD.t275 345.987
R420 VDD.t2435 VDD.t277 345.987
R421 VDD.t2419 VDD.t2435 345.987
R422 VDD.t2433 VDD.t1113 345.987
R423 VDD.t1113 VDD.t1039 345.987
R424 VDD.t1039 VDD.t1105 345.987
R425 VDD.t2292 VDD.t2298 345.987
R426 VDD.t2298 VDD.t2300 345.987
R427 VDD.t1342 VDD.t1350 345.987
R428 VDD.t1350 VDD.t454 345.987
R429 VDD.t842 VDD.t1064 345.987
R430 VDD.t611 VDD.t842 345.987
R431 VDD.t2306 VDD.t2308 345.987
R432 VDD.t2304 VDD.t2306 345.987
R433 VDD.t1701 VDD.t2304 345.987
R434 VDD.t1709 VDD.t1701 345.987
R435 VDD.t1693 VDD.t1070 345.987
R436 VDD.t1070 VDD.t840 345.987
R437 VDD.t840 VDD.t1076 345.987
R438 VDD.t2268 VDD.t2272 345.987
R439 VDD.t2270 VDD.t2268 345.987
R440 VDD.t609 VDD.t2270 345.987
R441 VDD.t1066 VDD.t609 345.987
R442 VDD.t1074 VDD.t1348 345.987
R443 VDD.t1348 VDD.t452 345.987
R444 VDD.t452 VDD.t1346 345.987
R445 VDD.n1093 VDD.t1638 343.055
R446 VDD.t782 VDD.t1880 312.28
R447 VDD.t1198 VDD.t1811 312.28
R448 VDD.t947 VDD.t1808 312.28
R449 VDD.t1604 VDD.t1815 312.28
R450 VDD.t1749 VDD.t1840 312.28
R451 VDD.t608 VDD.t1830 312.28
R452 VDD.t117 VDD.t1896 312.28
R453 VDD.t2078 VDD.t1845 312.28
R454 VDD.t765 VDD.t1303 312.28
R455 VDD.t2351 VDD.t1251 312.28
R456 VDD.t152 VDD.t183 312.28
R457 VDD.t527 VDD.t148 312.28
R458 VDD.t236 VDD.t474 312.28
R459 VDD.t847 VDD.t874 312.28
R460 VDD.t636 VDD.t2338 312.28
R461 VDD.t2285 VDD.t2292 312.28
R462 VDD.t1556 VDD.t2348 276.597
R463 VDD.t1482 VDD.t363 276.597
R464 VDD.t1490 VDD.t979 276.597
R465 VDD.t1512 VDD.t844 276.597
R466 VDD.t1476 VDD.t115 276.597
R467 VDD.t1558 VDD.t1607 276.597
R468 VDD.t1528 VDD.t969 276.597
R469 VDD.t1478 VDD.t633 276.597
R470 VDD.t1139 VDD.t1239 269.594
R471 VDD.t1088 VDD.t12 269.594
R472 VDD.t1047 VDD.t311 269.594
R473 VDD.t1091 VDD.t2558 269.594
R474 VDD.t1223 VDD.t1743 269.594
R475 VDD.t590 VDD.t552 269.594
R476 VDD.t861 VDD.t902 269.594
R477 VDD.t411 VDD.t522 269.594
R478 VDD.n1287 VDD.n1285 258.915
R479 VDD.n1305 VDD.n1303 258.915
R480 VDD.n1322 VDD.n1320 258.915
R481 VDD.n1339 VDD.n1337 258.915
R482 VDD.n1408 VDD.n1406 258.915
R483 VDD.n1425 VDD.n1423 258.915
R484 VDD.n375 VDD.n373 258.915
R485 VDD.n1270 VDD.n1268 258.915
R486 VDD.n1290 VDD.n1289 258.161
R487 VDD.n1308 VDD.n1307 258.161
R488 VDD.n1325 VDD.n1324 258.161
R489 VDD.n1342 VDD.n1341 258.161
R490 VDD.n1411 VDD.n1410 258.161
R491 VDD.n1428 VDD.n1427 258.161
R492 VDD.n378 VDD.n377 258.161
R493 VDD.n1273 VDD.n1272 258.161
R494 VDD.n1694 VDD.t1657 240.432
R495 VDD.n1101 VDD.t1691 240.432
R496 VDD.n1141 VDD.t936 240.432
R497 VDD.n1171 VDD.t2212 240.432
R498 VDD.n1195 VDD.t1337 240.432
R499 VDD.n754 VDD.t1768 240.432
R500 VDD.n731 VDD.t2389 240.432
R501 VDD.n641 VDD.t720 240.432
R502 VDD.n612 VDD.t1671 240.432
R503 VDD.n599 VDD.t976 240.432
R504 VDD.n693 VDD.t742 240.432
R505 VDD.n675 VDD.t790 240.432
R506 VDD.n534 VDD.t2387 240.432
R507 VDD.n522 VDD.t2522 240.432
R508 VDD.n468 VDD.t1762 240.432
R509 VDD.n452 VDD.t1229 240.432
R510 VDD.n843 VDD.t1321 240.432
R511 VDD.n840 VDD.t2247 240.432
R512 VDD.n909 VDD.t2216 240.432
R513 VDD.n901 VDD.t1725 240.432
R514 VDD.n973 VDD.t938 240.432
R515 VDD.n970 VDD.t2433 240.432
R516 VDD.n1037 VDD.t1693 240.432
R517 VDD.n1030 VDD.t1074 240.432
R518 VDD.t352 VDD.t1669 218.264
R519 VDD.t600 VDD.t740 218.264
R520 VDD.t1100 VDD.t2385 218.264
R521 VDD.t101 VDD.t1766 218.264
R522 VDD.t904 VDD.t1319 218.264
R523 VDD.t544 VDD.t2226 218.264
R524 VDD.t1152 VDD.t685 218.264
R525 VDD.t1655 VDD.t1705 218.264
R526 VDD.t989 VDD.t102 213.931
R527 VDD.t102 VDD.t2261 213.931
R528 VDD.t2261 VDD.t2259 213.931
R529 VDD.t2259 VDD.t2260 213.931
R530 VDD.t583 VDD.t585 213.931
R531 VDD.t585 VDD.t2289 213.931
R532 VDD.t2289 VDD.t2288 213.931
R533 VDD.t2288 VDD.t2290 213.931
R534 VDD.t2314 VDD.t2316 213.931
R535 VDD.t2316 VDD.t273 213.931
R536 VDD.t273 VDD.t219 213.931
R537 VDD.t219 VDD.t218 213.931
R538 VDD.t28 VDD.t30 213.931
R539 VDD.t30 VDD.t897 213.931
R540 VDD.t897 VDD.t898 213.931
R541 VDD.t898 VDD.t896 213.931
R542 VDD.t258 VDD.t254 213.931
R543 VDD.t254 VDD.t1034 213.931
R544 VDD.t1034 VDD.t1339 213.931
R545 VDD.t1339 VDD.t1033 213.931
R546 VDD.t1117 VDD.t1119 213.931
R547 VDD.t1119 VDD.t193 213.931
R548 VDD.t193 VDD.t905 213.931
R549 VDD.t905 VDD.t298 213.931
R550 VDD.t407 VDD.t250 213.931
R551 VDD.t250 VDD.t536 213.931
R552 VDD.t536 VDD.t189 213.931
R553 VDD.t189 VDD.t542 213.931
R554 VDD.t285 VDD.t1008 213.931
R555 VDD.t1008 VDD.t1057 213.931
R556 VDD.t1057 VDD.t1056 213.931
R557 VDD.t1056 VDD.t1055 213.931
R558 VDD.t892 VDD.t64 213.931
R559 VDD.t64 VDD.t603 213.931
R560 VDD.t603 VDD.t602 213.931
R561 VDD.t602 VDD.t601 213.931
R562 VDD.t170 VDD.t168 213.931
R563 VDD.t168 VDD.t1293 213.931
R564 VDD.t1293 VDD.t287 213.931
R565 VDD.t287 VDD.t1294 213.931
R566 VDD.t42 VDD.t191 213.931
R567 VDD.t191 VDD.t2350 213.931
R568 VDD.t2350 VDD.t2521 213.931
R569 VDD.t2521 VDD.t2520 213.931
R570 VDD.t1715 VDD.t1713 213.931
R571 VDD.t1713 VDD.t899 213.931
R572 VDD.t899 VDD.t503 213.931
R573 VDD.t503 VDD.t509 213.931
R574 VDD.t39 VDD.t999 213.931
R575 VDD.t999 VDD.t380 213.931
R576 VDD.t380 VDD.t984 213.931
R577 VDD.t984 VDD.t983 213.931
R578 VDD.t749 VDD.t747 213.931
R579 VDD.t747 VDD.t439 213.931
R580 VDD.t439 VDD.t438 213.931
R581 VDD.t438 VDD.t945 213.931
R582 VDD.t1006 VDD.t517 213.931
R583 VDD.t517 VDD.t763 213.931
R584 VDD.t763 VDD.t762 213.931
R585 VDD.t762 VDD.t761 213.931
R586 VDD.t1669 VDD.t1667 213.931
R587 VDD.t1667 VDD.t1665 213.931
R588 VDD.t2603 VDD.t2608 213.931
R589 VDD.t2608 VDD.t507 213.931
R590 VDD.t507 VDD.t161 213.931
R591 VDD.t161 VDD.t531 213.931
R592 VDD.t740 VDD.t738 213.931
R593 VDD.t738 VDD.t736 213.931
R594 VDD.t2385 VDD.t2383 213.931
R595 VDD.t2383 VDD.t2381 213.931
R596 VDD.t1766 VDD.t1764 213.931
R597 VDD.t1764 VDD.t1778 213.931
R598 VDD.t1319 VDD.t1333 213.931
R599 VDD.t1333 VDD.t1325 213.931
R600 VDD.t2226 VDD.t2210 213.931
R601 VDD.t2210 VDD.t2222 213.931
R602 VDD.t685 VDD.t932 213.931
R603 VDD.t932 VDD.t679 213.931
R604 VDD.t1705 VDD.t1687 213.931
R605 VDD.t1687 VDD.t1697 213.931
R606 VDD.t1789 VDD.t2189 205.749
R607 VDD.t2447 VDD.t519 205.749
R608 VDD.t106 VDD.t1216 205.749
R609 VDD.t136 VDD.t2550 205.749
R610 VDD.t2189 VDD.t2185 197.707
R611 VDD.t2185 VDD.t2183 197.707
R612 VDD.t519 VDD.t104 197.707
R613 VDD.t104 VDD.t376 197.707
R614 VDD.t2159 VDD.t2157 197.707
R615 VDD.t1216 VDD.t1178 197.707
R616 VDD.t1178 VDD.t1210 197.707
R617 VDD.t2579 VDD.t2571 197.707
R618 VDD.t2550 VDD.t2548 197.707
R619 VDD.t2548 VDD.t2546 197.707
R620 VDD.t1387 VDD.t1391 197.707
R621 VDD.t1966 VDD.t1960 197.707
R622 VDD.t1793 VDD.t1791 196.666
R623 VDD.t1929 VDD.t1793 196.666
R624 VDD.t1977 VDD.t1929 196.666
R625 VDD.t1991 VDD.t1977 196.666
R626 VDD.t2011 VDD.t1991 196.666
R627 VDD.t2135 VDD.t2027 196.666
R628 VDD.t2027 VDD.t2132 196.666
R629 VDD.t2067 VDD.t2069 196.666
R630 VDD.t2065 VDD.t2067 196.666
R631 VDD.t2125 VDD.t2065 196.666
R632 VDD.t2123 VDD.t2125 196.666
R633 VDD.t2025 VDD.t2123 196.666
R634 VDD.t800 VDD.t1462 196.666
R635 VDD.t1462 VDD.t1468 196.666
R636 VDD.t137 VDD.t210 196.666
R637 VDD.t208 VDD.t137 196.666
R638 VDD.t2009 VDD.t208 196.666
R639 VDD.t2007 VDD.t2009 196.666
R640 VDD.t2001 VDD.t2007 196.666
R641 VDD.t1633 VDD.t1631 196.666
R642 VDD.t1631 VDD.t1617 196.666
R643 VDD.t770 VDD.t857 196.666
R644 VDD.t855 VDD.t770 196.666
R645 VDD.t2477 VDD.t855 196.666
R646 VDD.t2486 VDD.t2477 196.666
R647 VDD.t2464 VDD.t2486 196.666
R648 VDD.t1464 VDD.t853 196.666
R649 VDD.t853 VDD.t851 196.666
R650 VDD.t1472 VDD.t1474 196.666
R651 VDD.t1470 VDD.t1472 196.666
R652 VDD.t2140 VDD.t1470 196.666
R653 VDD.t2033 VDD.t2140 196.666
R654 VDD.t2138 VDD.t2033 196.666
R655 VDD.t20 VDD.t757 196.666
R656 VDD.t757 VDD.t294 196.666
R657 VDD.t2230 VDD.t2228 196.666
R658 VDD.t2173 VDD.t2230 196.666
R659 VDD.t2471 VDD.t2173 196.666
R660 VDD.t2469 VDD.t2471 196.666
R661 VDD.t2493 VDD.t2469 196.666
R662 VDD.t2103 VDD.t2111 196.666
R663 VDD.t2111 VDD.t2085 196.666
R664 VDD.t2395 VDD.t2397 196.666
R665 VDD.t2393 VDD.t2395 196.666
R666 VDD.t2107 VDD.t2393 196.666
R667 VDD.t2101 VDD.t2107 196.666
R668 VDD.t2095 VDD.t2101 196.666
R669 VDD.t2501 VDD.t2499 196.666
R670 VDD.t2499 VDD.t2367 196.666
R671 VDD.t1147 VDD.t1145 196.666
R672 VDD.t1143 VDD.t1147 196.666
R673 VDD.t802 VDD.t1143 196.666
R674 VDD.t1358 VDD.t802 196.666
R675 VDD.t1460 VDD.t1358 196.666
R676 VDD.t1642 VDD.t1615 196.666
R677 VDD.t1615 VDD.t1629 196.666
R678 VDD.t1434 VDD.t866 196.666
R679 VDD.t864 VDD.t1434 196.666
R680 VDD.t16 VDD.t864 196.666
R681 VDD.t753 VDD.t16 196.666
R682 VDD.t290 VDD.t753 196.666
R683 VDD.t1611 VDD.t1627 196.666
R684 VDD.t1627 VDD.t1640 196.666
R685 VDD.t364 VDD.t108 196.666
R686 VDD.t313 VDD.t364 196.666
R687 VDD.t2508 VDD.t313 196.666
R688 VDD.t2355 VDD.t2508 196.666
R689 VDD.t2363 VDD.t2355 196.666
R690 VDD.t125 VDD.t426 196.666
R691 VDD.t426 VDD.t759 196.666
R692 VDD.t2073 VDD.t2075 196.666
R693 VDD.t2071 VDD.t2073 196.666
R694 VDD.t2093 VDD.t2071 196.666
R695 VDD.t2091 VDD.t2093 196.666
R696 VDD.t2081 VDD.t2091 196.666
R697 VDD.t2039 VDD.t2037 196.666
R698 VDD.t2037 VDD.t2035 196.666
R699 VDD.t337 VDD.t906 196.666
R700 VDD.t288 VDD.t337 196.666
R701 VDD.t123 VDD.t288 196.666
R702 VDD.t550 VDD.t123 196.666
R703 VDD.t548 VDD.t550 196.666
R704 VDD.t2495 VDD.t2491 196.666
R705 VDD.t2491 VDD.t2479 196.666
R706 VDD.t46 VDD.t267 196.666
R707 VDD.t350 VDD.t46 196.666
R708 VDD.t2497 VDD.t350 196.666
R709 VDD.t2483 VDD.t2497 196.666
R710 VDD.t2481 VDD.t2483 196.666
R711 VDD.t1985 VDD.t1995 196.666
R712 VDD.t1995 VDD.t1993 196.666
R713 VDD.t1206 VDD.t701 196.666
R714 VDD.t1204 VDD.t1206 196.666
R715 VDD.t2360 VDD.t1204 196.666
R716 VDD.t2515 VDD.t2360 196.666
R717 VDD.t2511 VDD.t2515 196.666
R718 VDD.t812 VDD.t810 196.666
R719 VDD.t810 VDD.t808 196.666
R720 VDD.t2121 VDD.t2119 196.666
R721 VDD.t2117 VDD.t2121 196.666
R722 VDD.t477 VDD.t2117 196.666
R723 VDD.t545 VDD.t477 196.666
R724 VDD.t993 VDD.t545 196.666
R725 VDD.t2155 VDD.t2143 196.666
R726 VDD.t2143 VDD.t2149 196.666
R727 VDD.t637 VDD.t397 196.666
R728 VDD.t395 VDD.t637 196.666
R729 VDD.t2358 VDD.t395 196.666
R730 VDD.t2506 VDD.t2358 196.666
R731 VDD.t2513 VDD.t2506 196.666
R732 VDD.t2005 VDD.t1981 196.666
R733 VDD.t1981 VDD.t1997 196.666
R734 VDD.t1164 VDD.t1092 196.666
R735 VDD.t1166 VDD.t1164 196.666
R736 VDD.t1176 VDD.t1166 196.666
R737 VDD.t1214 VDD.t1176 196.666
R738 VDD.t1101 VDD.t1214 196.666
R739 VDD.t2577 VDD.t2581 196.666
R740 VDD.t2581 VDD.t2565 196.666
R741 VDD.t2451 VDD.t2274 196.666
R742 VDD.t2449 VDD.t2451 196.666
R743 VDD.t2552 VDD.t2449 196.666
R744 VDD.t2461 VDD.t2552 196.666
R745 VDD.t2453 VDD.t2461 196.666
R746 VDD.t1399 VDD.t1397 196.666
R747 VDD.t1397 VDD.t1395 196.666
R748 VDD.t1182 VDD.t1184 196.666
R749 VDD.t1180 VDD.t1182 196.666
R750 VDD.t2187 VDD.t1180 196.666
R751 VDD.t2181 VDD.t2187 196.666
R752 VDD.t2179 VDD.t2181 196.666
R753 VDD.t1972 VDD.t1970 196.666
R754 VDD.t1970 VDD.t1968 196.666
R755 VDD.t661 VDD.t663 192.281
R756 VDD.t796 VDD.t355 192.281
R757 VDD.t796 VDD.t794 192.281
R758 VDD.t82 VDD.t84 192.281
R759 VDD.t88 VDD.t92 192.281
R760 VDD.t88 VDD.t90 192.281
R761 VDD.t1080 VDD.t1084 192.281
R762 VDD.t162 VDD.t8 192.281
R763 VDD.t162 VDD.t346 192.281
R764 VDD.t155 VDD.t113 192.281
R765 VDD.t1125 VDD.t1149 192.281
R766 VDD.t1125 VDD.t1123 192.281
R767 VDD.t341 VDD.t343 192.281
R768 VDD.t325 VDD.t321 192.281
R769 VDD.t325 VDD.t323 192.281
R770 VDD.t1753 VDD.t1755 192.281
R771 VDD.t25 VDD.t995 192.281
R772 VDD.t25 VDD.t110 192.281
R773 VDD.t2612 VDD.t2614 192.281
R774 VDD.t315 VDD.t393 192.281
R775 VDD.t1362 VDD.t1364 192.281
R776 VDD.t1362 VDD.t1360 192.281
R777 VDD.t68 VDD.t479 192.281
R778 VDD.t68 VDD.t303 192.281
R779 VDD.n1292 VDD.n1291 184.375
R780 VDD.n1310 VDD.n1309 184.375
R781 VDD.n1327 VDD.n1326 184.375
R782 VDD.n1344 VDD.n1343 184.375
R783 VDD.n1413 VDD.n1412 184.375
R784 VDD.n1430 VDD.n1429 184.375
R785 VDD.n380 VDD.n379 184.375
R786 VDD.n1275 VDD.n1274 184.375
R787 VDD.n1284 VDD.n1282 182.117
R788 VDD.n1302 VDD.n1300 182.117
R789 VDD.n1319 VDD.n1317 182.117
R790 VDD.n1336 VDD.n1334 182.117
R791 VDD.n1405 VDD.n1403 182.117
R792 VDD.n1422 VDD.n1420 182.117
R793 VDD.n372 VDD.n370 182.117
R794 VDD.n1267 VDD.n1265 182.117
R795 VDD.n1650 VDD.t1272 170.677
R796 VDD.n1616 VDD.t292 170.677
R797 VDD.n1591 VDD.t2099 170.677
R798 VDD.n1566 VDD.t2003 170.677
R799 VDD.n1541 VDD.t816 170.677
R800 VDD.n1516 VDD.t511 170.677
R801 VDD.n1500 VDD.t711 170.677
R802 VDD.n1466 VDD.t1158 170.677
R803 VDD.n1113 VDD.t659 169.468
R804 VDD.n1145 VDD.t80 169.468
R805 VDD.n1176 VDD.t1082 169.468
R806 VDD.n1208 VDD.t361 169.468
R807 VDD.n766 VDD.t339 169.468
R808 VDD.n740 VDD.t1751 169.468
R809 VDD.n654 VDD.t2610 169.468
R810 VDD.n1708 VDD.t299 169.468
R811 VDD.n1617 VDD.n1616 151.673
R812 VDD.n1592 VDD.n1591 151.673
R813 VDD.n1567 VDD.n1566 151.673
R814 VDD.n1542 VDD.n1541 151.673
R815 VDD.n1517 VDD.n1516 151.673
R816 VDD.n1467 VDD.n1466 151.673
R817 VDD.n1651 VDD.n1650 151.671
R818 VDD.n1501 VDD.n1500 151.671
R819 VDD.n637 VDD.n636 142.5
R820 VDD.n725 VDD.n724 142.5
R821 VDD.n554 VDD.n553 142.5
R822 VDD.n491 VDD.n490 142.5
R823 VDD.n868 VDD.n867 142.5
R824 VDD.n936 VDD.n935 142.5
R825 VDD.n999 VDD.n998 142.5
R826 VDD.n1063 VDD.n1062 142.5
R827 VDD.t1241 VDD.t1243 137.714
R828 VDD.t1239 VDD.t1241 137.714
R829 VDD.t1133 VDD.t1139 137.714
R830 VDD.t1494 VDD.t1556 137.714
R831 VDD.t2348 VDD.t2349 137.714
R832 VDD.t2349 VDD.t2347 137.714
R833 VDD.t2 VDD.t4 137.714
R834 VDD.t12 VDD.t2 137.714
R835 VDD.t1087 VDD.t1088 137.714
R836 VDD.t1530 VDD.t1482 137.714
R837 VDD.t363 VDD.t1005 137.714
R838 VDD.t1005 VDD.t508 137.714
R839 VDD.t269 VDD.t348 137.714
R840 VDD.t311 VDD.t269 137.714
R841 VDD.t883 VDD.t1047 137.714
R842 VDD.t1534 VDD.t1490 137.714
R843 VDD.t979 VDD.t262 137.714
R844 VDD.t262 VDD.t982 137.714
R845 VDD.t2554 VDD.t2556 137.714
R846 VDD.t2558 VDD.t2554 137.714
R847 VDD.t1169 VDD.t1091 137.714
R848 VDD.t1550 VDD.t1512 137.714
R849 VDD.t844 VDD.t846 137.714
R850 VDD.t846 VDD.t845 137.714
R851 VDD.t1745 VDD.t1747 137.714
R852 VDD.t1743 VDD.t1745 137.714
R853 VDD.t1222 VDD.t1223 137.714
R854 VDD.t1522 VDD.t1476 137.714
R855 VDD.t115 VDD.t253 137.714
R856 VDD.t253 VDD.t1010 137.714
R857 VDD.t554 VDD.t556 137.714
R858 VDD.t552 VDD.t554 137.714
R859 VDD.t589 VDD.t590 137.714
R860 VDD.t1562 VDD.t1558 137.714
R861 VDD.t1607 VDD.t1605 137.714
R862 VDD.t1605 VDD.t1606 137.714
R863 VDD.t35 VDD.t900 137.714
R864 VDD.t902 VDD.t35 137.714
R865 VDD.t621 VDD.t861 137.714
R866 VDD.t1566 VDD.t1528 137.714
R867 VDD.t969 VDD.t968 137.714
R868 VDD.t968 VDD.t967 137.714
R869 VDD.t497 VDD.t301 137.714
R870 VDD.t522 VDD.t497 137.714
R871 VDD.t160 VDD.t411 137.714
R872 VDD.t1524 VDD.t1478 137.714
R873 VDD.t633 VDD.t635 137.714
R874 VDD.t635 VDD.t634 137.714
R875 VDD.n1295 VDD.t1133 136.641
R876 VDD.n1313 VDD.t1087 136.641
R877 VDD.n1330 VDD.t883 136.641
R878 VDD.n1347 VDD.t1169 136.641
R879 VDD.n1416 VDD.t1222 136.641
R880 VDD.n1433 VDD.t589 136.641
R881 VDD.n383 VDD.t621 136.641
R882 VDD.n1278 VDD.t160 136.641
R883 VDD.t796 VDD.t583 135.973
R884 VDD.t88 VDD.t28 135.973
R885 VDD.t162 VDD.t1117 135.973
R886 VDD.t1125 VDD.t285 135.973
R887 VDD.t325 VDD.t170 135.973
R888 VDD.t25 VDD.t1715 135.973
R889 VDD.t1362 VDD.t1006 135.973
R890 VDD.t68 VDD.t2603 135.973
R891 VDD.n1296 VDD.t1494 121.615
R892 VDD.n1314 VDD.t1530 121.615
R893 VDD.n1331 VDD.t1534 121.615
R894 VDD.n1348 VDD.t1550 121.615
R895 VDD.n1417 VDD.t1522 121.615
R896 VDD.n1434 VDD.t1562 121.615
R897 VDD.n384 VDD.t1566 121.615
R898 VDD.n1279 VDD.t1524 121.615
R899 VDD.n1650 VDD.n1647 115.932
R900 VDD.n1616 VDD.n1613 115.932
R901 VDD.n1591 VDD.n1588 115.932
R902 VDD.n1566 VDD.n1563 115.932
R903 VDD.n1541 VDD.n1538 115.932
R904 VDD.n1516 VDD.n1513 115.932
R905 VDD.n1500 VDD.n1497 115.932
R906 VDD.n1466 VDD.n1463 115.932
R907 VDD.n1113 VDD.t989 110.591
R908 VDD.n1145 VDD.t2314 110.591
R909 VDD.n1176 VDD.t258 110.591
R910 VDD.n1208 VDD.t407 110.591
R911 VDD.n766 VDD.t892 110.591
R912 VDD.n740 VDD.t42 110.591
R913 VDD.n654 VDD.t39 110.591
R914 VDD.n1708 VDD.t749 110.591
R915 VDD.n1694 VDD.t1659 105.555
R916 VDD.n1101 VDD.t1703 105.555
R917 VDD.n1141 VDD.t687 105.555
R918 VDD.n1171 VDD.t2204 105.555
R919 VDD.n1195 VDD.t1329 105.555
R920 VDD.n754 VDD.t1772 105.555
R921 VDD.n731 VDD.t2377 105.555
R922 VDD.n641 VDD.t726 105.555
R923 VDD.n612 VDD.t1673 105.555
R924 VDD.n599 VDD.t461 105.555
R925 VDD.n693 VDD.t724 105.555
R926 VDD.n675 VDD.t1194 105.555
R927 VDD.n534 VDD.t2391 105.555
R928 VDD.n522 VDD.t2528 105.555
R929 VDD.n468 VDD.t1770 105.555
R930 VDD.n452 VDD.t1237 105.555
R931 VDD.n843 VDD.t1335 105.555
R932 VDD.n840 VDD.t2241 105.555
R933 VDD.n909 VDD.t2206 105.555
R934 VDD.n901 VDD.t1741 105.555
R935 VDD.n973 VDD.t928 105.555
R936 VDD.n970 VDD.t2419 105.555
R937 VDD.n1037 VDD.t1709 105.555
R938 VDD.n1030 VDD.t1066 105.555
R939 VDD.t985 VDD.n1113 103.339
R940 VDD.t2312 VDD.n1145 103.339
R941 VDD.t256 VDD.n1176 103.339
R942 VDD.t538 VDD.n1208 103.339
R943 VDD.t894 VDD.n766 103.339
R944 VDD.t263 VDD.n740 103.339
R945 VDD.t513 VDD.n654 103.339
R946 VDD.t751 VDD.n1708 103.339
R947 VDD.t796 VDD.t581 77.958
R948 VDD.t88 VDD.t32 77.958
R949 VDD.t162 VDD.t1121 77.958
R950 VDD.t1125 VDD.t849 77.958
R951 VDD.t325 VDD.t94 77.958
R952 VDD.t25 VDD.t1717 77.958
R953 VDD.t1362 VDD.t52 77.958
R954 VDD.t68 VDD.t2596 77.958
R955 VDD.t1842 VDD.t782 53.244
R956 VDD.t1874 VDD.t1198 53.244
R957 VDD.t1849 VDD.t947 53.244
R958 VDD.t1912 VDD.t1604 53.244
R959 VDD.t1822 VDD.t1749 53.244
R960 VDD.t1908 VDD.t608 53.244
R961 VDD.t1882 VDD.t117 53.244
R962 VDD.t1826 VDD.t2078 53.244
R963 VDD.t228 VDD.t515 53.244
R964 VDD.t1309 VDD.t765 53.244
R965 VDD.t641 VDD.t420 53.244
R966 VDD.t1253 VDD.t2351 53.244
R967 VDD.t1380 VDD.t2530 53.244
R968 VDD.t173 VDD.t152 53.244
R969 VDD.t1187 VDD.t1235 53.244
R970 VDD.t78 VDD.t527 53.244
R971 VDD.t1136 VDD.t2237 53.244
R972 VDD.t391 VDD.t236 53.244
R973 VDD.t745 VDD.t1735 53.244
R974 VDD.t868 VDD.t847 53.244
R975 VDD.t1601 VDD.t2415 53.244
R976 VDD.t2328 VDD.t636 53.244
R977 VDD.t15 VDD.t1072 53.244
R978 VDD.t2294 VDD.t2285 53.244
R979 VDD.t980 VDD.n632 47.617
R980 VDD.t515 VDD.n633 47.617
R981 VDD.n635 VDD.t1305 47.617
R982 VDD.n634 VDD.t1309 47.617
R983 VDD.t194 VDD.n720 47.617
R984 VDD.t420 VDD.n721 47.617
R985 VDD.n723 VDD.t98 47.617
R986 VDD.n722 VDD.t1253 47.617
R987 VDD.t2538 VDD.n549 47.617
R988 VDD.t2530 VDD.n550 47.617
R989 VDD.n552 VDD.t175 47.617
R990 VDD.n551 VDD.t173 47.617
R991 VDD.t1127 VDD.n486 47.617
R992 VDD.t1235 VDD.n487 47.617
R993 VDD.n489 VDD.t951 47.617
R994 VDD.n488 VDD.t78 47.617
R995 VDD.t2249 VDD.n863 47.617
R996 VDD.t2237 VDD.n864 47.617
R997 VDD.n866 VDD.t565 47.617
R998 VDD.n865 VDD.t391 47.617
R999 VDD.t1723 VDD.n931 47.617
R1000 VDD.t1735 VDD.n932 47.617
R1001 VDD.n934 VDD.t876 47.617
R1002 VDD.n933 VDD.t868 47.617
R1003 VDD.t2425 VDD.n994 47.617
R1004 VDD.t2415 VDD.n995 47.617
R1005 VDD.n997 VDD.t2336 47.617
R1006 VDD.n996 VDD.t2328 47.617
R1007 VDD.t1078 VDD.n1058 47.617
R1008 VDD.t1072 VDD.n1059 47.617
R1009 VDD.n1061 VDD.t2296 47.617
R1010 VDD.n1060 VDD.t2294 47.617
R1011 VDD.t433 VDD.t1448 47.617
R1012 VDD.t431 VDD.t1438 47.617
R1013 VDD.t432 VDD.t1679 47.617
R1014 VDD.t1012 VDD.t1677 47.617
R1015 VDD.t1013 VDD.t1675 47.617
R1016 VDD.t625 VDD.t2053 47.617
R1017 VDD.t626 VDD.t2061 47.617
R1018 VDD.t624 VDD.t734 47.617
R1019 VDD.t772 VDD.t732 47.617
R1020 VDD.t773 VDD.t722 47.617
R1021 VDD.t1269 VDD.t271 47.617
R1022 VDD.t1267 VDD.t405 47.617
R1023 VDD.t1268 VDD.t2375 47.617
R1024 VDD.t1297 VDD.t2373 47.617
R1025 VDD.t1296 VDD.t2371 47.617
R1026 VDD.t974 VDD.t499 47.617
R1027 VDD.t501 VDD.t525 47.617
R1028 VDD.t973 VDD.t1760 47.617
R1029 VDD.t328 VDD.t1776 47.617
R1030 VDD.t476 VDD.t1774 47.617
R1031 VDD.t1290 VDD.t1576 47.617
R1032 VDD.t1288 VDD.t1588 47.617
R1033 VDD.t1289 VDD.t1317 47.617
R1034 VDD.t249 VDD.t1327 47.617
R1035 VDD.t430 VDD.t1331 47.617
R1036 VDD.t27 VDD.t834 47.617
R1037 VDD.t1203 VDD.t824 47.617
R1038 VDD.t274 VDD.t2224 47.617
R1039 VDD.t167 VDD.t2208 47.617
R1040 VDD.t535 VDD.t2214 47.617
R1041 VDD.t2344 VDD.t1045 47.617
R1042 VDD.t2342 VDD.t1043 47.617
R1043 VDD.t2343 VDD.t934 47.617
R1044 VDD.t1153 VDD.t681 47.617
R1045 VDD.t1151 VDD.t930 47.617
R1046 VDD.t789 VDD.t1354 47.617
R1047 VDD.t787 VDD.t1340 47.617
R1048 VDD.t788 VDD.t1699 47.617
R1049 VDD.t1656 VDD.t1707 47.617
R1050 VDD.t1654 VDD.t1689 47.617
R1051 VDD.n1114 VDD.t985 47.137
R1052 VDD.n1146 VDD.t2312 47.137
R1053 VDD.n1177 VDD.t256 47.137
R1054 VDD.n1209 VDD.t538 47.137
R1055 VDD.n767 VDD.t894 47.137
R1056 VDD.n741 VDD.t263 47.137
R1057 VDD.n655 VDD.t513 47.137
R1058 VDD.n1709 VDD.t751 47.137
R1059 VDD.t2147 VDD.t284 45.992
R1060 VDD.t2151 VDD.t966 45.992
R1061 VDD.t2446 VDD.t715 45.992
R1062 VDD.t2448 VDD.t504 45.992
R1063 VDD.t2573 VDD.t231 45.992
R1064 VDD.t2569 VDD.t229 45.992
R1065 VDD.t215 VDD.t1174 45.992
R1066 VDD.t502 VDD.t141 45.992
R1067 VDD.t1385 VDD.t949 45.992
R1068 VDD.t1383 VDD.t950 45.992
R1069 VDD.t530 VDD.t2457 45.992
R1070 VDD.t248 VDD.t2455 45.992
R1071 VDD.t1962 VDD.t10 45.992
R1072 VDD.t1956 VDD.t100 45.992
R1073 VDD.t1790 VDD.t2175 45.992
R1074 VDD.t1788 VDD.t2191 45.992
R1075 VDD.n633 VDD.t980 44.495
R1076 VDD.t1307 VDD.n635 44.495
R1077 VDD.t1305 VDD.n634 44.495
R1078 VDD.n632 VDD.t143 44.495
R1079 VDD.n721 VDD.t194 44.495
R1080 VDD.t1245 VDD.n723 44.495
R1081 VDD.t98 VDD.n722 44.495
R1082 VDD.n720 VDD.t418 44.495
R1083 VDD.n550 VDD.t2538 44.495
R1084 VDD.t177 VDD.n552 44.495
R1085 VDD.t175 VDD.n551 44.495
R1086 VDD.n549 VDD.t2540 44.495
R1087 VDD.n487 VDD.t1127 44.495
R1088 VDD.t265 VDD.n489 44.495
R1089 VDD.t951 VDD.n488 44.495
R1090 VDD.n486 VDD.t1129 44.495
R1091 VDD.n864 VDD.t2249 44.495
R1092 VDD.t66 VDD.n866 44.495
R1093 VDD.t565 VDD.n865 44.495
R1094 VDD.n863 VDD.t2243 44.495
R1095 VDD.n932 VDD.t1723 44.495
R1096 VDD.t872 VDD.n934 44.495
R1097 VDD.t876 VDD.n933 44.495
R1098 VDD.n931 VDD.t1739 44.495
R1099 VDD.n995 VDD.t2425 44.495
R1100 VDD.t2332 VDD.n997 44.495
R1101 VDD.t2336 VDD.n996 44.495
R1102 VDD.n994 VDD.t2427 44.495
R1103 VDD.n1059 VDD.t1078 44.495
R1104 VDD.t2302 VDD.n1061 44.495
R1105 VDD.t2296 VDD.n1060 44.495
R1106 VDD.n1058 VDD.t1068 44.495
R1107 VDD.t1450 VDD.t433 44.494
R1108 VDD.t1448 VDD.t431 44.494
R1109 VDD.t1438 VDD.t432 44.494
R1110 VDD.t1679 VDD.t1012 44.494
R1111 VDD.t1677 VDD.t1013 44.494
R1112 VDD.t1675 VDD.t352 44.494
R1113 VDD.t2055 VDD.t625 44.494
R1114 VDD.t2053 VDD.t626 44.494
R1115 VDD.t2061 VDD.t624 44.494
R1116 VDD.t734 VDD.t772 44.494
R1117 VDD.t732 VDD.t773 44.494
R1118 VDD.t722 VDD.t600 44.494
R1119 VDD.t604 VDD.t1269 44.494
R1120 VDD.t271 VDD.t1267 44.494
R1121 VDD.t405 VDD.t1268 44.494
R1122 VDD.t2375 VDD.t1297 44.494
R1123 VDD.t2373 VDD.t1296 44.494
R1124 VDD.t2371 VDD.t1100 44.494
R1125 VDD.t997 VDD.t974 44.494
R1126 VDD.t499 VDD.t501 44.494
R1127 VDD.t525 VDD.t973 44.494
R1128 VDD.t1760 VDD.t328 44.494
R1129 VDD.t1776 VDD.t476 44.494
R1130 VDD.t1774 VDD.t101 44.494
R1131 VDD.t1594 VDD.t1290 44.494
R1132 VDD.t1576 VDD.t1288 44.494
R1133 VDD.t1588 VDD.t1289 44.494
R1134 VDD.t1317 VDD.t249 44.494
R1135 VDD.t1327 VDD.t430 44.494
R1136 VDD.t1331 VDD.t904 44.494
R1137 VDD.t828 VDD.t27 44.494
R1138 VDD.t834 VDD.t1203 44.494
R1139 VDD.t824 VDD.t274 44.494
R1140 VDD.t2224 VDD.t167 44.494
R1141 VDD.t2208 VDD.t535 44.494
R1142 VDD.t2214 VDD.t544 44.494
R1143 VDD.t1111 VDD.t2344 44.494
R1144 VDD.t1045 VDD.t2342 44.494
R1145 VDD.t1043 VDD.t2343 44.494
R1146 VDD.t934 VDD.t1153 44.494
R1147 VDD.t681 VDD.t1151 44.494
R1148 VDD.t930 VDD.t1152 44.494
R1149 VDD.t456 VDD.t789 44.494
R1150 VDD.t1354 VDD.t787 44.494
R1151 VDD.t1340 VDD.t788 44.494
R1152 VDD.t1699 VDD.t1656 44.494
R1153 VDD.t1707 VDD.t1654 44.494
R1154 VDD.t1689 VDD.t1655 44.494
R1155 VDD.n1645 VDD.t1842 44.17
R1156 VDD.n1646 VDD.t1906 44.17
R1157 VDD.t1272 VDD.n1649 44.17
R1158 VDD.t1280 VDD.n1648 44.17
R1159 VDD.n1611 VDD.t1874 44.17
R1160 VDD.n1612 VDD.t1835 44.17
R1161 VDD.t292 VDD.n1615 44.17
R1162 VDD.t424 VDD.n1614 44.17
R1163 VDD.n1586 VDD.t1849 44.17
R1164 VDD.n1587 VDD.t1910 44.17
R1165 VDD.t2099 VDD.n1590 44.17
R1166 VDD.t2089 VDD.n1589 44.17
R1167 VDD.n1561 VDD.t1912 44.17
R1168 VDD.n1562 VDD.t1865 44.17
R1169 VDD.t2003 VDD.n1565 44.17
R1170 VDD.t1989 VDD.n1564 44.17
R1171 VDD.n1536 VDD.t1822 44.17
R1172 VDD.n1537 VDD.t1888 44.17
R1173 VDD.t816 VDD.n1540 44.17
R1174 VDD.t806 VDD.n1539 44.17
R1175 VDD.n1511 VDD.t1908 44.17
R1176 VDD.n1512 VDD.t1890 44.17
R1177 VDD.t511 VDD.n1515 44.17
R1178 VDD.t458 VDD.n1514 44.17
R1179 VDD.n1495 VDD.t1882 44.17
R1180 VDD.n1496 VDD.t1847 44.17
R1181 VDD.t711 VDD.n1499 44.17
R1182 VDD.t707 VDD.n1498 44.17
R1183 VDD.n1461 VDD.t1826 44.17
R1184 VDD.n1462 VDD.t1894 44.17
R1185 VDD.t1158 VDD.n1465 44.17
R1186 VDD.t1156 VDD.n1464 44.17
R1187 VDD.t284 VDD.t2153 42.976
R1188 VDD.t966 VDD.t2147 42.976
R1189 VDD.t283 VDD.t2151 42.976
R1190 VDD.t403 VDD.t2446 42.976
R1191 VDD.t715 VDD.t2448 42.976
R1192 VDD.t504 VDD.t2447 42.976
R1193 VDD.t231 VDD.t2567 42.976
R1194 VDD.t229 VDD.t2573 42.976
R1195 VDD.t230 VDD.t2569 42.976
R1196 VDD.t1212 VDD.t215 42.976
R1197 VDD.t1174 VDD.t502 42.976
R1198 VDD.t141 VDD.t106 42.976
R1199 VDD.t949 VDD.t1393 42.976
R1200 VDD.t950 VDD.t1385 42.976
R1201 VDD.t948 VDD.t1383 42.976
R1202 VDD.t2459 VDD.t530 42.976
R1203 VDD.t2457 VDD.t248 42.976
R1204 VDD.t2455 VDD.t136 42.976
R1205 VDD.t10 VDD.t1964 42.976
R1206 VDD.t100 VDD.t1962 42.976
R1207 VDD.t172 VDD.t1956 42.976
R1208 VDD.t2177 VDD.t1790 42.976
R1209 VDD.t2175 VDD.t1788 42.976
R1210 VDD.t2191 VDD.t1789 42.976
R1211 VDD.t1906 VDD.n1645 41.273
R1212 VDD.t1884 VDD.n1646 41.273
R1213 VDD.n1649 VDD.t1280 41.273
R1214 VDD.n1648 VDD.t1278 41.273
R1215 VDD.t1835 VDD.n1611 41.273
R1216 VDD.t1902 VDD.n1612 41.273
R1217 VDD.n1615 VDD.t424 41.273
R1218 VDD.n1614 VDD.t755 41.273
R1219 VDD.t1910 VDD.n1586 41.273
R1220 VDD.t1892 VDD.n1587 41.273
R1221 VDD.n1590 VDD.t2089 41.273
R1222 VDD.n1589 VDD.t2115 41.273
R1223 VDD.t1865 VDD.n1561 41.273
R1224 VDD.t1824 VDD.n1562 41.273
R1225 VDD.n1565 VDD.t1989 41.273
R1226 VDD.n1564 VDD.t1983 41.273
R1227 VDD.t1888 VDD.n1536 41.273
R1228 VDD.t1852 VDD.n1537 41.273
R1229 VDD.n1540 VDD.t806 41.273
R1230 VDD.n1539 VDD.t1466 41.273
R1231 VDD.t1890 VDD.n1511 41.273
R1232 VDD.t1869 VDD.n1512 41.273
R1233 VDD.n1515 VDD.t458 41.273
R1234 VDD.n1514 VDD.t242 41.273
R1235 VDD.t1847 VDD.n1495 41.273
R1236 VDD.t1828 VDD.n1496 41.273
R1237 VDD.n1499 VDD.t707 41.273
R1238 VDD.n1498 VDD.t703 41.273
R1239 VDD.t1894 VDD.n1461 41.273
R1240 VDD.t1855 VDD.n1462 41.273
R1241 VDD.n1465 VDD.t1156 41.273
R1242 VDD.n1464 VDD.t1160 41.273
R1243 VDD.n1253 VDD.t403 37.698
R1244 VDD.n1239 VDD.t1212 37.698
R1245 VDD.n398 VDD.t2459 37.698
R1246 VDD.n1390 VDD.t2177 37.698
R1247 VDD.n1483 VDD.t1897 30.726
R1248 VDD.n1717 VDD.t1445 30.238
R1249 VDD.n1731 VDD.t1618 30.238
R1250 VDD.n1203 VDD.t1591 30.238
R1251 VDD.n811 VDD.t295 30.238
R1252 VDD.n821 VDD.t2086 30.238
R1253 VDD.n649 VDD.t2058 30.238
R1254 VDD.n418 VDD.t2566 30.238
R1255 VDD.n407 VDD.t1396 30.238
R1256 VDD.n837 VDD.t1585 30.238
R1257 VDD.n898 VDD.t837 30.238
R1258 VDD.n967 VDD.t1106 30.238
R1259 VDD.n1027 VDD.t1347 30.238
R1260 VDD.n11 VDD.t488 30.163
R1261 VDD.n3 VDD.t2165 30.163
R1262 VDD.n1832 VDD.t2171 30.163
R1263 VDD.n47 VDD.t653 30.163
R1264 VDD.n1784 VDD.t1810 30.163
R1265 VDD.n51 VDD.t652 30.163
R1266 VDD.n1690 VDD.t2133 30.163
R1267 VDD.n1680 VDD.t1469 30.163
R1268 VDD.n1083 VDD.t852 30.163
R1269 VDD.n1104 VDD.t1353 30.163
R1270 VDD.n1138 VDD.t1110 30.163
R1271 VDD.n1167 VDD.t62 30.163
R1272 VDD.n1091 VDD.t2114 30.163
R1273 VDD.n445 VDD.t2368 30.163
R1274 VDD.n436 VDD.t1630 30.163
R1275 VDD.n794 VDD.t1641 30.163
R1276 VDD.n803 VDD.t760 30.163
R1277 VDD.n757 VDD.t384 30.163
R1278 VDD.n734 VDD.t23 30.163
R1279 VDD.n615 VDD.t297 30.163
R1280 VDD.n606 VDD.t1447 30.163
R1281 VDD.n690 VDD.t1189 30.163
R1282 VDD.n678 VDD.t2046 30.163
R1283 VDD.n531 VDD.t2537 30.163
R1284 VDD.n519 VDD.t261 30.163
R1285 VDD.n1374 VDD.t2036 30.163
R1286 VDD.n1366 VDD.t2480 30.163
R1287 VDD.n1671 VDD.t1994 30.163
R1288 VDD.n1358 VDD.t809 30.163
R1289 VDD.n1393 VDD.t1969 30.163
R1290 VDD.n1262 VDD.t2150 30.163
R1291 VDD.n428 VDD.t1998 30.163
R1292 VDD.n69 VDD.t644 30.163
R1293 VDD.n126 VDD.t2467 30.163
R1294 VDD.n183 VDD.t2127 30.163
R1295 VDD.n240 VDD.t1614 30.163
R1296 VDD.n87 VDD.t2583 30.163
R1297 VDD.n97 VDD.t2488 30.163
R1298 VDD.n144 VDD.t2193 30.163
R1299 VDD.n154 VDD.t2137 30.163
R1300 VDD.n201 VDD.t916 30.163
R1301 VDD.n211 VDD.t1637 30.163
R1302 VDD.n338 VDD.t448 30.163
R1303 VDD.n330 VDD.t2518 30.163
R1304 VDD.n309 VDD.t2365 30.163
R1305 VDD.n288 VDD.t74 30.163
R1306 VDD.n255 VDD.t1955 30.163
R1307 VDD.n247 VDD.t618 30.163
R1308 VDD.n461 VDD.t1232 30.163
R1309 VDD.n449 VDD.t234 30.163
R1310 VDD.n846 VDD.t2254 30.163
R1311 VDD.n906 VDD.t1720 30.163
R1312 VDD.n976 VDD.t2418 30.163
R1313 VDD.n1041 VDD.t1077 30.163
R1314 VDD.n1763 VDD.t1422 30.163
R1315 VDD.n1773 VDD.t564 30.163
R1316 VDD.n1647 VDD.t1951 29.891
R1317 VDD.n1613 VDD.t463 29.891
R1318 VDD.n1588 VDD.t1054 29.891
R1319 VDD.n1563 VDD.t308 29.891
R1320 VDD.n1538 VDD.t1134 29.891
R1321 VDD.n1513 VDD.t336 29.891
R1322 VDD.n1497 VDD.t767 29.891
R1323 VDD.n1463 VDD.t943 29.891
R1324 VDD.n636 VDD.t228 28.957
R1325 VDD.n724 VDD.t641 28.957
R1326 VDD.n553 VDD.t1380 28.957
R1327 VDD.n490 VDD.t1187 28.957
R1328 VDD.n867 VDD.t1136 28.957
R1329 VDD.n935 VDD.t745 28.957
R1330 VDD.n998 VDD.t1601 28.957
R1331 VDD.n1062 VDD.t15 28.957
R1332 VDD.n1556 VDD.t1980 28.913
R1333 VDD.n31 VDD.t164 28.664
R1334 VDD.n36 VDD.t885 28.664
R1335 VDD.n19 VDD.t665 28.664
R1336 VDD.n24 VDD.t2170 28.664
R1337 VDD.n1791 VDD.t2445 28.664
R1338 VDD.n1796 VDD.t1096 28.664
R1339 VDD.n1802 VDD.t2264 28.664
R1340 VDD.n1807 VDD.t1821 28.664
R1341 VDD.n1638 VDD.t1277 28.664
R1342 VDD.n1633 VDD.t1881 28.664
R1343 VDD.n1620 VDD.t1812 28.664
R1344 VDD.n1606 VDD.t19 28.664
R1345 VDD.n1595 VDD.t1809 28.664
R1346 VDD.n1581 VDD.t2110 28.664
R1347 VDD.n1570 VDD.t1816 28.664
R1348 VDD.n1545 VDD.t1841 28.664
R1349 VDD.n1531 VDD.t799 28.664
R1350 VDD.n1520 VDD.t1831 28.664
R1351 VDD.n1506 VDD.t225 28.664
R1352 VDD.n1488 VDD.t714 28.664
R1353 VDD.n1470 VDD.t1846 28.664
R1354 VDD.n1456 VDD.t1155 28.664
R1355 VDD.n586 VDD.t1304 28.664
R1356 VDD.n591 VDD.t128 28.664
R1357 VDD.n621 VDD.t1670 28.664
R1358 VDD.n626 VDD.t1437 28.664
R1359 VDD.n710 VDD.t1252 28.664
R1360 VDD.n715 VDD.t793 28.664
R1361 VDD.n697 VDD.t741 28.664
R1362 VDD.n702 VDD.t2050 28.664
R1363 VDD.n557 VDD.t184 28.664
R1364 VDD.n562 VDD.t2527 28.664
R1365 VDD.n538 VDD.t2386 28.664
R1366 VDD.n543 VDD.t55 28.664
R1367 VDD.n1385 VDD.t2190 28.664
R1368 VDD.n1380 VDD.t1959 28.664
R1369 VDD.n1248 VDD.t520 28.664
R1370 VDD.n1243 VDD.t2146 28.664
R1371 VDD.n1234 VDD.t1217 28.664
R1372 VDD.n1229 VDD.t2576 28.664
R1373 VDD.n393 VDD.t2551 28.664
R1374 VDD.n388 VDD.t1390 28.664
R1375 VDD.n80 VDD.t2485 28.664
R1376 VDD.n75 VDD.t567 28.664
R1377 VDD.n108 VDD.t2562 28.664
R1378 VDD.n103 VDD.t472 28.664
R1379 VDD.n137 VDD.t2134 28.664
R1380 VDD.n132 VDD.t1377 28.664
R1381 VDD.n165 VDD.t2201 28.664
R1382 VDD.n160 VDD.t560 28.664
R1383 VDD.n194 VDD.t1623 28.664
R1384 VDD.n189 VDD.t1403 28.664
R1385 VDD.n222 VDD.t920 28.664
R1386 VDD.n217 VDD.t1926 28.664
R1387 VDD.n358 VDD.t1019 28.664
R1388 VDD.n363 VDD.t464 28.664
R1389 VDD.n346 VDD.t1795 28.664
R1390 VDD.n351 VDD.t2517 28.664
R1391 VDD.n275 VDD.t1417 28.664
R1392 VDD.n280 VDD.t1917 28.664
R1393 VDD.n263 VDD.t569 28.664
R1394 VDD.n268 VDD.t71 28.664
R1395 VDD.n493 VDD.t149 28.664
R1396 VDD.n498 VDD.t1262 28.664
R1397 VDD.n475 VDD.t1767 28.664
R1398 VDD.n480 VDD.t400 28.664
R1399 VDD.n871 VDD.t475 28.664
R1400 VDD.n876 VDD.t2258 28.664
R1401 VDD.n852 VDD.t1320 28.664
R1402 VDD.n857 VDD.t1579 28.664
R1403 VDD.n883 VDD.t875 28.664
R1404 VDD.n888 VDD.t1728 28.664
R1405 VDD.n920 VDD.t2227 28.664
R1406 VDD.n925 VDD.t831 28.664
R1407 VDD.n949 VDD.t2339 28.664
R1408 VDD.n954 VDD.t2438 28.664
R1409 VDD.n983 VDD.t686 28.664
R1410 VDD.n988 VDD.t1042 28.664
R1411 VDD.n1012 VDD.t2293 28.664
R1412 VDD.n1017 VDD.t612 28.664
R1413 VDD.n1047 VDD.t1706 28.664
R1414 VDD.n1052 VDD.t455 28.664
R1415 VDD.n1756 VDD.t1945 28.664
R1416 VDD.n1751 VDD.t1314 28.664
R1417 VDD.n1745 VDD.t2593 28.664
R1418 VDD.n1740 VDD.t1430 28.664
R1419 VDD.n1841 VDD.t49 28.57
R1420 VDD.n1847 VDD.t1758 28.57
R1421 VDD.n1819 VDD.t247 28.57
R1422 VDD.n1825 VDD.t51 28.57
R1423 VDD.n59 VDD.t334 28.57
R1424 VDD.n1068 VDD.t664 28.57
R1425 VDD.n1123 VDD.t356 28.57
R1426 VDD.n1004 VDD.t85 28.57
R1427 VDD.n1153 VDD.t93 28.57
R1428 VDD.n941 VDD.t1085 28.57
R1429 VDD.n1183 VDD.t9 28.57
R1430 VDD.n1212 VDD.t114 28.57
R1431 VDD.n1219 VDD.t1150 28.57
R1432 VDD.n506 VDD.t344 28.57
R1433 VDD.n777 VDD.t322 28.57
R1434 VDD.n577 VDD.t1756 28.57
R1435 VDD.n570 VDD.t996 28.57
R1436 VDD.n659 VDD.t2615 28.57
R1437 VDD.n1704 VDD.t394 28.57
R1438 VDD.n1697 VDD.t1365 28.57
R1439 VDD.n667 VDD.t480 28.57
R1440 VDD.n173 VDD.t1089 28.57
R1441 VDD.n178 VDD.t2439 28.57
R1442 VDD.n121 VDD.t534 28.57
R1443 VDD.n116 VDD.t779 28.57
R1444 VDD.n235 VDD.t443 28.57
R1445 VDD.n230 VDD.t14 28.57
R1446 VDD.n64 VDD.t2311 28.57
R1447 VDD.n318 VDD.t972 28.57
R1448 VDD.n324 VDD.t1021 28.57
R1449 VDD.n302 VDD.t1142 28.57
R1450 VDD.n296 VDD.t1300 28.57
R1451 VDD.n1292 VDD.t533 28.568
R1452 VDD.n1310 VDD.t1283 28.568
R1453 VDD.n1327 VDD.t959 28.568
R1454 VDD.n1344 VDD.t122 28.568
R1455 VDD.n1413 VDD.t133 28.568
R1456 VDD.n1430 VDD.t630 28.568
R1457 VDD.n380 VDD.t1937 28.568
R1458 VDD.n1275 VDD.t1260 28.568
R1459 VDD.n32 VDD.t537 28.565
R1460 VDD.n32 VDD.t56 28.565
R1461 VDD.n37 VDD.t696 28.565
R1462 VDD.n37 VDD.t694 28.565
R1463 VDD.n20 VDD.t676 28.565
R1464 VDD.n20 VDD.t675 28.565
R1465 VDD.n25 VDD.t2164 28.565
R1466 VDD.n25 VDD.t2162 28.565
R1467 VDD.n10 VDD.t490 28.565
R1468 VDD.n10 VDD.t489 28.565
R1469 VDD.n13 VDD.t1644 28.565
R1470 VDD.n13 VDD.t1646 28.565
R1471 VDD.n14 VDD.t1645 28.565
R1472 VDD.n14 VDD.t674 28.565
R1473 VDD.n9 VDD.t672 28.565
R1474 VDD.n9 VDD.t671 28.565
R1475 VDD.n2 VDD.t2169 28.565
R1476 VDD.n2 VDD.t2168 28.565
R1477 VDD.n5 VDD.t2234 28.565
R1478 VDD.n5 VDD.t2233 28.565
R1479 VDD.n6 VDD.t2232 28.565
R1480 VDD.n6 VDD.t717 28.565
R1481 VDD.n1 VDD.t887 28.565
R1482 VDD.n1 VDD.t886 28.565
R1483 VDD.n1831 VDD.t2167 28.565
R1484 VDD.n1831 VDD.t2166 28.565
R1485 VDD.n1834 VDD.t187 28.565
R1486 VDD.n1834 VDD.t543 28.565
R1487 VDD.n1835 VDD.t205 28.565
R1488 VDD.n1835 VDD.t668 28.565
R1489 VDD.n1830 VDD.t667 28.565
R1490 VDD.n1830 VDD.t666 28.565
R1491 VDD.n1840 VDD.t188 28.565
R1492 VDD.n1840 VDD.t1011 28.565
R1493 VDD.n1846 VDD.t1757 28.565
R1494 VDD.n1846 VDD.t1759 28.565
R1495 VDD.n1818 VDD.t506 28.565
R1496 VDD.n1818 VDD.t374 28.565
R1497 VDD.n1824 VDD.t320 28.565
R1498 VDD.n1824 VDD.t317 28.565
R1499 VDD.n46 VDD.t1095 28.565
R1500 VDD.n46 VDD.t1094 28.565
R1501 VDD.n42 VDD.t648 28.565
R1502 VDD.n42 VDD.t640 28.565
R1503 VDD.n43 VDD.t639 28.565
R1504 VDD.n43 VDD.t2408 28.565
R1505 VDD.n45 VDD.t2402 28.565
R1506 VDD.n45 VDD.t2401 28.565
R1507 VDD.n1792 VDD.t2410 28.565
R1508 VDD.n1792 VDD.t2409 28.565
R1509 VDD.n1797 VDD.t651 28.565
R1510 VDD.n1797 VDD.t650 28.565
R1511 VDD.n1803 VDD.t2263 28.565
R1512 VDD.n1803 VDD.t2262 28.565
R1513 VDD.n1808 VDD.t1864 28.565
R1514 VDD.n1808 VDD.t1863 28.565
R1515 VDD.n1783 VDD.t1834 28.565
R1516 VDD.n1783 VDD.t1914 28.565
R1517 VDD.n1786 VDD.t2284 28.565
R1518 VDD.n1786 VDD.t2283 28.565
R1519 VDD.n1787 VDD.t2282 28.565
R1520 VDD.n1787 VDD.t2407 28.565
R1521 VDD.n1782 VDD.t2406 28.565
R1522 VDD.n1782 VDD.t2405 28.565
R1523 VDD.n50 VDD.t655 28.565
R1524 VDD.n50 VDD.t654 28.565
R1525 VDD.n53 VDD.t1786 28.565
R1526 VDD.n53 VDD.t1785 28.565
R1527 VDD.n54 VDD.t1784 28.565
R1528 VDD.n54 VDD.t1844 28.565
R1529 VDD.n49 VDD.t1839 28.565
R1530 VDD.n49 VDD.t1807 28.565
R1531 VDD.n58 VDD.t333 28.565
R1532 VDD.n58 VDD.t335 28.565
R1533 VDD.n1716 VDD.t1457 28.565
R1534 VDD.n1716 VDD.t1455 28.565
R1535 VDD.n1715 VDD.t1660 28.565
R1536 VDD.n1715 VDD.t1658 28.565
R1537 VDD.n1712 VDD.t1648 28.565
R1538 VDD.n1712 VDD.t1664 28.565
R1539 VDD.n1713 VDD.t1652 28.565
R1540 VDD.n1713 VDD.t1650 28.565
R1541 VDD.n1689 VDD.t2136 28.565
R1542 VDD.n1689 VDD.t2028 28.565
R1543 VDD.n1684 VDD.t1792 28.565
R1544 VDD.n1684 VDD.t1794 28.565
R1545 VDD.n1685 VDD.t1930 28.565
R1546 VDD.n1685 VDD.t1978 28.565
R1547 VDD.n1687 VDD.t1992 28.565
R1548 VDD.n1687 VDD.t2012 28.565
R1549 VDD.n1679 VDD.t801 28.565
R1550 VDD.n1679 VDD.t1463 28.565
R1551 VDD.n1674 VDD.t2070 28.565
R1552 VDD.n1674 VDD.t2068 28.565
R1553 VDD.n1675 VDD.t2066 28.565
R1554 VDD.n1675 VDD.t2126 28.565
R1555 VDD.n1677 VDD.t2124 28.565
R1556 VDD.n1677 VDD.t2026 28.565
R1557 VDD.n1730 VDD.t1634 28.565
R1558 VDD.n1730 VDD.t1632 28.565
R1559 VDD.n1725 VDD.t2008 28.565
R1560 VDD.n1725 VDD.t2002 28.565
R1561 VDD.n1726 VDD.t209 28.565
R1562 VDD.n1726 VDD.t2010 28.565
R1563 VDD.n1727 VDD.t211 28.565
R1564 VDD.n1727 VDD.t138 28.565
R1565 VDD.n1639 VDD.t1275 28.565
R1566 VDD.n1639 VDD.t1271 28.565
R1567 VDD.n1634 VDD.t1862 28.565
R1568 VDD.n1634 VDD.t1818 28.565
R1569 VDD.n1621 VDD.t1868 28.565
R1570 VDD.n1621 VDD.t1858 28.565
R1571 VDD.n1607 VDD.t429 28.565
R1572 VDD.n1607 VDD.t423 28.565
R1573 VDD.n1596 VDD.t1838 28.565
R1574 VDD.n1596 VDD.t1820 28.565
R1575 VDD.n1582 VDD.t2098 28.565
R1576 VDD.n1582 VDD.t2088 28.565
R1577 VDD.n1571 VDD.t1905 28.565
R1578 VDD.n1571 VDD.t1860 28.565
R1579 VDD.n1557 VDD.t2000 28.565
R1580 VDD.n1557 VDD.t1988 28.565
R1581 VDD.n1546 VDD.t1814 28.565
R1582 VDD.n1546 VDD.t1877 28.565
R1583 VDD.n1532 VDD.t815 28.565
R1584 VDD.n1532 VDD.t805 28.565
R1585 VDD.n1521 VDD.t1899 28.565
R1586 VDD.n1521 VDD.t1872 28.565
R1587 VDD.n1507 VDD.t487 28.565
R1588 VDD.n1507 VDD.t607 28.565
R1589 VDD.n1487 VDD.t710 28.565
R1590 VDD.n1487 VDD.t706 28.565
R1591 VDD.n1482 VDD.t1879 28.565
R1592 VDD.n1482 VDD.t1833 28.565
R1593 VDD.n1471 VDD.t1901 28.565
R1594 VDD.n1471 VDD.t1887 28.565
R1595 VDD.n1457 VDD.t775 28.565
R1596 VDD.n1457 VDD.t1163 28.565
R1597 VDD.n1082 VDD.t1465 28.565
R1598 VDD.n1082 VDD.t854 28.565
R1599 VDD.n1077 VDD.t858 28.565
R1600 VDD.n1077 VDD.t771 28.565
R1601 VDD.n1078 VDD.t856 28.565
R1602 VDD.n1078 VDD.t2478 28.565
R1603 VDD.n1080 VDD.t2487 28.565
R1604 VDD.n1080 VDD.t2465 28.565
R1605 VDD.n1067 VDD.t662 28.565
R1606 VDD.n1067 VDD.t660 28.565
R1607 VDD.n1122 VDD.t797 28.565
R1608 VDD.n1122 VDD.t795 28.565
R1609 VDD.n1103 VDD.t1357 28.565
R1610 VDD.n1103 VDD.t1345 28.565
R1611 VDD.n1073 VDD.t1200 28.565
R1612 VDD.n1073 VDD.t1221 28.565
R1613 VDD.n1074 VDD.t1202 28.565
R1614 VDD.n1074 VDD.t1696 28.565
R1615 VDD.n1102 VDD.t1704 28.565
R1616 VDD.n1102 VDD.t1692 28.565
R1617 VDD.n1003 VDD.t83 28.565
R1618 VDD.n1003 VDD.t81 28.565
R1619 VDD.n1152 VDD.t89 28.565
R1620 VDD.n1152 VDD.t91 28.565
R1621 VDD.n1137 VDD.t1038 28.565
R1622 VDD.n1137 VDD.t1104 28.565
R1623 VDD.n1008 VDD.t2320 28.565
R1624 VDD.n1008 VDD.t2322 28.565
R1625 VDD.n1009 VDD.t2324 28.565
R1626 VDD.n1009 VDD.t941 28.565
R1627 VDD.n1136 VDD.t688 28.565
R1628 VDD.n1136 VDD.t937 28.565
R1629 VDD.n940 VDD.t1081 28.565
R1630 VDD.n940 VDD.t1083 28.565
R1631 VDD.n1182 VDD.t163 28.565
R1632 VDD.n1182 VDD.t347 28.565
R1633 VDD.n1166 VDD.t839 28.565
R1634 VDD.n1166 VDD.t827 28.565
R1635 VDD.n945 VDD.t595 28.565
R1636 VDD.n945 VDD.t597 28.565
R1637 VDD.n946 VDD.t593 28.565
R1638 VDD.n946 VDD.t2219 28.565
R1639 VDD.n1165 VDD.t2205 28.565
R1640 VDD.n1165 VDD.t2213 28.565
R1641 VDD.n1202 VDD.t1583 28.565
R1642 VDD.n1202 VDD.t1593 28.565
R1643 VDD.n1201 VDD.t1330 28.565
R1644 VDD.n1201 VDD.t1338 28.565
R1645 VDD.n1198 VDD.t319 28.565
R1646 VDD.n1198 VDD.t1324 28.565
R1647 VDD.n1199 VDD.t437 28.565
R1648 VDD.n1199 VDD.t371 28.565
R1649 VDD.n1211 VDD.t156 28.565
R1650 VDD.n1211 VDD.t362 28.565
R1651 VDD.n1218 VDD.t1126 28.565
R1652 VDD.n1218 VDD.t1124 28.565
R1653 VDD.n1090 VDD.t2084 28.565
R1654 VDD.n1090 VDD.t2106 28.565
R1655 VDD.n1085 VDD.t2016 28.565
R1656 VDD.n1085 VDD.t2018 28.565
R1657 VDD.n1086 VDD.t2014 28.565
R1658 VDD.n1086 VDD.t1609 28.565
R1659 VDD.n1088 VDD.t1626 28.565
R1660 VDD.n1088 VDD.t1639 28.565
R1661 VDD.n807 VDD.t1475 28.565
R1662 VDD.n807 VDD.t1473 28.565
R1663 VDD.n806 VDD.t1471 28.565
R1664 VDD.n806 VDD.t2141 28.565
R1665 VDD.n805 VDD.t2034 28.565
R1666 VDD.n805 VDD.t2139 28.565
R1667 VDD.n810 VDD.t21 28.565
R1668 VDD.n810 VDD.t758 28.565
R1669 VDD.n817 VDD.t2229 28.565
R1670 VDD.n817 VDD.t2231 28.565
R1671 VDD.n816 VDD.t2174 28.565
R1672 VDD.n816 VDD.t2472 28.565
R1673 VDD.n815 VDD.t2470 28.565
R1674 VDD.n815 VDD.t2494 28.565
R1675 VDD.n820 VDD.t2104 28.565
R1676 VDD.n820 VDD.t2112 28.565
R1677 VDD.n444 VDD.t2502 28.565
R1678 VDD.n444 VDD.t2500 28.565
R1679 VDD.n439 VDD.t2398 28.565
R1680 VDD.n439 VDD.t2396 28.565
R1681 VDD.n440 VDD.t2394 28.565
R1682 VDD.n440 VDD.t2108 28.565
R1683 VDD.n442 VDD.t2102 28.565
R1684 VDD.n442 VDD.t2096 28.565
R1685 VDD.n435 VDD.t1643 28.565
R1686 VDD.n435 VDD.t1616 28.565
R1687 VDD.n430 VDD.t1146 28.565
R1688 VDD.n430 VDD.t1148 28.565
R1689 VDD.n431 VDD.t1144 28.565
R1690 VDD.n431 VDD.t803 28.565
R1691 VDD.n433 VDD.t1359 28.565
R1692 VDD.n433 VDD.t1461 28.565
R1693 VDD.n793 VDD.t1612 28.565
R1694 VDD.n793 VDD.t1628 28.565
R1695 VDD.n788 VDD.t867 28.565
R1696 VDD.n788 VDD.t1435 28.565
R1697 VDD.n789 VDD.t865 28.565
R1698 VDD.n789 VDD.t17 28.565
R1699 VDD.n791 VDD.t754 28.565
R1700 VDD.n791 VDD.t291 28.565
R1701 VDD.n802 VDD.t126 28.565
R1702 VDD.n802 VDD.t427 28.565
R1703 VDD.n797 VDD.t109 28.565
R1704 VDD.n797 VDD.t365 28.565
R1705 VDD.n798 VDD.t314 28.565
R1706 VDD.n798 VDD.t2509 28.565
R1707 VDD.n800 VDD.t2356 28.565
R1708 VDD.n800 VDD.t2364 28.565
R1709 VDD.n505 VDD.t342 28.565
R1710 VDD.n505 VDD.t340 28.565
R1711 VDD.n776 VDD.t326 28.565
R1712 VDD.n776 VDD.t324 28.565
R1713 VDD.n756 VDD.t382 28.565
R1714 VDD.n756 VDD.t386 28.565
R1715 VDD.n511 VDD.t246 28.565
R1716 VDD.n511 VDD.t496 28.565
R1717 VDD.n512 VDD.t373 28.565
R1718 VDD.n512 VDD.t1783 28.565
R1719 VDD.n755 VDD.t1773 28.565
R1720 VDD.n755 VDD.t1769 28.565
R1721 VDD.n576 VDD.t1754 28.565
R1722 VDD.n576 VDD.t1752 28.565
R1723 VDD.n569 VDD.t26 28.565
R1724 VDD.n569 VDD.t111 28.565
R1725 VDD.n733 VDD.t186 28.565
R1726 VDD.n733 VDD.t417 28.565
R1727 VDD.n582 VDD.t227 28.565
R1728 VDD.n582 VDD.t166 28.565
R1729 VDD.n583 VDD.t482 28.565
R1730 VDD.n583 VDD.t2380 28.565
R1731 VDD.n732 VDD.t2378 28.565
R1732 VDD.n732 VDD.t2390 28.565
R1733 VDD.n658 VDD.t2613 28.565
R1734 VDD.n658 VDD.t2611 28.565
R1735 VDD.n648 VDD.t2042 28.565
R1736 VDD.n648 VDD.t2060 28.565
R1737 VDD.n647 VDD.t727 28.565
R1738 VDD.n647 VDD.t721 28.565
R1739 VDD.n644 VDD.t2020 28.565
R1740 VDD.n644 VDD.t731 28.565
R1741 VDD.n645 VDD.t2024 28.565
R1742 VDD.n645 VDD.t2022 28.565
R1743 VDD.n1703 VDD.t316 28.565
R1744 VDD.n1703 VDD.t300 28.565
R1745 VDD.n1696 VDD.t1363 28.565
R1746 VDD.n1696 VDD.t1361 28.565
R1747 VDD.n587 VDD.t1302 28.565
R1748 VDD.n587 VDD.t1312 28.565
R1749 VDD.n592 VDD.t700 28.565
R1750 VDD.n592 VDD.t992 28.565
R1751 VDD.n622 VDD.t1668 28.565
R1752 VDD.n622 VDD.t1666 28.565
R1753 VDD.n627 VDD.t1453 28.565
R1754 VDD.n627 VDD.t1441 28.565
R1755 VDD.n614 VDD.t367 28.565
R1756 VDD.n614 VDD.t1003 28.565
R1757 VDD.n596 VDD.t1024 28.565
R1758 VDD.n596 VDD.t1028 28.565
R1759 VDD.n597 VDD.t1026 28.565
R1760 VDD.n597 VDD.t1662 28.565
R1761 VDD.n613 VDD.t1674 28.565
R1762 VDD.n613 VDD.t1672 28.565
R1763 VDD.n605 VDD.t1443 28.565
R1764 VDD.n605 VDD.t1459 28.565
R1765 VDD.n600 VDD.t146 28.565
R1766 VDD.n600 VDD.t402 28.565
R1767 VDD.n601 VDD.t678 28.565
R1768 VDD.n601 VDD.t925 28.565
R1769 VDD.n604 VDD.t462 28.565
R1770 VDD.n604 VDD.t977 28.565
R1771 VDD.n666 VDD.t69 28.565
R1772 VDD.n666 VDD.t304 28.565
R1773 VDD.n711 VDD.t1250 28.565
R1774 VDD.n711 VDD.t1248 28.565
R1775 VDD.n716 VDD.t199 28.565
R1776 VDD.n716 VDD.t197 28.565
R1777 VDD.n698 VDD.t739 28.565
R1778 VDD.n698 VDD.t737 28.565
R1779 VDD.n703 VDD.t2064 28.565
R1780 VDD.n703 VDD.t2052 28.565
R1781 VDD.n689 VDD.t1193 28.565
R1782 VDD.n689 VDD.t1191 28.565
R1783 VDD.n672 VDD.t435 28.565
R1784 VDD.n672 VDD.t379 28.565
R1785 VDD.n673 VDD.t159 28.565
R1786 VDD.n673 VDD.t729 28.565
R1787 VDD.n688 VDD.t725 28.565
R1788 VDD.n688 VDD.t743 28.565
R1789 VDD.n677 VDD.t2048 28.565
R1790 VDD.n677 VDD.t2044 28.565
R1791 VDD.n682 VDD.t1051 28.565
R1792 VDD.n682 VDD.t1053 28.565
R1793 VDD.n683 VDD.t1049 28.565
R1794 VDD.n683 VDD.t201 28.565
R1795 VDD.n676 VDD.t1195 28.565
R1796 VDD.n676 VDD.t791 28.565
R1797 VDD.n558 VDD.t182 28.565
R1798 VDD.n558 VDD.t180 28.565
R1799 VDD.n563 VDD.t2535 28.565
R1800 VDD.n563 VDD.t2533 28.565
R1801 VDD.n539 VDD.t2384 28.565
R1802 VDD.n539 VDD.t2382 28.565
R1803 VDD.n544 VDD.t358 28.565
R1804 VDD.n544 VDD.t97 28.565
R1805 VDD.n530 VDD.t2545 28.565
R1806 VDD.n530 VDD.t2543 28.565
R1807 VDD.n514 VDD.t2281 28.565
R1808 VDD.n514 VDD.t2279 28.565
R1809 VDD.n515 VDD.t2277 28.565
R1810 VDD.n515 VDD.t2370 28.565
R1811 VDD.n529 VDD.t2392 28.565
R1812 VDD.n529 VDD.t2388 28.565
R1813 VDD.n518 VDD.t354 28.565
R1814 VDD.n518 VDD.t860 28.565
R1815 VDD.n523 VDD.t2606 28.565
R1816 VDD.n523 VDD.t2599 28.565
R1817 VDD.n524 VDD.t2601 28.565
R1818 VDD.n524 VDD.t2525 28.565
R1819 VDD.n517 VDD.t2529 28.565
R1820 VDD.n517 VDD.t2523 28.565
R1821 VDD.n1373 VDD.t2040 28.565
R1822 VDD.n1373 VDD.t2038 28.565
R1823 VDD.n1368 VDD.t2076 28.565
R1824 VDD.n1368 VDD.t2074 28.565
R1825 VDD.n1369 VDD.t2072 28.565
R1826 VDD.n1369 VDD.t2094 28.565
R1827 VDD.n1371 VDD.t2092 28.565
R1828 VDD.n1371 VDD.t2082 28.565
R1829 VDD.n1365 VDD.t2496 28.565
R1830 VDD.n1365 VDD.t2492 28.565
R1831 VDD.n1360 VDD.t907 28.565
R1832 VDD.n1360 VDD.t338 28.565
R1833 VDD.n1361 VDD.t289 28.565
R1834 VDD.n1361 VDD.t124 28.565
R1835 VDD.n1363 VDD.t551 28.565
R1836 VDD.n1363 VDD.t549 28.565
R1837 VDD.n1670 VDD.t1986 28.565
R1838 VDD.n1670 VDD.t1996 28.565
R1839 VDD.n1665 VDD.t268 28.565
R1840 VDD.n1665 VDD.t47 28.565
R1841 VDD.n1666 VDD.t351 28.565
R1842 VDD.n1666 VDD.t2498 28.565
R1843 VDD.n1668 VDD.t2484 28.565
R1844 VDD.n1668 VDD.t2482 28.565
R1845 VDD.n1357 VDD.t813 28.565
R1846 VDD.n1357 VDD.t811 28.565
R1847 VDD.n1352 VDD.t702 28.565
R1848 VDD.n1352 VDD.t1207 28.565
R1849 VDD.n1353 VDD.t1205 28.565
R1850 VDD.n1353 VDD.t2361 28.565
R1851 VDD.n1355 VDD.t2516 28.565
R1852 VDD.n1355 VDD.t2512 28.565
R1853 VDD.n1386 VDD.t2186 28.565
R1854 VDD.n1386 VDD.t2184 28.565
R1855 VDD.n1381 VDD.t1967 28.565
R1856 VDD.n1381 VDD.t1961 28.565
R1857 VDD.n1392 VDD.t1973 28.565
R1858 VDD.n1392 VDD.t1971 28.565
R1859 VDD.n1394 VDD.t1185 28.565
R1860 VDD.n1394 VDD.t1183 28.565
R1861 VDD.n1395 VDD.t1181 28.565
R1862 VDD.n1395 VDD.t2188 28.565
R1863 VDD.n1397 VDD.t2182 28.565
R1864 VDD.n1397 VDD.t2180 28.565
R1865 VDD.n1291 VDD.t410 28.565
R1866 VDD.n1291 VDD.t45 28.565
R1867 VDD.n1283 VDD.t1503 28.565
R1868 VDD.n1282 VDD.t1481 28.565
R1869 VDD.n1282 VDD.t1547 28.565
R1870 VDD.n1309 VDD.t1287 28.565
R1871 VDD.n1309 VDD.t1285 28.565
R1872 VDD.n1301 VDD.t1569 28.565
R1873 VDD.n1300 VDD.t1521 28.565
R1874 VDD.n1300 VDD.t1571 28.565
R1875 VDD.n1326 VDD.t957 28.565
R1876 VDD.n1326 VDD.t955 28.565
R1877 VDD.n1318 VDD.t1497 28.565
R1878 VDD.n1317 VDD.t1553 28.565
R1879 VDD.n1317 VDD.t1517 28.565
R1880 VDD.n1343 VDD.t140 28.565
R1881 VDD.n1343 VDD.t988 28.565
R1882 VDD.n1335 VDD.t1515 28.565
R1883 VDD.n1334 VDD.t1565 28.565
R1884 VDD.n1334 VDD.t1527 28.565
R1885 VDD.n1249 VDD.t105 28.565
R1886 VDD.n1249 VDD.t377 28.565
R1887 VDD.n1244 VDD.t2160 28.565
R1888 VDD.n1244 VDD.t2158 28.565
R1889 VDD.n1261 VDD.t2156 28.565
R1890 VDD.n1261 VDD.t2144 28.565
R1891 VDD.n1256 VDD.t2120 28.565
R1892 VDD.n1256 VDD.t2122 28.565
R1893 VDD.n1257 VDD.t2118 28.565
R1894 VDD.n1257 VDD.t478 28.565
R1895 VDD.n1259 VDD.t546 28.565
R1896 VDD.n1259 VDD.t994 28.565
R1897 VDD.n1235 VDD.t1179 28.565
R1898 VDD.n1235 VDD.t1211 28.565
R1899 VDD.n1230 VDD.t2580 28.565
R1900 VDD.n1230 VDD.t2572 28.565
R1901 VDD.n427 VDD.t2006 28.565
R1902 VDD.n427 VDD.t1982 28.565
R1903 VDD.n422 VDD.t398 28.565
R1904 VDD.n422 VDD.t638 28.565
R1905 VDD.n423 VDD.t396 28.565
R1906 VDD.n423 VDD.t2359 28.565
R1907 VDD.n425 VDD.t2507 28.565
R1908 VDD.n425 VDD.t2514 28.565
R1909 VDD.n417 VDD.t2578 28.565
R1910 VDD.n417 VDD.t2582 28.565
R1911 VDD.n412 VDD.t1215 28.565
R1912 VDD.n412 VDD.t1102 28.565
R1913 VDD.n413 VDD.t1167 28.565
R1914 VDD.n413 VDD.t1177 28.565
R1915 VDD.n414 VDD.t1093 28.565
R1916 VDD.n414 VDD.t1165 28.565
R1917 VDD.n394 VDD.t2549 28.565
R1918 VDD.n394 VDD.t2547 28.565
R1919 VDD.n389 VDD.t1388 28.565
R1920 VDD.n389 VDD.t1392 28.565
R1921 VDD.n406 VDD.t1400 28.565
R1922 VDD.n406 VDD.t1398 28.565
R1923 VDD.n401 VDD.t2462 28.565
R1924 VDD.n401 VDD.t2454 28.565
R1925 VDD.n402 VDD.t2450 28.565
R1926 VDD.n402 VDD.t2553 28.565
R1927 VDD.n403 VDD.t2275 28.565
R1928 VDD.n403 VDD.t2452 28.565
R1929 VDD.n1412 VDD.t131 28.565
R1930 VDD.n1412 VDD.t135 28.565
R1931 VDD.n1404 VDD.t1485 28.565
R1932 VDD.n1403 VDD.t1541 28.565
R1933 VDD.n1403 VDD.t1501 28.565
R1934 VDD.n1429 VDD.t628 28.565
R1935 VDD.n1429 VDD.t632 28.565
R1936 VDD.n1421 VDD.t1561 28.565
R1937 VDD.n1420 VDD.t1509 28.565
R1938 VDD.n1420 VDD.t1499 28.565
R1939 VDD.n379 VDD.t1935 28.565
R1940 VDD.n379 VDD.t1933 28.565
R1941 VDD.n371 VDD.t1505 28.565
R1942 VDD.n370 VDD.t1487 28.565
R1943 VDD.n370 VDD.t1543 28.565
R1944 VDD.n172 VDD.t483 28.565
R1945 VDD.n172 VDD.t926 28.565
R1946 VDD.n177 VDD.t2441 28.565
R1947 VDD.n177 VDD.t2440 28.565
R1948 VDD.n120 VDD.t129 28.565
R1949 VDD.n120 VDD.t359 28.565
R1950 VDD.n115 VDD.t781 28.565
R1951 VDD.n115 VDD.t780 28.565
R1952 VDD.n71 VDD.t77 28.565
R1953 VDD.n71 VDD.t76 28.565
R1954 VDD.n72 VDD.t1941 28.565
R1955 VDD.n72 VDD.t642 28.565
R1956 VDD.n68 VDD.t910 28.565
R1957 VDD.n68 VDD.t147 28.565
R1958 VDD.n67 VDD.t1947 28.565
R1959 VDD.n67 VDD.t1942 28.565
R1960 VDD.n128 VDD.t2443 28.565
R1961 VDD.n128 VDD.t2442 28.565
R1962 VDD.n129 VDD.t819 28.565
R1963 VDD.n129 VDD.t2444 28.565
R1964 VDD.n125 VDD.t2490 28.565
R1965 VDD.n125 VDD.t2489 28.565
R1966 VDD.n124 VDD.t818 28.565
R1967 VDD.n124 VDD.t1255 28.565
R1968 VDD.n185 VDD.t657 28.565
R1969 VDD.n185 VDD.t656 28.565
R1970 VDD.n186 VDD.t1371 28.565
R1971 VDD.n186 VDD.t658 28.565
R1972 VDD.n182 VDD.t2030 28.565
R1973 VDD.n182 VDD.t2029 28.565
R1974 VDD.n181 VDD.t1373 28.565
R1975 VDD.n181 VDD.t1372 28.565
R1976 VDD.n242 VDD.t777 28.565
R1977 VDD.n242 VDD.t776 28.565
R1978 VDD.n243 VDD.t1407 28.565
R1979 VDD.n243 VDD.t778 28.565
R1980 VDD.n239 VDD.t1613 28.565
R1981 VDD.n239 VDD.t1610 28.565
R1982 VDD.n238 VDD.t1401 28.565
R1983 VDD.n238 VDD.t1409 28.565
R1984 VDD.n234 VDD.t445 28.565
R1985 VDD.n234 VDD.t444 28.565
R1986 VDD.n229 VDD.t524 28.565
R1987 VDD.n229 VDD.t460 28.565
R1988 VDD.n63 VDD.t2291 28.565
R1989 VDD.n63 VDD.t2310 28.565
R1990 VDD.n81 VDD.t2473 28.565
R1991 VDD.n81 VDD.t2468 28.565
R1992 VDD.n76 VDD.t568 28.565
R1993 VDD.n76 VDD.t1256 28.565
R1994 VDD.n109 VDD.t2584 28.565
R1995 VDD.n109 VDD.t2586 28.565
R1996 VDD.n104 VDD.t473 28.565
R1997 VDD.n104 VDD.t471 28.565
R1998 VDD.n89 VDD.t2607 28.565
R1999 VDD.n89 VDD.t2318 28.565
R2000 VDD.n90 VDD.t1208 28.565
R2001 VDD.n90 VDD.t2602 28.565
R2002 VDD.n86 VDD.t2563 28.565
R2003 VDD.n86 VDD.t2585 28.565
R2004 VDD.n85 VDD.t588 28.565
R2005 VDD.n85 VDD.t587 28.565
R2006 VDD.n92 VDD.t280 28.565
R2007 VDD.n92 VDD.t279 28.565
R2008 VDD.n93 VDD.t2564 28.565
R2009 VDD.n93 VDD.t281 28.565
R2010 VDD.n96 VDD.t2476 28.565
R2011 VDD.n96 VDD.t2475 28.565
R2012 VDD.n95 VDD.t2560 28.565
R2013 VDD.n95 VDD.t2561 28.565
R2014 VDD.n138 VDD.t2032 28.565
R2015 VDD.n138 VDD.t2031 28.565
R2016 VDD.n133 VDD.t1379 28.565
R2017 VDD.n133 VDD.t1378 28.565
R2018 VDD.n166 VDD.t2200 28.565
R2019 VDD.n166 VDD.t2199 28.565
R2020 VDD.n161 VDD.t562 28.565
R2021 VDD.n161 VDD.t561 28.565
R2022 VDD.n146 VDD.t862 28.565
R2023 VDD.n146 VDD.t118 28.565
R2024 VDD.n147 VDD.t1374 28.565
R2025 VDD.n147 VDD.t863 28.565
R2026 VDD.n143 VDD.t2194 28.565
R2027 VDD.n143 VDD.t2202 28.565
R2028 VDD.n142 VDD.t1376 28.565
R2029 VDD.n142 VDD.t1375 28.565
R2030 VDD.n149 VDD.t690 28.565
R2031 VDD.n149 VDD.t689 28.565
R2032 VDD.n150 VDD.t2196 28.565
R2033 VDD.n150 VDD.t691 28.565
R2034 VDD.n153 VDD.t2131 28.565
R2035 VDD.n153 VDD.t2130 28.565
R2036 VDD.n152 VDD.t2198 28.565
R2037 VDD.n152 VDD.t2197 28.565
R2038 VDD.n195 VDD.t1621 28.565
R2039 VDD.n195 VDD.t1619 28.565
R2040 VDD.n190 VDD.t1402 28.565
R2041 VDD.n190 VDD.t1404 28.565
R2042 VDD.n223 VDD.t918 28.565
R2043 VDD.n223 VDD.t917 28.565
R2044 VDD.n218 VDD.t1925 28.565
R2045 VDD.n218 VDD.t1924 28.565
R2046 VDD.n203 VDD.t786 28.565
R2047 VDD.n203 VDD.t785 28.565
R2048 VDD.n204 VDD.t1412 28.565
R2049 VDD.n204 VDD.t1173 28.565
R2050 VDD.n200 VDD.t915 28.565
R2051 VDD.n200 VDD.t912 28.565
R2052 VDD.n199 VDD.t1411 28.565
R2053 VDD.n199 VDD.t1410 28.565
R2054 VDD.n206 VDD.t1974 28.565
R2055 VDD.n206 VDD.t1976 28.565
R2056 VDD.n207 VDD.t911 28.565
R2057 VDD.n207 VDD.t1975 28.565
R2058 VDD.n210 VDD.t1636 28.565
R2059 VDD.n210 VDD.t1635 28.565
R2060 VDD.n209 VDD.t913 28.565
R2061 VDD.n209 VDD.t922 28.565
R2062 VDD.n359 VDD.t1018 28.565
R2063 VDD.n359 VDD.t1017 28.565
R2064 VDD.n364 VDD.t447 28.565
R2065 VDD.n364 VDD.t446 28.565
R2066 VDD.n347 VDD.t1806 28.565
R2067 VDD.n347 VDD.t1803 28.565
R2068 VDD.n352 VDD.t2505 28.565
R2069 VDD.n352 VDD.t2362 28.565
R2070 VDD.n337 VDD.t450 28.565
R2071 VDD.n337 VDD.t449 28.565
R2072 VDD.n340 VDD.t1172 28.565
R2073 VDD.n340 VDD.t1171 28.565
R2074 VDD.n341 VDD.t1170 28.565
R2075 VDD.n341 VDD.t1804 28.565
R2076 VDD.n336 VDD.t1805 28.565
R2077 VDD.n336 VDD.t1799 28.565
R2078 VDD.n329 VDD.t2357 28.565
R2079 VDD.n329 VDD.t2519 28.565
R2080 VDD.n332 VDD.t415 28.565
R2081 VDD.n332 VDD.t414 28.565
R2082 VDD.n333 VDD.t413 28.565
R2083 VDD.n333 VDD.t468 28.565
R2084 VDD.n328 VDD.t470 28.565
R2085 VDD.n328 VDD.t469 28.565
R2086 VDD.n317 VDD.t971 28.565
R2087 VDD.n317 VDD.t970 28.565
R2088 VDD.n323 VDD.t1020 28.565
R2089 VDD.n323 VDD.t1022 28.565
R2090 VDD.n308 VDD.t2354 28.565
R2091 VDD.n308 VDD.t2510 28.565
R2092 VDD.n311 VDD.t212 28.565
R2093 VDD.n311 VDD.t232 28.565
R2094 VDD.n312 VDD.t927 28.565
R2095 VDD.n312 VDD.t1800 28.565
R2096 VDD.n307 VDD.t1802 28.565
R2097 VDD.n307 VDD.t1801 28.565
R2098 VDD.n301 VDD.t1140 28.565
R2099 VDD.n301 VDD.t1141 28.565
R2100 VDD.n295 VDD.t1299 28.565
R2101 VDD.n295 VDD.t1298 28.565
R2102 VDD.n287 VDD.t70 28.565
R2103 VDD.n287 VDD.t619 28.565
R2104 VDD.n290 VDD.t50 28.565
R2105 VDD.n290 VDD.t213 28.565
R2106 VDD.n291 VDD.t48 28.565
R2107 VDD.n291 VDD.t574 28.565
R2108 VDD.n286 VDD.t573 28.565
R2109 VDD.n286 VDD.t580 28.565
R2110 VDD.n276 VDD.t1416 28.565
R2111 VDD.n276 VDD.t1415 28.565
R2112 VDD.n281 VDD.t1922 28.565
R2113 VDD.n281 VDD.t1918 28.565
R2114 VDD.n264 VDD.t579 28.565
R2115 VDD.n264 VDD.t578 28.565
R2116 VDD.n269 VDD.t73 28.565
R2117 VDD.n269 VDD.t72 28.565
R2118 VDD.n254 VDD.t1954 28.565
R2119 VDD.n254 VDD.t1952 28.565
R2120 VDD.n257 VDD.t63 28.565
R2121 VDD.n257 VDD.t34 28.565
R2122 VDD.n258 VDD.t345 28.565
R2123 VDD.n258 VDD.t575 28.565
R2124 VDD.n253 VDD.t571 28.565
R2125 VDD.n253 VDD.t570 28.565
R2126 VDD.n246 VDD.t617 28.565
R2127 VDD.n246 VDD.t616 28.565
R2128 VDD.n249 VDD.t252 28.565
R2129 VDD.n249 VDD.t964 28.565
R2130 VDD.n250 VDD.t963 28.565
R2131 VDD.n250 VDD.t1916 28.565
R2132 VDD.n245 VDD.t1915 28.565
R2133 VDD.n245 VDD.t1953 28.565
R2134 VDD.n1274 VDD.t1258 28.565
R2135 VDD.n1274 VDD.t1219 28.565
R2136 VDD.n1266 VDD.t1555 28.565
R2137 VDD.n1265 VDD.t1519 28.565
R2138 VDD.n1265 VDD.t1493 28.565
R2139 VDD.n494 VDD.t221 28.565
R2140 VDD.n494 VDD.t541 28.565
R2141 VDD.n499 VDD.t1266 28.565
R2142 VDD.n499 VDD.t1264 28.565
R2143 VDD.n476 VDD.t1765 28.565
R2144 VDD.n476 VDD.t1779 28.565
R2145 VDD.n481 VDD.t217 28.565
R2146 VDD.n481 VDD.t529 28.565
R2147 VDD.n460 VDD.t1228 28.565
R2148 VDD.n460 VDD.t1226 28.565
R2149 VDD.n464 VDD.t7 28.565
R2150 VDD.n464 VDD.t494 28.565
R2151 VDD.n465 VDD.t492 28.565
R2152 VDD.n465 VDD.t1781 28.565
R2153 VDD.n459 VDD.t1771 28.565
R2154 VDD.n459 VDD.t1763 28.565
R2155 VDD.n448 VDD.t154 28.565
R2156 VDD.n448 VDD.t369 28.565
R2157 VDD.n453 VDD.t485 28.565
R2158 VDD.n453 VDD.t330 28.565
R2159 VDD.n454 VDD.t332 28.565
R2160 VDD.n454 VDD.t1234 28.565
R2161 VDD.n447 VDD.t1238 28.565
R2162 VDD.n447 VDD.t1230 28.565
R2163 VDD.n872 VDD.t599 28.565
R2164 VDD.n872 VDD.t961 28.565
R2165 VDD.n877 VDD.t2236 28.565
R2166 VDD.n877 VDD.t2240 28.565
R2167 VDD.n853 VDD.t1334 28.565
R2168 VDD.n853 VDD.t1326 28.565
R2169 VDD.n858 VDD.t1581 28.565
R2170 VDD.n858 VDD.t1575 28.565
R2171 VDD.n845 VDD.t2246 28.565
R2172 VDD.n845 VDD.t2256 28.565
R2173 VDD.n829 VDD.t1059 28.565
R2174 VDD.n829 VDD.t1061 28.565
R2175 VDD.n830 VDD.t1063 28.565
R2176 VDD.n830 VDD.t1316 28.565
R2177 VDD.n844 VDD.t1336 28.565
R2178 VDD.n844 VDD.t1322 28.565
R2179 VDD.n836 VDD.t1573 28.565
R2180 VDD.n836 VDD.t1587 28.565
R2181 VDD.n835 VDD.t2242 28.565
R2182 VDD.n835 VDD.t2248 28.565
R2183 VDD.n832 VDD.t889 28.565
R2184 VDD.n832 VDD.t2252 28.565
R2185 VDD.n833 VDD.t891 28.565
R2186 VDD.n833 VDD.t223 28.565
R2187 VDD.n884 VDD.t879 28.565
R2188 VDD.n884 VDD.t871 28.565
R2189 VDD.n889 VDD.t1738 28.565
R2190 VDD.n889 VDD.t1730 28.565
R2191 VDD.n921 VDD.t2211 28.565
R2192 VDD.n921 VDD.t2223 28.565
R2193 VDD.n926 VDD.t823 28.565
R2194 VDD.n926 VDD.t58 28.565
R2195 VDD.n905 VDD.t1722 28.565
R2196 VDD.n905 VDD.t1732 28.565
R2197 VDD.n910 VDD.t1712 28.565
R2198 VDD.n910 VDD.t1684 28.565
R2199 VDD.n911 VDD.t1686 28.565
R2200 VDD.n911 VDD.t2221 28.565
R2201 VDD.n904 VDD.t2207 28.565
R2202 VDD.n904 VDD.t2217 28.565
R2203 VDD.n897 VDD.t833 28.565
R2204 VDD.n897 VDD.t60 28.565
R2205 VDD.n896 VDD.t1742 28.565
R2206 VDD.n896 VDD.t1726 28.565
R2207 VDD.n893 VDD.t1030 28.565
R2208 VDD.n893 VDD.t1734 28.565
R2209 VDD.n894 VDD.t1032 28.565
R2210 VDD.n894 VDD.t1116 28.565
R2211 VDD.n950 VDD.t2331 28.565
R2212 VDD.n950 VDD.t2335 28.565
R2213 VDD.n955 VDD.t2424 28.565
R2214 VDD.n955 VDD.t2432 28.565
R2215 VDD.n984 VDD.t933 28.565
R2216 VDD.n984 VDD.t680 28.565
R2217 VDD.n989 VDD.t1108 28.565
R2218 VDD.n989 VDD.t1036 28.565
R2219 VDD.n975 VDD.t2422 28.565
R2220 VDD.n975 VDD.t2430 28.565
R2221 VDD.n959 VDD.t1292 28.565
R2222 VDD.n959 VDD.t388 28.565
R2223 VDD.n960 VDD.t390 28.565
R2224 VDD.n960 VDD.t684 28.565
R2225 VDD.n974 VDD.t929 28.565
R2226 VDD.n974 VDD.t939 28.565
R2227 VDD.n966 VDD.t1114 28.565
R2228 VDD.n966 VDD.t1040 28.565
R2229 VDD.n965 VDD.t2420 28.565
R2230 VDD.n965 VDD.t2434 28.565
R2231 VDD.n962 VDD.t278 28.565
R2232 VDD.n962 VDD.t2436 28.565
R2233 VDD.n963 VDD.t698 28.565
R2234 VDD.n963 VDD.t276 28.565
R2235 VDD.n1013 VDD.t2299 28.565
R2236 VDD.n1013 VDD.t2301 28.565
R2237 VDD.n1018 VDD.t1065 28.565
R2238 VDD.n1018 VDD.t843 28.565
R2239 VDD.n1048 VDD.t1688 28.565
R2240 VDD.n1048 VDD.t1698 28.565
R2241 VDD.n1053 VDD.t1343 28.565
R2242 VDD.n1053 VDD.t1351 28.565
R2243 VDD.n1040 VDD.t1071 28.565
R2244 VDD.n1040 VDD.t841 28.565
R2245 VDD.n1033 VDD.t2309 28.565
R2246 VDD.n1033 VDD.t2307 28.565
R2247 VDD.n1034 VDD.t2305 28.565
R2248 VDD.n1034 VDD.t1702 28.565
R2249 VDD.n1039 VDD.t1710 28.565
R2250 VDD.n1039 VDD.t1694 28.565
R2251 VDD.n1026 VDD.t1349 28.565
R2252 VDD.n1026 VDD.t453 28.565
R2253 VDD.n1025 VDD.t1067 28.565
R2254 VDD.n1025 VDD.t1075 28.565
R2255 VDD.n1022 VDD.t2271 28.565
R2256 VDD.n1022 VDD.t610 28.565
R2257 VDD.n1023 VDD.t2273 28.565
R2258 VDD.n1023 VDD.t2269 28.565
R2259 VDD.n1757 VDD.t1949 28.565
R2260 VDD.n1757 VDD.t1946 28.565
R2261 VDD.n1752 VDD.t451 28.565
R2262 VDD.n1752 VDD.t965 28.565
R2263 VDD.n1746 VDD.t2590 28.565
R2264 VDD.n1746 VDD.t2592 28.565
R2265 VDD.n1741 VDD.t1428 28.565
R2266 VDD.n1741 VDD.t1429 28.565
R2267 VDD.n1765 VDD.t1432 28.565
R2268 VDD.n1765 VDD.t1433 28.565
R2269 VDD.n1766 VDD.t1943 28.565
R2270 VDD.n1766 VDD.t1431 28.565
R2271 VDD.n1762 VDD.t1423 28.565
R2272 VDD.n1762 VDD.t1424 28.565
R2273 VDD.n1761 VDD.t1948 28.565
R2274 VDD.n1761 VDD.t1944 28.565
R2275 VDD.n1768 VDD.t116 28.565
R2276 VDD.n1768 VDD.t978 28.565
R2277 VDD.n1769 VDD.t1420 28.565
R2278 VDD.n1769 VDD.t975 28.565
R2279 VDD.n1772 VDD.t206 28.565
R2280 VDD.n1772 VDD.t909 28.565
R2281 VDD.n1771 VDD.t1419 28.565
R2282 VDD.n1771 VDD.t1421 28.565
R2283 VDD.n636 VDD.t1307 23.418
R2284 VDD.n724 VDD.t1245 23.418
R2285 VDD.n553 VDD.t177 23.418
R2286 VDD.n490 VDD.t265 23.418
R2287 VDD.n867 VDD.t66 23.418
R2288 VDD.n935 VDD.t872 23.418
R2289 VDD.n998 VDD.t2332 23.418
R2290 VDD.n1062 VDD.t2302 23.418
R2291 VDD.n1683 VDD.t2135 23.317
R2292 VDD.n1673 VDD.t800 23.317
R2293 VDD.n1724 VDD.t1633 23.317
R2294 VDD.n1076 VDD.t1464 23.317
R2295 VDD.n813 VDD.t20 23.317
R2296 VDD.n823 VDD.t2103 23.317
R2297 VDD.n438 VDD.t2501 23.317
R2298 VDD.n429 VDD.t1642 23.317
R2299 VDD.n787 VDD.t1611 23.317
R2300 VDD.n796 VDD.t125 23.317
R2301 VDD.n1367 VDD.t2039 23.317
R2302 VDD.n1359 VDD.t2495 23.317
R2303 VDD.n1664 VDD.t1985 23.317
R2304 VDD.n1351 VDD.t812 23.317
R2305 VDD.n421 VDD.t2005 23.317
R2306 VDD.n411 VDD.t2577 23.317
R2307 VDD.n400 VDD.t1399 23.317
R2308 VDD.n1255 VDD.t2155 23.316
R2309 VDD.n1399 VDD.t1972 23.316
R2310 VDD.n1113 VDD.t661 22.813
R2311 VDD.n1145 VDD.t82 22.813
R2312 VDD.n1176 VDD.t1080 22.813
R2313 VDD.n1208 VDD.t155 22.813
R2314 VDD.n766 VDD.t341 22.813
R2315 VDD.n740 VDD.t1753 22.813
R2316 VDD.n654 VDD.t2612 22.813
R2317 VDD.n1708 VDD.t315 22.813
R2318 VDD.n1647 VDD.t1884 20.998
R2319 VDD.n1613 VDD.t1902 20.998
R2320 VDD.n1588 VDD.t1892 20.998
R2321 VDD.n1563 VDD.t1824 20.998
R2322 VDD.n1538 VDD.t1852 20.998
R2323 VDD.n1513 VDD.t1869 20.998
R2324 VDD.n1497 VDD.t1828 20.998
R2325 VDD.n1463 VDD.t1855 20.998
R2326 VDD.n1255 VDD.t993 20.186
R2327 VDD.n1399 VDD.t2179 20.186
R2328 VDD.n1683 VDD.t2011 20.183
R2329 VDD.n1673 VDD.t2025 20.183
R2330 VDD.n1724 VDD.t2001 20.183
R2331 VDD.n1076 VDD.t2464 20.183
R2332 VDD.n813 VDD.t2138 20.183
R2333 VDD.n823 VDD.t2493 20.183
R2334 VDD.n438 VDD.t2095 20.183
R2335 VDD.n429 VDD.t1460 20.183
R2336 VDD.n787 VDD.t290 20.183
R2337 VDD.n796 VDD.t2363 20.183
R2338 VDD.n1367 VDD.t2081 20.183
R2339 VDD.n1359 VDD.t548 20.183
R2340 VDD.n1664 VDD.t2481 20.183
R2341 VDD.n1351 VDD.t2511 20.183
R2342 VDD.n421 VDD.t2513 20.183
R2343 VDD.n411 VDD.t1101 20.183
R2344 VDD.n400 VDD.t2453 20.183
R2345 VDD.n1693 VDD.n1682 15.439
R2346 VDD.n31 VDD.t360 14.284
R2347 VDD.n36 VDD.t695 14.284
R2348 VDD.n19 VDD.t669 14.284
R2349 VDD.n24 VDD.t2163 14.284
R2350 VDD.n1842 VDD.t1597 14.284
R2351 VDD.n1848 VDD.t239 14.284
R2352 VDD.n1820 VDD.t884 14.284
R2353 VDD.n1826 VDD.t2341 14.284
R2354 VDD.n1791 VDD.t2400 14.284
R2355 VDD.n1796 VDD.t1099 14.284
R2356 VDD.n1802 VDD.t2265 14.284
R2357 VDD.n1807 VDD.t1873 14.284
R2358 VDD.n60 VDD.t2327 14.284
R2359 VDD.n1638 VDD.t1279 14.284
R2360 VDD.n1633 VDD.t1843 14.284
R2361 VDD.n1620 VDD.t1875 14.284
R2362 VDD.n1606 VDD.t756 14.284
R2363 VDD.n1595 VDD.t1850 14.284
R2364 VDD.n1581 VDD.t2116 14.284
R2365 VDD.n1570 VDD.t1913 14.284
R2366 VDD.n1556 VDD.t1984 14.284
R2367 VDD.n1545 VDD.t1823 14.284
R2368 VDD.n1531 VDD.t1467 14.284
R2369 VDD.n1520 VDD.t1909 14.284
R2370 VDD.n1506 VDD.t243 14.284
R2371 VDD.n1488 VDD.t704 14.284
R2372 VDD.n1483 VDD.t1883 14.284
R2373 VDD.n1470 VDD.t1827 14.284
R2374 VDD.n1456 VDD.t1161 14.284
R2375 VDD.n1069 VDD.t986 14.284
R2376 VDD.n1124 VDD.t582 14.284
R2377 VDD.n1005 VDD.t2313 14.284
R2378 VDD.n1154 VDD.t33 14.284
R2379 VDD.n942 VDD.t257 14.284
R2380 VDD.n1184 VDD.t1122 14.284
R2381 VDD.n1213 VDD.t539 14.284
R2382 VDD.n1220 VDD.t850 14.284
R2383 VDD.n507 VDD.t895 14.284
R2384 VDD.n778 VDD.t95 14.284
R2385 VDD.n578 VDD.t264 14.284
R2386 VDD.n571 VDD.t1718 14.284
R2387 VDD.n660 VDD.t514 14.284
R2388 VDD.n1705 VDD.t752 14.284
R2389 VDD.n1698 VDD.t53 14.284
R2390 VDD.n586 VDD.t1310 14.284
R2391 VDD.n591 VDD.t144 14.284
R2392 VDD.n621 VDD.t1676 14.284
R2393 VDD.n626 VDD.t1451 14.284
R2394 VDD.n668 VDD.t2597 14.284
R2395 VDD.n710 VDD.t1254 14.284
R2396 VDD.n715 VDD.t419 14.284
R2397 VDD.n697 VDD.t723 14.284
R2398 VDD.n702 VDD.t2056 14.284
R2399 VDD.n557 VDD.t174 14.284
R2400 VDD.n562 VDD.t2541 14.284
R2401 VDD.n538 VDD.t2372 14.284
R2402 VDD.n543 VDD.t605 14.284
R2403 VDD.n1385 VDD.t2192 14.284
R2404 VDD.n1380 VDD.t1965 14.284
R2405 VDD.n1248 VDD.t505 14.284
R2406 VDD.n1243 VDD.t2154 14.284
R2407 VDD.n1234 VDD.t142 14.284
R2408 VDD.n1229 VDD.t2568 14.284
R2409 VDD.n393 VDD.t2456 14.284
R2410 VDD.n388 VDD.t1394 14.284
R2411 VDD.n174 VDD.t2413 14.284
R2412 VDD.n179 VDD.t86 14.284
R2413 VDD.n122 VDD.t1653 14.284
R2414 VDD.n117 VDD.t235 14.284
R2415 VDD.n236 VDD.t622 14.284
R2416 VDD.n231 VDD.t440 14.284
R2417 VDD.n65 VDD.t244 14.284
R2418 VDD.n80 VDD.t2466 14.284
R2419 VDD.n75 VDD.t1209 14.284
R2420 VDD.n108 VDD.t2587 14.284
R2421 VDD.n103 VDD.t647 14.284
R2422 VDD.n137 VDD.t2142 14.284
R2423 VDD.n132 VDD.t1369 14.284
R2424 VDD.n165 VDD.t2195 14.284
R2425 VDD.n160 VDD.t559 14.284
R2426 VDD.n194 VDD.t1620 14.284
R2427 VDD.n189 VDD.t1408 14.284
R2428 VDD.n222 VDD.t914 14.284
R2429 VDD.n217 VDD.t1923 14.284
R2430 VDD.n358 VDD.t1014 14.284
R2431 VDD.n363 VDD.t467 14.284
R2432 VDD.n346 VDD.t1796 14.284
R2433 VDD.n351 VDD.t2366 14.284
R2434 VDD.n319 VDD.t649 14.284
R2435 VDD.n325 VDD.t202 14.284
R2436 VDD.n303 VDD.t2346 14.284
R2437 VDD.n297 VDD.t375 14.284
R2438 VDD.n275 VDD.t1418 14.284
R2439 VDD.n280 VDD.t1921 14.284
R2440 VDD.n263 VDD.t572 14.284
R2441 VDD.n268 VDD.t718 14.284
R2442 VDD.n493 VDD.t79 14.284
R2443 VDD.n498 VDD.t1130 14.284
R2444 VDD.n475 VDD.t1775 14.284
R2445 VDD.n480 VDD.t998 14.284
R2446 VDD.n871 VDD.t392 14.284
R2447 VDD.n876 VDD.t2244 14.284
R2448 VDD.n852 VDD.t1332 14.284
R2449 VDD.n857 VDD.t1595 14.284
R2450 VDD.n883 VDD.t869 14.284
R2451 VDD.n888 VDD.t1740 14.284
R2452 VDD.n920 VDD.t2215 14.284
R2453 VDD.n925 VDD.t829 14.284
R2454 VDD.n949 VDD.t2329 14.284
R2455 VDD.n954 VDD.t2428 14.284
R2456 VDD.n983 VDD.t931 14.284
R2457 VDD.n988 VDD.t1112 14.284
R2458 VDD.n1012 VDD.t2295 14.284
R2459 VDD.n1017 VDD.t1069 14.284
R2460 VDD.n1047 VDD.t1690 14.284
R2461 VDD.n1052 VDD.t457 14.284
R2462 VDD.n1756 VDD.t1940 14.284
R2463 VDD.n1751 VDD.t962 14.284
R2464 VDD.n1745 VDD.t2595 14.284
R2465 VDD.n1740 VDD.t1427 14.284
R2466 VDD.n1290 VDD.t1557 14.283
R2467 VDD.n1308 VDD.t1483 14.283
R2468 VDD.n1325 VDD.t1491 14.283
R2469 VDD.n1342 VDD.t1513 14.283
R2470 VDD.n1411 VDD.t1477 14.283
R2471 VDD.n1428 VDD.t1559 14.283
R2472 VDD.n378 VDD.t1529 14.283
R2473 VDD.n1273 VDD.t1479 14.283
R2474 VDD.n1286 VDD.t1244 14.283
R2475 VDD.n1304 VDD.t5 14.283
R2476 VDD.n1321 VDD.t349 14.283
R2477 VDD.n1338 VDD.t2557 14.283
R2478 VDD.n1407 VDD.t1748 14.283
R2479 VDD.n1424 VDD.t557 14.283
R2480 VDD.n374 VDD.t901 14.283
R2481 VDD.n1269 VDD.t302 14.283
R2482 VDD.n30 VDD.t37 14.282
R2483 VDD.n30 VDD.t38 14.282
R2484 VDD.n35 VDD.t693 14.282
R2485 VDD.n35 VDD.t692 14.282
R2486 VDD.n18 VDD.t673 14.282
R2487 VDD.n18 VDD.t670 14.282
R2488 VDD.n23 VDD.t2161 14.282
R2489 VDD.n23 VDD.t2172 14.282
R2490 VDD.n1839 VDD.t1596 14.282
R2491 VDD.n1839 VDD.t1598 14.282
R2492 VDD.n1845 VDD.t238 14.282
R2493 VDD.n1845 VDD.t237 14.282
R2494 VDD.n1817 VDD.t190 14.282
R2495 VDD.n1817 VDD.t282 14.282
R2496 VDD.n1823 VDD.t2340 14.282
R2497 VDD.n1823 VDD.t2399 14.282
R2498 VDD.n1790 VDD.t2403 14.282
R2499 VDD.n1790 VDD.t2404 14.282
R2500 VDD.n1795 VDD.t1098 14.282
R2501 VDD.n1795 VDD.t1097 14.282
R2502 VDD.n1801 VDD.t2267 14.282
R2503 VDD.n1801 VDD.t2266 14.282
R2504 VDD.n1806 VDD.t1854 14.282
R2505 VDD.n1806 VDD.t1851 14.282
R2506 VDD.n57 VDD.t2326 14.282
R2507 VDD.n57 VDD.t2325 14.282
R2508 VDD.n1637 VDD.t1273 14.282
R2509 VDD.n1637 VDD.t1281 14.282
R2510 VDD.n1632 VDD.t1907 14.282
R2511 VDD.n1632 VDD.t1885 14.282
R2512 VDD.n1619 VDD.t1836 14.282
R2513 VDD.n1619 VDD.t1903 14.282
R2514 VDD.n1605 VDD.t293 14.282
R2515 VDD.n1605 VDD.t425 14.282
R2516 VDD.n1594 VDD.t1911 14.282
R2517 VDD.n1594 VDD.t1893 14.282
R2518 VDD.n1580 VDD.t2100 14.282
R2519 VDD.n1580 VDD.t2090 14.282
R2520 VDD.n1569 VDD.t1866 14.282
R2521 VDD.n1569 VDD.t1825 14.282
R2522 VDD.n1555 VDD.t2004 14.282
R2523 VDD.n1555 VDD.t1990 14.282
R2524 VDD.n1544 VDD.t1889 14.282
R2525 VDD.n1544 VDD.t1853 14.282
R2526 VDD.n1530 VDD.t817 14.282
R2527 VDD.n1530 VDD.t807 14.282
R2528 VDD.n1519 VDD.t1891 14.282
R2529 VDD.n1519 VDD.t1870 14.282
R2530 VDD.n1505 VDD.t512 14.282
R2531 VDD.n1505 VDD.t459 14.282
R2532 VDD.n1490 VDD.t712 14.282
R2533 VDD.n1490 VDD.t708 14.282
R2534 VDD.n1485 VDD.t1848 14.282
R2535 VDD.n1485 VDD.t1829 14.282
R2536 VDD.n1469 VDD.t1895 14.282
R2537 VDD.n1469 VDD.t1856 14.282
R2538 VDD.n1455 VDD.t1159 14.282
R2539 VDD.n1455 VDD.t1157 14.282
R2540 VDD.n1066 VDD.t990 14.282
R2541 VDD.n1066 VDD.t103 14.282
R2542 VDD.n1121 VDD.t584 14.282
R2543 VDD.n1121 VDD.t586 14.282
R2544 VDD.n1002 VDD.t2315 14.282
R2545 VDD.n1002 VDD.t2317 14.282
R2546 VDD.n1151 VDD.t29 14.282
R2547 VDD.n1151 VDD.t31 14.282
R2548 VDD.n939 VDD.t259 14.282
R2549 VDD.n939 VDD.t255 14.282
R2550 VDD.n1181 VDD.t1118 14.282
R2551 VDD.n1181 VDD.t1120 14.282
R2552 VDD.n1214 VDD.t408 14.282
R2553 VDD.n1214 VDD.t251 14.282
R2554 VDD.n1221 VDD.t286 14.282
R2555 VDD.n1221 VDD.t1009 14.282
R2556 VDD.n504 VDD.t893 14.282
R2557 VDD.n504 VDD.t65 14.282
R2558 VDD.n775 VDD.t171 14.282
R2559 VDD.n775 VDD.t169 14.282
R2560 VDD.n575 VDD.t43 14.282
R2561 VDD.n575 VDD.t192 14.282
R2562 VDD.n568 VDD.t1716 14.282
R2563 VDD.n568 VDD.t1714 14.282
R2564 VDD.n661 VDD.t40 14.282
R2565 VDD.n661 VDD.t1000 14.282
R2566 VDD.n1706 VDD.t750 14.282
R2567 VDD.n1706 VDD.t748 14.282
R2568 VDD.n1699 VDD.t1007 14.282
R2569 VDD.n1699 VDD.t518 14.282
R2570 VDD.n585 VDD.t1308 14.282
R2571 VDD.n585 VDD.t1306 14.282
R2572 VDD.n590 VDD.t981 14.282
R2573 VDD.n590 VDD.t516 14.282
R2574 VDD.n620 VDD.t1680 14.282
R2575 VDD.n620 VDD.t1678 14.282
R2576 VDD.n625 VDD.t1449 14.282
R2577 VDD.n625 VDD.t1439 14.282
R2578 VDD.n669 VDD.t2604 14.282
R2579 VDD.n669 VDD.t2609 14.282
R2580 VDD.n709 VDD.t1246 14.282
R2581 VDD.n709 VDD.t99 14.282
R2582 VDD.n714 VDD.t195 14.282
R2583 VDD.n714 VDD.t421 14.282
R2584 VDD.n696 VDD.t735 14.282
R2585 VDD.n696 VDD.t733 14.282
R2586 VDD.n701 VDD.t2054 14.282
R2587 VDD.n701 VDD.t2062 14.282
R2588 VDD.n556 VDD.t178 14.282
R2589 VDD.n556 VDD.t176 14.282
R2590 VDD.n561 VDD.t2539 14.282
R2591 VDD.n561 VDD.t2531 14.282
R2592 VDD.n537 VDD.t2376 14.282
R2593 VDD.n537 VDD.t2374 14.282
R2594 VDD.n542 VDD.t272 14.282
R2595 VDD.n542 VDD.t406 14.282
R2596 VDD.n1384 VDD.t2178 14.282
R2597 VDD.n1384 VDD.t2176 14.282
R2598 VDD.n1379 VDD.t1963 14.282
R2599 VDD.n1379 VDD.t1957 14.282
R2600 VDD.n1289 VDD.t1537 14.282
R2601 VDD.n1289 VDD.t1495 14.282
R2602 VDD.n1285 VDD.t1242 14.282
R2603 VDD.n1285 VDD.t1240 14.282
R2604 VDD.n1307 VDD.t1549 14.282
R2605 VDD.n1307 VDD.t1531 14.282
R2606 VDD.n1303 VDD.t3 14.282
R2607 VDD.n1303 VDD.t13 14.282
R2608 VDD.n1324 VDD.t1545 14.282
R2609 VDD.n1324 VDD.t1535 14.282
R2610 VDD.n1320 VDD.t270 14.282
R2611 VDD.n1320 VDD.t312 14.282
R2612 VDD.n1341 VDD.t1489 14.282
R2613 VDD.n1341 VDD.t1551 14.282
R2614 VDD.n1337 VDD.t2555 14.282
R2615 VDD.n1337 VDD.t2559 14.282
R2616 VDD.n1247 VDD.t404 14.282
R2617 VDD.n1247 VDD.t716 14.282
R2618 VDD.n1242 VDD.t2148 14.282
R2619 VDD.n1242 VDD.t2152 14.282
R2620 VDD.n1233 VDD.t1213 14.282
R2621 VDD.n1233 VDD.t1175 14.282
R2622 VDD.n1228 VDD.t2574 14.282
R2623 VDD.n1228 VDD.t2570 14.282
R2624 VDD.n392 VDD.t2460 14.282
R2625 VDD.n392 VDD.t2458 14.282
R2626 VDD.n387 VDD.t1386 14.282
R2627 VDD.n387 VDD.t1384 14.282
R2628 VDD.n1410 VDD.t1539 14.282
R2629 VDD.n1410 VDD.t1523 14.282
R2630 VDD.n1406 VDD.t1746 14.282
R2631 VDD.n1406 VDD.t1744 14.282
R2632 VDD.n1427 VDD.t1507 14.282
R2633 VDD.n1427 VDD.t1563 14.282
R2634 VDD.n1423 VDD.t555 14.282
R2635 VDD.n1423 VDD.t553 14.282
R2636 VDD.n377 VDD.t1511 14.282
R2637 VDD.n377 VDD.t1567 14.282
R2638 VDD.n373 VDD.t36 14.282
R2639 VDD.n373 VDD.t903 14.282
R2640 VDD.n171 VDD.t2411 14.282
R2641 VDD.n171 VDD.t2412 14.282
R2642 VDD.n176 VDD.t953 14.282
R2643 VDD.n176 VDD.t87 14.282
R2644 VDD.n119 VDD.t1681 14.282
R2645 VDD.n119 VDD.t1682 14.282
R2646 VDD.n114 VDD.t613 14.282
R2647 VDD.n114 VDD.t614 14.282
R2648 VDD.n233 VDD.t306 14.282
R2649 VDD.n233 VDD.t305 14.282
R2650 VDD.n228 VDD.t442 14.282
R2651 VDD.n228 VDD.t441 14.282
R2652 VDD.n62 VDD.t24 14.282
R2653 VDD.n62 VDD.t214 14.282
R2654 VDD.n79 VDD.t2474 14.282
R2655 VDD.n79 VDD.t2463 14.282
R2656 VDD.n74 VDD.t151 14.282
R2657 VDD.n74 VDD.t150 14.282
R2658 VDD.n107 VDD.t2589 14.282
R2659 VDD.n107 VDD.t2588 14.282
R2660 VDD.n102 VDD.t646 14.282
R2661 VDD.n102 VDD.t645 14.282
R2662 VDD.n136 VDD.t2129 14.282
R2663 VDD.n136 VDD.t2128 14.282
R2664 VDD.n131 VDD.t1370 14.282
R2665 VDD.n131 VDD.t1368 14.282
R2666 VDD.n164 VDD.t2080 14.282
R2667 VDD.n164 VDD.t2203 14.282
R2668 VDD.n159 VDD.t563 14.282
R2669 VDD.n159 VDD.t558 14.282
R2670 VDD.n193 VDD.t1624 14.282
R2671 VDD.n193 VDD.t1622 14.282
R2672 VDD.n188 VDD.t1406 14.282
R2673 VDD.n188 VDD.t1405 14.282
R2674 VDD.n221 VDD.t921 14.282
R2675 VDD.n221 VDD.t919 14.282
R2676 VDD.n216 VDD.t1928 14.282
R2677 VDD.n216 VDD.t1927 14.282
R2678 VDD.n357 VDD.t1016 14.282
R2679 VDD.n357 VDD.t1015 14.282
R2680 VDD.n362 VDD.t466 14.282
R2681 VDD.n362 VDD.t465 14.282
R2682 VDD.n345 VDD.t1798 14.282
R2683 VDD.n345 VDD.t1797 14.282
R2684 VDD.n350 VDD.t2504 14.282
R2685 VDD.n350 VDD.t2503 14.282
R2686 VDD.n316 VDD.t241 14.282
R2687 VDD.n316 VDD.t240 14.282
R2688 VDD.n322 VDD.t1 14.282
R2689 VDD.n322 VDD.t0 14.282
R2690 VDD.n300 VDD.t2345 14.282
R2691 VDD.n300 VDD.t2414 14.282
R2692 VDD.n294 VDD.t41 14.282
R2693 VDD.n294 VDD.t157 14.282
R2694 VDD.n274 VDD.t1413 14.282
R2695 VDD.n274 VDD.t1414 14.282
R2696 VDD.n279 VDD.t1920 14.282
R2697 VDD.n279 VDD.t1919 14.282
R2698 VDD.n262 VDD.t577 14.282
R2699 VDD.n262 VDD.t576 14.282
R2700 VDD.n267 VDD.t75 14.282
R2701 VDD.n267 VDD.t615 14.282
R2702 VDD.n1272 VDD.t1533 14.282
R2703 VDD.n1272 VDD.t1525 14.282
R2704 VDD.n1268 VDD.t498 14.282
R2705 VDD.n1268 VDD.t523 14.282
R2706 VDD.n492 VDD.t266 14.282
R2707 VDD.n492 VDD.t952 14.282
R2708 VDD.n497 VDD.t1128 14.282
R2709 VDD.n497 VDD.t1236 14.282
R2710 VDD.n474 VDD.t1761 14.282
R2711 VDD.n474 VDD.t1777 14.282
R2712 VDD.n479 VDD.t500 14.282
R2713 VDD.n479 VDD.t526 14.282
R2714 VDD.n870 VDD.t67 14.282
R2715 VDD.n870 VDD.t566 14.282
R2716 VDD.n875 VDD.t2250 14.282
R2717 VDD.n875 VDD.t2238 14.282
R2718 VDD.n851 VDD.t1318 14.282
R2719 VDD.n851 VDD.t1328 14.282
R2720 VDD.n856 VDD.t1577 14.282
R2721 VDD.n856 VDD.t1589 14.282
R2722 VDD.n882 VDD.t873 14.282
R2723 VDD.n882 VDD.t877 14.282
R2724 VDD.n887 VDD.t1724 14.282
R2725 VDD.n887 VDD.t1736 14.282
R2726 VDD.n919 VDD.t2225 14.282
R2727 VDD.n919 VDD.t2209 14.282
R2728 VDD.n924 VDD.t835 14.282
R2729 VDD.n924 VDD.t825 14.282
R2730 VDD.n948 VDD.t2333 14.282
R2731 VDD.n948 VDD.t2337 14.282
R2732 VDD.n953 VDD.t2426 14.282
R2733 VDD.n953 VDD.t2416 14.282
R2734 VDD.n982 VDD.t935 14.282
R2735 VDD.n982 VDD.t682 14.282
R2736 VDD.n987 VDD.t1046 14.282
R2737 VDD.n987 VDD.t1044 14.282
R2738 VDD.n1011 VDD.t2303 14.282
R2739 VDD.n1011 VDD.t2297 14.282
R2740 VDD.n1016 VDD.t1079 14.282
R2741 VDD.n1016 VDD.t1073 14.282
R2742 VDD.n1046 VDD.t1700 14.282
R2743 VDD.n1046 VDD.t1708 14.282
R2744 VDD.n1051 VDD.t1355 14.282
R2745 VDD.n1051 VDD.t1341 14.282
R2746 VDD.n1755 VDD.t1939 14.282
R2747 VDD.n1755 VDD.t1938 14.282
R2748 VDD.n1750 VDD.t643 14.282
R2749 VDD.n1750 VDD.t719 14.282
R2750 VDD.n1744 VDD.t2594 14.282
R2751 VDD.n1744 VDD.t2591 14.282
R2752 VDD.n1739 VDD.t1425 14.282
R2753 VDD.n1739 VDD.t1426 14.282
R2754 VDD.n1296 VDD.t1536 12.385
R2755 VDD.n1314 VDD.t1548 12.385
R2756 VDD.n1331 VDD.t1544 12.385
R2757 VDD.n1348 VDD.t1488 12.385
R2758 VDD.n1417 VDD.t1538 12.385
R2759 VDD.n1434 VDD.t1506 12.385
R2760 VDD.n384 VDD.t1510 12.385
R2761 VDD.n1279 VDD.t1532 12.385
R2762 VDD.n1693 VDD.n1692 10.379
R2763 VDD.n1734 VDD.n1733 9.353
R2764 VDD.n1253 VDD.t283 8.293
R2765 VDD.n1239 VDD.t230 8.293
R2766 VDD.n398 VDD.t948 8.293
R2767 VDD.n1390 VDD.t172 8.293
R2768 VDD.n1297 VDD.n1295 6.376
R2769 VDD.n1315 VDD.n1313 6.376
R2770 VDD.n1332 VDD.n1330 6.376
R2771 VDD.n1349 VDD.n1347 6.376
R2772 VDD.n1418 VDD.n1416 6.376
R2773 VDD.n1435 VDD.n1433 6.376
R2774 VDD.n385 VDD.n383 6.376
R2775 VDD.n1280 VDD.n1278 6.376
R2776 VDD.n1645 VDD.t784 6.189
R2777 VDD.n1646 VDD.t783 6.189
R2778 VDD.n1649 VDD.t1950 6.189
R2779 VDD.n1648 VDD.t1931 6.189
R2780 VDD.n1611 VDD.t1197 6.189
R2781 VDD.n1612 VDD.t1196 6.189
R2782 VDD.n1615 VDD.t1004 6.189
R2783 VDD.n1614 VDD.t203 6.189
R2784 VDD.n1586 VDD.t946 6.189
R2785 VDD.n1587 VDD.t1313 6.189
R2786 VDD.n1590 VDD.t1366 6.189
R2787 VDD.n1589 VDD.t1367 6.189
R2788 VDD.n1561 VDD.t1603 6.189
R2789 VDD.n1562 VDD.t1602 6.189
R2790 VDD.n1565 VDD.t310 6.189
R2791 VDD.n1564 VDD.t309 6.189
R2792 VDD.n1536 VDD.t1750 6.189
R2793 VDD.n1537 VDD.t1787 6.189
R2794 VDD.n1540 VDD.t623 6.189
R2795 VDD.n1539 VDD.t1135 6.189
R2796 VDD.n1511 VDD.t821 6.189
R2797 VDD.n1512 VDD.t820 6.189
R2798 VDD.n1515 VDD.t923 6.189
R2799 VDD.n1514 VDD.t908 6.189
R2800 VDD.n1495 VDD.t1090 6.189
R2801 VDD.n1496 VDD.t1295 6.189
R2802 VDD.n1499 VDD.t769 6.189
R2803 VDD.n1498 VDD.t768 6.189
R2804 VDD.n1461 VDD.t2077 6.189
R2805 VDD.n1462 VDD.t2079 6.189
R2806 VDD.n1465 VDD.t942 6.189
R2807 VDD.n1464 VDD.t944 6.189
R2808 VDD.n1281 VDD.n1280 4.897
R2809 VDD.n1297 VDD.n1296 4.688
R2810 VDD.n1315 VDD.n1314 4.688
R2811 VDD.n1332 VDD.n1331 4.688
R2812 VDD.n1349 VDD.n1348 4.688
R2813 VDD.n1418 VDD.n1417 4.688
R2814 VDD.n1435 VDD.n1434 4.688
R2815 VDD.n385 VDD.n384 4.688
R2816 VDD.n1280 VDD.n1279 4.688
R2817 VDD.n632 VDD.t307 4.524
R2818 VDD.n633 VDD.t327 4.524
R2819 VDD.n635 VDD.t766 4.524
R2820 VDD.n634 VDD.t764 4.524
R2821 VDD.n720 VDD.t120 4.524
R2822 VDD.n721 VDD.t119 4.524
R2823 VDD.n723 VDD.t2353 4.524
R2824 VDD.n722 VDD.t2352 4.524
R2825 VDD.n549 VDD.t1381 4.524
R2826 VDD.n550 VDD.t1382 4.524
R2827 VDD.n552 VDD.t207 4.524
R2828 VDD.n551 VDD.t510 4.524
R2829 VDD.n486 VDD.t1131 4.524
R2830 VDD.n487 VDD.t1186 4.524
R2831 VDD.n489 VDD.t547 4.524
R2832 VDD.n488 VDD.t1001 4.524
R2833 VDD.n863 VDD.t1137 4.524
R2834 VDD.n864 VDD.t1138 4.524
R2835 VDD.n866 VDD.t204 4.524
R2836 VDD.n865 VDD.t107 4.524
R2837 VDD.n931 VDD.t746 4.524
R2838 VDD.n932 VDD.t744 4.524
R2839 VDD.n934 VDD.t848 4.524
R2840 VDD.n933 VDD.t11 4.524
R2841 VDD.n994 VDD.t1600 4.524
R2842 VDD.n995 VDD.t1599 4.524
R2843 VDD.n997 VDD.t880 4.524
R2844 VDD.n996 VDD.t881 4.524
R2845 VDD.n1058 VDD.t521 4.524
R2846 VDD.n1059 VDD.t112 4.524
R2847 VDD.n1061 VDD.t2286 4.524
R2848 VDD.n1060 VDD.t2287 4.524
R2849 VDD.n1389 VDD.n1388 4.331
R2850 VDD.n1252 VDD.n1251 4.331
R2851 VDD.n397 VDD.n396 4.331
R2852 VDD.n40 VDD.n34 4.276
R2853 VDD.n28 VDD.n22 4.276
R2854 VDD.n1800 VDD.n1794 4.276
R2855 VDD.n1811 VDD.n1805 4.276
R2856 VDD.n595 VDD.n589 4.276
R2857 VDD.n630 VDD.n624 4.276
R2858 VDD.n719 VDD.n713 4.276
R2859 VDD.n706 VDD.n700 4.276
R2860 VDD.n566 VDD.n560 4.276
R2861 VDD.n547 VDD.n541 4.276
R2862 VDD.n367 VDD.n361 4.276
R2863 VDD.n355 VDD.n349 4.276
R2864 VDD.n284 VDD.n278 4.276
R2865 VDD.n272 VDD.n266 4.276
R2866 VDD.n502 VDD.n496 4.276
R2867 VDD.n484 VDD.n478 4.276
R2868 VDD.n880 VDD.n874 4.276
R2869 VDD.n861 VDD.n855 4.276
R2870 VDD.n892 VDD.n886 4.276
R2871 VDD.n929 VDD.n923 4.276
R2872 VDD.n958 VDD.n952 4.276
R2873 VDD.n992 VDD.n986 4.276
R2874 VDD.n1021 VDD.n1015 4.276
R2875 VDD.n1056 VDD.n1050 4.276
R2876 VDD.n1093 VDD.t1625 2.932
R2877 VDD.n1294 VDD.n1288 2.572
R2878 VDD.n1312 VDD.n1306 2.572
R2879 VDD.n1329 VDD.n1323 2.572
R2880 VDD.n1346 VDD.n1340 2.572
R2881 VDD.n1415 VDD.n1409 2.572
R2882 VDD.n1432 VDD.n1426 2.572
R2883 VDD.n382 VDD.n376 2.572
R2884 VDD.n1277 VDD.n1271 2.572
R2885 VDD.n1583 VDD.n1582 2.546
R2886 VDD.n1558 VDD.n1557 2.546
R2887 VDD.n1293 VDD.n1292 2.542
R2888 VDD.n1311 VDD.n1310 2.542
R2889 VDD.n1328 VDD.n1327 2.542
R2890 VDD.n1345 VDD.n1344 2.542
R2891 VDD.n1414 VDD.n1413 2.542
R2892 VDD.n1431 VDD.n1430 2.542
R2893 VDD.n381 VDD.n380 2.542
R2894 VDD.n1276 VDD.n1275 2.542
R2895 VDD.n1484 VDD.n1482 2.531
R2896 VDD.n33 VDD.n32 2.451
R2897 VDD.n21 VDD.n20 2.451
R2898 VDD.n1793 VDD.n1792 2.451
R2899 VDD.n1804 VDD.n1803 2.451
R2900 VDD.n1635 VDD.n1634 2.451
R2901 VDD.n1622 VDD.n1621 2.451
R2902 VDD.n1597 VDD.n1596 2.451
R2903 VDD.n1572 VDD.n1571 2.451
R2904 VDD.n1547 VDD.n1546 2.451
R2905 VDD.n1522 VDD.n1521 2.451
R2906 VDD.n1472 VDD.n1471 2.451
R2907 VDD.n588 VDD.n587 2.451
R2908 VDD.n623 VDD.n622 2.451
R2909 VDD.n712 VDD.n711 2.451
R2910 VDD.n699 VDD.n698 2.451
R2911 VDD.n559 VDD.n558 2.451
R2912 VDD.n540 VDD.n539 2.451
R2913 VDD.n1387 VDD.n1386 2.451
R2914 VDD.n1250 VDD.n1249 2.451
R2915 VDD.n1236 VDD.n1235 2.451
R2916 VDD.n395 VDD.n394 2.451
R2917 VDD.n77 VDD.n76 2.451
R2918 VDD.n105 VDD.n104 2.451
R2919 VDD.n134 VDD.n133 2.451
R2920 VDD.n162 VDD.n161 2.451
R2921 VDD.n191 VDD.n190 2.451
R2922 VDD.n219 VDD.n218 2.451
R2923 VDD.n360 VDD.n359 2.451
R2924 VDD.n348 VDD.n347 2.451
R2925 VDD.n277 VDD.n276 2.451
R2926 VDD.n265 VDD.n264 2.451
R2927 VDD.n495 VDD.n494 2.451
R2928 VDD.n477 VDD.n476 2.451
R2929 VDD.n873 VDD.n872 2.451
R2930 VDD.n854 VDD.n853 2.451
R2931 VDD.n885 VDD.n884 2.451
R2932 VDD.n922 VDD.n921 2.451
R2933 VDD.n951 VDD.n950 2.451
R2934 VDD.n985 VDD.n984 2.451
R2935 VDD.n1014 VDD.n1013 2.451
R2936 VDD.n1049 VDD.n1048 2.451
R2937 VDD.n1758 VDD.n1757 2.451
R2938 VDD.n1747 VDD.n1746 2.451
R2939 VDD.n38 VDD.n37 2.449
R2940 VDD.n26 VDD.n25 2.449
R2941 VDD.n1798 VDD.n1797 2.449
R2942 VDD.n1809 VDD.n1808 2.449
R2943 VDD.n1640 VDD.n1639 2.449
R2944 VDD.n1608 VDD.n1607 2.449
R2945 VDD.n1533 VDD.n1532 2.449
R2946 VDD.n1508 VDD.n1507 2.449
R2947 VDD.n1458 VDD.n1457 2.449
R2948 VDD.n593 VDD.n592 2.449
R2949 VDD.n628 VDD.n627 2.449
R2950 VDD.n717 VDD.n716 2.449
R2951 VDD.n704 VDD.n703 2.449
R2952 VDD.n564 VDD.n563 2.449
R2953 VDD.n545 VDD.n544 2.449
R2954 VDD.n1382 VDD.n1381 2.449
R2955 VDD.n1245 VDD.n1244 2.449
R2956 VDD.n1231 VDD.n1230 2.449
R2957 VDD.n390 VDD.n389 2.449
R2958 VDD.n82 VDD.n81 2.449
R2959 VDD.n110 VDD.n109 2.449
R2960 VDD.n139 VDD.n138 2.449
R2961 VDD.n167 VDD.n166 2.449
R2962 VDD.n196 VDD.n195 2.449
R2963 VDD.n224 VDD.n223 2.449
R2964 VDD.n365 VDD.n364 2.449
R2965 VDD.n353 VDD.n352 2.449
R2966 VDD.n282 VDD.n281 2.449
R2967 VDD.n270 VDD.n269 2.449
R2968 VDD.n500 VDD.n499 2.449
R2969 VDD.n482 VDD.n481 2.449
R2970 VDD.n878 VDD.n877 2.449
R2971 VDD.n859 VDD.n858 2.449
R2972 VDD.n890 VDD.n889 2.449
R2973 VDD.n927 VDD.n926 2.449
R2974 VDD.n956 VDD.n955 2.449
R2975 VDD.n990 VDD.n989 2.449
R2976 VDD.n1019 VDD.n1018 2.449
R2977 VDD.n1054 VDD.n1053 2.449
R2978 VDD.n1753 VDD.n1752 2.449
R2979 VDD.n1742 VDD.n1741 2.449
R2980 VDD.n1489 VDD.n1487 2.399
R2981 VDD.n1842 VDD.n1841 2.195
R2982 VDD.n1848 VDD.n1847 2.195
R2983 VDD.n1820 VDD.n1819 2.195
R2984 VDD.n1826 VDD.n1825 2.195
R2985 VDD.n60 VDD.n59 2.195
R2986 VDD.n1069 VDD.n1068 2.195
R2987 VDD.n1124 VDD.n1123 2.195
R2988 VDD.n1005 VDD.n1004 2.195
R2989 VDD.n1154 VDD.n1153 2.195
R2990 VDD.n942 VDD.n941 2.195
R2991 VDD.n1184 VDD.n1183 2.195
R2992 VDD.n1213 VDD.n1212 2.195
R2993 VDD.n1220 VDD.n1219 2.195
R2994 VDD.n507 VDD.n506 2.195
R2995 VDD.n778 VDD.n777 2.195
R2996 VDD.n578 VDD.n577 2.195
R2997 VDD.n571 VDD.n570 2.195
R2998 VDD.n660 VDD.n659 2.195
R2999 VDD.n1705 VDD.n1704 2.195
R3000 VDD.n1698 VDD.n1697 2.195
R3001 VDD.n668 VDD.n667 2.195
R3002 VDD.n174 VDD.n173 2.195
R3003 VDD.n179 VDD.n178 2.195
R3004 VDD.n122 VDD.n121 2.195
R3005 VDD.n117 VDD.n116 2.195
R3006 VDD.n236 VDD.n235 2.195
R3007 VDD.n231 VDD.n230 2.195
R3008 VDD.n65 VDD.n64 2.195
R3009 VDD.n319 VDD.n318 2.195
R3010 VDD.n325 VDD.n324 2.195
R3011 VDD.n303 VDD.n302 2.195
R3012 VDD.n297 VDD.n296 2.195
R3013 VDD.n1222 VDD.n1221 1.833
R3014 VDD.n1700 VDD.n1699 1.833
R3015 VDD.n670 VDD.n669 1.833
R3016 VDD.n1215 VDD.n1214 1.811
R3017 VDD.n662 VDD.n661 1.811
R3018 VDD.n1707 VDD.n1706 1.811
R3019 VDD.n1849 VDD.n1845 1.72
R3020 VDD.n1827 VDD.n1823 1.72
R3021 VDD.n61 VDD.n57 1.72
R3022 VDD.n1125 VDD.n1121 1.72
R3023 VDD.n1155 VDD.n1151 1.72
R3024 VDD.n1185 VDD.n1181 1.72
R3025 VDD.n779 VDD.n775 1.72
R3026 VDD.n572 VDD.n568 1.72
R3027 VDD.n175 VDD.n171 1.72
R3028 VDD.n118 VDD.n114 1.72
R3029 VDD.n232 VDD.n228 1.72
R3030 VDD.n326 VDD.n322 1.72
R3031 VDD.n304 VDD.n300 1.72
R3032 VDD.n1843 VDD.n1839 1.698
R3033 VDD.n1821 VDD.n1817 1.698
R3034 VDD.n1070 VDD.n1066 1.698
R3035 VDD.n1006 VDD.n1002 1.698
R3036 VDD.n943 VDD.n939 1.698
R3037 VDD.n508 VDD.n504 1.698
R3038 VDD.n579 VDD.n575 1.698
R3039 VDD.n180 VDD.n176 1.698
R3040 VDD.n123 VDD.n119 1.698
R3041 VDD.n237 VDD.n233 1.698
R3042 VDD.n66 VDD.n62 1.698
R3043 VDD.n320 VDD.n316 1.698
R3044 VDD.n298 VDD.n294 1.698
R3045 VDD.n1841 VDD.n1840 1.651
R3046 VDD.n1847 VDD.n1846 1.651
R3047 VDD.n1819 VDD.n1818 1.651
R3048 VDD.n1825 VDD.n1824 1.651
R3049 VDD.n59 VDD.n58 1.651
R3050 VDD.n1068 VDD.n1067 1.651
R3051 VDD.n1123 VDD.n1122 1.651
R3052 VDD.n1004 VDD.n1003 1.651
R3053 VDD.n1153 VDD.n1152 1.651
R3054 VDD.n941 VDD.n940 1.651
R3055 VDD.n1183 VDD.n1182 1.651
R3056 VDD.n1212 VDD.n1211 1.651
R3057 VDD.n1219 VDD.n1218 1.651
R3058 VDD.n506 VDD.n505 1.651
R3059 VDD.n777 VDD.n776 1.651
R3060 VDD.n577 VDD.n576 1.651
R3061 VDD.n570 VDD.n569 1.651
R3062 VDD.n659 VDD.n658 1.651
R3063 VDD.n1704 VDD.n1703 1.651
R3064 VDD.n1697 VDD.n1696 1.651
R3065 VDD.n667 VDD.n666 1.651
R3066 VDD.n173 VDD.n172 1.651
R3067 VDD.n178 VDD.n177 1.651
R3068 VDD.n121 VDD.n120 1.651
R3069 VDD.n116 VDD.n115 1.651
R3070 VDD.n235 VDD.n234 1.651
R3071 VDD.n230 VDD.n229 1.651
R3072 VDD.n64 VDD.n63 1.651
R3073 VDD.n318 VDD.n317 1.651
R3074 VDD.n324 VDD.n323 1.651
R3075 VDD.n302 VDD.n301 1.651
R3076 VDD.n296 VDD.n295 1.651
R3077 VDD.n1714 VDD.n1713 1.647
R3078 VDD.n1728 VDD.n1727 1.647
R3079 VDD.n1200 VDD.n1199 1.647
R3080 VDD.n808 VDD.n807 1.647
R3081 VDD.n818 VDD.n817 1.647
R3082 VDD.n646 VDD.n645 1.647
R3083 VDD.n415 VDD.n414 1.647
R3084 VDD.n404 VDD.n403 1.647
R3085 VDD.n834 VDD.n833 1.647
R3086 VDD.n895 VDD.n894 1.647
R3087 VDD.n964 VDD.n963 1.647
R3088 VDD.n1024 VDD.n1023 1.647
R3089 VDD.n15 VDD.n13 1.564
R3090 VDD.n7 VDD.n5 1.564
R3091 VDD.n1836 VDD.n1834 1.564
R3092 VDD.n44 VDD.n42 1.564
R3093 VDD.n1788 VDD.n1786 1.564
R3094 VDD.n55 VDD.n53 1.564
R3095 VDD.n1686 VDD.n1684 1.564
R3096 VDD.n1676 VDD.n1674 1.564
R3097 VDD.n1079 VDD.n1077 1.564
R3098 VDD.n1075 VDD.n1073 1.564
R3099 VDD.n1010 VDD.n1008 1.564
R3100 VDD.n947 VDD.n945 1.564
R3101 VDD.n1087 VDD.n1085 1.564
R3102 VDD.n441 VDD.n439 1.564
R3103 VDD.n432 VDD.n430 1.564
R3104 VDD.n790 VDD.n788 1.564
R3105 VDD.n799 VDD.n797 1.564
R3106 VDD.n513 VDD.n511 1.564
R3107 VDD.n584 VDD.n582 1.564
R3108 VDD.n598 VDD.n596 1.564
R3109 VDD.n602 VDD.n600 1.564
R3110 VDD.n674 VDD.n672 1.564
R3111 VDD.n684 VDD.n682 1.564
R3112 VDD.n516 VDD.n514 1.564
R3113 VDD.n525 VDD.n523 1.564
R3114 VDD.n1370 VDD.n1368 1.564
R3115 VDD.n1362 VDD.n1360 1.564
R3116 VDD.n1667 VDD.n1665 1.564
R3117 VDD.n1354 VDD.n1352 1.564
R3118 VDD.n1396 VDD.n1394 1.564
R3119 VDD.n1258 VDD.n1256 1.564
R3120 VDD.n424 VDD.n422 1.564
R3121 VDD.n73 VDD.n71 1.564
R3122 VDD.n130 VDD.n128 1.564
R3123 VDD.n187 VDD.n185 1.564
R3124 VDD.n244 VDD.n242 1.564
R3125 VDD.n91 VDD.n89 1.564
R3126 VDD.n94 VDD.n92 1.564
R3127 VDD.n148 VDD.n146 1.564
R3128 VDD.n151 VDD.n149 1.564
R3129 VDD.n205 VDD.n203 1.564
R3130 VDD.n208 VDD.n206 1.564
R3131 VDD.n342 VDD.n340 1.564
R3132 VDD.n334 VDD.n332 1.564
R3133 VDD.n313 VDD.n311 1.564
R3134 VDD.n292 VDD.n290 1.564
R3135 VDD.n259 VDD.n257 1.564
R3136 VDD.n251 VDD.n249 1.564
R3137 VDD.n466 VDD.n464 1.564
R3138 VDD.n455 VDD.n453 1.564
R3139 VDD.n831 VDD.n829 1.564
R3140 VDD.n912 VDD.n910 1.564
R3141 VDD.n961 VDD.n959 1.564
R3142 VDD.n1035 VDD.n1033 1.564
R3143 VDD.n1767 VDD.n1765 1.564
R3144 VDD.n1770 VDD.n1768 1.564
R3145 VDD.n827 VDD.n826 1.496
R3146 VDD.n826 VDD.n825 1.232
R3147 VDD.n1097 VDD.n1096 1.223
R3148 VDD.n1377 VDD.n1376 1.212
R3149 VDD.n1491 VDD.n1490 1.195
R3150 VDD.n1486 VDD.n1485 1.195
R3151 VDD.n1484 VDD.n1483 1.194
R3152 VDD.n1636 VDD.n1632 1.114
R3153 VDD.n1295 VDD.t1132 1.057
R3154 VDD.n1313 VDD.t1086 1.057
R3155 VDD.n1330 VDD.t882 1.057
R3156 VDD.n1347 VDD.t1168 1.057
R3157 VDD.n1416 VDD.t1224 1.057
R3158 VDD.n1433 VDD.t591 1.057
R3159 VDD.n383 VDD.t620 1.057
R3160 VDD.n1278 VDD.t412 1.057
R3161 VDD.n1376 VDD.n1375 1.025
R3162 VDD.n1489 VDD.n1488 1.002
R3163 VDD.n1718 VDD.n1717 0.983
R3164 VDD.n1729 VDD.n1728 0.983
R3165 VDD.n1204 VDD.n1203 0.983
R3166 VDD.n809 VDD.n808 0.983
R3167 VDD.n819 VDD.n818 0.983
R3168 VDD.n650 VDD.n649 0.983
R3169 VDD.n416 VDD.n415 0.983
R3170 VDD.n405 VDD.n404 0.983
R3171 VDD.n838 VDD.n837 0.983
R3172 VDD.n899 VDD.n898 0.983
R3173 VDD.n968 VDD.n967 0.983
R3174 VDD.n1028 VDD.n1027 0.983
R3175 VDD.n34 VDD.n30 0.922
R3176 VDD.n39 VDD.n35 0.922
R3177 VDD.n22 VDD.n18 0.922
R3178 VDD.n27 VDD.n23 0.922
R3179 VDD.n1794 VDD.n1790 0.922
R3180 VDD.n1799 VDD.n1795 0.922
R3181 VDD.n1805 VDD.n1801 0.922
R3182 VDD.n1810 VDD.n1806 0.922
R3183 VDD.n1641 VDD.n1637 0.922
R3184 VDD.n1623 VDD.n1619 0.922
R3185 VDD.n1609 VDD.n1605 0.922
R3186 VDD.n1598 VDD.n1594 0.922
R3187 VDD.n1584 VDD.n1580 0.922
R3188 VDD.n1573 VDD.n1569 0.922
R3189 VDD.n1559 VDD.n1555 0.922
R3190 VDD.n1548 VDD.n1544 0.922
R3191 VDD.n1534 VDD.n1530 0.922
R3192 VDD.n1523 VDD.n1519 0.922
R3193 VDD.n1509 VDD.n1505 0.922
R3194 VDD.n1473 VDD.n1469 0.922
R3195 VDD.n1459 VDD.n1455 0.922
R3196 VDD.n589 VDD.n585 0.922
R3197 VDD.n594 VDD.n590 0.922
R3198 VDD.n624 VDD.n620 0.922
R3199 VDD.n629 VDD.n625 0.922
R3200 VDD.n713 VDD.n709 0.922
R3201 VDD.n718 VDD.n714 0.922
R3202 VDD.n700 VDD.n696 0.922
R3203 VDD.n705 VDD.n701 0.922
R3204 VDD.n560 VDD.n556 0.922
R3205 VDD.n565 VDD.n561 0.922
R3206 VDD.n541 VDD.n537 0.922
R3207 VDD.n546 VDD.n542 0.922
R3208 VDD.n1388 VDD.n1384 0.922
R3209 VDD.n1383 VDD.n1379 0.922
R3210 VDD.n1251 VDD.n1247 0.922
R3211 VDD.n1246 VDD.n1242 0.922
R3212 VDD.n1237 VDD.n1233 0.922
R3213 VDD.n1232 VDD.n1228 0.922
R3214 VDD.n396 VDD.n392 0.922
R3215 VDD.n391 VDD.n387 0.922
R3216 VDD.n83 VDD.n79 0.922
R3217 VDD.n78 VDD.n74 0.922
R3218 VDD.n111 VDD.n107 0.922
R3219 VDD.n106 VDD.n102 0.922
R3220 VDD.n140 VDD.n136 0.922
R3221 VDD.n135 VDD.n131 0.922
R3222 VDD.n168 VDD.n164 0.922
R3223 VDD.n163 VDD.n159 0.922
R3224 VDD.n197 VDD.n193 0.922
R3225 VDD.n192 VDD.n188 0.922
R3226 VDD.n225 VDD.n221 0.922
R3227 VDD.n220 VDD.n216 0.922
R3228 VDD.n361 VDD.n357 0.922
R3229 VDD.n366 VDD.n362 0.922
R3230 VDD.n349 VDD.n345 0.922
R3231 VDD.n354 VDD.n350 0.922
R3232 VDD.n278 VDD.n274 0.922
R3233 VDD.n283 VDD.n279 0.922
R3234 VDD.n266 VDD.n262 0.922
R3235 VDD.n271 VDD.n267 0.922
R3236 VDD.n496 VDD.n492 0.922
R3237 VDD.n501 VDD.n497 0.922
R3238 VDD.n478 VDD.n474 0.922
R3239 VDD.n483 VDD.n479 0.922
R3240 VDD.n874 VDD.n870 0.922
R3241 VDD.n879 VDD.n875 0.922
R3242 VDD.n855 VDD.n851 0.922
R3243 VDD.n860 VDD.n856 0.922
R3244 VDD.n886 VDD.n882 0.922
R3245 VDD.n891 VDD.n887 0.922
R3246 VDD.n923 VDD.n919 0.922
R3247 VDD.n928 VDD.n924 0.922
R3248 VDD.n952 VDD.n948 0.922
R3249 VDD.n957 VDD.n953 0.922
R3250 VDD.n986 VDD.n982 0.922
R3251 VDD.n991 VDD.n987 0.922
R3252 VDD.n1015 VDD.n1011 0.922
R3253 VDD.n1020 VDD.n1016 0.922
R3254 VDD.n1050 VDD.n1046 0.922
R3255 VDD.n1055 VDD.n1051 0.922
R3256 VDD.n1759 VDD.n1755 0.922
R3257 VDD.n1754 VDD.n1750 0.922
R3258 VDD.n1748 VDD.n1744 0.922
R3259 VDD.n1743 VDD.n1739 0.922
R3260 VDD.n33 VDD.n31 0.921
R3261 VDD.n38 VDD.n36 0.921
R3262 VDD.n21 VDD.n19 0.921
R3263 VDD.n26 VDD.n24 0.921
R3264 VDD.n1793 VDD.n1791 0.921
R3265 VDD.n1798 VDD.n1796 0.921
R3266 VDD.n1804 VDD.n1802 0.921
R3267 VDD.n1809 VDD.n1807 0.921
R3268 VDD.n1640 VDD.n1638 0.921
R3269 VDD.n1635 VDD.n1633 0.921
R3270 VDD.n1622 VDD.n1620 0.921
R3271 VDD.n1608 VDD.n1606 0.921
R3272 VDD.n1597 VDD.n1595 0.921
R3273 VDD.n1583 VDD.n1581 0.921
R3274 VDD.n1572 VDD.n1570 0.921
R3275 VDD.n1558 VDD.n1556 0.921
R3276 VDD.n1547 VDD.n1545 0.921
R3277 VDD.n1533 VDD.n1531 0.921
R3278 VDD.n1522 VDD.n1520 0.921
R3279 VDD.n1508 VDD.n1506 0.921
R3280 VDD.n1472 VDD.n1470 0.921
R3281 VDD.n1458 VDD.n1456 0.921
R3282 VDD.n588 VDD.n586 0.921
R3283 VDD.n593 VDD.n591 0.921
R3284 VDD.n623 VDD.n621 0.921
R3285 VDD.n628 VDD.n626 0.921
R3286 VDD.n712 VDD.n710 0.921
R3287 VDD.n717 VDD.n715 0.921
R3288 VDD.n699 VDD.n697 0.921
R3289 VDD.n704 VDD.n702 0.921
R3290 VDD.n559 VDD.n557 0.921
R3291 VDD.n564 VDD.n562 0.921
R3292 VDD.n540 VDD.n538 0.921
R3293 VDD.n545 VDD.n543 0.921
R3294 VDD.n1387 VDD.n1385 0.921
R3295 VDD.n1382 VDD.n1380 0.921
R3296 VDD.n1250 VDD.n1248 0.921
R3297 VDD.n1245 VDD.n1243 0.921
R3298 VDD.n1236 VDD.n1234 0.921
R3299 VDD.n1231 VDD.n1229 0.921
R3300 VDD.n395 VDD.n393 0.921
R3301 VDD.n390 VDD.n388 0.921
R3302 VDD.n82 VDD.n80 0.921
R3303 VDD.n77 VDD.n75 0.921
R3304 VDD.n110 VDD.n108 0.921
R3305 VDD.n105 VDD.n103 0.921
R3306 VDD.n139 VDD.n137 0.921
R3307 VDD.n134 VDD.n132 0.921
R3308 VDD.n167 VDD.n165 0.921
R3309 VDD.n162 VDD.n160 0.921
R3310 VDD.n196 VDD.n194 0.921
R3311 VDD.n191 VDD.n189 0.921
R3312 VDD.n224 VDD.n222 0.921
R3313 VDD.n219 VDD.n217 0.921
R3314 VDD.n360 VDD.n358 0.921
R3315 VDD.n365 VDD.n363 0.921
R3316 VDD.n348 VDD.n346 0.921
R3317 VDD.n353 VDD.n351 0.921
R3318 VDD.n277 VDD.n275 0.921
R3319 VDD.n282 VDD.n280 0.921
R3320 VDD.n265 VDD.n263 0.921
R3321 VDD.n270 VDD.n268 0.921
R3322 VDD.n495 VDD.n493 0.921
R3323 VDD.n500 VDD.n498 0.921
R3324 VDD.n477 VDD.n475 0.921
R3325 VDD.n482 VDD.n480 0.921
R3326 VDD.n873 VDD.n871 0.921
R3327 VDD.n878 VDD.n876 0.921
R3328 VDD.n854 VDD.n852 0.921
R3329 VDD.n859 VDD.n857 0.921
R3330 VDD.n885 VDD.n883 0.921
R3331 VDD.n890 VDD.n888 0.921
R3332 VDD.n922 VDD.n920 0.921
R3333 VDD.n927 VDD.n925 0.921
R3334 VDD.n951 VDD.n949 0.921
R3335 VDD.n956 VDD.n954 0.921
R3336 VDD.n985 VDD.n983 0.921
R3337 VDD.n990 VDD.n988 0.921
R3338 VDD.n1014 VDD.n1012 0.921
R3339 VDD.n1019 VDD.n1017 0.921
R3340 VDD.n1049 VDD.n1047 0.921
R3341 VDD.n1054 VDD.n1052 0.921
R3342 VDD.n1758 VDD.n1756 0.921
R3343 VDD.n1753 VDD.n1751 0.921
R3344 VDD.n1747 VDD.n1745 0.921
R3345 VDD.n1742 VDD.n1740 0.921
R3346 VDD.n1719 VDD.n1714 0.908
R3347 VDD.n1205 VDD.n1200 0.908
R3348 VDD.n651 VDD.n646 0.908
R3349 VDD.n839 VDD.n834 0.908
R3350 VDD.n900 VDD.n895 0.908
R3351 VDD.n969 VDD.n964 0.908
R3352 VDD.n1029 VDD.n1024 0.908
R3353 VDD.n1293 VDD.n1290 0.863
R3354 VDD.n1311 VDD.n1308 0.863
R3355 VDD.n1328 VDD.n1325 0.863
R3356 VDD.n1345 VDD.n1342 0.863
R3357 VDD.n1414 VDD.n1411 0.863
R3358 VDD.n1431 VDD.n1428 0.863
R3359 VDD.n381 VDD.n378 0.863
R3360 VDD.n1276 VDD.n1273 0.863
R3361 VDD.n1688 VDD.n1686 0.85
R3362 VDD.n1678 VDD.n1676 0.85
R3363 VDD.n1081 VDD.n1079 0.85
R3364 VDD.n1089 VDD.n1087 0.85
R3365 VDD.n443 VDD.n441 0.85
R3366 VDD.n434 VDD.n432 0.85
R3367 VDD.n792 VDD.n790 0.85
R3368 VDD.n801 VDD.n799 0.85
R3369 VDD.n1372 VDD.n1370 0.85
R3370 VDD.n1364 VDD.n1362 0.85
R3371 VDD.n1669 VDD.n1667 0.85
R3372 VDD.n1356 VDD.n1354 0.85
R3373 VDD.n1398 VDD.n1396 0.85
R3374 VDD.n1260 VDD.n1258 0.85
R3375 VDD.n426 VDD.n424 0.85
R3376 VDD.n1843 VDD.n1842 0.806
R3377 VDD.n1821 VDD.n1820 0.806
R3378 VDD.n1070 VDD.n1069 0.806
R3379 VDD.n1006 VDD.n1005 0.806
R3380 VDD.n943 VDD.n942 0.806
R3381 VDD.n508 VDD.n507 0.806
R3382 VDD.n579 VDD.n578 0.806
R3383 VDD.n180 VDD.n179 0.806
R3384 VDD.n123 VDD.n122 0.806
R3385 VDD.n237 VDD.n236 0.806
R3386 VDD.n66 VDD.n65 0.806
R3387 VDD.n320 VDD.n319 0.806
R3388 VDD.n298 VDD.n297 0.806
R3389 VDD.n1849 VDD.n1848 0.778
R3390 VDD.n1827 VDD.n1826 0.778
R3391 VDD.n61 VDD.n60 0.778
R3392 VDD.n1125 VDD.n1124 0.778
R3393 VDD.n1155 VDD.n1154 0.778
R3394 VDD.n1185 VDD.n1184 0.778
R3395 VDD.n779 VDD.n778 0.778
R3396 VDD.n572 VDD.n571 0.778
R3397 VDD.n175 VDD.n174 0.778
R3398 VDD.n118 VDD.n117 0.778
R3399 VDD.n232 VDD.n231 0.778
R3400 VDD.n326 VDD.n325 0.778
R3401 VDD.n304 VDD.n303 0.778
R3402 VDD.n1215 VDD.n1213 0.777
R3403 VDD.n662 VDD.n660 0.777
R3404 VDD.n1707 VDD.n1705 0.777
R3405 VDD.n11 VDD.n10 0.747
R3406 VDD.n15 VDD.n14 0.747
R3407 VDD.n3 VDD.n2 0.747
R3408 VDD.n7 VDD.n6 0.747
R3409 VDD.n1832 VDD.n1831 0.747
R3410 VDD.n1836 VDD.n1835 0.747
R3411 VDD.n47 VDD.n46 0.747
R3412 VDD.n44 VDD.n43 0.747
R3413 VDD.n1784 VDD.n1783 0.747
R3414 VDD.n1788 VDD.n1787 0.747
R3415 VDD.n51 VDD.n50 0.747
R3416 VDD.n55 VDD.n54 0.747
R3417 VDD.n1690 VDD.n1689 0.747
R3418 VDD.n1686 VDD.n1685 0.747
R3419 VDD.n1688 VDD.n1687 0.747
R3420 VDD.n1680 VDD.n1679 0.747
R3421 VDD.n1676 VDD.n1675 0.747
R3422 VDD.n1678 VDD.n1677 0.747
R3423 VDD.n1083 VDD.n1082 0.747
R3424 VDD.n1079 VDD.n1078 0.747
R3425 VDD.n1081 VDD.n1080 0.747
R3426 VDD.n1104 VDD.n1103 0.747
R3427 VDD.n1075 VDD.n1074 0.747
R3428 VDD.n1138 VDD.n1137 0.747
R3429 VDD.n1010 VDD.n1009 0.747
R3430 VDD.n1167 VDD.n1166 0.747
R3431 VDD.n947 VDD.n946 0.747
R3432 VDD.n1091 VDD.n1090 0.747
R3433 VDD.n1087 VDD.n1086 0.747
R3434 VDD.n1089 VDD.n1088 0.747
R3435 VDD.n445 VDD.n444 0.747
R3436 VDD.n441 VDD.n440 0.747
R3437 VDD.n443 VDD.n442 0.747
R3438 VDD.n436 VDD.n435 0.747
R3439 VDD.n432 VDD.n431 0.747
R3440 VDD.n434 VDD.n433 0.747
R3441 VDD.n794 VDD.n793 0.747
R3442 VDD.n790 VDD.n789 0.747
R3443 VDD.n792 VDD.n791 0.747
R3444 VDD.n803 VDD.n802 0.747
R3445 VDD.n799 VDD.n798 0.747
R3446 VDD.n801 VDD.n800 0.747
R3447 VDD.n757 VDD.n756 0.747
R3448 VDD.n513 VDD.n512 0.747
R3449 VDD.n734 VDD.n733 0.747
R3450 VDD.n584 VDD.n583 0.747
R3451 VDD.n615 VDD.n614 0.747
R3452 VDD.n598 VDD.n597 0.747
R3453 VDD.n606 VDD.n605 0.747
R3454 VDD.n602 VDD.n601 0.747
R3455 VDD.n690 VDD.n689 0.747
R3456 VDD.n674 VDD.n673 0.747
R3457 VDD.n678 VDD.n677 0.747
R3458 VDD.n684 VDD.n683 0.747
R3459 VDD.n531 VDD.n530 0.747
R3460 VDD.n516 VDD.n515 0.747
R3461 VDD.n519 VDD.n518 0.747
R3462 VDD.n525 VDD.n524 0.747
R3463 VDD.n1374 VDD.n1373 0.747
R3464 VDD.n1370 VDD.n1369 0.747
R3465 VDD.n1372 VDD.n1371 0.747
R3466 VDD.n1366 VDD.n1365 0.747
R3467 VDD.n1362 VDD.n1361 0.747
R3468 VDD.n1364 VDD.n1363 0.747
R3469 VDD.n1671 VDD.n1670 0.747
R3470 VDD.n1667 VDD.n1666 0.747
R3471 VDD.n1669 VDD.n1668 0.747
R3472 VDD.n1358 VDD.n1357 0.747
R3473 VDD.n1354 VDD.n1353 0.747
R3474 VDD.n1356 VDD.n1355 0.747
R3475 VDD.n1393 VDD.n1392 0.747
R3476 VDD.n1396 VDD.n1395 0.747
R3477 VDD.n1398 VDD.n1397 0.747
R3478 VDD.n1262 VDD.n1261 0.747
R3479 VDD.n1258 VDD.n1257 0.747
R3480 VDD.n1260 VDD.n1259 0.747
R3481 VDD.n428 VDD.n427 0.747
R3482 VDD.n424 VDD.n423 0.747
R3483 VDD.n426 VDD.n425 0.747
R3484 VDD.n73 VDD.n72 0.747
R3485 VDD.n69 VDD.n68 0.747
R3486 VDD.n130 VDD.n129 0.747
R3487 VDD.n126 VDD.n125 0.747
R3488 VDD.n187 VDD.n186 0.747
R3489 VDD.n183 VDD.n182 0.747
R3490 VDD.n244 VDD.n243 0.747
R3491 VDD.n240 VDD.n239 0.747
R3492 VDD.n91 VDD.n90 0.747
R3493 VDD.n87 VDD.n86 0.747
R3494 VDD.n94 VDD.n93 0.747
R3495 VDD.n97 VDD.n96 0.747
R3496 VDD.n148 VDD.n147 0.747
R3497 VDD.n144 VDD.n143 0.747
R3498 VDD.n151 VDD.n150 0.747
R3499 VDD.n154 VDD.n153 0.747
R3500 VDD.n205 VDD.n204 0.747
R3501 VDD.n201 VDD.n200 0.747
R3502 VDD.n208 VDD.n207 0.747
R3503 VDD.n211 VDD.n210 0.747
R3504 VDD.n338 VDD.n337 0.747
R3505 VDD.n342 VDD.n341 0.747
R3506 VDD.n330 VDD.n329 0.747
R3507 VDD.n334 VDD.n333 0.747
R3508 VDD.n309 VDD.n308 0.747
R3509 VDD.n313 VDD.n312 0.747
R3510 VDD.n288 VDD.n287 0.747
R3511 VDD.n292 VDD.n291 0.747
R3512 VDD.n255 VDD.n254 0.747
R3513 VDD.n259 VDD.n258 0.747
R3514 VDD.n247 VDD.n246 0.747
R3515 VDD.n251 VDD.n250 0.747
R3516 VDD.n461 VDD.n460 0.747
R3517 VDD.n466 VDD.n465 0.747
R3518 VDD.n449 VDD.n448 0.747
R3519 VDD.n455 VDD.n454 0.747
R3520 VDD.n846 VDD.n845 0.747
R3521 VDD.n831 VDD.n830 0.747
R3522 VDD.n906 VDD.n905 0.747
R3523 VDD.n912 VDD.n911 0.747
R3524 VDD.n976 VDD.n975 0.747
R3525 VDD.n961 VDD.n960 0.747
R3526 VDD.n1041 VDD.n1040 0.747
R3527 VDD.n1035 VDD.n1034 0.747
R3528 VDD.n1767 VDD.n1766 0.747
R3529 VDD.n1763 VDD.n1762 0.747
R3530 VDD.n1770 VDD.n1769 0.747
R3531 VDD.n1773 VDD.n1772 0.747
R3532 VDD.n1222 VDD.n1220 0.74
R3533 VDD.n1700 VDD.n1698 0.74
R3534 VDD.n670 VDD.n668 0.74
R3535 VDD.n12 VDD.n9 0.689
R3536 VDD.n4 VDD.n1 0.689
R3537 VDD.n1833 VDD.n1830 0.689
R3538 VDD.n48 VDD.n45 0.689
R3539 VDD.n1785 VDD.n1782 0.689
R3540 VDD.n52 VDD.n49 0.689
R3541 VDD.n1717 VDD.n1716 0.689
R3542 VDD.n1718 VDD.n1715 0.689
R3543 VDD.n1714 VDD.n1712 0.689
R3544 VDD.n1731 VDD.n1730 0.689
R3545 VDD.n1729 VDD.n1725 0.689
R3546 VDD.n1728 VDD.n1726 0.689
R3547 VDD.n1106 VDD.n1102 0.689
R3548 VDD.n1140 VDD.n1136 0.689
R3549 VDD.n1169 VDD.n1165 0.689
R3550 VDD.n1203 VDD.n1202 0.689
R3551 VDD.n1204 VDD.n1201 0.689
R3552 VDD.n1200 VDD.n1198 0.689
R3553 VDD.n808 VDD.n806 0.689
R3554 VDD.n809 VDD.n805 0.689
R3555 VDD.n811 VDD.n810 0.689
R3556 VDD.n818 VDD.n816 0.689
R3557 VDD.n819 VDD.n815 0.689
R3558 VDD.n821 VDD.n820 0.689
R3559 VDD.n759 VDD.n755 0.689
R3560 VDD.n736 VDD.n732 0.689
R3561 VDD.n649 VDD.n648 0.689
R3562 VDD.n650 VDD.n647 0.689
R3563 VDD.n646 VDD.n644 0.689
R3564 VDD.n617 VDD.n613 0.689
R3565 VDD.n608 VDD.n604 0.689
R3566 VDD.n692 VDD.n688 0.689
R3567 VDD.n680 VDD.n676 0.689
R3568 VDD.n533 VDD.n529 0.689
R3569 VDD.n521 VDD.n517 0.689
R3570 VDD.n418 VDD.n417 0.689
R3571 VDD.n416 VDD.n412 0.689
R3572 VDD.n415 VDD.n413 0.689
R3573 VDD.n407 VDD.n406 0.689
R3574 VDD.n405 VDD.n401 0.689
R3575 VDD.n404 VDD.n402 0.689
R3576 VDD.n70 VDD.n67 0.689
R3577 VDD.n127 VDD.n124 0.689
R3578 VDD.n184 VDD.n181 0.689
R3579 VDD.n241 VDD.n238 0.689
R3580 VDD.n88 VDD.n85 0.689
R3581 VDD.n98 VDD.n95 0.689
R3582 VDD.n145 VDD.n142 0.689
R3583 VDD.n155 VDD.n152 0.689
R3584 VDD.n202 VDD.n199 0.689
R3585 VDD.n212 VDD.n209 0.689
R3586 VDD.n339 VDD.n336 0.689
R3587 VDD.n331 VDD.n328 0.689
R3588 VDD.n310 VDD.n307 0.689
R3589 VDD.n289 VDD.n286 0.689
R3590 VDD.n256 VDD.n253 0.689
R3591 VDD.n248 VDD.n245 0.689
R3592 VDD.n463 VDD.n459 0.689
R3593 VDD.n451 VDD.n447 0.689
R3594 VDD.n848 VDD.n844 0.689
R3595 VDD.n837 VDD.n836 0.689
R3596 VDD.n838 VDD.n835 0.689
R3597 VDD.n834 VDD.n832 0.689
R3598 VDD.n908 VDD.n904 0.689
R3599 VDD.n898 VDD.n897 0.689
R3600 VDD.n899 VDD.n896 0.689
R3601 VDD.n895 VDD.n893 0.689
R3602 VDD.n978 VDD.n974 0.689
R3603 VDD.n967 VDD.n966 0.689
R3604 VDD.n968 VDD.n965 0.689
R3605 VDD.n964 VDD.n962 0.689
R3606 VDD.n1043 VDD.n1039 0.689
R3607 VDD.n1027 VDD.n1026 0.689
R3608 VDD.n1028 VDD.n1025 0.689
R3609 VDD.n1024 VDD.n1022 0.689
R3610 VDD.n1764 VDD.n1761 0.689
R3611 VDD.n1774 VDD.n1771 0.689
R3612 VDD.n34 VDD.n33 0.686
R3613 VDD.n39 VDD.n38 0.686
R3614 VDD.n22 VDD.n21 0.686
R3615 VDD.n27 VDD.n26 0.686
R3616 VDD.n1794 VDD.n1793 0.686
R3617 VDD.n1799 VDD.n1798 0.686
R3618 VDD.n1805 VDD.n1804 0.686
R3619 VDD.n1810 VDD.n1809 0.686
R3620 VDD.n1641 VDD.n1640 0.686
R3621 VDD.n1636 VDD.n1635 0.686
R3622 VDD.n1623 VDD.n1622 0.686
R3623 VDD.n1609 VDD.n1608 0.686
R3624 VDD.n1598 VDD.n1597 0.686
R3625 VDD.n1584 VDD.n1583 0.686
R3626 VDD.n1573 VDD.n1572 0.686
R3627 VDD.n1559 VDD.n1558 0.686
R3628 VDD.n1548 VDD.n1547 0.686
R3629 VDD.n1534 VDD.n1533 0.686
R3630 VDD.n1523 VDD.n1522 0.686
R3631 VDD.n1509 VDD.n1508 0.686
R3632 VDD.n1473 VDD.n1472 0.686
R3633 VDD.n1459 VDD.n1458 0.686
R3634 VDD.n589 VDD.n588 0.686
R3635 VDD.n594 VDD.n593 0.686
R3636 VDD.n624 VDD.n623 0.686
R3637 VDD.n629 VDD.n628 0.686
R3638 VDD.n713 VDD.n712 0.686
R3639 VDD.n718 VDD.n717 0.686
R3640 VDD.n700 VDD.n699 0.686
R3641 VDD.n705 VDD.n704 0.686
R3642 VDD.n560 VDD.n559 0.686
R3643 VDD.n565 VDD.n564 0.686
R3644 VDD.n541 VDD.n540 0.686
R3645 VDD.n546 VDD.n545 0.686
R3646 VDD.n1388 VDD.n1387 0.686
R3647 VDD.n1383 VDD.n1382 0.686
R3648 VDD.n1251 VDD.n1250 0.686
R3649 VDD.n1246 VDD.n1245 0.686
R3650 VDD.n1232 VDD.n1231 0.686
R3651 VDD.n1237 VDD.n1236 0.686
R3652 VDD.n396 VDD.n395 0.686
R3653 VDD.n391 VDD.n390 0.686
R3654 VDD.n78 VDD.n77 0.686
R3655 VDD.n83 VDD.n82 0.686
R3656 VDD.n106 VDD.n105 0.686
R3657 VDD.n111 VDD.n110 0.686
R3658 VDD.n135 VDD.n134 0.686
R3659 VDD.n140 VDD.n139 0.686
R3660 VDD.n163 VDD.n162 0.686
R3661 VDD.n168 VDD.n167 0.686
R3662 VDD.n192 VDD.n191 0.686
R3663 VDD.n197 VDD.n196 0.686
R3664 VDD.n220 VDD.n219 0.686
R3665 VDD.n225 VDD.n224 0.686
R3666 VDD.n361 VDD.n360 0.686
R3667 VDD.n366 VDD.n365 0.686
R3668 VDD.n349 VDD.n348 0.686
R3669 VDD.n354 VDD.n353 0.686
R3670 VDD.n278 VDD.n277 0.686
R3671 VDD.n283 VDD.n282 0.686
R3672 VDD.n266 VDD.n265 0.686
R3673 VDD.n271 VDD.n270 0.686
R3674 VDD.n496 VDD.n495 0.686
R3675 VDD.n501 VDD.n500 0.686
R3676 VDD.n478 VDD.n477 0.686
R3677 VDD.n483 VDD.n482 0.686
R3678 VDD.n874 VDD.n873 0.686
R3679 VDD.n879 VDD.n878 0.686
R3680 VDD.n855 VDD.n854 0.686
R3681 VDD.n860 VDD.n859 0.686
R3682 VDD.n886 VDD.n885 0.686
R3683 VDD.n891 VDD.n890 0.686
R3684 VDD.n923 VDD.n922 0.686
R3685 VDD.n928 VDD.n927 0.686
R3686 VDD.n952 VDD.n951 0.686
R3687 VDD.n957 VDD.n956 0.686
R3688 VDD.n986 VDD.n985 0.686
R3689 VDD.n991 VDD.n990 0.686
R3690 VDD.n1015 VDD.n1014 0.686
R3691 VDD.n1020 VDD.n1019 0.686
R3692 VDD.n1050 VDD.n1049 0.686
R3693 VDD.n1055 VDD.n1054 0.686
R3694 VDD.n1759 VDD.n1758 0.686
R3695 VDD.n1754 VDD.n1753 0.686
R3696 VDD.n1748 VDD.n1747 0.686
R3697 VDD.n1743 VDD.n1742 0.686
R3698 VDD.n1735 VDD.n1672 0.675
R3699 VDD.n1294 VDD.n1293 0.646
R3700 VDD.n1312 VDD.n1311 0.646
R3701 VDD.n1329 VDD.n1328 0.646
R3702 VDD.n1346 VDD.n1345 0.646
R3703 VDD.n1415 VDD.n1414 0.646
R3704 VDD.n1432 VDD.n1431 0.646
R3705 VDD.n382 VDD.n381 0.646
R3706 VDD.n1277 VDD.n1276 0.646
R3707 VDD.n12 VDD.n11 0.59
R3708 VDD.n4 VDD.n3 0.59
R3709 VDD.n1833 VDD.n1832 0.59
R3710 VDD.n48 VDD.n47 0.59
R3711 VDD.n1785 VDD.n1784 0.59
R3712 VDD.n52 VDD.n51 0.59
R3713 VDD.n70 VDD.n69 0.59
R3714 VDD.n127 VDD.n126 0.59
R3715 VDD.n184 VDD.n183 0.59
R3716 VDD.n241 VDD.n240 0.59
R3717 VDD.n88 VDD.n87 0.59
R3718 VDD.n98 VDD.n97 0.59
R3719 VDD.n145 VDD.n144 0.59
R3720 VDD.n155 VDD.n154 0.59
R3721 VDD.n202 VDD.n201 0.59
R3722 VDD.n212 VDD.n211 0.59
R3723 VDD.n339 VDD.n338 0.59
R3724 VDD.n331 VDD.n330 0.59
R3725 VDD.n310 VDD.n309 0.59
R3726 VDD.n289 VDD.n288 0.59
R3727 VDD.n256 VDD.n255 0.59
R3728 VDD.n248 VDD.n247 0.59
R3729 VDD.n1764 VDD.n1763 0.59
R3730 VDD.n1774 VDD.n1773 0.59
R3731 VDD.n1491 VDD.n1489 0.587
R3732 VDD.n1486 VDD.n1484 0.587
R3733 VDD.n1139 VDD.n1138 0.571
R3734 VDD.n607 VDD.n606 0.571
R3735 VDD.n691 VDD.n690 0.571
R3736 VDD.n532 VDD.n531 0.571
R3737 VDD.n520 VDD.n519 0.571
R3738 VDD.n462 VDD.n461 0.571
R3739 VDD.n450 VDD.n449 0.571
R3740 VDD.n907 VDD.n906 0.571
R3741 VDD.n1042 VDD.n1041 0.571
R3742 VDD.n735 VDD.n734 0.57
R3743 VDD.n616 VDD.n615 0.57
R3744 VDD.n847 VDD.n846 0.57
R3745 VDD.n1105 VDD.n1104 0.569
R3746 VDD.n1168 VDD.n1167 0.569
R3747 VDD.n758 VDD.n757 0.569
R3748 VDD.n679 VDD.n678 0.569
R3749 VDD.n977 VDD.n976 0.569
R3750 VDD.n1732 VDD.n1731 0.5
R3751 VDD.n812 VDD.n811 0.5
R3752 VDD.n822 VDD.n821 0.5
R3753 VDD.n419 VDD.n418 0.5
R3754 VDD.n408 VDD.n407 0.5
R3755 VDD.n1732 VDD.n1729 0.483
R3756 VDD.n812 VDD.n809 0.483
R3757 VDD.n822 VDD.n819 0.483
R3758 VDD.n419 VDD.n416 0.483
R3759 VDD.n408 VDD.n405 0.483
R3760 VDD.n763 VDD.n513 0.452
R3761 VDD.n619 VDD.n598 0.452
R3762 VDD.n981 VDD.n961 0.452
R3763 VDD.n1110 VDD.n1075 0.452
R3764 VDD.n1174 VDD.n947 0.452
R3765 VDD.n738 VDD.n584 0.452
R3766 VDD.n850 VDD.n831 0.452
R3767 VDD.n685 VDD.n684 0.452
R3768 VDD.n1143 VDD.n1010 0.451
R3769 VDD.n695 VDD.n674 0.451
R3770 VDD.n536 VDD.n516 0.451
R3771 VDD.n16 VDD.n15 0.451
R3772 VDD.n8 VDD.n7 0.451
R3773 VDD.n1837 VDD.n1836 0.451
R3774 VDD.n1816 VDD.n44 0.451
R3775 VDD.n1789 VDD.n1788 0.451
R3776 VDD.n56 VDD.n55 0.451
R3777 VDD.n1450 VDD.n73 0.451
R3778 VDD.n1446 VDD.n130 0.451
R3779 VDD.n1442 VDD.n187 0.451
R3780 VDD.n1438 VDD.n244 0.451
R3781 VDD.n100 VDD.n91 0.451
R3782 VDD.n99 VDD.n94 0.451
R3783 VDD.n157 VDD.n148 0.451
R3784 VDD.n156 VDD.n151 0.451
R3785 VDD.n214 VDD.n205 0.451
R3786 VDD.n213 VDD.n208 0.451
R3787 VDD.n343 VDD.n342 0.451
R3788 VDD.n335 VDD.n334 0.451
R3789 VDD.n314 VDD.n313 0.451
R3790 VDD.n293 VDD.n292 0.451
R3791 VDD.n260 VDD.n259 0.451
R3792 VDD.n252 VDD.n251 0.451
R3793 VDD.n1776 VDD.n1767 0.451
R3794 VDD.n1775 VDD.n1770 0.451
R3795 VDD.n526 VDD.n525 0.451
R3796 VDD.n456 VDD.n455 0.451
R3797 VDD.n603 VDD.n602 0.45
R3798 VDD.n1036 VDD.n1035 0.449
R3799 VDD.n1092 VDD.n1091 0.433
R3800 VDD.n467 VDD.n466 0.419
R3801 VDD.n913 VDD.n912 0.419
R3802 VDD.n1092 VDD.n1089 0.416
R3803 VDD.n1072 VDD.n1071 0.4
R3804 VDD.n1157 VDD.n1156 0.4
R3805 VDD.n510 VDD.n509 0.4
R3806 VDD.n781 VDD.n780 0.4
R3807 VDD.n581 VDD.n580 0.4
R3808 VDD.n574 VDD.n573 0.4
R3809 VDD.n1662 VDD.n1661 0.398
R3810 VDD.n1661 VDD.n1660 0.398
R3811 VDD.n1660 VDD.n1659 0.398
R3812 VDD.n1659 VDD.n1658 0.398
R3813 VDD.n1658 VDD.n1657 0.398
R3814 VDD.n1657 VDD.n1656 0.398
R3815 VDD.n1656 VDD.n1655 0.398
R3816 VDD.n84 VDD.n78 0.345
R3817 VDD.n112 VDD.n106 0.345
R3818 VDD.n141 VDD.n135 0.345
R3819 VDD.n169 VDD.n163 0.345
R3820 VDD.n198 VDD.n192 0.345
R3821 VDD.n226 VDD.n220 0.345
R3822 VDD.n1238 VDD.n1232 0.343
R3823 VDD.n1238 VDD.n1237 0.343
R3824 VDD.n1760 VDD.n1754 0.342
R3825 VDD.n1749 VDD.n1743 0.342
R3826 VDD.n84 VDD.n83 0.34
R3827 VDD.n112 VDD.n111 0.34
R3828 VDD.n141 VDD.n140 0.34
R3829 VDD.n169 VDD.n168 0.34
R3830 VDD.n198 VDD.n197 0.34
R3831 VDD.n226 VDD.n225 0.34
R3832 VDD.n1760 VDD.n1759 0.336
R3833 VDD.n1749 VDD.n1748 0.336
R3834 VDD.n1642 VDD.n1636 0.334
R3835 VDD.n1438 VDD.n1437 0.326
R3836 VDD.n1642 VDD.n1641 0.305
R3837 VDD.n786 VDD.n785 0.303
R3838 VDD.n663 VDD.n662 0.296
R3839 VDD.n1710 VDD.n1707 0.296
R3840 VDD.n1216 VDD.n1215 0.295
R3841 VDD.n1223 VDD.n1222 0.286
R3842 VDD.n1225 VDD.n828 0.286
R3843 VDD.n1701 VDD.n1700 0.285
R3844 VDD.n671 VDD.n670 0.285
R3845 VDD.n1492 VDD.n1486 0.284
R3846 VDD.n828 VDD.n827 0.283
R3847 VDD.n1663 VDD.n1662 0.28
R3848 VDD.n1722 VDD.n1693 0.277
R3849 VDD.n17 VDD.n8 0.276
R3850 VDD.n344 VDD.n335 0.276
R3851 VDD.n261 VDD.n252 0.276
R3852 VDD.n903 VDD.n902 0.272
R3853 VDD.n842 VDD.n841 0.272
R3854 VDD.n100 VDD.n99 0.272
R3855 VDD.n157 VDD.n156 0.272
R3856 VDD.n214 VDD.n213 0.272
R3857 VDD.n1776 VDD.n1775 0.272
R3858 VDD.n972 VDD.n971 0.271
R3859 VDD.n1032 VDD.n1031 0.271
R3860 VDD.n528 VDD.n527 0.271
R3861 VDD.n458 VDD.n457 0.271
R3862 VDD.n611 VDD.n610 0.271
R3863 VDD.n687 VDD.n686 0.271
R3864 VDD.n1492 VDD.n1491 0.255
R3865 VDD.n1443 VDD.n180 0.254
R3866 VDD.n1447 VDD.n123 0.254
R3867 VDD.n1439 VDD.n237 0.254
R3868 VDD.n1451 VDD.n66 0.254
R3869 VDD.n1844 VDD.n1843 0.253
R3870 VDD.n1822 VDD.n1821 0.253
R3871 VDD.n321 VDD.n320 0.253
R3872 VDD.n299 VDD.n298 0.253
R3873 VDD.n1264 VDD.n1254 0.252
R3874 VDD.n729 VDD.n728 0.244
R3875 VDD.n1452 VDD.n61 0.242
R3876 VDD.n1444 VDD.n175 0.242
R3877 VDD.n1448 VDD.n118 0.242
R3878 VDD.n1440 VDD.n232 0.242
R3879 VDD.n1850 VDD.n1849 0.241
R3880 VDD.n1828 VDD.n1827 0.241
R3881 VDD.n327 VDD.n326 0.241
R3882 VDD.n305 VDD.n304 0.241
R3883 VDD.n1391 VDD.n1378 0.233
R3884 VDD.n1072 VDD.n1070 0.23
R3885 VDD.n1007 VDD.n1006 0.23
R3886 VDD.n944 VDD.n943 0.23
R3887 VDD.n510 VDD.n508 0.23
R3888 VDD.n581 VDD.n579 0.23
R3889 VDD.n1126 VDD.n1125 0.218
R3890 VDD.n1157 VDD.n1155 0.218
R3891 VDD.n1186 VDD.n1185 0.218
R3892 VDD.n781 VDD.n779 0.218
R3893 VDD.n574 VDD.n572 0.218
R3894 VDD.n386 VDD.n369 0.215
R3895 VDD.n1691 VDD.n1690 0.208
R3896 VDD.n1681 VDD.n1680 0.208
R3897 VDD.n1084 VDD.n1083 0.208
R3898 VDD.n446 VDD.n445 0.208
R3899 VDD.n437 VDD.n436 0.208
R3900 VDD.n795 VDD.n794 0.208
R3901 VDD.n804 VDD.n803 0.208
R3902 VDD.n1375 VDD.n1374 0.208
R3903 VDD.n1376 VDD.n1366 0.208
R3904 VDD.n1672 VDD.n1671 0.208
R3905 VDD.n1378 VDD.n1358 0.208
R3906 VDD.n1400 VDD.n1393 0.208
R3907 VDD.n1263 VDD.n1262 0.208
R3908 VDD.n1227 VDD.n428 0.208
R3909 VDD.n1389 VDD.n1383 0.203
R3910 VDD.n1252 VDD.n1246 0.203
R3911 VDD.n397 VDD.n391 0.203
R3912 VDD.n1691 VDD.n1688 0.195
R3913 VDD.n1681 VDD.n1678 0.195
R3914 VDD.n1084 VDD.n1081 0.195
R3915 VDD.n446 VDD.n443 0.195
R3916 VDD.n437 VDD.n434 0.195
R3917 VDD.n795 VDD.n792 0.195
R3918 VDD.n804 VDD.n801 0.195
R3919 VDD.n1375 VDD.n1372 0.195
R3920 VDD.n1376 VDD.n1364 0.195
R3921 VDD.n1672 VDD.n1669 0.195
R3922 VDD.n1378 VDD.n1356 0.195
R3923 VDD.n1400 VDD.n1398 0.195
R3924 VDD.n1263 VDD.n1260 0.195
R3925 VDD.n1227 VDD.n426 0.195
R3926 VDD.n410 VDD.n399 0.195
R3927 VDD.n1240 VDD.n1227 0.194
R3928 VDD.n1624 VDD.n1623 0.193
R3929 VDD.n1599 VDD.n1598 0.193
R3930 VDD.n1574 VDD.n1573 0.193
R3931 VDD.n1549 VDD.n1548 0.193
R3932 VDD.n1524 VDD.n1523 0.193
R3933 VDD.n1474 VDD.n1473 0.193
R3934 VDD.n1610 VDD.n1609 0.189
R3935 VDD.n1585 VDD.n1584 0.189
R3936 VDD.n1560 VDD.n1559 0.189
R3937 VDD.n1535 VDD.n1534 0.189
R3938 VDD.n1510 VDD.n1509 0.189
R3939 VDD.n1460 VDD.n1459 0.189
R3940 VDD.n643 VDD.n640 0.186
R3941 VDD.n1164 VDD.n1163 0.186
R3942 VDD.n1226 VDD.n786 0.185
R3943 VDD.n730 VDD.n729 0.185
R3944 VDD.n1197 VDD.n1194 0.184
R3945 VDD.n752 VDD.n751 0.182
R3946 VDD.n657 VDD.n653 0.182
R3947 VDD.n764 VDD.n763 0.182
R3948 VDD.n1851 VDD.n41 0.182
R3949 VDD.n1135 VDD.n1134 0.18
R3950 VDD.n1098 VDD.n1097 0.18
R3951 VDD.n40 VDD.n39 0.179
R3952 VDD.n28 VDD.n27 0.179
R3953 VDD.n1800 VDD.n1799 0.179
R3954 VDD.n1811 VDD.n1810 0.179
R3955 VDD.n595 VDD.n594 0.179
R3956 VDD.n630 VDD.n629 0.179
R3957 VDD.n719 VDD.n718 0.179
R3958 VDD.n706 VDD.n705 0.179
R3959 VDD.n566 VDD.n565 0.179
R3960 VDD.n547 VDD.n546 0.179
R3961 VDD.n367 VDD.n366 0.179
R3962 VDD.n355 VDD.n354 0.179
R3963 VDD.n284 VDD.n283 0.179
R3964 VDD.n272 VDD.n271 0.179
R3965 VDD.n502 VDD.n501 0.179
R3966 VDD.n484 VDD.n483 0.179
R3967 VDD.n880 VDD.n879 0.179
R3968 VDD.n861 VDD.n860 0.179
R3969 VDD.n892 VDD.n891 0.179
R3970 VDD.n929 VDD.n928 0.179
R3971 VDD.n958 VDD.n957 0.179
R3972 VDD.n992 VDD.n991 0.179
R3973 VDD.n1021 VDD.n1020 0.179
R3974 VDD.n1056 VDD.n1055 0.179
R3975 VDD.n1778 VDD.n1777 0.177
R3976 VDD.n1111 VDD.n1110 0.177
R3977 VDD.n1144 VDD.n1143 0.176
R3978 VDD.n869 VDD.n862 0.175
R3979 VDD.n937 VDD.n930 0.175
R3980 VDD.n1000 VDD.n993 0.175
R3981 VDD.n638 VDD.n631 0.175
R3982 VDD.n1064 VDD.n1057 0.175
R3983 VDD.n503 VDD.n485 0.175
R3984 VDD.n555 VDD.n548 0.174
R3985 VDD.n1175 VDD.n1174 0.174
R3986 VDD.n113 VDD.n101 0.174
R3987 VDD.n170 VDD.n158 0.174
R3988 VDD.n227 VDD.n215 0.174
R3989 VDD.n368 VDD.n356 0.174
R3990 VDD.n285 VDD.n273 0.174
R3991 VDD.n1813 VDD.n1812 0.174
R3992 VDD.n41 VDD.n29 0.174
R3993 VDD.n1210 VDD.n1207 0.173
R3994 VDD.n1814 VDD.n1813 0.172
R3995 VDD.n1692 VDD.n1691 0.17
R3996 VDD.n751 VDD.n567 0.168
R3997 VDD.n1097 VDD.n1084 0.168
R3998 VDD.n708 VDD.n707 0.168
R3999 VDD.n1682 VDD.n1681 0.166
R4000 VDD.n315 VDD.n306 0.164
R4001 VDD.n739 VDD.n738 0.164
R4002 VDD.n321 VDD.n315 0.163
R4003 VDD.n1838 VDD.n1829 0.162
R4004 VDD.n1450 VDD.n1449 0.162
R4005 VDD.n631 VDD.n619 0.162
R4006 VDD.n707 VDD.n695 0.162
R4007 VDD.n548 VDD.n536 0.162
R4008 VDD.n862 VDD.n850 0.162
R4009 VDD.n993 VDD.n981 0.162
R4010 VDD.n29 VDD.n17 0.161
R4011 VDD.n356 VDD.n344 0.161
R4012 VDD.n273 VDD.n261 0.161
R4013 VDD.n1446 VDD.n1445 0.161
R4014 VDD.n1822 VDD.n1816 0.161
R4015 VDD.n1451 VDD.n1450 0.161
R4016 VDD.n485 VDD.n473 0.161
R4017 VDD.n930 VDD.n918 0.161
R4018 VDD.n1057 VDD.n1045 0.161
R4019 VDD.n1844 VDD.n1838 0.16
R4020 VDD.n1442 VDD.n1441 0.16
R4021 VDD.n1711 VDD.n1710 0.159
R4022 VDD.n101 VDD.n100 0.159
R4023 VDD.n158 VDD.n157 0.159
R4024 VDD.n215 VDD.n214 0.159
R4025 VDD.n1777 VDD.n1776 0.159
R4026 VDD.n1439 VDD.n1438 0.158
R4027 VDD.n1443 VDD.n1442 0.158
R4028 VDD.n1447 VDD.n1446 0.158
R4029 VDD.n1779 VDD.n1778 0.158
R4030 VDD.n640 VDD.n639 0.155
R4031 VDD.n1777 VDD.n1760 0.15
R4032 VDD.n1778 VDD.n1749 0.15
R4033 VDD.n299 VDD.n293 0.145
R4034 VDD.n41 VDD.n40 0.143
R4035 VDD.n29 VDD.n28 0.142
R4036 VDD.n1813 VDD.n1800 0.142
R4037 VDD.n631 VDD.n630 0.142
R4038 VDD.n707 VDD.n706 0.142
R4039 VDD.n548 VDD.n547 0.142
R4040 VDD.n356 VDD.n355 0.142
R4041 VDD.n273 VDD.n272 0.142
R4042 VDD.n485 VDD.n484 0.142
R4043 VDD.n862 VDD.n861 0.142
R4044 VDD.n930 VDD.n929 0.142
R4045 VDD.n993 VDD.n992 0.142
R4046 VDD.n1057 VDD.n1056 0.142
R4047 VDD.n1812 VDD.n1811 0.141
R4048 VDD.n368 VDD.n367 0.141
R4049 VDD.n285 VDD.n284 0.141
R4050 VDD.n1401 VDD.n1391 0.131
R4051 VDD.n1240 VDD.n1238 0.129
R4052 VDD.n1449 VDD.n113 0.129
R4053 VDD.n306 VDD.n285 0.129
R4054 VDD.n1445 VDD.n170 0.128
R4055 VDD.n1441 VDD.n227 0.128
R4056 VDD.n783 VDD.n503 0.128
R4057 VDD.n1224 VDD.n881 0.128
R4058 VDD.n1194 VDD.n938 0.128
R4059 VDD.n1163 VDD.n1001 0.128
R4060 VDD.n1134 VDD.n1065 0.128
R4061 VDD.n639 VDD.n595 0.125
R4062 VDD.n727 VDD.n719 0.125
R4063 VDD.n881 VDD.n880 0.125
R4064 VDD.n938 VDD.n892 0.125
R4065 VDD.n1001 VDD.n958 0.125
R4066 VDD.n1065 VDD.n1021 0.125
R4067 VDD.n503 VDD.n502 0.124
R4068 VDD.n567 VDD.n566 0.123
R4069 VDD.n1297 VDD.n1294 0.118
R4070 VDD.n1315 VDD.n1312 0.118
R4071 VDD.n1332 VDD.n1329 0.118
R4072 VDD.n1349 VDD.n1346 0.118
R4073 VDD.n1418 VDD.n1415 0.118
R4074 VDD.n1435 VDD.n1432 0.118
R4075 VDD.n385 VDD.n382 0.118
R4076 VDD.n1280 VDD.n1277 0.118
R4077 VDD.n1722 VDD.n1721 0.117
R4078 VDD.n369 VDD.n368 0.117
R4079 VDD.n827 VDD.n804 0.114
R4080 VDD.n1241 VDD.n1240 0.113
R4081 VDD.n828 VDD.n795 0.113
R4082 VDD.n369 VDD.n327 0.111
R4083 VDD.n1099 VDD.n1098 0.105
R4084 VDD.n1281 VDD.n1264 0.104
R4085 VDD.n1815 VDD.n1814 0.102
R4086 VDD.n785 VDD.n446 0.1
R4087 VDD.n786 VDD.n437 0.1
R4088 VDD.n1734 VDD.n1723 0.098
R4089 VDD.n1779 VDD.n1738 0.098
R4090 VDD.n1160 VDD.n1150 0.098
R4091 VDD.n773 VDD.n772 0.097
R4092 VDD.n743 VDD.n742 0.097
R4093 VDD.n748 VDD.n747 0.097
R4094 VDD.n1735 VDD.n1734 0.097
R4095 VDD.n1288 VDD.n1284 0.095
R4096 VDD.n1306 VDD.n1302 0.095
R4097 VDD.n1323 VDD.n1319 0.095
R4098 VDD.n1340 VDD.n1336 0.095
R4099 VDD.n1409 VDD.n1405 0.095
R4100 VDD.n1426 VDD.n1422 0.095
R4101 VDD.n376 VDD.n372 0.095
R4102 VDD.n1271 VDD.n1267 0.095
R4103 VDD.n1116 VDD.n1115 0.093
R4104 VDD.n1738 VDD.n1737 0.088
R4105 VDD.n1781 VDD.n1780 0.088
R4106 VDD.n771 VDD.n770 0.086
R4107 VDD.n665 VDD.n664 0.085
R4108 VDD.n1736 VDD.n1735 0.083
R4109 VDD.n1814 VDD.n1781 0.082
R4110 VDD.n1120 VDD.n1119 0.082
R4111 VDD.n1149 VDD.n1148 0.082
R4112 VDD.n1217 VDD.n1216 0.081
R4113 VDD.n1180 VDD.n1179 0.081
R4114 VDD.n327 VDD.n321 0.078
R4115 VDD.n746 VDD.n745 0.077
R4116 VDD.n1710 VDD.n1702 0.076
R4117 VDD.n1452 VDD.n1451 0.075
R4118 VDD.n1850 VDD.n1844 0.075
R4119 VDD.n1828 VDD.n1822 0.075
R4120 VDD.n305 VDD.n299 0.075
R4121 VDD.n1719 VDD.n1718 0.075
R4122 VDD.n1205 VDD.n1204 0.075
R4123 VDD.n651 VDD.n650 0.075
R4124 VDD.n839 VDD.n838 0.075
R4125 VDD.n900 VDD.n899 0.075
R4126 VDD.n969 VDD.n968 0.075
R4127 VDD.n1029 VDD.n1028 0.075
R4128 VDD.n1436 VDD.n1419 0.073
R4129 VDD.n1440 VDD.n1439 0.073
R4130 VDD.n1444 VDD.n1443 0.073
R4131 VDD.n1448 VDD.n1447 0.073
R4132 VDD.n1736 VDD.n1663 0.062
R4133 VDD.n101 VDD.n84 0.062
R4134 VDD.n113 VDD.n112 0.062
R4135 VDD.n158 VDD.n141 0.062
R4136 VDD.n170 VDD.n169 0.062
R4137 VDD.n215 VDD.n198 0.062
R4138 VDD.n227 VDD.n226 0.062
R4139 VDD.n1333 VDD.n410 0.061
R4140 VDD.n1350 VDD.n1333 0.061
R4141 VDD.n1333 VDD.n1316 0.06
R4142 VDD.n1643 VDD.n1642 0.059
R4143 VDD.n1493 VDD.n1492 0.059
R4144 VDD.n785 VDD.n784 0.057
R4145 VDD.n1299 VDD.n1298 0.055
R4146 VDD.n410 VDD.n409 0.055
R4147 VDD.n1733 VDD.n1732 0.054
R4148 VDD.n1095 VDD.n1092 0.054
R4149 VDD.n814 VDD.n812 0.054
R4150 VDD.n824 VDD.n822 0.054
R4151 VDD.n420 VDD.n419 0.054
R4152 VDD.n409 VDD.n408 0.054
R4153 VDD.n1402 VDD.n1401 0.054
R4154 VDD.n1378 VDD.n1377 0.053
R4155 VDD.n1264 VDD.n1263 0.053
R4156 VDD.n1227 VDD.n1226 0.051
R4157 VDD.n1419 VDD.n1402 0.049
R4158 VDD.n1225 VDD.n1224 0.048
R4159 VDD.n1737 VDD.n1454 0.047
R4160 VDD.n1031 VDD.n1029 0.047
R4161 VDD.n1299 VDD.n1241 0.046
R4162 VDD.n902 VDD.n900 0.045
R4163 VDD.n1720 VDD.n1719 0.045
R4164 VDD.n1206 VDD.n1205 0.045
R4165 VDD.n652 VDD.n651 0.045
R4166 VDD.n971 VDD.n969 0.045
R4167 VDD.n841 VDD.n839 0.044
R4168 VDD.n784 VDD.n783 0.044
R4169 VDD.n1738 VDD.n1453 0.043
R4170 VDD.n471 VDD.n470 0.043
R4171 VDD.n916 VDD.n915 0.042
R4172 VDD.n761 VDD.n753 0.042
R4173 VDD.n1117 VDD.n1112 0.042
R4174 VDD.n1108 VDD.n1100 0.041
R4175 VDD.n1191 VDD.n1190 0.041
R4176 VDD.n1131 VDD.n1130 0.04
R4177 VDD.n1172 VDD.n1170 0.04
R4178 VDD.n1401 VDD.n1400 0.039
R4179 VDD.n1737 VDD.n1736 0.038
R4180 VDD.n1437 VDD.n1436 0.037
R4181 VDD.n1241 VDD.n420 0.037
R4182 VDD.n1437 VDD.n386 0.036
R4183 VDD.n1226 VDD.n1225 0.032
R4184 VDD.n1631 VDD.n1630 0.03
R4185 VDD.n1627 VDD.n1626 0.03
R4186 VDD.n1602 VDD.n1601 0.03
R4187 VDD.n1577 VDD.n1576 0.03
R4188 VDD.n1552 VDD.n1551 0.03
R4189 VDD.n1527 VDD.n1526 0.03
R4190 VDD.n1481 VDD.n1480 0.03
R4191 VDD.n1477 VDD.n1476 0.03
R4192 VDD.n1391 VDD.n1389 0.03
R4193 VDD.n1254 VDD.n1252 0.03
R4194 VDD.n399 VDD.n397 0.03
R4195 VDD.n1298 VDD.n1281 0.03
R4196 VDD.n469 VDD.n467 0.03
R4197 VDD.n914 VDD.n913 0.03
R4198 VDD.n1224 VDD.n1223 0.027
R4199 VDD.n1163 VDD.n1162 0.026
R4200 VDD.n1134 VDD.n1133 0.026
R4201 VDD.n783 VDD.n782 0.025
R4202 VDD.n1194 VDD.n1193 0.025
R4203 VDD.n1721 VDD.n1695 0.023
R4204 VDD.n643 VDD.n642 0.023
R4205 VDD.n1197 VDD.n1196 0.023
R4206 VDD.n1653 VDD.n1644 0.023
R4207 VDD.n1503 VDD.n1494 0.023
R4208 VDD.n1441 VDD.n1440 0.023
R4209 VDD.n1445 VDD.n1444 0.023
R4210 VDD.n1449 VDD.n1448 0.023
R4211 VDD.n306 VDD.n305 0.023
R4212 VDD.n1829 VDD.n1828 0.023
R4213 VDD.n0 VDD 0.022
R4214 VDD VDD.n0 0.022
R4215 VDD.n751 VDD.n750 0.022
R4216 VDD.n782 VDD.n781 0.021
R4217 VDD.n1625 VDD.n1624 0.021
R4218 VDD.n1617 VDD.n1610 0.021
R4219 VDD.n1600 VDD.n1599 0.021
R4220 VDD.n1592 VDD.n1585 0.021
R4221 VDD.n1575 VDD.n1574 0.021
R4222 VDD.n1567 VDD.n1560 0.021
R4223 VDD.n1550 VDD.n1549 0.021
R4224 VDD.n1542 VDD.n1535 0.021
R4225 VDD.n1525 VDD.n1524 0.021
R4226 VDD.n1517 VDD.n1510 0.021
R4227 VDD.n1475 VDD.n1474 0.021
R4228 VDD.n1467 VDD.n1460 0.021
R4229 VDD.n759 VDD.n758 0.021
R4230 VDD.n1851 VDD.n1850 0.02
R4231 VDD.n1148 VDD.n1007 0.02
R4232 VDD.n1179 VDD.n944 0.02
R4233 VDD.n745 VDD.n581 0.02
R4234 VDD.n750 VDD.n574 0.02
R4235 VDD.n770 VDD.n510 0.02
R4236 VDD.n1119 VDD.n1072 0.02
R4237 VDD.n1106 VDD.n1105 0.02
R4238 VDD.n1169 VDD.n1168 0.02
R4239 VDD.n736 VDD.n735 0.02
R4240 VDD.n617 VDD.n616 0.02
R4241 VDD.n680 VDD.n679 0.02
R4242 VDD.n848 VDD.n847 0.02
R4243 VDD.n978 VDD.n977 0.02
R4244 VDD.n1814 VDD.n1789 0.019
R4245 VDD.n1140 VDD.n1139 0.019
R4246 VDD.n608 VDD.n607 0.019
R4247 VDD.n692 VDD.n691 0.019
R4248 VDD.n533 VDD.n532 0.019
R4249 VDD.n521 VDD.n520 0.019
R4250 VDD.n451 VDD.n450 0.019
R4251 VDD.n1402 VDD.n1350 0.018
R4252 VDD.n463 VDD.n462 0.018
R4253 VDD.n908 VDD.n907 0.018
R4254 VDD.n1043 VDD.n1042 0.018
R4255 VDD.n729 VDD.n671 0.016
R4256 VDD.n1644 VDD.n1643 0.015
R4257 VDD.n1494 VDD.n1493 0.015
R4258 VDD.n1780 VDD.n1779 0.012
R4259 VDD VDD.n1851 0.011
R4260 VDD.n16 VDD.n12 0.011
R4261 VDD.n8 VDD.n4 0.011
R4262 VDD.n1837 VDD.n1833 0.011
R4263 VDD.n1816 VDD.n48 0.011
R4264 VDD.n1789 VDD.n1785 0.011
R4265 VDD.n56 VDD.n52 0.011
R4266 VDD.n1127 VDD.n1126 0.011
R4267 VDD.n1158 VDD.n1157 0.011
R4268 VDD.n1142 VDD.n1140 0.011
R4269 VDD.n1187 VDD.n1186 0.011
R4270 VDD.n737 VDD.n736 0.011
R4271 VDD.n609 VDD.n608 0.011
R4272 VDD.n694 VDD.n692 0.011
R4273 VDD.n535 VDD.n533 0.011
R4274 VDD.n526 VDD.n521 0.011
R4275 VDD.n1450 VDD.n70 0.011
R4276 VDD.n1446 VDD.n127 0.011
R4277 VDD.n1442 VDD.n184 0.011
R4278 VDD.n1438 VDD.n241 0.011
R4279 VDD.n100 VDD.n88 0.011
R4280 VDD.n99 VDD.n98 0.011
R4281 VDD.n157 VDD.n145 0.011
R4282 VDD.n156 VDD.n155 0.011
R4283 VDD.n214 VDD.n202 0.011
R4284 VDD.n213 VDD.n212 0.011
R4285 VDD.n343 VDD.n339 0.011
R4286 VDD.n335 VDD.n331 0.011
R4287 VDD.n314 VDD.n310 0.011
R4288 VDD.n293 VDD.n289 0.011
R4289 VDD.n260 VDD.n256 0.011
R4290 VDD.n252 VDD.n248 0.011
R4291 VDD.n472 VDD.n463 0.011
R4292 VDD.n456 VDD.n451 0.011
R4293 VDD.n849 VDD.n848 0.011
R4294 VDD.n917 VDD.n908 0.011
R4295 VDD.n1044 VDD.n1043 0.011
R4296 VDD.n1776 VDD.n1764 0.011
R4297 VDD.n1775 VDD.n1774 0.011
R4298 VDD.n1781 VDD.n56 0.011
R4299 VDD.n618 VDD.n617 0.01
R4300 VDD.n681 VDD.n680 0.01
R4301 VDD.n979 VDD.n978 0.01
R4302 VDD.n1117 VDD.n1116 0.009
R4303 VDD.n1107 VDD.n1106 0.009
R4304 VDD.n1172 VDD.n1169 0.009
R4305 VDD.n1723 VDD.n1722 0.009
R4306 VDD.n760 VDD.n759 0.008
R4307 VDD.n1780 VDD.n1452 0.007
R4308 VDD.n1159 VDD.n1158 0.007
R4309 VDD.n1816 VDD.n1815 0.007
R4310 VDD.n1132 VDD.n1129 0.007
R4311 VDD.n728 VDD.n708 0.006
R4312 VDD.n657 VDD.n656 0.005
R4313 VDD.n1189 VDD.n1187 0.005
R4314 VDD.n1655 VDD.n1654 0.005
R4315 VDD.n1661 VDD.n1504 0.005
R4316 VDD.n1316 VDD.n1299 0.004
R4317 VDD.n761 VDD.n760 0.003
R4318 VDD.n1298 VDD.n1297 0.003
R4319 VDD.n1316 VDD.n1315 0.003
R4320 VDD.n1333 VDD.n1332 0.003
R4321 VDD.n1350 VDD.n1349 0.003
R4322 VDD.n1419 VDD.n1418 0.003
R4323 VDD.n1436 VDD.n1435 0.003
R4324 VDD.n386 VDD.n385 0.003
R4325 VDD.n1192 VDD.n1189 0.003
R4326 VDD.n1132 VDD.n1131 0.003
R4327 VDD.n1284 VDD.n1283 0.003
R4328 VDD.n1302 VDD.n1301 0.003
R4329 VDD.n1319 VDD.n1318 0.003
R4330 VDD.n1336 VDD.n1335 0.003
R4331 VDD.n1405 VDD.n1404 0.003
R4332 VDD.n1422 VDD.n1421 0.003
R4333 VDD.n372 VDD.n371 0.003
R4334 VDD.n1267 VDD.n1266 0.003
R4335 VDD.n1628 VDD.n1627 0.002
R4336 VDD.n1603 VDD.n1602 0.002
R4337 VDD.n1578 VDD.n1577 0.002
R4338 VDD.n1553 VDD.n1552 0.002
R4339 VDD.n1528 VDD.n1527 0.002
R4340 VDD.n1478 VDD.n1477 0.002
R4341 VDD.n293 VDD.n0 0.002
R4342 VDD.n471 VDD.n469 0.002
R4343 VDD.n1044 VDD.n1038 0.002
R4344 VDD.n1629 VDD.n1628 0.002
R4345 VDD.n1604 VDD.n1603 0.002
R4346 VDD.n1579 VDD.n1578 0.002
R4347 VDD.n1554 VDD.n1553 0.002
R4348 VDD.n1529 VDD.n1528 0.002
R4349 VDD.n1479 VDD.n1478 0.002
R4350 VDD.n609 VDD.n603 0.002
R4351 VDD.n1654 VDD.n1631 0.002
R4352 VDD.n1504 VDD.n1481 0.002
R4353 VDD.n1160 VDD.n1159 0.001
R4354 VDD.n1625 VDD.n1618 0.001
R4355 VDD.n1600 VDD.n1593 0.001
R4356 VDD.n1575 VDD.n1568 0.001
R4357 VDD.n1550 VDD.n1543 0.001
R4358 VDD.n1525 VDD.n1518 0.001
R4359 VDD.n1475 VDD.n1468 0.001
R4360 VDD.n1108 VDD.n1107 0.001
R4361 VDD.n916 VDD.n914 0.001
R4362 VDD.n1652 VDD.n1651 0.001
R4363 VDD.n1502 VDD.n1501 0.001
R4364 VDD.n728 VDD.n727 0.001
R4365 VDD.n1129 VDD.n1127 0.001
R4366 VDD.n1654 VDD.n1653 0.001
R4367 VDD.n1504 VDD.n1503 0.001
R4368 VDD.n1628 VDD.n1625 0.001
R4369 VDD.n1603 VDD.n1600 0.001
R4370 VDD.n1578 VDD.n1575 0.001
R4371 VDD.n1553 VDD.n1550 0.001
R4372 VDD.n1528 VDD.n1525 0.001
R4373 VDD.n1478 VDD.n1475 0.001
R4374 VDD.n1192 VDD.n1191 0.001
R4375 VDD.n774 VDD.n773 0.001
R4376 VDD.n744 VDD.n743 0.001
R4377 VDD.n749 VDD.n748 0.001
R4378 VDD.n685 VDD.n681 0.001
R4379 VDD.n980 VDD.n979 0.001
R4380 VDD.n17 VDD.n16 0.001
R4381 VDD.n344 VDD.n343 0.001
R4382 VDD.n261 VDD.n260 0.001
R4383 VDD.n727 VDD.n726 0.001
R4384 VDD.n1838 VDD.n1837 0.001
R4385 VDD.n315 VDD.n314 0.001
R4386 VDD.n825 VDD.n824 0.001
R4387 VDD.n826 VDD.n814 0.001
R4388 VDD.n1096 VDD.n1095 0.001
R4389 VDD.n1065 VDD.n1064 0.001
R4390 VDD.n639 VDD.n638 0.001
R4391 VDD.n1001 VDD.n1000 0.001
R4392 VDD.n938 VDD.n937 0.001
R4393 VDD.n1287 VDD.n1286 0.001
R4394 VDD.n1305 VDD.n1304 0.001
R4395 VDD.n1322 VDD.n1321 0.001
R4396 VDD.n1339 VDD.n1338 0.001
R4397 VDD.n1408 VDD.n1407 0.001
R4398 VDD.n1425 VDD.n1424 0.001
R4399 VDD.n375 VDD.n374 0.001
R4400 VDD.n1270 VDD.n1269 0.001
R4401 VDD.n768 VDD.n765 0.001
R4402 VDD.n769 VDD.n768 0.001
R4403 VDD.n472 VDD.n471 0.001
R4404 VDD.n1189 VDD.n1188 0.001
R4405 VDD.n1656 VDD.n1629 0.001
R4406 VDD.n1657 VDD.n1604 0.001
R4407 VDD.n1658 VDD.n1579 0.001
R4408 VDD.n1659 VDD.n1554 0.001
R4409 VDD.n1660 VDD.n1529 0.001
R4410 VDD.n1662 VDD.n1479 0.001
R4411 VDD.n1691 VDD.n1683 0.001
R4412 VDD.n1681 VDD.n1673 0.001
R4413 VDD.n1733 VDD.n1724 0.001
R4414 VDD.n1084 VDD.n1076 0.001
R4415 VDD.n814 VDD.n813 0.001
R4416 VDD.n824 VDD.n823 0.001
R4417 VDD.n446 VDD.n438 0.001
R4418 VDD.n437 VDD.n429 0.001
R4419 VDD.n795 VDD.n787 0.001
R4420 VDD.n804 VDD.n796 0.001
R4421 VDD.n1375 VDD.n1367 0.001
R4422 VDD.n1376 VDD.n1359 0.001
R4423 VDD.n1672 VDD.n1664 0.001
R4424 VDD.n1378 VDD.n1351 0.001
R4425 VDD.n1227 VDD.n421 0.001
R4426 VDD.n420 VDD.n411 0.001
R4427 VDD.n409 VDD.n400 0.001
R4428 VDD.n1263 VDD.n1255 0.001
R4429 VDD.n1400 VDD.n1399 0.001
R4430 VDD.n1095 VDD.n1094 0.001
R4431 VDD.n1038 VDD.n1036 0.001
R4432 VDD.n1129 VDD.n1128 0.001
R4433 VDD.n664 VDD.n663 0.001
R4434 VDD.n762 VDD.n752 0.001
R4435 VDD.n769 VDD.n764 0.001
R4436 VDD.n1193 VDD.n1192 0.001
R4437 VDD.n1173 VDD.n1164 0.001
R4438 VDD.n1133 VDD.n1132 0.001
R4439 VDD.n1118 VDD.n1111 0.001
R4440 VDD.n1109 VDD.n1099 0.001
R4441 VDD.n473 VDD.n472 0.001
R4442 VDD.n918 VDD.n917 0.001
R4443 VDD.n1045 VDD.n1044 0.001
R4444 VDD.n1207 VDD.n1206 0.001
R4445 VDD.n653 VDD.n652 0.001
R4446 VDD.n1720 VDD.n1711 0.001
R4447 VDD.n1118 VDD.n1117 0.001
R4448 VDD.n686 VDD.n685 0.001
R4449 VDD.n774 VDD.n771 0.001
R4450 VDD.n610 VDD.n609 0.001
R4451 VDD.n527 VDD.n526 0.001
R4452 VDD.n457 VDD.n456 0.001
R4453 VDD.n1161 VDD.n1149 0.001
R4454 VDD.n1142 VDD.n1135 0.001
R4455 VDD.n737 VDD.n730 0.001
R4456 VDD.n749 VDD.n746 0.001
R4457 VDD.n744 VDD.n739 0.001
R4458 VDD.n762 VDD.n761 0.001
R4459 VDD.n1216 VDD.n1210 0.001
R4460 VDD.n1178 VDD.n1175 0.001
R4461 VDD.n1147 VDD.n1144 0.001
R4462 VDD.n1192 VDD.n1180 0.001
R4463 VDD.n1132 VDD.n1120 0.001
R4464 VDD.n1206 VDD.n1197 0.001
R4465 VDD.n652 VDD.n643 0.001
R4466 VDD.n1223 VDD.n1217 0.001
R4467 VDD.n671 VDD.n665 0.001
R4468 VDD.n663 VDD.n657 0.001
R4469 VDD.n1653 VDD.n1652 0.001
R4470 VDD.n1503 VDD.n1502 0.001
R4471 VDD.n980 VDD.n972 0.001
R4472 VDD.n618 VDD.n611 0.001
R4473 VDD.n849 VDD.n842 0.001
R4474 VDD.n694 VDD.n687 0.001
R4475 VDD.n535 VDD.n528 0.001
R4476 VDD.n472 VDD.n458 0.001
R4477 VDD.n917 VDD.n903 0.001
R4478 VDD.n1044 VDD.n1032 0.001
R4479 VDD.n1702 VDD.n1701 0.001
R4480 VDD.n1721 VDD.n1720 0.001
R4481 VDD.n782 VDD.n774 0.001
R4482 VDD.n881 VDD.n869 0.001
R4483 VDD.n567 VDD.n555 0.001
R4484 VDD.n917 VDD.n916 0.001
R4485 VDD.n1162 VDD.n1161 0.001
R4486 VDD.n1109 VDD.n1108 0.001
R4487 VDD.n1618 VDD.n1617 0.001
R4488 VDD.n1593 VDD.n1592 0.001
R4489 VDD.n1568 VDD.n1567 0.001
R4490 VDD.n1543 VDD.n1542 0.001
R4491 VDD.n1518 VDD.n1517 0.001
R4492 VDD.n1468 VDD.n1467 0.001
R4493 VDD.n1143 VDD.n1142 0.001
R4494 VDD.n738 VDD.n737 0.001
R4495 VDD.n1174 VDD.n1173 0.001
R4496 VDD.n1110 VDD.n1109 0.001
R4497 VDD.n850 VDD.n849 0.001
R4498 VDD.n763 VDD.n762 0.001
R4499 VDD.n695 VDD.n694 0.001
R4500 VDD.n536 VDD.n535 0.001
R4501 VDD.n619 VDD.n618 0.001
R4502 VDD.n981 VDD.n980 0.001
R4503 VDD.n1179 VDD.n1178 0.001
R4504 VDD.n1148 VDD.n1147 0.001
R4505 VDD.n770 VDD.n769 0.001
R4506 VDD.n1119 VDD.n1118 0.001
R4507 VDD.n750 VDD.n749 0.001
R4508 VDD.n745 VDD.n744 0.001
R4509 VDD.n1161 VDD.n1160 0.001
R4510 VDD.n1173 VDD.n1172 0.001
R4511 VDD.n1288 VDD.n1287 0.001
R4512 VDD.n1306 VDD.n1305 0.001
R4513 VDD.n1323 VDD.n1322 0.001
R4514 VDD.n1340 VDD.n1339 0.001
R4515 VDD.n1409 VDD.n1408 0.001
R4516 VDD.n1426 VDD.n1425 0.001
R4517 VDD.n376 VDD.n375 0.001
R4518 VDD.n1271 VDD.n1270 0.001
R4519 a_11521_19244.n6 a_11521_19244.n5 501.28
R4520 a_11521_19244.t10 a_11521_19244.t19 437.233
R4521 a_11521_19244.t16 a_11521_19244.t7 415.315
R4522 a_11521_19244.t5 a_11521_19244.n3 313.873
R4523 a_11521_19244.n5 a_11521_19244.t15 294.986
R4524 a_11521_19244.n2 a_11521_19244.t18 272.288
R4525 a_11521_19244.n6 a_11521_19244.t17 236.009
R4526 a_11521_19244.n9 a_11521_19244.t10 216.627
R4527 a_11521_19244.n7 a_11521_19244.t16 216.111
R4528 a_11521_19244.n8 a_11521_19244.t11 214.686
R4529 a_11521_19244.t19 a_11521_19244.n8 214.686
R4530 a_11521_19244.n1 a_11521_19244.t9 214.335
R4531 a_11521_19244.t7 a_11521_19244.n1 214.335
R4532 a_11521_19244.n4 a_11521_19244.t12 190.152
R4533 a_11521_19244.n4 a_11521_19244.t5 190.152
R4534 a_11521_19244.n2 a_11521_19244.t14 160.666
R4535 a_11521_19244.n3 a_11521_19244.t13 160.666
R4536 a_11521_19244.n7 a_11521_19244.n6 148.428
R4537 a_11521_19244.n5 a_11521_19244.t8 110.859
R4538 a_11521_19244.n3 a_11521_19244.n2 96.129
R4539 a_11521_19244.n8 a_11521_19244.t4 80.333
R4540 a_11521_19244.n1 a_11521_19244.t6 80.333
R4541 a_11521_19244.t17 a_11521_19244.n4 80.333
R4542 a_11521_19244.t0 a_11521_19244.n11 28.57
R4543 a_11521_19244.n0 a_11521_19244.t1 28.565
R4544 a_11521_19244.n0 a_11521_19244.t2 28.565
R4545 a_11521_19244.n11 a_11521_19244.t3 17.638
R4546 a_11521_19244.n10 a_11521_19244.n9 5.589
R4547 a_11521_19244.n9 a_11521_19244.n7 2.923
R4548 a_11521_19244.n10 a_11521_19244.n0 0.693
R4549 a_11521_19244.n11 a_11521_19244.n10 0.597
R4550 a_15556_20132.n0 a_15556_20132.t8 214.335
R4551 a_15556_20132.t10 a_15556_20132.n0 214.335
R4552 a_15556_20132.n1 a_15556_20132.t10 143.851
R4553 a_15556_20132.n1 a_15556_20132.t7 135.658
R4554 a_15556_20132.n0 a_15556_20132.t9 80.333
R4555 a_15556_20132.n2 a_15556_20132.t5 28.565
R4556 a_15556_20132.n2 a_15556_20132.t6 28.565
R4557 a_15556_20132.n4 a_15556_20132.t4 28.565
R4558 a_15556_20132.n4 a_15556_20132.t1 28.565
R4559 a_15556_20132.t0 a_15556_20132.n7 28.565
R4560 a_15556_20132.n7 a_15556_20132.t2 28.565
R4561 a_15556_20132.n3 a_15556_20132.t3 9.714
R4562 a_15556_20132.n3 a_15556_20132.n2 1.003
R4563 a_15556_20132.n6 a_15556_20132.n5 0.833
R4564 a_15556_20132.n5 a_15556_20132.n4 0.653
R4565 a_15556_20132.n7 a_15556_20132.n6 0.653
R4566 a_15556_20132.n5 a_15556_20132.n3 0.341
R4567 a_15556_20132.n6 a_15556_20132.n1 0.032
R4568 a_5860_19519.n0 a_5860_19519.t3 14.282
R4569 a_5860_19519.t0 a_5860_19519.n0 14.282
R4570 a_5860_19519.n0 a_5860_19519.n12 122.747
R4571 a_5860_19519.n8 a_5860_19519.n10 74.302
R4572 a_5860_19519.n12 a_5860_19519.n8 50.575
R4573 a_5860_19519.n12 a_5860_19519.n11 157.665
R4574 a_5860_19519.n11 a_5860_19519.t7 8.7
R4575 a_5860_19519.n11 a_5860_19519.t1 8.7
R4576 a_5860_19519.n10 a_5860_19519.n9 90.436
R4577 a_5860_19519.n9 a_5860_19519.t4 14.282
R4578 a_5860_19519.n9 a_5860_19519.t5 14.282
R4579 a_5860_19519.n8 a_5860_19519.n7 90.416
R4580 a_5860_19519.n7 a_5860_19519.t6 14.282
R4581 a_5860_19519.n7 a_5860_19519.t2 14.282
R4582 a_5860_19519.n10 a_5860_19519.n1 342.688
R4583 a_5860_19519.n1 a_5860_19519.n6 126.566
R4584 a_5860_19519.n6 a_5860_19519.t13 294.653
R4585 a_5860_19519.n6 a_5860_19519.t9 111.663
R4586 a_5860_19519.n1 a_5860_19519.n5 552.333
R4587 a_5860_19519.n5 a_5860_19519.n4 6.615
R4588 a_5860_19519.n4 a_5860_19519.t15 93.989
R4589 a_5860_19519.n4 a_5860_19519.t8 198.043
R4590 a_5860_19519.n5 a_5860_19519.n3 97.816
R4591 a_5860_19519.n3 a_5860_19519.t14 80.333
R4592 a_5860_19519.n3 a_5860_19519.t11 394.151
R4593 a_5860_19519.t11 a_5860_19519.n2 269.523
R4594 a_5860_19519.n2 a_5860_19519.t12 160.666
R4595 a_5860_19519.n2 a_5860_19519.t10 269.523
R4596 a_5917_18826.n2 a_5917_18826.t6 318.922
R4597 a_5917_18826.n1 a_5917_18826.t4 273.935
R4598 a_5917_18826.n1 a_5917_18826.t7 273.935
R4599 a_5917_18826.n2 a_5917_18826.t5 269.116
R4600 a_5917_18826.n4 a_5917_18826.n0 193.227
R4601 a_5917_18826.t6 a_5917_18826.n1 179.142
R4602 a_5917_18826.n3 a_5917_18826.n2 106.999
R4603 a_5917_18826.t2 a_5917_18826.n4 28.568
R4604 a_5917_18826.n0 a_5917_18826.t0 28.565
R4605 a_5917_18826.n0 a_5917_18826.t1 28.565
R4606 a_5917_18826.n3 a_5917_18826.t3 18.149
R4607 a_5917_18826.n4 a_5917_18826.n3 3.726
R4608 a_21150_9929.n0 a_21150_9929.n13 122.999
R4609 a_21150_9929.t0 a_21150_9929.n0 14.282
R4610 a_21150_9929.n0 a_21150_9929.t3 14.282
R4611 a_21150_9929.n13 a_21150_9929.n11 50.575
R4612 a_21150_9929.n11 a_21150_9929.n9 74.302
R4613 a_21150_9929.n13 a_21150_9929.n12 157.665
R4614 a_21150_9929.n12 a_21150_9929.t4 8.7
R4615 a_21150_9929.n12 a_21150_9929.t1 8.7
R4616 a_21150_9929.n11 a_21150_9929.n10 90.416
R4617 a_21150_9929.n10 a_21150_9929.t2 14.282
R4618 a_21150_9929.n10 a_21150_9929.t5 14.282
R4619 a_21150_9929.n9 a_21150_9929.n8 90.436
R4620 a_21150_9929.n8 a_21150_9929.t7 14.282
R4621 a_21150_9929.n8 a_21150_9929.t6 14.282
R4622 a_21150_9929.n1 a_21150_9929.t15 217.826
R4623 a_21150_9929.n9 a_21150_9929.n1 277.579
R4624 a_21150_9929.n1 a_21150_9929.n6 133.839
R4625 a_21150_9929.t15 a_21150_9929.t14 437.233
R4626 a_21150_9929.t14 a_21150_9929.n7 214.686
R4627 a_21150_9929.n7 a_21150_9929.t19 80.333
R4628 a_21150_9929.n7 a_21150_9929.t10 214.686
R4629 a_21150_9929.n6 a_21150_9929.n2 563.136
R4630 a_21150_9929.n6 a_21150_9929.t11 178.973
R4631 a_21150_9929.t11 a_21150_9929.n5 80.333
R4632 a_21150_9929.n5 a_21150_9929.t12 190.152
R4633 a_21150_9929.n5 a_21150_9929.t16 190.152
R4634 a_21150_9929.t16 a_21150_9929.n4 313.873
R4635 a_21150_9929.n4 a_21150_9929.t9 160.666
R4636 a_21150_9929.n4 a_21150_9929.n3 96.129
R4637 a_21150_9929.n3 a_21150_9929.t18 160.666
R4638 a_21150_9929.n3 a_21150_9929.t8 272.288
R4639 a_21150_9929.n2 a_21150_9929.t13 294.986
R4640 a_21150_9929.n2 a_21150_9929.t17 110.859
R4641 a_31893_6205.t0 a_31893_6205.n7 16.058
R4642 a_31893_6205.n7 a_31893_6205.n5 0.575
R4643 a_31893_6205.n5 a_31893_6205.n9 0.2
R4644 a_31893_6205.n9 a_31893_6205.t5 16.058
R4645 a_31893_6205.n9 a_31893_6205.n8 0.999
R4646 a_31893_6205.n8 a_31893_6205.t4 14.282
R4647 a_31893_6205.n8 a_31893_6205.t3 14.282
R4648 a_31893_6205.n7 a_31893_6205.n6 0.999
R4649 a_31893_6205.n6 a_31893_6205.t6 14.282
R4650 a_31893_6205.n6 a_31893_6205.t2 14.282
R4651 a_31893_6205.n5 a_31893_6205.n3 0.227
R4652 a_31893_6205.n3 a_31893_6205.n4 1.511
R4653 a_31893_6205.n4 a_31893_6205.t1 14.282
R4654 a_31893_6205.n4 a_31893_6205.t10 14.282
R4655 a_31893_6205.n3 a_31893_6205.n0 0.669
R4656 a_31893_6205.n0 a_31893_6205.n1 0.001
R4657 a_31893_6205.n0 a_31893_6205.n2 267.767
R4658 a_31893_6205.n2 a_31893_6205.t7 14.282
R4659 a_31893_6205.n2 a_31893_6205.t8 14.282
R4660 a_31893_6205.n1 a_31893_6205.t11 14.282
R4661 a_31893_6205.n1 a_31893_6205.t9 14.282
R4662 a_12900_12829.t8 a_12900_12829.n2 404.877
R4663 a_12900_12829.n1 a_12900_12829.t6 210.902
R4664 a_12900_12829.n3 a_12900_12829.t8 136.943
R4665 a_12900_12829.n2 a_12900_12829.n1 107.801
R4666 a_12900_12829.n1 a_12900_12829.t5 80.333
R4667 a_12900_12829.n2 a_12900_12829.t7 80.333
R4668 a_12900_12829.n0 a_12900_12829.t1 17.4
R4669 a_12900_12829.n0 a_12900_12829.t0 17.4
R4670 a_12900_12829.n4 a_12900_12829.t3 15.032
R4671 a_12900_12829.t2 a_12900_12829.n5 14.282
R4672 a_12900_12829.n5 a_12900_12829.t4 14.282
R4673 a_12900_12829.n5 a_12900_12829.n4 1.65
R4674 a_12900_12829.n3 a_12900_12829.n0 0.672
R4675 a_12900_12829.n4 a_12900_12829.n3 0.665
R4676 a_13164_12246.t4 a_13164_12246.t7 800.071
R4677 a_13164_12246.n3 a_13164_12246.n2 672.951
R4678 a_13164_12246.n1 a_13164_12246.t6 285.109
R4679 a_13164_12246.n2 a_13164_12246.t4 193.602
R4680 a_13164_12246.n1 a_13164_12246.t5 160.666
R4681 a_13164_12246.n2 a_13164_12246.n1 91.507
R4682 a_13164_12246.n0 a_13164_12246.t0 28.57
R4683 a_13164_12246.n4 a_13164_12246.t1 28.565
R4684 a_13164_12246.t2 a_13164_12246.n4 28.565
R4685 a_13164_12246.n0 a_13164_12246.t3 17.638
R4686 a_13164_12246.n4 a_13164_12246.n3 0.69
R4687 a_13164_12246.n3 a_13164_12246.n0 0.6
R4688 a_17356_9635.n0 a_17356_9635.t8 214.335
R4689 a_17356_9635.t10 a_17356_9635.n0 214.335
R4690 a_17356_9635.n1 a_17356_9635.t10 143.851
R4691 a_17356_9635.n1 a_17356_9635.t7 135.658
R4692 a_17356_9635.n0 a_17356_9635.t9 80.333
R4693 a_17356_9635.n2 a_17356_9635.t5 28.565
R4694 a_17356_9635.n2 a_17356_9635.t6 28.565
R4695 a_17356_9635.n4 a_17356_9635.t4 28.565
R4696 a_17356_9635.n4 a_17356_9635.t2 28.565
R4697 a_17356_9635.n7 a_17356_9635.t3 28.565
R4698 a_17356_9635.t0 a_17356_9635.n7 28.565
R4699 a_17356_9635.n6 a_17356_9635.t1 9.714
R4700 a_17356_9635.n7 a_17356_9635.n6 1.003
R4701 a_17356_9635.n5 a_17356_9635.n3 0.833
R4702 a_17356_9635.n3 a_17356_9635.n2 0.653
R4703 a_17356_9635.n5 a_17356_9635.n4 0.653
R4704 a_17356_9635.n6 a_17356_9635.n5 0.341
R4705 a_17356_9635.n3 a_17356_9635.n1 0.032
R4706 VSS.n380 VSS.t389 20.872
R4707 VSS.n383 VSS.t423 20.872
R4708 VSS.n123 VSS.t103 20.872
R4709 VSS.n48 VSS.t140 20.872
R4710 VSS.n379 VSS.t335 20.83
R4711 VSS.n382 VSS.t218 20.83
R4712 VSS.n122 VSS.t95 20.83
R4713 VSS.n47 VSS.t374 20.83
R4714 VSS.n426 VSS.t260 20.763
R4715 VSS.n385 VSS.t124 20.763
R4716 VSS.n226 VSS.t386 20.763
R4717 VSS.n211 VSS.t293 20.763
R4718 VSS.n388 VSS.t66 20.763
R4719 VSS.n421 VSS.t281 20.763
R4720 VSS.n223 VSS.t242 20.763
R4721 VSS.n347 VSS.t10 20.763
R4722 VSS.n429 VSS.t272 20.763
R4723 VSS.n400 VSS.t104 20.763
R4724 VSS.n180 VSS.t177 20.763
R4725 VSS.n322 VSS.t301 20.763
R4726 VSS.n233 VSS.t90 20.763
R4727 VSS.n317 VSS.t432 20.763
R4728 VSS.n461 VSS.t247 20.763
R4729 VSS.n464 VSS.t26 20.763
R4730 VSS.n459 VSS.t365 20.763
R4731 VSS.n457 VSS.t353 20.763
R4732 VSS.n472 VSS.t163 20.763
R4733 VSS.n476 VSS.t111 20.763
R4734 VSS.n480 VSS.t145 20.763
R4735 VSS.n454 VSS.t155 20.763
R4736 VSS.n161 VSS.t419 20.763
R4737 VSS.n358 VSS.t210 20.763
R4738 VSS.n30 VSS.t277 20.763
R4739 VSS.n152 VSS.t428 20.763
R4740 VSS.n140 VSS.t39 20.763
R4741 VSS.n34 VSS.t361 20.763
R4742 VSS.n175 VSS.t340 20.763
R4743 VSS.n53 VSS.t17 20.763
R4744 VSS.n147 VSS.t435 20.763
R4745 VSS.n96 VSS.t204 20.763
R4746 VSS.n144 VSS.t315 20.763
R4747 VSS.n93 VSS.t164 20.763
R4748 VSS.n90 VSS.t379 20.763
R4749 VSS.n131 VSS.t371 20.763
R4750 VSS.n455 VSS.t330 20.677
R4751 VSS.n466 VSS.t334 20.677
R4752 VSS.n474 VSS.t336 20.677
R4753 VSS.n478 VSS.t328 20.677
R4754 VSS.n482 VSS.t331 20.677
R4755 VSS.n462 VSS.t329 20.676
R4756 VSS.n468 VSS.t333 20.676
R4757 VSS.n470 VSS.t327 20.676
R4758 VSS.n54 VSS.t120 20.614
R4759 VSS.n427 VSS.t311 20.606
R4760 VSS.n386 VSS.t397 20.606
R4761 VSS.n227 VSS.t171 20.606
R4762 VSS.n212 VSS.t258 20.606
R4763 VSS.n389 VSS.t254 20.606
R4764 VSS.n422 VSS.t305 20.606
R4765 VSS.n224 VSS.t89 20.606
R4766 VSS.n348 VSS.t319 20.606
R4767 VSS.n430 VSS.t197 20.606
R4768 VSS.n401 VSS.t346 20.606
R4769 VSS.n181 VSS.t341 20.606
R4770 VSS.n323 VSS.t268 20.606
R4771 VSS.n234 VSS.t203 20.606
R4772 VSS.n318 VSS.t324 20.606
R4773 VSS.n162 VSS.t403 20.606
R4774 VSS.n359 VSS.t181 20.606
R4775 VSS.n31 VSS.t135 20.606
R4776 VSS.n153 VSS.t3 20.606
R4777 VSS.n141 VSS.t58 20.606
R4778 VSS.n35 VSS.t150 20.606
R4779 VSS.n176 VSS.t271 20.606
R4780 VSS.n148 VSS.t38 20.606
R4781 VSS.n97 VSS.t410 20.606
R4782 VSS.n145 VSS.t170 20.606
R4783 VSS.n94 VSS.t382 20.606
R4784 VSS.n91 VSS.t118 20.606
R4785 VSS.n132 VSS.t264 20.606
R4786 VSS.n236 VSS.t373 20.5
R4787 VSS.n243 VSS.t106 20.5
R4788 VSS.n241 VSS.t266 20.5
R4789 VSS.n239 VSS.t350 20.5
R4790 VSS.n237 VSS.t112 20.224
R4791 VSS.n307 VSS.t234 20.223
R4792 VSS.n307 VSS.t437 20.223
R4793 VSS.n307 VSS.t377 20.223
R4794 VSS.n404 VSS.t322 18.354
R4795 VSS.n39 VSS.t384 18.354
R4796 VSS.n73 VSS.t229 18.354
R4797 VSS.n335 VSS.t174 18.185
R4798 VSS.n437 VSS.t390 18.185
R4799 VSS.n206 VSS.t47 18.185
R4800 VSS.n415 VSS.t398 18.185
R4801 VSS.n183 VSS.t214 18.185
R4802 VSS.n182 VSS.t34 18.185
R4803 VSS.n444 VSS.t240 18.185
R4804 VSS.n409 VSS.t33 18.185
R4805 VSS.n193 VSS.t71 18.185
R4806 VSS.n433 VSS.t207 18.185
R4807 VSS.n199 VSS.t96 18.185
R4808 VSS.n442 VSS.t304 18.185
R4809 VSS.n187 VSS.t93 18.185
R4810 VSS.n394 VSS.t30 18.185
R4811 VSS.n230 VSS.t351 18.185
R4812 VSS.n231 VSS.t233 18.185
R4813 VSS.n391 VSS.t134 18.185
R4814 VSS.n229 VSS.t156 18.185
R4815 VSS.n334 VSS.t84 18.185
R4816 VSS.n333 VSS.t219 18.185
R4817 VSS.n405 VSS.t393 18.185
R4818 VSS.n493 VSS.t132 18.185
R4819 VSS.n13 VSS.t61 18.185
R4820 VSS.n367 VSS.t80 18.185
R4821 VSS.n20 VSS.t211 18.185
R4822 VSS.n361 VSS.t8 18.185
R4823 VSS.n5 VSS.t401 18.185
R4824 VSS.n373 VSS.t357 18.185
R4825 VSS.n178 VSS.t303 18.185
R4826 VSS.n350 VSS.t55 18.185
R4827 VSS.n165 VSS.t148 18.185
R4828 VSS.n164 VSS.t25 18.185
R4829 VSS.n166 VSS.t137 18.185
R4830 VSS.n62 VSS.t278 18.185
R4831 VSS.n63 VSS.t230 18.185
R4832 VSS.n64 VSS.t422 18.185
R4833 VSS.n65 VSS.t31 18.185
R4834 VSS.n116 VSS.t113 18.185
R4835 VSS.n112 VSS.t221 18.185
R4836 VSS.n105 VSS.t308 18.185
R4837 VSS.n75 VSS.t196 18.185
R4838 VSS.n99 VSS.t391 18.185
R4839 VSS.n67 VSS.t123 18.185
R4840 VSS.n1 VSS.t105 18.185
R4841 VSS.n313 VSS.t27 18.178
R4842 VSS.n244 VSS.t368 18.178
R4843 VSS.n311 VSS.t169 18.178
R4844 VSS.n452 VSS.t168 18.178
R4845 VSS.n451 VSS.t323 18.178
R4846 VSS.n245 VSS.t217 18.178
R4847 VSS.n312 VSS.t82 18.178
R4848 VSS.n308 VSS.t228 18.178
R4849 VSS.n246 VSS.t421 18.178
R4850 VSS.n450 VSS.t363 18.178
R4851 VSS.n309 VSS.t413 18.178
R4852 VSS.n449 VSS.t44 18.178
R4853 VSS.n247 VSS.t235 18.178
R4854 VSS.n395 VSS.t187 18.178
R4855 VSS.n310 VSS.t236 18.178
R4856 VSS.n44 VSS.t76 18.178
R4857 VSS.n55 VSS.t359 18.178
R4858 VSS.n396 VSS.t356 18.176
R4859 VSS.n155 VSS.t283 18.176
R4860 VSS.n134 VSS.t376 18.176
R4861 VSS.n390 VSS.t279 18.089
R4862 VSS.n214 VSS.t45 17.959
R4863 VSS.n332 VSS.t342 17.959
R4864 VSS.n38 VSS.t180 17.959
R4865 VSS.n158 VSS.t100 17.959
R4866 VSS.n59 VSS.t176 17.959
R4867 VSS.n61 VSS.t0 17.959
R4868 VSS.n221 VSS.t188 17.929
R4869 VSS.n500 VSS.t395 17.929
R4870 VSS.n327 VSS.t213 17.929
R4871 VSS.n496 VSS.t153 17.929
R4872 VSS.n320 VSS.t251 17.929
R4873 VSS.n393 VSS.t392 17.929
R4874 VSS.n171 VSS.t173 17.929
R4875 VSS.n168 VSS.t28 17.929
R4876 VSS.n41 VSS.t49 17.929
R4877 VSS.n129 VSS.t299 17.929
R4878 VSS.n127 VSS.t199 17.929
R4879 VSS.n125 VSS.t108 17.929
R4880 VSS.n398 VSS.t42 17.925
R4881 VSS.n315 VSS.t253 17.925
R4882 VSS.n343 VSS.t114 17.925
R4883 VSS.n424 VSS.t388 17.925
R4884 VSS.n487 VSS.t183 17.925
R4885 VSS.n338 VSS.t83 17.925
R4886 VSS.n355 VSS.t59 17.925
R4887 VSS.n352 VSS.t7 17.925
R4888 VSS.n150 VSS.t396 17.925
R4889 VSS.n137 VSS.t60 17.925
R4890 VSS.n82 VSS.t433 17.925
R4891 VSS.n84 VSS.t208 17.925
R4892 VSS.n407 VSS.t191 17.888
R4893 VSS.n403 VSS.t394 17.884
R4894 VSS.n301 VSS.t288 17.508
R4895 VSS.n250 VSS.t286 17.508
R4896 VSS.n257 VSS.t289 17.508
R4897 VSS.n280 VSS.t291 17.508
R4898 VSS.n286 VSS.t285 17.508
R4899 VSS.n293 VSS.t290 17.508
R4900 VSS.n273 VSS.t287 17.508
R4901 VSS.n266 VSS.t284 17.508
R4902 VSS.n302 VSS.t239 17.504
R4903 VSS.n251 VSS.t78 17.504
R4904 VSS.n258 VSS.t249 17.504
R4905 VSS.n281 VSS.t190 17.504
R4906 VSS.n287 VSS.t194 17.504
R4907 VSS.n294 VSS.t126 17.504
R4908 VSS.n274 VSS.t130 17.504
R4909 VSS.n267 VSS.t343 17.504
R4910 VSS.n397 VSS.t81 17.4
R4911 VSS.n397 VSS.t43 17.4
R4912 VSS.n314 VSS.t193 17.4
R4913 VSS.n314 VSS.t54 17.4
R4914 VSS.n220 VSS.t205 17.4
R4915 VSS.n220 VSS.t40 17.4
R4916 VSS.n499 VSS.t162 17.4
R4917 VSS.n499 VSS.t122 17.4
R4918 VSS.n342 VSS.t16 17.4
R4919 VSS.n342 VSS.t115 17.4
R4920 VSS.n423 VSS.t138 17.4
R4921 VSS.n423 VSS.t200 17.4
R4922 VSS.n326 VSS.t223 17.4
R4923 VSS.n326 VSS.t201 17.4
R4924 VSS.n486 VSS.t50 17.4
R4925 VSS.n486 VSS.t152 17.4
R4926 VSS.n495 VSS.t261 17.4
R4927 VSS.n495 VSS.t36 17.4
R4928 VSS.n337 VSS.t74 17.4
R4929 VSS.n337 VSS.t189 17.4
R4930 VSS.n319 VSS.t139 17.4
R4931 VSS.n319 VSS.t21 17.4
R4932 VSS.n213 VSS.t87 17.4
R4933 VSS.n213 VSS.t110 17.4
R4934 VSS.n406 VSS.t402 17.4
R4935 VSS.n406 VSS.t72 17.4
R4936 VSS.n402 VSS.t46 17.4
R4937 VSS.n402 VSS.t399 17.4
R4938 VSS.n331 VSS.t128 17.4
R4939 VSS.n331 VSS.t88 17.4
R4940 VSS.n392 VSS.t98 17.4
R4941 VSS.n392 VSS.t404 17.4
R4942 VSS.n354 VSS.t18 17.4
R4943 VSS.n354 VSS.t400 17.4
R4944 VSS.n351 VSS.t41 17.4
R4945 VSS.n351 VSS.t75 17.4
R4946 VSS.n37 VSS.t13 17.4
R4947 VSS.n37 VSS.t157 17.4
R4948 VSS.n170 VSS.t20 17.4
R4949 VSS.n170 VSS.t11 17.4
R4950 VSS.n167 VSS.t65 17.4
R4951 VSS.n167 VSS.t19 17.4
R4952 VSS.n40 VSS.t227 17.4
R4953 VSS.n40 VSS.t407 17.4
R4954 VSS.n157 VSS.t297 17.4
R4955 VSS.n157 VSS.t12 17.4
R4956 VSS.n149 VSS.t97 17.4
R4957 VSS.n149 VSS.t295 17.4
R4958 VSS.n136 VSS.t252 17.4
R4959 VSS.n136 VSS.t24 17.4
R4960 VSS.n58 VSS.t185 17.4
R4961 VSS.n58 VSS.t420 17.4
R4962 VSS.n128 VSS.t338 17.4
R4963 VSS.n128 VSS.t52 17.4
R4964 VSS.n126 VSS.t79 17.4
R4965 VSS.n126 VSS.t312 17.4
R4966 VSS.n124 VSS.t69 17.4
R4967 VSS.n124 VSS.t222 17.4
R4968 VSS.n60 VSS.t416 17.4
R4969 VSS.n60 VSS.t216 17.4
R4970 VSS.n81 VSS.t317 17.4
R4971 VSS.n81 VSS.t5 17.4
R4972 VSS.n83 VSS.t215 17.4
R4973 VSS.n83 VSS.t57 17.4
R4974 VSS.n404 VSS.t337 9.906
R4975 VSS.n39 VSS.t172 9.906
R4976 VSS.n73 VSS.t339 9.906
R4977 VSS.n437 VSS.t125 9.568
R4978 VSS.n206 VSS.t385 9.568
R4979 VSS.n415 VSS.t310 9.568
R4980 VSS.n183 VSS.t257 9.568
R4981 VSS.n182 VSS.t256 9.568
R4982 VSS.n444 VSS.t309 9.568
R4983 VSS.n409 VSS.t70 9.568
R4984 VSS.n193 VSS.t243 9.568
R4985 VSS.n433 VSS.t306 9.568
R4986 VSS.n199 VSS.t320 9.568
R4987 VSS.n442 VSS.t307 9.568
R4988 VSS.n187 VSS.t321 9.568
R4989 VSS.n13 VSS.t418 9.568
R4990 VSS.n367 VSS.t144 9.568
R4991 VSS.n20 VSS.t86 9.568
R4992 VSS.n361 VSS.t151 9.568
R4993 VSS.n5 VSS.t143 9.568
R4994 VSS.n373 VSS.t149 9.568
R4995 VSS.n112 VSS.t314 9.568
R4996 VSS.n105 VSS.t318 9.568
R4997 VSS.n75 VSS.t434 9.568
R4998 VSS.n99 VSS.t411 9.568
R4999 VSS.n67 VSS.t383 9.568
R5000 VSS.n1 VSS.t412 9.568
R5001 VSS.n335 VSS.t326 9.487
R5002 VSS.n394 VSS.t273 9.487
R5003 VSS.n230 VSS.t179 9.487
R5004 VSS.n231 VSS.t269 9.487
R5005 VSS.n391 VSS.t344 9.487
R5006 VSS.n229 VSS.t270 9.487
R5007 VSS.n334 VSS.t91 9.487
R5008 VSS.n333 VSS.t325 9.487
R5009 VSS.n405 VSS.t414 9.487
R5010 VSS.n493 VSS.t415 9.487
R5011 VSS.n178 VSS.t141 9.487
R5012 VSS.n350 VSS.t142 9.487
R5013 VSS.n165 VSS.t380 9.487
R5014 VSS.n164 VSS.t263 9.487
R5015 VSS.n166 VSS.t262 9.487
R5016 VSS.n62 VSS.t35 9.487
R5017 VSS.n63 VSS.t275 9.487
R5018 VSS.n64 VSS.t248 9.487
R5019 VSS.n65 VSS.t119 9.487
R5020 VSS.n116 VSS.t121 9.487
R5021 VSS.n390 VSS.t345 9.46
R5022 VSS.n313 VSS.t430 9.319
R5023 VSS.n244 VSS.t186 9.319
R5024 VSS.n311 VSS.t64 9.319
R5025 VSS.n452 VSS.t425 9.319
R5026 VSS.n451 VSS.t354 9.319
R5027 VSS.n245 VSS.t238 9.319
R5028 VSS.n312 VSS.t431 9.319
R5029 VSS.n308 VSS.t282 9.319
R5030 VSS.n246 VSS.t438 9.319
R5031 VSS.n450 VSS.t370 9.319
R5032 VSS.n309 VSS.t367 9.319
R5033 VSS.n449 VSS.t355 9.319
R5034 VSS.n247 VSS.t378 9.319
R5035 VSS.n395 VSS.t427 9.319
R5036 VSS.n310 VSS.t409 9.319
R5037 VSS.n44 VSS.t116 9.319
R5038 VSS.n55 VSS.t364 9.319
R5039 VSS.n396 VSS.t302 9.317
R5040 VSS.n155 VSS.t358 9.317
R5041 VSS.n134 VSS.t426 9.317
R5042 VSS.n302 VSS.t131 8.702
R5043 VSS.n251 VSS.t408 8.702
R5044 VSS.n258 VSS.t99 8.702
R5045 VSS.n281 VSS.t4 8.702
R5046 VSS.n287 VSS.t166 8.702
R5047 VSS.n294 VSS.t198 8.702
R5048 VSS.n274 VSS.t298 8.702
R5049 VSS.n267 VSS.t192 8.702
R5050 VSS.n301 VSS.t102 8.702
R5051 VSS.n250 VSS.t244 8.702
R5052 VSS.n257 VSS.t1 8.702
R5053 VSS.n280 VSS.t63 8.702
R5054 VSS.n286 VSS.t439 8.702
R5055 VSS.n293 VSS.t316 8.702
R5056 VSS.n273 VSS.t117 8.702
R5057 VSS.n266 VSS.t175 8.702
R5058 VSS.n235 VSS.t62 8.7
R5059 VSS.n235 VSS.t372 8.7
R5060 VSS.n425 VSS.t159 8.7
R5061 VSS.n425 VSS.t259 8.7
R5062 VSS.n384 VSS.t32 8.7
R5063 VSS.n384 VSS.t165 8.7
R5064 VSS.n225 VSS.t226 8.7
R5065 VSS.n225 VSS.t387 8.7
R5066 VSS.n210 VSS.t250 8.7
R5067 VSS.n210 VSS.t294 8.7
R5068 VSS.n242 VSS.t48 8.7
R5069 VSS.n242 VSS.t107 8.7
R5070 VSS.n387 VSS.t23 8.7
R5071 VSS.n387 VSS.t195 8.7
R5072 VSS.n420 VSS.t206 8.7
R5073 VSS.n420 VSS.t280 8.7
R5074 VSS.n240 VSS.t184 8.7
R5075 VSS.n240 VSS.t267 8.7
R5076 VSS.n222 VSS.t224 8.7
R5077 VSS.n222 VSS.t241 8.7
R5078 VSS.n346 VSS.t77 8.7
R5079 VSS.n346 VSS.t53 8.7
R5080 VSS.n238 VSS.t56 8.7
R5081 VSS.n238 VSS.t349 8.7
R5082 VSS.n428 VSS.t274 8.7
R5083 VSS.n428 VSS.t360 8.7
R5084 VSS.n399 VSS.t94 8.7
R5085 VSS.n399 VSS.t160 8.7
R5086 VSS.n179 VSS.t178 8.7
R5087 VSS.n179 VSS.t255 8.7
R5088 VSS.n321 VSS.t300 8.7
R5089 VSS.n321 VSS.t161 8.7
R5090 VSS.n378 VSS.t51 8.7
R5091 VSS.n378 VSS.t332 8.7
R5092 VSS.n381 VSS.t237 8.7
R5093 VSS.n381 VSS.t136 8.7
R5094 VSS.n232 VSS.t6 8.7
R5095 VSS.n232 VSS.t92 8.7
R5096 VSS.n316 VSS.t232 8.7
R5097 VSS.n316 VSS.t429 8.7
R5098 VSS.n460 VSS.t246 8.7
R5099 VSS.n460 VSS.t347 8.7
R5100 VSS.n463 VSS.t2 8.7
R5101 VSS.n463 VSS.t109 8.7
R5102 VSS.n458 VSS.t366 8.7
R5103 VSS.n458 VSS.t212 8.7
R5104 VSS.n456 VSS.t352 8.7
R5105 VSS.n456 VSS.t68 8.7
R5106 VSS.n471 VSS.t167 8.7
R5107 VSS.n471 VSS.t225 8.7
R5108 VSS.n475 VSS.t67 8.7
R5109 VSS.n475 VSS.t73 8.7
R5110 VSS.n479 VSS.t146 8.7
R5111 VSS.n479 VSS.t154 8.7
R5112 VSS.n453 VSS.t231 8.7
R5113 VSS.n453 VSS.t182 8.7
R5114 VSS.n160 VSS.t296 8.7
R5115 VSS.n160 VSS.t417 8.7
R5116 VSS.n357 VSS.t405 8.7
R5117 VSS.n357 VSS.t209 8.7
R5118 VSS.n29 VSS.t276 8.7
R5119 VSS.n29 VSS.t406 8.7
R5120 VSS.n151 VSS.t424 8.7
R5121 VSS.n151 VSS.t29 8.7
R5122 VSS.n139 VSS.t133 8.7
R5123 VSS.n139 VSS.t85 8.7
R5124 VSS.n33 VSS.t129 8.7
R5125 VSS.n33 VSS.t362 8.7
R5126 VSS.n174 VSS.t220 8.7
R5127 VSS.n174 VSS.t348 8.7
R5128 VSS.n52 VSS.t101 8.7
R5129 VSS.n52 VSS.t127 8.7
R5130 VSS.n121 VSS.t158 8.7
R5131 VSS.n121 VSS.t147 8.7
R5132 VSS.n46 VSS.t202 8.7
R5133 VSS.n46 VSS.t375 8.7
R5134 VSS.n146 VSS.t265 8.7
R5135 VSS.n146 VSS.t436 8.7
R5136 VSS.n95 VSS.t245 8.7
R5137 VSS.n95 VSS.t37 8.7
R5138 VSS.n143 VSS.t292 8.7
R5139 VSS.n143 VSS.t313 8.7
R5140 VSS.n92 VSS.t9 8.7
R5141 VSS.n92 VSS.t15 8.7
R5142 VSS.n89 VSS.t381 8.7
R5143 VSS.n89 VSS.t14 8.7
R5144 VSS.n130 VSS.t369 8.7
R5145 VSS.n130 VSS.t22 8.7
R5146 VSS.n303 VSS.n301 2.025
R5147 VSS.n252 VSS.n250 2.025
R5148 VSS.n259 VSS.n257 2.025
R5149 VSS.n282 VSS.n280 2.025
R5150 VSS.n288 VSS.n286 2.025
R5151 VSS.n295 VSS.n293 2.025
R5152 VSS.n275 VSS.n273 2.025
R5153 VSS.n268 VSS.n266 2.025
R5154 VSS.n303 VSS.n302 1.953
R5155 VSS.n252 VSS.n251 1.953
R5156 VSS.n259 VSS.n258 1.953
R5157 VSS.n282 VSS.n281 1.953
R5158 VSS.n288 VSS.n287 1.953
R5159 VSS.n295 VSS.n294 1.953
R5160 VSS.n275 VSS.n274 1.953
R5161 VSS.n268 VSS.n267 1.953
R5162 VSS.n426 VSS.n425 0.948
R5163 VSS.n385 VSS.n384 0.948
R5164 VSS.n226 VSS.n225 0.948
R5165 VSS.n211 VSS.n210 0.948
R5166 VSS.n388 VSS.n387 0.948
R5167 VSS.n421 VSS.n420 0.948
R5168 VSS.n223 VSS.n222 0.948
R5169 VSS.n347 VSS.n346 0.948
R5170 VSS.n429 VSS.n428 0.948
R5171 VSS.n400 VSS.n399 0.948
R5172 VSS.n180 VSS.n179 0.948
R5173 VSS.n322 VSS.n321 0.948
R5174 VSS.n233 VSS.n232 0.948
R5175 VSS.n317 VSS.n316 0.948
R5176 VSS.n461 VSS.n460 0.948
R5177 VSS.n464 VSS.n463 0.948
R5178 VSS.n459 VSS.n458 0.948
R5179 VSS.n457 VSS.n456 0.948
R5180 VSS.n472 VSS.n471 0.948
R5181 VSS.n476 VSS.n475 0.948
R5182 VSS.n480 VSS.n479 0.948
R5183 VSS.n454 VSS.n453 0.948
R5184 VSS.n161 VSS.n160 0.948
R5185 VSS.n358 VSS.n357 0.948
R5186 VSS.n30 VSS.n29 0.948
R5187 VSS.n152 VSS.n151 0.948
R5188 VSS.n140 VSS.n139 0.948
R5189 VSS.n34 VSS.n33 0.948
R5190 VSS.n175 VSS.n174 0.948
R5191 VSS.n53 VSS.n52 0.948
R5192 VSS.n147 VSS.n146 0.948
R5193 VSS.n96 VSS.n95 0.948
R5194 VSS.n144 VSS.n143 0.948
R5195 VSS.n93 VSS.n92 0.948
R5196 VSS.n90 VSS.n89 0.948
R5197 VSS.n131 VSS.n130 0.948
R5198 VSS.n236 VSS.n235 0.889
R5199 VSS.n243 VSS.n242 0.889
R5200 VSS.n241 VSS.n240 0.889
R5201 VSS.n239 VSS.n238 0.889
R5202 VSS.n379 VSS.n378 0.889
R5203 VSS.n382 VSS.n381 0.889
R5204 VSS.n122 VSS.n121 0.889
R5205 VSS.n47 VSS.n46 0.889
R5206 VSS.n332 VSS.n331 0.795
R5207 VSS.n158 VSS.n157 0.795
R5208 VSS.n59 VSS.n58 0.795
R5209 VSS.n214 VSS.n213 0.791
R5210 VSS.n38 VSS.n37 0.791
R5211 VSS.n61 VSS.n60 0.791
R5212 VSS.n398 VSS.n397 0.72
R5213 VSS.n315 VSS.n314 0.72
R5214 VSS.n221 VSS.n220 0.72
R5215 VSS.n500 VSS.n499 0.72
R5216 VSS.n343 VSS.n342 0.72
R5217 VSS.n424 VSS.n423 0.72
R5218 VSS.n327 VSS.n326 0.72
R5219 VSS.n487 VSS.n486 0.72
R5220 VSS.n496 VSS.n495 0.72
R5221 VSS.n338 VSS.n337 0.72
R5222 VSS.n320 VSS.n319 0.72
R5223 VSS.n407 VSS.n406 0.72
R5224 VSS.n403 VSS.n402 0.72
R5225 VSS.n393 VSS.n392 0.72
R5226 VSS.n355 VSS.n354 0.72
R5227 VSS.n352 VSS.n351 0.72
R5228 VSS.n171 VSS.n170 0.72
R5229 VSS.n168 VSS.n167 0.72
R5230 VSS.n41 VSS.n40 0.72
R5231 VSS.n150 VSS.n149 0.72
R5232 VSS.n137 VSS.n136 0.72
R5233 VSS.n129 VSS.n128 0.72
R5234 VSS.n127 VSS.n126 0.72
R5235 VSS.n125 VSS.n124 0.72
R5236 VSS.n82 VSS.n81 0.72
R5237 VSS.n84 VSS.n83 0.72
R5238 VSS.n380 VSS.n379 0.449
R5239 VSS.n383 VSS.n382 0.449
R5240 VSS.n123 VSS.n122 0.449
R5241 VSS.n48 VSS.n47 0.449
R5242 VSS.n503 VSS.n396 0.311
R5243 VSS.n325 VSS.n313 0.309
R5244 VSS.n306 VSS.n244 0.309
R5245 VSS.n325 VSS.n311 0.309
R5246 VSS.n484 VSS.n452 0.309
R5247 VSS.n484 VSS.n451 0.309
R5248 VSS.n306 VSS.n245 0.309
R5249 VSS.n325 VSS.n312 0.309
R5250 VSS.n325 VSS.n308 0.309
R5251 VSS.n306 VSS.n246 0.309
R5252 VSS.n484 VSS.n450 0.309
R5253 VSS.n484 VSS.n449 0.309
R5254 VSS.n306 VSS.n247 0.309
R5255 VSS.n503 VSS.n395 0.309
R5256 VSS.n325 VSS.n310 0.309
R5257 VSS.n156 VSS.n155 0.266
R5258 VSS.n135 VSS.n134 0.266
R5259 VSS.n45 VSS.n44 0.264
R5260 VSS.n56 VSS.n55 0.264
R5261 VSS.n325 VSS.n309 0.259
R5262 VSS.n503 VSS.n390 0.239
R5263 VSS.n494 VSS.n404 0.229
R5264 VSS VSS.n39 0.229
R5265 VSS VSS.n73 0.229
R5266 VSS.n462 VSS.n461 0.198
R5267 VSS.n477 VSS.n476 0.198
R5268 VSS.n481 VSS.n480 0.198
R5269 VSS.n465 VSS.n464 0.198
R5270 VSS.n473 VSS.n472 0.198
R5271 VSS.n467 VSS.n459 0.197
R5272 VSS.n469 VSS.n457 0.197
R5273 VSS.n455 VSS.n454 0.197
R5274 VSS.n228 VSS.n227 0.147
R5275 VSS.n503 VSS.n386 0.146
R5276 VSS.n503 VSS.n389 0.146
R5277 VSS.n325 VSS.n224 0.146
R5278 VSS.n485 VSS.n430 0.146
R5279 VSS.n503 VSS.n401 0.146
R5280 VSS.n349 VSS.n181 0.146
R5281 VSS.n325 VSS.n323 0.146
R5282 VSS.n325 VSS.n234 0.146
R5283 VSS.n325 VSS.n318 0.146
R5284 VSS VSS.n162 0.146
R5285 VSS VSS.n31 0.146
R5286 VSS VSS.n153 0.146
R5287 VSS VSS.n141 0.146
R5288 VSS VSS.n176 0.146
R5289 VSS VSS.n54 0.146
R5290 VSS VSS.n148 0.146
R5291 VSS VSS.n145 0.146
R5292 VSS VSS.n91 0.146
R5293 VSS VSS.n132 0.146
R5294 VSS.n325 VSS.n320 0.143
R5295 VSS.n325 VSS.n221 0.142
R5296 VSS.n485 VSS.n427 0.142
R5297 VSS.n349 VSS.n348 0.142
R5298 VSS.n494 VSS.n407 0.142
R5299 VSS.n503 VSS.n393 0.142
R5300 VSS VSS.n41 0.142
R5301 VSS VSS.n359 0.142
R5302 VSS VSS.n35 0.142
R5303 VSS VSS.n129 0.142
R5304 VSS VSS.n94 0.142
R5305 VSS VSS.n171 0.141
R5306 VSS VSS.n97 0.141
R5307 VSS.n349 VSS.n212 0.14
R5308 VSS.n485 VSS.n422 0.14
R5309 VSS VSS.n127 0.138
R5310 VSS VSS.n125 0.138
R5311 VSS.n503 VSS.n398 0.138
R5312 VSS.n325 VSS.n315 0.138
R5313 VSS.n501 VSS.n500 0.138
R5314 VSS.n503 VSS.n403 0.138
R5315 VSS VSS.n150 0.138
R5316 VSS VSS.n137 0.138
R5317 VSS.n328 VSS.n327 0.137
R5318 VSS VSS.n168 0.137
R5319 VSS VSS.n82 0.136
R5320 VSS.n497 VSS.n496 0.136
R5321 VSS.n485 VSS.n424 0.135
R5322 VSS VSS.n84 0.135
R5323 VSS.n339 VSS.n338 0.135
R5324 VSS.n488 VSS.n487 0.133
R5325 VSS VSS.n355 0.132
R5326 VSS.n344 VSS.n343 0.129
R5327 VSS VSS.n352 0.129
R5328 VSS.n504 VSS.n383 0.126
R5329 VSS.n427 VSS.n426 0.125
R5330 VSS.n386 VSS.n385 0.125
R5331 VSS.n227 VSS.n226 0.125
R5332 VSS.n212 VSS.n211 0.125
R5333 VSS.n389 VSS.n388 0.125
R5334 VSS.n422 VSS.n421 0.125
R5335 VSS.n224 VSS.n223 0.125
R5336 VSS.n348 VSS.n347 0.125
R5337 VSS.n430 VSS.n429 0.125
R5338 VSS.n401 VSS.n400 0.125
R5339 VSS.n181 VSS.n180 0.125
R5340 VSS.n323 VSS.n322 0.125
R5341 VSS.n234 VSS.n233 0.125
R5342 VSS.n318 VSS.n317 0.125
R5343 VSS.n162 VSS.n161 0.125
R5344 VSS.n359 VSS.n358 0.125
R5345 VSS.n31 VSS.n30 0.125
R5346 VSS.n153 VSS.n152 0.125
R5347 VSS.n141 VSS.n140 0.125
R5348 VSS.n35 VSS.n34 0.125
R5349 VSS.n176 VSS.n175 0.125
R5350 VSS.n54 VSS.n53 0.125
R5351 VSS.n148 VSS.n147 0.125
R5352 VSS.n97 VSS.n96 0.125
R5353 VSS.n145 VSS.n144 0.125
R5354 VSS.n94 VSS.n93 0.125
R5355 VSS.n91 VSS.n90 0.125
R5356 VSS.n132 VSS.n131 0.125
R5357 VSS.n49 VSS.n48 0.125
R5358 VSS.n505 VSS.n380 0.124
R5359 VSS VSS.n123 0.124
R5360 VSS.n349 VSS.n183 0.119
R5361 VSS.n485 VSS.n433 0.119
R5362 VSS.n113 VSS.n112 0.118
R5363 VSS.n485 VSS.n442 0.118
R5364 VSS.n349 VSS.n182 0.117
R5365 VSS.n410 VSS.n409 0.116
R5366 VSS.n21 VSS.n20 0.116
R5367 VSS.n76 VSS.n75 0.116
R5368 VSS.n68 VSS.n67 0.116
R5369 VSS.n194 VSS.n193 0.115
R5370 VSS.n362 VSS.n361 0.115
R5371 VSS.n188 VSS.n187 0.114
R5372 VSS.n368 VSS.n367 0.114
R5373 VSS.n106 VSS.n105 0.114
R5374 VSS.n438 VSS.n437 0.113
R5375 VSS.n207 VSS.n206 0.113
R5376 VSS.n445 VSS.n444 0.113
R5377 VSS.n6 VSS.n5 0.113
R5378 VSS.n374 VSS.n373 0.113
R5379 VSS.n100 VSS.n99 0.112
R5380 VSS.n14 VSS.n13 0.111
R5381 VSS.n2 VSS.n1 0.111
R5382 VSS.n416 VSS.n415 0.11
R5383 VSS.n200 VSS.n199 0.11
R5384 VSS.n304 VSS.n303 0.095
R5385 VSS.n253 VSS.n252 0.095
R5386 VSS.n260 VSS.n259 0.095
R5387 VSS.n283 VSS.n282 0.095
R5388 VSS.n289 VSS.n288 0.095
R5389 VSS.n296 VSS.n295 0.095
R5390 VSS.n276 VSS.n275 0.095
R5391 VSS.n269 VSS.n268 0.095
R5392 VSS VSS.n138 0.067
R5393 VSS.n307 VSS.n243 0.062
R5394 VSS.n307 VSS.n241 0.062
R5395 VSS.n307 VSS.n239 0.062
R5396 VSS.n237 VSS.n236 0.061
R5397 VSS VSS.n156 0.045
R5398 VSS VSS.n45 0.045
R5399 VSS VSS.n56 0.045
R5400 VSS VSS.n135 0.045
R5401 VSS.n349 VSS.n214 0.044
R5402 VSS.n336 VSS.n332 0.044
R5403 VSS VSS.n38 0.044
R5404 VSS VSS.n158 0.044
R5405 VSS VSS.n59 0.044
R5406 VSS VSS.n61 0.044
R5407 VSS.n438 VSS.n436 0.04
R5408 VSS.n188 VSS.n186 0.04
R5409 VSS VSS.n32 0.034
R5410 VSS.n469 VSS.n468 0.028
R5411 VSS.n467 VSS.n466 0.028
R5412 VSS.n481 VSS.n478 0.028
R5413 VSS.n465 VSS.n462 0.028
R5414 VSS.n477 VSS.n474 0.028
R5415 VSS.n473 VSS.n470 0.028
R5416 VSS.n483 VSS.n455 0.023
R5417 VSS.n485 VSS.n432 0.022
R5418 VSS.n325 VSS.n324 0.022
R5419 VSS.n503 VSS.n394 0.02
R5420 VSS.n447 VSS.n446 0.018
R5421 VSS.n196 VSS.n195 0.018
R5422 VSS.n202 VSS.n201 0.018
R5423 VSS.n16 VSS.n15 0.018
R5424 VSS.n370 VSS.n369 0.018
R5425 VSS.n23 VSS.n22 0.018
R5426 VSS.n364 VSS.n363 0.018
R5427 VSS.n8 VSS.n7 0.018
R5428 VSS.n376 VSS.n375 0.018
R5429 VSS VSS.n36 0.018
R5430 VSS VSS.n159 0.018
R5431 VSS VSS.n142 0.018
R5432 VSS.n111 VSS.n110 0.018
R5433 VSS.n108 VSS.n107 0.018
R5434 VSS.n78 VSS.n77 0.018
R5435 VSS.n102 VSS.n101 0.018
R5436 VSS.n70 VSS.n69 0.018
R5437 VSS.n4 VSS.n3 0.018
R5438 VSS.n503 VSS.n391 0.018
R5439 VSS.n325 VSS.n229 0.018
R5440 VSS.n325 VSS.n230 0.018
R5441 VSS.n325 VSS.n231 0.018
R5442 VSS.n494 VSS.n493 0.017
R5443 VSS VSS.n166 0.017
R5444 VSS VSS.n64 0.017
R5445 VSS VSS.n165 0.017
R5446 VSS VSS.n63 0.017
R5447 VSS VSS.n164 0.017
R5448 VSS VSS.n62 0.017
R5449 VSS.n217 VSS.n216 0.016
R5450 VSS.n336 VSS.n335 0.015
R5451 VSS.n336 VSS.n334 0.015
R5452 VSS.n336 VSS.n333 0.015
R5453 VSS.n494 VSS.n405 0.015
R5454 VSS VSS.n178 0.015
R5455 VSS VSS.n350 0.015
R5456 VSS VSS.n65 0.015
R5457 VSS VSS.n116 0.015
R5458 VSS VSS.n154 0.014
R5459 VSS VSS.n43 0.014
R5460 VSS VSS.n57 0.014
R5461 VSS VSS.n133 0.014
R5462 VSS.n485 VSS.n431 0.011
R5463 VSS.n494 VSS.n491 0.011
R5464 VSS.n336 VSS.n330 0.011
R5465 VSS.n209 VSS.n208 0.011
R5466 VSS.n10 VSS.n9 0.011
R5467 VSS.n8 VSS.n6 0.01
R5468 VSS VSS.n120 0.009
R5469 VSS.n196 VSS.n194 0.007
R5470 VSS.n329 VSS.n328 0.007
R5471 VSS.n418 VSS.n416 0.006
R5472 VSS.n447 VSS.n445 0.006
R5473 VSS.n202 VSS.n200 0.006
R5474 VSS.n494 VSS.n492 0.006
R5475 VSS.n115 VSS.n114 0.006
R5476 VSS.n502 VSS.n501 0.005
R5477 VSS.n341 VSS.n217 0.005
R5478 VSS.n370 VSS.n368 0.005
R5479 VSS.n364 VSS.n362 0.005
R5480 VSS.n376 VSS.n374 0.005
R5481 VSS VSS.n42 0.005
R5482 VSS VSS.n50 0.005
R5483 VSS VSS.n119 0.005
R5484 VSS.n78 VSS.n76 0.005
R5485 VSS.n102 VSS.n100 0.005
R5486 VSS.n306 VSS.n305 0.005
R5487 VSS.n483 VSS.n482 0.004
R5488 VSS.n345 VSS.n344 0.004
R5489 VSS.n412 VSS.n410 0.004
R5490 VSS.n108 VSS.n106 0.004
R5491 VSS.n4 VSS.n2 0.004
R5492 VSS.n349 VSS.n215 0.004
R5493 VSS.n489 VSS.n488 0.004
R5494 VSS.n498 VSS.n497 0.004
R5495 VSS.n340 VSS.n339 0.004
R5496 VSS.n505 VSS.n504 0.003
R5497 VSS.n325 VSS.n228 0.003
R5498 VSS.n23 VSS.n21 0.003
R5499 VSS.n70 VSS.n68 0.003
R5500 VSS.n418 VSS.n417 0.003
R5501 VSS.n412 VSS.n411 0.003
R5502 VSS.n439 VSS.n438 0.003
R5503 VSS.n264 VSS.n263 0.002
R5504 VSS.n205 VSS.n204 0.002
R5505 VSS.n16 VSS.n14 0.002
R5506 VSS VSS.n173 0.002
R5507 VSS VSS.n118 0.002
R5508 VSS VSS.n117 0.002
R5509 VSS.n485 VSS.n484 0.002
R5510 VSS.n484 VSS.n483 0.002
R5511 VSS.n189 VSS.n188 0.002
R5512 VSS VSS.n18 0.002
R5513 VSS VSS.n25 0.002
R5514 VSS VSS.n80 0.002
R5515 VSS VSS.n11 0.002
R5516 VSS VSS.n72 0.002
R5517 VSS.n197 VSS.n196 0.001
R5518 VSS.n349 VSS.n197 0.001
R5519 VSS.n203 VSS.n202 0.001
R5520 VSS.n349 VSS.n203 0.001
R5521 VSS.n485 VSS.n448 0.001
R5522 VSS.n448 VSS.n447 0.001
R5523 VSS.n191 VSS.n190 0.001
R5524 VSS.n349 VSS.n191 0.001
R5525 VSS.n307 VSS.n237 0.001
R5526 VSS VSS.n49 0.001
R5527 VSS VSS.n28 0.001
R5528 VSS VSS.n88 0.001
R5529 VSS.n474 VSS.n473 0.001
R5530 VSS.n466 VSS.n465 0.001
R5531 VSS.n482 VSS.n481 0.001
R5532 VSS.n478 VSS.n477 0.001
R5533 VSS.n470 VSS.n469 0.001
R5534 VSS.n468 VSS.n467 0.001
R5535 VSS.n307 VSS.n306 0.001
R5536 VSS.n325 VSS.n307 0.001
R5537 VSS VSS.n349 0.001
R5538 VSS VSS.n505 0.001
R5539 VSS.n441 VSS.n440 0.001
R5540 VSS.n485 VSS.n441 0.001
R5541 VSS.n336 VSS.n219 0.001
R5542 VSS.n341 VSS.n218 0.001
R5543 VSS.n494 VSS.n490 0.001
R5544 VSS.n345 VSS.n341 0.001
R5545 VSS.n349 VSS.n345 0.001
R5546 VSS.n305 VSS.n304 0.001
R5547 VSS.n305 VSS.n253 0.001
R5548 VSS.n305 VSS.n260 0.001
R5549 VSS.n305 VSS.n283 0.001
R5550 VSS.n305 VSS.n289 0.001
R5551 VSS.n305 VSS.n296 0.001
R5552 VSS.n305 VSS.n276 0.001
R5553 VSS.n305 VSS.n269 0.001
R5554 VSS.n304 VSS.n300 0.001
R5555 VSS.n253 VSS.n249 0.001
R5556 VSS.n260 VSS.n256 0.001
R5557 VSS.n283 VSS.n279 0.001
R5558 VSS.n289 VSS.n285 0.001
R5559 VSS.n296 VSS.n292 0.001
R5560 VSS.n276 VSS.n272 0.001
R5561 VSS.n269 VSS.n265 0.001
R5562 VSS VSS.n26 0.001
R5563 VSS VSS.n27 0.001
R5564 VSS VSS.n85 0.001
R5565 VSS VSS.n86 0.001
R5566 VSS VSS.n87 0.001
R5567 VSS.n190 VSS.n184 0.001
R5568 VSS.n440 VSS.n434 0.001
R5569 VSS.n416 VSS.n414 0.001
R5570 VSS.n200 VSS.n198 0.001
R5571 VSS.n305 VSS.n277 0.001
R5572 VSS.n14 VSS.n12 0.001
R5573 VSS.n2 VSS.n0 0.001
R5574 VSS.n305 VSS.n297 0.001
R5575 VSS.n100 VSS.n98 0.001
R5576 VSS.n305 VSS.n270 0.001
R5577 VSS.n305 VSS.n254 0.001
R5578 VSS.n445 VSS.n443 0.001
R5579 VSS.n374 VSS.n372 0.001
R5580 VSS.n208 VSS.n207 0.001
R5581 VSS.n106 VSS.n104 0.001
R5582 VSS.n368 VSS.n366 0.001
R5583 VSS.n362 VSS.n360 0.001
R5584 VSS.n194 VSS.n192 0.001
R5585 VSS.n305 VSS.n261 0.001
R5586 VSS.n305 VSS.n262 0.001
R5587 VSS.n21 VSS.n19 0.001
R5588 VSS.n68 VSS.n66 0.001
R5589 VSS.n305 VSS.n298 0.001
R5590 VSS.n410 VSS.n408 0.001
R5591 VSS.n76 VSS.n74 0.001
R5592 VSS.n305 VSS.n290 0.001
R5593 VSS.n114 VSS.n113 0.001
R5594 VSS.n305 VSS.n248 0.001
R5595 VSS.n305 VSS.n255 0.001
R5596 VSS.n305 VSS.n284 0.001
R5597 VSS.n305 VSS.n291 0.001
R5598 VSS.n305 VSS.n271 0.001
R5599 VSS.n305 VSS.n299 0.001
R5600 VSS.n305 VSS.n278 0.001
R5601 VSS.n305 VSS.n264 0.001
R5602 VSS VSS.n172 0.001
R5603 VSS VSS.n356 0.001
R5604 VSS VSS.n353 0.001
R5605 VSS VSS.n169 0.001
R5606 VSS.n504 VSS.n503 0.001
R5607 VSS.n439 VSS.n435 0.001
R5608 VSS.n440 VSS.n439 0.001
R5609 VSS.n349 VSS.n209 0.001
R5610 VSS.n485 VSS.n419 0.001
R5611 VSS.n503 VSS.n502 0.001
R5612 VSS.n329 VSS.n325 0.001
R5613 VSS.n485 VSS.n413 0.001
R5614 VSS.n494 VSS.n489 0.001
R5615 VSS.n503 VSS.n498 0.001
R5616 VSS.n340 VSS.n336 0.001
R5617 VSS.n189 VSS.n185 0.001
R5618 VSS.n190 VSS.n189 0.001
R5619 VSS VSS.n17 0.001
R5620 VSS VSS.n371 0.001
R5621 VSS VSS.n24 0.001
R5622 VSS VSS.n365 0.001
R5623 VSS VSS.n10 0.001
R5624 VSS VSS.n377 0.001
R5625 VSS VSS.n177 0.001
R5626 VSS VSS.n163 0.001
R5627 VSS VSS.n51 0.001
R5628 VSS VSS.n115 0.001
R5629 VSS VSS.n109 0.001
R5630 VSS VSS.n79 0.001
R5631 VSS VSS.n103 0.001
R5632 VSS VSS.n71 0.001
R5633 VSS.n506 VSS 0.001
R5634 VSS.n341 VSS.n340 0.001
R5635 VSS.n489 VSS.n485 0.001
R5636 VSS.n377 VSS.n376 0.001
R5637 VSS.n498 VSS.n494 0.001
R5638 VSS.n506 VSS.n4 0.001
R5639 VSS.n365 VSS.n364 0.001
R5640 VSS.n103 VSS.n102 0.001
R5641 VSS.n413 VSS.n412 0.001
R5642 VSS.n24 VSS.n23 0.001
R5643 VSS.n79 VSS.n78 0.001
R5644 VSS.n336 VSS.n329 0.001
R5645 VSS.n71 VSS.n70 0.001
R5646 VSS.n10 VSS.n8 0.001
R5647 VSS.n109 VSS.n108 0.001
R5648 VSS.n371 VSS.n370 0.001
R5649 VSS.n419 VSS.n418 0.001
R5650 VSS.n209 VSS.n205 0.001
R5651 VSS.n115 VSS.n111 0.001
R5652 VSS.n17 VSS.n16 0.001
R5653 a_17946_9198.t5 a_17946_9198.t4 574.43
R5654 a_17946_9198.n1 a_17946_9198.t7 285.109
R5655 a_17946_9198.n3 a_17946_9198.n2 197.217
R5656 a_17946_9198.n4 a_17946_9198.n0 192.754
R5657 a_17946_9198.n1 a_17946_9198.t6 160.666
R5658 a_17946_9198.n2 a_17946_9198.t5 160.666
R5659 a_17946_9198.n2 a_17946_9198.n1 114.829
R5660 a_17946_9198.t3 a_17946_9198.n4 28.568
R5661 a_17946_9198.n0 a_17946_9198.t2 28.565
R5662 a_17946_9198.n0 a_17946_9198.t1 28.565
R5663 a_17946_9198.n3 a_17946_9198.t0 18.838
R5664 a_17946_9198.n4 a_17946_9198.n3 1.129
R5665 a_n3111_15192.n0 a_n3111_15192.t2 14.282
R5666 a_n3111_15192.t0 a_n3111_15192.n0 14.282
R5667 a_n3111_15192.n0 a_n3111_15192.n16 90.436
R5668 a_n3111_15192.n16 a_n3111_15192.n2 74.302
R5669 a_n3111_15192.n2 a_n3111_15192.n4 50.575
R5670 a_n3111_15192.n4 a_n3111_15192.n5 110.084
R5671 a_n3111_15192.n16 a_n3111_15192.n6 201.691
R5672 a_n3111_15192.n6 a_n3111_15192.n8 16.411
R5673 a_n3111_15192.n8 a_n3111_15192.t13 198.921
R5674 a_n3111_15192.t13 a_n3111_15192.t14 415.315
R5675 a_n3111_15192.t14 a_n3111_15192.n15 214.335
R5676 a_n3111_15192.n15 a_n3111_15192.t16 80.333
R5677 a_n3111_15192.n15 a_n3111_15192.t17 214.335
R5678 a_n3111_15192.n8 a_n3111_15192.n14 861.987
R5679 a_n3111_15192.n14 a_n3111_15192.n9 560.726
R5680 a_n3111_15192.n14 a_n3111_15192.n13 65.07
R5681 a_n3111_15192.n13 a_n3111_15192.n12 6.615
R5682 a_n3111_15192.n12 a_n3111_15192.t20 93.989
R5683 a_n3111_15192.n13 a_n3111_15192.n11 97.816
R5684 a_n3111_15192.n11 a_n3111_15192.t23 80.333
R5685 a_n3111_15192.n11 a_n3111_15192.t8 394.151
R5686 a_n3111_15192.t8 a_n3111_15192.n10 269.523
R5687 a_n3111_15192.n10 a_n3111_15192.t12 160.666
R5688 a_n3111_15192.n10 a_n3111_15192.t11 269.523
R5689 a_n3111_15192.n12 a_n3111_15192.t19 198.043
R5690 a_n3111_15192.n9 a_n3111_15192.t22 294.653
R5691 a_n3111_15192.n9 a_n3111_15192.t21 111.663
R5692 a_n3111_15192.n6 a_n3111_15192.t15 217.716
R5693 a_n3111_15192.t15 a_n3111_15192.t9 415.315
R5694 a_n3111_15192.t9 a_n3111_15192.n7 214.335
R5695 a_n3111_15192.n7 a_n3111_15192.t10 80.333
R5696 a_n3111_15192.n7 a_n3111_15192.t18 214.335
R5697 a_n3111_15192.n5 a_n3111_15192.t4 14.282
R5698 a_n3111_15192.n5 a_n3111_15192.t6 14.282
R5699 a_n3111_15192.n4 a_n3111_15192.n3 157.665
R5700 a_n3111_15192.n3 a_n3111_15192.t3 8.7
R5701 a_n3111_15192.n3 a_n3111_15192.t5 8.7
R5702 a_n3111_15192.n2 a_n3111_15192.n1 90.416
R5703 a_n3111_15192.n1 a_n3111_15192.t1 14.282
R5704 a_n3111_15192.n1 a_n3111_15192.t7 14.282
R5705 a_7735_24460.n0 a_7735_24460.n1 0.001
R5706 a_7735_24460.n0 a_7735_24460.t1 14.282
R5707 a_7735_24460.t3 a_7735_24460.n0 14.282
R5708 a_7735_24460.n1 a_7735_24460.n9 267.767
R5709 a_7735_24460.n9 a_7735_24460.t4 14.282
R5710 a_7735_24460.n9 a_7735_24460.t5 14.282
R5711 a_7735_24460.n1 a_7735_24460.n7 0.669
R5712 a_7735_24460.n7 a_7735_24460.n8 1.511
R5713 a_7735_24460.n8 a_7735_24460.t2 14.282
R5714 a_7735_24460.n8 a_7735_24460.t0 14.282
R5715 a_7735_24460.n7 a_7735_24460.n6 0.227
R5716 a_7735_24460.n6 a_7735_24460.n3 0.575
R5717 a_7735_24460.n6 a_7735_24460.n5 0.2
R5718 a_7735_24460.n5 a_7735_24460.t8 16.058
R5719 a_7735_24460.n5 a_7735_24460.n4 0.999
R5720 a_7735_24460.n4 a_7735_24460.t6 14.282
R5721 a_7735_24460.n4 a_7735_24460.t7 14.282
R5722 a_7735_24460.n3 a_7735_24460.n2 0.999
R5723 a_7735_24460.n2 a_7735_24460.t9 14.282
R5724 a_7735_24460.n2 a_7735_24460.t10 14.282
R5725 a_7735_24460.n3 a_7735_24460.t11 16.058
R5726 a_8419_26709.t7 a_8419_26709.t6 800.071
R5727 a_8419_26709.n3 a_8419_26709.n2 672.951
R5728 a_8419_26709.n1 a_8419_26709.t5 285.109
R5729 a_8419_26709.n2 a_8419_26709.t7 193.602
R5730 a_8419_26709.n1 a_8419_26709.t4 160.666
R5731 a_8419_26709.n2 a_8419_26709.n1 91.507
R5732 a_8419_26709.n0 a_8419_26709.t1 28.57
R5733 a_8419_26709.t0 a_8419_26709.n4 28.565
R5734 a_8419_26709.n4 a_8419_26709.t3 28.565
R5735 a_8419_26709.n0 a_8419_26709.t2 17.638
R5736 a_8419_26709.n4 a_8419_26709.n3 0.69
R5737 a_8419_26709.n3 a_8419_26709.n0 0.6
R5738 a_9415_27296.n0 a_9415_27296.t0 14.282
R5739 a_9415_27296.n0 a_9415_27296.t5 14.282
R5740 a_9415_27296.n1 a_9415_27296.t1 14.282
R5741 a_9415_27296.n1 a_9415_27296.t2 14.282
R5742 a_9415_27296.n3 a_9415_27296.t4 14.282
R5743 a_9415_27296.t3 a_9415_27296.n3 14.282
R5744 a_9415_27296.n3 a_9415_27296.n2 2.546
R5745 a_9415_27296.n2 a_9415_27296.n1 2.367
R5746 a_9415_27296.n2 a_9415_27296.n0 0.001
R5747 A[3].n16 A[3].n6 2170.52
R5748 A[3].n11 A[3].n10 535.449
R5749 A[3].t17 A[3].t1 437.233
R5750 A[3].t19 A[3].t20 437.233
R5751 A[3].t23 A[3].t24 437.233
R5752 A[3].t22 A[3].t10 415.315
R5753 A[3].t11 A[3].t12 415.315
R5754 A[3].t9 A[3].t28 415.315
R5755 A[3].t14 A[3].n8 313.873
R5756 A[3].n10 A[3].t8 294.986
R5757 A[3].n7 A[3].t2 272.288
R5758 A[3].n11 A[3].t27 245.184
R5759 A[3].n5 A[3].t11 221.468
R5760 A[3].n2 A[3].t17 219.798
R5761 A[3].n13 A[3].t23 218.628
R5762 A[3].n2 A[3].t22 217.276
R5763 A[3].n5 A[3].t9 217.129
R5764 A[3].n15 A[3].t19 217.024
R5765 A[3].n1 A[3].t31 214.686
R5766 A[3].t1 A[3].n1 214.686
R5767 A[3].n14 A[3].t29 214.686
R5768 A[3].t20 A[3].n14 214.686
R5769 A[3].n12 A[3].t16 214.686
R5770 A[3].t24 A[3].n12 214.686
R5771 A[3].n0 A[3].t26 214.335
R5772 A[3].t10 A[3].n0 214.335
R5773 A[3].n3 A[3].t25 214.335
R5774 A[3].t12 A[3].n3 214.335
R5775 A[3].n4 A[3].t6 214.335
R5776 A[3].t28 A[3].n4 214.335
R5777 A[3].n9 A[3].t14 190.152
R5778 A[3].n9 A[3].t4 190.152
R5779 A[3].n7 A[3].t3 160.666
R5780 A[3].n8 A[3].t30 160.666
R5781 A[3].n10 A[3].t15 110.859
R5782 A[3].n8 A[3].n7 96.129
R5783 A[3].n1 A[3].t0 80.333
R5784 A[3].n0 A[3].t13 80.333
R5785 A[3].n3 A[3].t5 80.333
R5786 A[3].n4 A[3].t21 80.333
R5787 A[3].n14 A[3].t7 80.333
R5788 A[3].t27 A[3].n9 80.333
R5789 A[3].n12 A[3].t18 80.333
R5790 A[3].n6 A[3].n5 54.612
R5791 A[3].n6 A[3].n2 49.781
R5792 A[3].n16 A[3].n15 28.756
R5793 A[3].n13 A[3].n11 14.9
R5794 A[3] A[3].n16 2.747
R5795 A[3].n15 A[3].n13 2.599
R5796 a_29769_12318.n2 a_29769_12318.t9 214.335
R5797 a_29769_12318.t7 a_29769_12318.n2 214.335
R5798 a_29769_12318.n3 a_29769_12318.t7 143.851
R5799 a_29769_12318.n3 a_29769_12318.t10 135.658
R5800 a_29769_12318.n2 a_29769_12318.t8 80.333
R5801 a_29769_12318.n4 a_29769_12318.t6 28.565
R5802 a_29769_12318.n4 a_29769_12318.t5 28.565
R5803 a_29769_12318.n0 a_29769_12318.t3 28.565
R5804 a_29769_12318.n0 a_29769_12318.t1 28.565
R5805 a_29769_12318.t4 a_29769_12318.n7 28.565
R5806 a_29769_12318.n7 a_29769_12318.t2 28.565
R5807 a_29769_12318.n1 a_29769_12318.t0 9.714
R5808 a_29769_12318.n1 a_29769_12318.n0 1.003
R5809 a_29769_12318.n6 a_29769_12318.n5 0.833
R5810 a_29769_12318.n5 a_29769_12318.n4 0.653
R5811 a_29769_12318.n7 a_29769_12318.n6 0.653
R5812 a_29769_12318.n6 a_29769_12318.n1 0.341
R5813 a_29769_12318.n5 a_29769_12318.n3 0.032
R5814 a_21466_26701.t7 a_21466_26701.t6 800.071
R5815 a_21466_26701.n3 a_21466_26701.n2 672.951
R5816 a_21466_26701.n1 a_21466_26701.t5 285.109
R5817 a_21466_26701.n2 a_21466_26701.t7 193.602
R5818 a_21466_26701.n1 a_21466_26701.t4 160.666
R5819 a_21466_26701.n2 a_21466_26701.n1 91.507
R5820 a_21466_26701.t0 a_21466_26701.n4 28.57
R5821 a_21466_26701.n0 a_21466_26701.t3 28.565
R5822 a_21466_26701.n0 a_21466_26701.t2 28.565
R5823 a_21466_26701.n4 a_21466_26701.t1 17.638
R5824 a_21466_26701.n3 a_21466_26701.n0 0.69
R5825 a_21466_26701.n4 a_21466_26701.n3 0.6
R5826 a_22462_27288.n0 a_22462_27288.t1 14.282
R5827 a_22462_27288.n0 a_22462_27288.t2 14.282
R5828 a_22462_27288.n1 a_22462_27288.t4 14.282
R5829 a_22462_27288.n1 a_22462_27288.t5 14.282
R5830 a_22462_27288.n3 a_22462_27288.t3 14.282
R5831 a_22462_27288.t0 a_22462_27288.n3 14.282
R5832 a_22462_27288.n2 a_22462_27288.n0 2.546
R5833 a_22462_27288.n2 a_22462_27288.n1 2.367
R5834 a_22462_27288.n3 a_22462_27288.n2 0.001
R5835 a_30430_6928.n5 a_30430_6928.n4 465.933
R5836 a_30430_6928.t15 a_30430_6928.t4 415.315
R5837 a_30430_6928.n1 a_30430_6928.t5 394.151
R5838 a_30430_6928.n4 a_30430_6928.t10 294.653
R5839 a_30430_6928.n0 a_30430_6928.t7 269.523
R5840 a_30430_6928.t5 a_30430_6928.n0 269.523
R5841 a_30430_6928.n7 a_30430_6928.t15 220.285
R5842 a_30430_6928.n6 a_30430_6928.t14 214.335
R5843 a_30430_6928.t4 a_30430_6928.n6 214.335
R5844 a_30430_6928.n2 a_30430_6928.t11 198.043
R5845 a_30430_6928.n10 a_30430_6928.n9 192.754
R5846 a_30430_6928.n5 a_30430_6928.n3 163.88
R5847 a_30430_6928.n0 a_30430_6928.t6 160.666
R5848 a_30430_6928.n4 a_30430_6928.t9 111.663
R5849 a_30430_6928.n3 a_30430_6928.n1 97.816
R5850 a_30430_6928.n2 a_30430_6928.t12 93.989
R5851 a_30430_6928.n6 a_30430_6928.t8 80.333
R5852 a_30430_6928.n1 a_30430_6928.t13 80.333
R5853 a_30430_6928.n7 a_30430_6928.n5 61.538
R5854 a_30430_6928.n9 a_30430_6928.t1 28.568
R5855 a_30430_6928.n10 a_30430_6928.t3 28.565
R5856 a_30430_6928.t0 a_30430_6928.n10 28.565
R5857 a_30430_6928.n8 a_30430_6928.t2 18.824
R5858 a_30430_6928.n3 a_30430_6928.n2 6.615
R5859 a_30430_6928.n8 a_30430_6928.n7 5.5
R5860 a_30430_6928.n9 a_30430_6928.n8 1.105
R5861 a_33377_10390.n0 a_33377_10390.t10 214.335
R5862 a_33377_10390.t8 a_33377_10390.n0 214.335
R5863 a_33377_10390.n1 a_33377_10390.t8 143.851
R5864 a_33377_10390.n1 a_33377_10390.t7 135.658
R5865 a_33377_10390.n0 a_33377_10390.t9 80.333
R5866 a_33377_10390.n2 a_33377_10390.t0 28.565
R5867 a_33377_10390.n2 a_33377_10390.t1 28.565
R5868 a_33377_10390.n4 a_33377_10390.t2 28.565
R5869 a_33377_10390.n4 a_33377_10390.t6 28.565
R5870 a_33377_10390.n7 a_33377_10390.t5 28.565
R5871 a_33377_10390.t4 a_33377_10390.n7 28.565
R5872 a_33377_10390.n6 a_33377_10390.t3 9.714
R5873 a_33377_10390.n7 a_33377_10390.n6 1.003
R5874 a_33377_10390.n5 a_33377_10390.n3 0.833
R5875 a_33377_10390.n3 a_33377_10390.n2 0.653
R5876 a_33377_10390.n5 a_33377_10390.n4 0.653
R5877 a_33377_10390.n6 a_33377_10390.n5 0.341
R5878 a_33377_10390.n3 a_33377_10390.n1 0.032
R5879 a_31466_2550.n1 a_31466_2550.t4 318.922
R5880 a_31466_2550.n0 a_31466_2550.t5 273.935
R5881 a_31466_2550.n0 a_31466_2550.t7 273.935
R5882 a_31466_2550.n1 a_31466_2550.t6 269.116
R5883 a_31466_2550.n4 a_31466_2550.n3 193.227
R5884 a_31466_2550.t4 a_31466_2550.n0 179.142
R5885 a_31466_2550.n2 a_31466_2550.n1 106.999
R5886 a_31466_2550.n3 a_31466_2550.t1 28.568
R5887 a_31466_2550.n4 a_31466_2550.t2 28.565
R5888 a_31466_2550.t0 a_31466_2550.n4 28.565
R5889 a_31466_2550.n2 a_31466_2550.t3 18.149
R5890 a_31466_2550.n3 a_31466_2550.n2 3.726
R5891 a_32011_1857.n0 a_32011_1857.t7 14.282
R5892 a_32011_1857.t1 a_32011_1857.n0 14.282
R5893 a_32011_1857.n0 a_32011_1857.n8 90.416
R5894 a_32011_1857.n8 a_32011_1857.n7 50.575
R5895 a_32011_1857.n8 a_32011_1857.n4 74.302
R5896 a_32011_1857.n7 a_32011_1857.n6 157.665
R5897 a_32011_1857.n6 a_32011_1857.t4 8.7
R5898 a_32011_1857.n6 a_32011_1857.t0 8.7
R5899 a_32011_1857.n7 a_32011_1857.n5 122.999
R5900 a_32011_1857.n5 a_32011_1857.t5 14.282
R5901 a_32011_1857.n5 a_32011_1857.t6 14.282
R5902 a_32011_1857.n4 a_32011_1857.n3 90.436
R5903 a_32011_1857.n3 a_32011_1857.t3 14.282
R5904 a_32011_1857.n3 a_32011_1857.t2 14.282
R5905 a_32011_1857.n4 a_32011_1857.n1 154.155
R5906 a_32011_1857.n1 a_32011_1857.t11 408.806
R5907 a_32011_1857.t8 a_32011_1857.n2 160.666
R5908 a_32011_1857.n1 a_32011_1857.t8 989.744
R5909 a_32011_1857.n2 a_32011_1857.t10 287.241
R5910 a_32011_1857.n2 a_32011_1857.t9 287.241
R5911 a_31893_1857.t0 a_31893_1857.n0 14.282
R5912 a_31893_1857.n0 a_31893_1857.t5 14.282
R5913 a_31893_1857.n0 a_31893_1857.n9 0.999
R5914 a_31893_1857.n6 a_31893_1857.n8 0.575
R5915 a_31893_1857.n9 a_31893_1857.n6 0.2
R5916 a_31893_1857.n9 a_31893_1857.t1 16.058
R5917 a_31893_1857.n8 a_31893_1857.n7 0.999
R5918 a_31893_1857.n7 a_31893_1857.t8 14.282
R5919 a_31893_1857.n7 a_31893_1857.t6 14.282
R5920 a_31893_1857.n8 a_31893_1857.t7 16.058
R5921 a_31893_1857.n6 a_31893_1857.n4 0.227
R5922 a_31893_1857.n4 a_31893_1857.n5 1.511
R5923 a_31893_1857.n5 a_31893_1857.t3 14.282
R5924 a_31893_1857.n5 a_31893_1857.t4 14.282
R5925 a_31893_1857.n4 a_31893_1857.n1 0.669
R5926 a_31893_1857.n1 a_31893_1857.n2 0.001
R5927 a_31893_1857.n1 a_31893_1857.n3 267.767
R5928 a_31893_1857.n3 a_31893_1857.t9 14.282
R5929 a_31893_1857.n3 a_31893_1857.t11 14.282
R5930 a_31893_1857.n2 a_31893_1857.t2 14.282
R5931 a_31893_1857.n2 a_31893_1857.t10 14.282
R5932 a_17301_11213.n17 a_17301_11213.n16 538.835
R5933 a_17301_11213.n9 a_17301_11213.n8 501.28
R5934 a_17301_11213.t6 a_17301_11213.t19 437.233
R5935 a_17301_11213.t7 a_17301_11213.t4 415.315
R5936 a_17301_11213.t8 a_17301_11213.n6 313.873
R5937 a_17301_11213.n8 a_17301_11213.t17 294.986
R5938 a_17301_11213.n5 a_17301_11213.t11 272.288
R5939 a_17301_11213.n9 a_17301_11213.t12 236.01
R5940 a_17301_11213.n12 a_17301_11213.t6 216.627
R5941 a_17301_11213.n10 a_17301_11213.t7 216.111
R5942 a_17301_11213.n11 a_17301_11213.t14 214.686
R5943 a_17301_11213.t19 a_17301_11213.n11 214.686
R5944 a_17301_11213.n4 a_17301_11213.t5 214.335
R5945 a_17301_11213.t4 a_17301_11213.n4 214.335
R5946 a_17301_11213.n19 a_17301_11213.n18 192.754
R5947 a_17301_11213.n7 a_17301_11213.t8 190.152
R5948 a_17301_11213.n7 a_17301_11213.t13 190.152
R5949 a_17301_11213.n5 a_17301_11213.t15 160.666
R5950 a_17301_11213.n6 a_17301_11213.t16 160.666
R5951 a_17301_11213.n10 a_17301_11213.n9 148.428
R5952 a_17301_11213.n8 a_17301_11213.t10 110.859
R5953 a_17301_11213.n6 a_17301_11213.n5 96.129
R5954 a_17301_11213.n11 a_17301_11213.t18 80.333
R5955 a_17301_11213.n4 a_17301_11213.t9 80.333
R5956 a_17301_11213.t12 a_17301_11213.n7 80.333
R5957 a_17301_11213.n18 a_17301_11213.t2 28.568
R5958 a_17301_11213.n19 a_17301_11213.t3 28.565
R5959 a_17301_11213.t1 a_17301_11213.n19 28.565
R5960 a_17301_11213.n17 a_17301_11213.t0 18.514
R5961 a_17301_11213.n16 a_17301_11213.n15 4.161
R5962 a_17301_11213.n12 a_17301_11213.n10 2.923
R5963 a_17301_11213.n18 a_17301_11213.n17 1.177
R5964 a_17301_11213.n13 a_17301_11213.n12 0.707
R5965 a_17301_11213.n15 a_17301_11213.n14 0.078
R5966 a_17301_11213.n1 a_17301_11213.n0 0.045
R5967 a_17301_11213.n3 a_17301_11213.n2 0.006
R5968 a_17301_11213.n15 a_17301_11213.n1 0.003
R5969 a_17301_11213.n13 a_17301_11213.n3 0.002
R5970 a_17301_11213.n15 a_17301_11213.n13 0.001
R5971 A[6].n16 A[6].n6 2865.54
R5972 A[6].n2 A[6].t25 2858.78
R5973 A[6].n6 A[6].n2 2573.2
R5974 A[6].n11 A[6].n10 535.449
R5975 A[6].t25 A[6].t29 437.233
R5976 A[6].t0 A[6].t24 437.233
R5977 A[6].t31 A[6].t13 437.233
R5978 A[6].t22 A[6].t17 415.315
R5979 A[6].t10 A[6].t2 415.315
R5980 A[6].t11 A[6].t28 415.315
R5981 A[6].t19 A[6].n8 313.873
R5982 A[6].n10 A[6].t4 294.986
R5983 A[6].n7 A[6].t12 272.288
R5984 A[6].n11 A[6].t9 245.184
R5985 A[6].n5 A[6].t11 238.523
R5986 A[6].n13 A[6].t31 218.627
R5987 A[6].n5 A[6].t10 217.897
R5988 A[6].n2 A[6].t22 217.528
R5989 A[6].n15 A[6].t0 217.023
R5990 A[6].n1 A[6].t16 214.686
R5991 A[6].t29 A[6].n1 214.686
R5992 A[6].n14 A[6].t5 214.686
R5993 A[6].t24 A[6].n14 214.686
R5994 A[6].n12 A[6].t21 214.686
R5995 A[6].t13 A[6].n12 214.686
R5996 A[6].n0 A[6].t30 214.335
R5997 A[6].t17 A[6].n0 214.335
R5998 A[6].n3 A[6].t15 214.335
R5999 A[6].t2 A[6].n3 214.335
R6000 A[6].n4 A[6].t8 214.335
R6001 A[6].t28 A[6].n4 214.335
R6002 A[6].n9 A[6].t6 190.152
R6003 A[6].n9 A[6].t19 190.152
R6004 A[6].n7 A[6].t1 160.666
R6005 A[6].n8 A[6].t3 160.666
R6006 A[6].n10 A[6].t23 110.859
R6007 A[6].n8 A[6].n7 96.129
R6008 A[6].n0 A[6].t18 80.333
R6009 A[6].n1 A[6].t27 80.333
R6010 A[6].n3 A[6].t20 80.333
R6011 A[6].n4 A[6].t7 80.333
R6012 A[6].n14 A[6].t26 80.333
R6013 A[6].t9 A[6].n9 80.333
R6014 A[6].n12 A[6].t14 80.333
R6015 A[6].n16 A[6].n15 37.965
R6016 A[6].n13 A[6].n11 14.9
R6017 A[6].n15 A[6].n13 2.599
R6018 A[6] A[6].n16 2.485
R6019 A[6].n6 A[6].n5 0.274
R6020 a_16219_21171.t0 a_16219_21171.t1 17.4
R6021 a_15570_21782.n0 a_15570_21782.t7 214.335
R6022 a_15570_21782.t9 a_15570_21782.n0 214.335
R6023 a_15570_21782.n1 a_15570_21782.t9 143.851
R6024 a_15570_21782.n1 a_15570_21782.t10 135.658
R6025 a_15570_21782.n0 a_15570_21782.t8 80.333
R6026 a_15570_21782.n4 a_15570_21782.t3 28.565
R6027 a_15570_21782.n4 a_15570_21782.t1 28.565
R6028 a_15570_21782.n2 a_15570_21782.t6 28.565
R6029 a_15570_21782.n2 a_15570_21782.t5 28.565
R6030 a_15570_21782.n7 a_15570_21782.t2 28.565
R6031 a_15570_21782.t4 a_15570_21782.n7 28.565
R6032 a_15570_21782.n5 a_15570_21782.t0 9.714
R6033 a_15570_21782.n5 a_15570_21782.n4 1.003
R6034 a_15570_21782.n6 a_15570_21782.n3 0.833
R6035 a_15570_21782.n3 a_15570_21782.n2 0.653
R6036 a_15570_21782.n7 a_15570_21782.n6 0.653
R6037 a_15570_21782.n6 a_15570_21782.n5 0.341
R6038 a_15570_21782.n3 a_15570_21782.n1 0.032
R6039 a_20058_21029.t8 a_20058_21029.n2 404.877
R6040 a_20058_21029.n1 a_20058_21029.t5 210.902
R6041 a_20058_21029.n3 a_20058_21029.t8 136.949
R6042 a_20058_21029.n2 a_20058_21029.n1 107.801
R6043 a_20058_21029.n1 a_20058_21029.t6 80.333
R6044 a_20058_21029.n2 a_20058_21029.t7 80.333
R6045 a_20058_21029.n0 a_20058_21029.t3 17.4
R6046 a_20058_21029.n0 a_20058_21029.t4 17.4
R6047 a_20058_21029.n4 a_20058_21029.t2 15.032
R6048 a_20058_21029.n5 a_20058_21029.t1 14.282
R6049 a_20058_21029.t0 a_20058_21029.n5 14.282
R6050 a_20058_21029.n5 a_20058_21029.n4 1.65
R6051 a_20058_21029.n3 a_20058_21029.n0 0.657
R6052 a_20058_21029.n4 a_20058_21029.n3 0.614
R6053 a_18991_21663.t7 a_18991_21663.t4 800.071
R6054 a_18991_21663.n3 a_18991_21663.n2 672.95
R6055 a_18991_21663.n1 a_18991_21663.t5 285.109
R6056 a_18991_21663.n2 a_18991_21663.t7 193.602
R6057 a_18991_21663.n1 a_18991_21663.t6 160.666
R6058 a_18991_21663.n2 a_18991_21663.n1 91.507
R6059 a_18991_21663.n0 a_18991_21663.t1 28.57
R6060 a_18991_21663.n4 a_18991_21663.t2 28.565
R6061 a_18991_21663.t3 a_18991_21663.n4 28.565
R6062 a_18991_21663.n0 a_18991_21663.t0 17.638
R6063 a_18991_21663.n4 a_18991_21663.n3 0.693
R6064 a_18991_21663.n3 a_18991_21663.n0 0.597
R6065 a_10641_5411.n5 a_10641_5411.n4 501.28
R6066 a_10641_5411.t11 a_10641_5411.t7 437.233
R6067 a_10641_5411.t17 a_10641_5411.t15 415.315
R6068 a_10641_5411.t19 a_10641_5411.n2 313.873
R6069 a_10641_5411.n4 a_10641_5411.t13 294.986
R6070 a_10641_5411.n1 a_10641_5411.t4 272.288
R6071 a_10641_5411.n5 a_10641_5411.t14 236.01
R6072 a_10641_5411.n8 a_10641_5411.t11 216.627
R6073 a_10641_5411.n6 a_10641_5411.t17 216.111
R6074 a_10641_5411.n7 a_10641_5411.t5 214.686
R6075 a_10641_5411.t7 a_10641_5411.n7 214.686
R6076 a_10641_5411.n0 a_10641_5411.t16 214.335
R6077 a_10641_5411.t15 a_10641_5411.n0 214.335
R6078 a_10641_5411.n11 a_10641_5411.n10 192.754
R6079 a_10641_5411.n3 a_10641_5411.t19 190.152
R6080 a_10641_5411.n3 a_10641_5411.t8 190.152
R6081 a_10641_5411.n1 a_10641_5411.t9 160.666
R6082 a_10641_5411.n2 a_10641_5411.t10 160.666
R6083 a_10641_5411.n6 a_10641_5411.n5 148.428
R6084 a_10641_5411.n4 a_10641_5411.t18 110.859
R6085 a_10641_5411.n9 a_10641_5411.n8 102.569
R6086 a_10641_5411.n2 a_10641_5411.n1 96.129
R6087 a_10641_5411.n7 a_10641_5411.t12 80.333
R6088 a_10641_5411.n0 a_10641_5411.t6 80.333
R6089 a_10641_5411.t14 a_10641_5411.n3 80.333
R6090 a_10641_5411.n10 a_10641_5411.t3 28.568
R6091 a_10641_5411.n11 a_10641_5411.t2 28.565
R6092 a_10641_5411.t1 a_10641_5411.n11 28.565
R6093 a_10641_5411.n9 a_10641_5411.t0 18.523
R6094 a_10641_5411.n8 a_10641_5411.n6 2.923
R6095 a_10641_5411.n10 a_10641_5411.n9 1.167
R6096 a_14372_4127.t3 a_14372_4127.n7 16.058
R6097 a_14372_4127.n7 a_14372_4127.n5 0.575
R6098 a_14372_4127.n5 a_14372_4127.n9 0.2
R6099 a_14372_4127.n9 a_14372_4127.t7 16.058
R6100 a_14372_4127.n9 a_14372_4127.n8 0.999
R6101 a_14372_4127.n8 a_14372_4127.t8 14.282
R6102 a_14372_4127.n8 a_14372_4127.t6 14.282
R6103 a_14372_4127.n7 a_14372_4127.n6 0.999
R6104 a_14372_4127.n6 a_14372_4127.t5 14.282
R6105 a_14372_4127.n6 a_14372_4127.t4 14.282
R6106 a_14372_4127.n5 a_14372_4127.n3 0.227
R6107 a_14372_4127.n3 a_14372_4127.n4 1.511
R6108 a_14372_4127.n4 a_14372_4127.t9 14.282
R6109 a_14372_4127.n4 a_14372_4127.t11 14.282
R6110 a_14372_4127.n3 a_14372_4127.n0 0.669
R6111 a_14372_4127.n0 a_14372_4127.n1 0.001
R6112 a_14372_4127.n0 a_14372_4127.n2 267.767
R6113 a_14372_4127.n2 a_14372_4127.t1 14.282
R6114 a_14372_4127.n2 a_14372_4127.t0 14.282
R6115 a_14372_4127.n1 a_14372_4127.t10 14.282
R6116 a_14372_4127.n1 a_14372_4127.t2 14.282
R6117 a_13951_10690.n2 a_13951_10690.t6 318.922
R6118 a_13951_10690.n1 a_13951_10690.t7 273.935
R6119 a_13951_10690.n1 a_13951_10690.t5 273.935
R6120 a_13951_10690.n2 a_13951_10690.t4 269.116
R6121 a_13951_10690.n4 a_13951_10690.n0 193.227
R6122 a_13951_10690.t6 a_13951_10690.n1 179.142
R6123 a_13951_10690.n3 a_13951_10690.n2 106.999
R6124 a_13951_10690.t1 a_13951_10690.n4 28.568
R6125 a_13951_10690.n0 a_13951_10690.t3 28.565
R6126 a_13951_10690.n0 a_13951_10690.t2 28.565
R6127 a_13951_10690.n3 a_13951_10690.t0 18.149
R6128 a_13951_10690.n4 a_13951_10690.n3 3.726
R6129 a_14496_9265.t0 a_14496_9265.t1 380.209
R6130 a_14496_9997.t0 a_14496_9997.n0 14.282
R6131 a_14496_9997.n0 a_14496_9997.t1 14.282
R6132 a_14496_9997.n0 a_14496_9997.n16 90.436
R6133 a_14496_9997.n12 a_14496_9997.n15 50.575
R6134 a_14496_9997.n16 a_14496_9997.n12 74.302
R6135 a_14496_9997.n15 a_14496_9997.n14 157.665
R6136 a_14496_9997.n14 a_14496_9997.t6 8.7
R6137 a_14496_9997.n14 a_14496_9997.t7 8.7
R6138 a_14496_9997.n15 a_14496_9997.n13 122.999
R6139 a_14496_9997.n13 a_14496_9997.t3 14.282
R6140 a_14496_9997.n13 a_14496_9997.t4 14.282
R6141 a_14496_9997.n12 a_14496_9997.n11 90.416
R6142 a_14496_9997.n11 a_14496_9997.t5 14.282
R6143 a_14496_9997.n11 a_14496_9997.t2 14.282
R6144 a_14496_9997.n16 a_14496_9997.n1 216.635
R6145 a_14496_9997.n1 a_14496_9997.n3 16.411
R6146 a_14496_9997.n3 a_14496_9997.t13 198.921
R6147 a_14496_9997.t13 a_14496_9997.t21 415.315
R6148 a_14496_9997.t21 a_14496_9997.n10 214.335
R6149 a_14496_9997.n10 a_14496_9997.t23 80.333
R6150 a_14496_9997.n10 a_14496_9997.t8 214.335
R6151 a_14496_9997.n3 a_14496_9997.n9 861.987
R6152 a_14496_9997.n9 a_14496_9997.n4 560.726
R6153 a_14496_9997.n9 a_14496_9997.n8 65.07
R6154 a_14496_9997.n8 a_14496_9997.n7 6.615
R6155 a_14496_9997.n7 a_14496_9997.t18 93.989
R6156 a_14496_9997.n8 a_14496_9997.n6 97.816
R6157 a_14496_9997.n6 a_14496_9997.t19 80.333
R6158 a_14496_9997.n6 a_14496_9997.t9 394.151
R6159 a_14496_9997.t9 a_14496_9997.n5 269.523
R6160 a_14496_9997.n5 a_14496_9997.t10 160.666
R6161 a_14496_9997.n5 a_14496_9997.t11 269.523
R6162 a_14496_9997.n7 a_14496_9997.t17 198.043
R6163 a_14496_9997.n4 a_14496_9997.t20 294.653
R6164 a_14496_9997.n4 a_14496_9997.t12 111.663
R6165 a_14496_9997.n1 a_14496_9997.t15 217.716
R6166 a_14496_9997.t15 a_14496_9997.t22 415.315
R6167 a_14496_9997.t22 a_14496_9997.n2 214.335
R6168 a_14496_9997.n2 a_14496_9997.t14 80.333
R6169 a_14496_9997.n2 a_14496_9997.t16 214.335
R6170 a_9647_19525.t0 a_9647_19525.t1 17.4
R6171 a_11523_19541.n1 a_11523_19541.t7 318.922
R6172 a_11523_19541.n0 a_11523_19541.t6 274.739
R6173 a_11523_19541.n0 a_11523_19541.t4 274.739
R6174 a_11523_19541.n1 a_11523_19541.t5 269.116
R6175 a_11523_19541.t7 a_11523_19541.n0 179.946
R6176 a_11523_19541.n2 a_11523_19541.n1 105.178
R6177 a_11523_19541.n3 a_11523_19541.t2 29.444
R6178 a_11523_19541.t3 a_11523_19541.n4 28.565
R6179 a_11523_19541.n4 a_11523_19541.t1 28.565
R6180 a_11523_19541.n2 a_11523_19541.t0 18.145
R6181 a_11523_19541.n3 a_11523_19541.n2 2.878
R6182 a_11523_19541.n4 a_11523_19541.n3 0.764
R6183 a_12063_18848.n0 a_12063_18848.n1 0.001
R6184 a_12063_18848.n0 a_12063_18848.t9 14.282
R6185 a_12063_18848.t0 a_12063_18848.n0 14.282
R6186 a_12063_18848.n1 a_12063_18848.n9 267.767
R6187 a_12063_18848.n9 a_12063_18848.t11 14.282
R6188 a_12063_18848.n9 a_12063_18848.t10 14.282
R6189 a_12063_18848.n1 a_12063_18848.n7 0.669
R6190 a_12063_18848.n7 a_12063_18848.n8 1.511
R6191 a_12063_18848.n8 a_12063_18848.t1 14.282
R6192 a_12063_18848.n8 a_12063_18848.t2 14.282
R6193 a_12063_18848.n7 a_12063_18848.n6 0.227
R6194 a_12063_18848.n6 a_12063_18848.n3 0.2
R6195 a_12063_18848.n6 a_12063_18848.n5 0.575
R6196 a_12063_18848.n5 a_12063_18848.t6 16.058
R6197 a_12063_18848.n5 a_12063_18848.n4 0.999
R6198 a_12063_18848.n4 a_12063_18848.t8 14.282
R6199 a_12063_18848.n4 a_12063_18848.t7 14.282
R6200 a_12063_18848.n3 a_12063_18848.n2 0.999
R6201 a_12063_18848.n2 a_12063_18848.t5 14.282
R6202 a_12063_18848.n2 a_12063_18848.t3 14.282
R6203 a_12063_18848.n3 a_12063_18848.t4 16.058
R6204 a_12181_18848.n0 a_12181_18848.t6 14.282
R6205 a_12181_18848.t5 a_12181_18848.n0 14.282
R6206 a_12181_18848.n0 a_12181_18848.n8 122.747
R6207 a_12181_18848.n4 a_12181_18848.n6 74.302
R6208 a_12181_18848.n8 a_12181_18848.n4 50.575
R6209 a_12181_18848.n8 a_12181_18848.n7 157.665
R6210 a_12181_18848.n7 a_12181_18848.t0 8.7
R6211 a_12181_18848.n7 a_12181_18848.t4 8.7
R6212 a_12181_18848.n6 a_12181_18848.n5 90.436
R6213 a_12181_18848.n5 a_12181_18848.t2 14.282
R6214 a_12181_18848.n5 a_12181_18848.t1 14.282
R6215 a_12181_18848.n4 a_12181_18848.n3 90.416
R6216 a_12181_18848.n3 a_12181_18848.t3 14.282
R6217 a_12181_18848.n3 a_12181_18848.t7 14.282
R6218 a_12181_18848.n6 a_12181_18848.n1 294.955
R6219 a_12181_18848.t11 a_12181_18848.n2 160.666
R6220 a_12181_18848.n1 a_12181_18848.t11 867.393
R6221 a_12181_18848.n2 a_12181_18848.t9 287.241
R6222 a_12181_18848.n2 a_12181_18848.t10 287.241
R6223 a_12181_18848.n1 a_12181_18848.t8 545.094
R6224 a_12886_4101.n1 a_12886_4101.t4 318.922
R6225 a_12886_4101.n0 a_12886_4101.t5 274.739
R6226 a_12886_4101.n0 a_12886_4101.t6 274.739
R6227 a_12886_4101.n1 a_12886_4101.t7 269.116
R6228 a_12886_4101.t4 a_12886_4101.n0 179.946
R6229 a_12886_4101.n2 a_12886_4101.n1 107.263
R6230 a_12886_4101.n3 a_12886_4101.t3 29.444
R6231 a_12886_4101.t0 a_12886_4101.n4 28.565
R6232 a_12886_4101.n4 a_12886_4101.t2 28.565
R6233 a_12886_4101.n2 a_12886_4101.t1 18.145
R6234 a_12886_4101.n3 a_12886_4101.n2 2.878
R6235 a_12886_4101.n4 a_12886_4101.n3 0.764
R6236 a_12474_4127.n0 a_12474_4127.n9 1.511
R6237 a_12474_4127.n0 a_12474_4127.t1 14.282
R6238 a_12474_4127.t0 a_12474_4127.n0 14.282
R6239 a_12474_4127.n9 a_12474_4127.n5 0.227
R6240 a_12474_4127.n9 a_12474_4127.n6 0.669
R6241 a_12474_4127.n6 a_12474_4127.n7 0.001
R6242 a_12474_4127.n6 a_12474_4127.n8 267.767
R6243 a_12474_4127.n8 a_12474_4127.t7 14.282
R6244 a_12474_4127.n8 a_12474_4127.t8 14.282
R6245 a_12474_4127.n7 a_12474_4127.t2 14.282
R6246 a_12474_4127.n7 a_12474_4127.t6 14.282
R6247 a_12474_4127.n5 a_12474_4127.n2 0.575
R6248 a_12474_4127.n5 a_12474_4127.n4 0.2
R6249 a_12474_4127.n4 a_12474_4127.t3 16.058
R6250 a_12474_4127.n4 a_12474_4127.n3 0.999
R6251 a_12474_4127.n3 a_12474_4127.t4 14.282
R6252 a_12474_4127.n3 a_12474_4127.t5 14.282
R6253 a_12474_4127.n2 a_12474_4127.n1 0.999
R6254 a_12474_4127.n1 a_12474_4127.t9 14.282
R6255 a_12474_4127.n1 a_12474_4127.t11 14.282
R6256 a_12474_4127.n2 a_12474_4127.t10 16.058
R6257 a_12592_4127.n0 a_12592_4127.n12 122.999
R6258 a_12592_4127.n0 a_12592_4127.t5 14.282
R6259 a_12592_4127.t4 a_12592_4127.n0 14.282
R6260 a_12592_4127.n12 a_12592_4127.n10 50.575
R6261 a_12592_4127.n10 a_12592_4127.n8 74.302
R6262 a_12592_4127.n12 a_12592_4127.n11 157.665
R6263 a_12592_4127.n11 a_12592_4127.t7 8.7
R6264 a_12592_4127.n11 a_12592_4127.t0 8.7
R6265 a_12592_4127.n10 a_12592_4127.n9 90.416
R6266 a_12592_4127.n9 a_12592_4127.t6 14.282
R6267 a_12592_4127.n9 a_12592_4127.t2 14.282
R6268 a_12592_4127.n8 a_12592_4127.n7 90.436
R6269 a_12592_4127.n7 a_12592_4127.t3 14.282
R6270 a_12592_4127.n7 a_12592_4127.t1 14.282
R6271 a_12592_4127.n8 a_12592_4127.n1 342.688
R6272 a_12592_4127.n1 a_12592_4127.n6 126.566
R6273 a_12592_4127.n6 a_12592_4127.t15 294.653
R6274 a_12592_4127.n6 a_12592_4127.t8 111.663
R6275 a_12592_4127.n1 a_12592_4127.n5 552.333
R6276 a_12592_4127.n5 a_12592_4127.n4 6.615
R6277 a_12592_4127.n4 a_12592_4127.t10 93.989
R6278 a_12592_4127.n5 a_12592_4127.n3 97.816
R6279 a_12592_4127.n3 a_12592_4127.t14 80.333
R6280 a_12592_4127.n3 a_12592_4127.t9 394.151
R6281 a_12592_4127.t9 a_12592_4127.n2 269.523
R6282 a_12592_4127.n2 a_12592_4127.t13 160.666
R6283 a_12592_4127.n2 a_12592_4127.t11 269.523
R6284 a_12592_4127.n4 a_12592_4127.t12 198.043
R6285 a_5899_21662.t5 a_5899_21662.t6 800.071
R6286 a_5899_21662.n3 a_5899_21662.n2 672.95
R6287 a_5899_21662.n1 a_5899_21662.t7 285.109
R6288 a_5899_21662.n2 a_5899_21662.t5 193.602
R6289 a_5899_21662.n1 a_5899_21662.t4 160.666
R6290 a_5899_21662.n2 a_5899_21662.n1 91.507
R6291 a_5899_21662.t0 a_5899_21662.n4 28.57
R6292 a_5899_21662.n0 a_5899_21662.t2 28.565
R6293 a_5899_21662.n0 a_5899_21662.t3 28.565
R6294 a_5899_21662.n4 a_5899_21662.t1 17.638
R6295 a_5899_21662.n3 a_5899_21662.n0 0.693
R6296 a_5899_21662.n4 a_5899_21662.n3 0.597
R6297 a_5959_21688.n0 a_5959_21688.t5 14.282
R6298 a_5959_21688.n0 a_5959_21688.t4 14.282
R6299 a_5959_21688.n1 a_5959_21688.t2 14.282
R6300 a_5959_21688.n1 a_5959_21688.t0 14.282
R6301 a_5959_21688.t3 a_5959_21688.n3 14.282
R6302 a_5959_21688.n3 a_5959_21688.t1 14.282
R6303 a_5959_21688.n2 a_5959_21688.n0 2.546
R6304 a_5959_21688.n2 a_5959_21688.n1 2.367
R6305 a_5959_21688.n3 a_5959_21688.n2 0.001
R6306 a_10687_7087.n4 a_10687_7087.t7 214.335
R6307 a_10687_7087.t9 a_10687_7087.n4 214.335
R6308 a_10687_7087.n5 a_10687_7087.t9 143.851
R6309 a_10687_7087.n5 a_10687_7087.t10 135.658
R6310 a_10687_7087.n4 a_10687_7087.t8 80.333
R6311 a_10687_7087.n0 a_10687_7087.t5 28.565
R6312 a_10687_7087.n0 a_10687_7087.t6 28.565
R6313 a_10687_7087.n2 a_10687_7087.t1 28.565
R6314 a_10687_7087.n2 a_10687_7087.t3 28.565
R6315 a_10687_7087.n7 a_10687_7087.t2 28.565
R6316 a_10687_7087.t0 a_10687_7087.n7 28.565
R6317 a_10687_7087.n1 a_10687_7087.t4 9.714
R6318 a_10687_7087.n1 a_10687_7087.n0 1.003
R6319 a_10687_7087.n6 a_10687_7087.n3 0.833
R6320 a_10687_7087.n3 a_10687_7087.n2 0.653
R6321 a_10687_7087.n7 a_10687_7087.n6 0.653
R6322 a_10687_7087.n3 a_10687_7087.n1 0.341
R6323 a_10687_7087.n6 a_10687_7087.n5 0.032
R6324 a_11277_6650.t7 a_11277_6650.t4 800.071
R6325 a_11277_6650.n3 a_11277_6650.n2 659.097
R6326 a_11277_6650.n1 a_11277_6650.t5 285.109
R6327 a_11277_6650.n2 a_11277_6650.t7 193.602
R6328 a_11277_6650.n4 a_11277_6650.n0 192.754
R6329 a_11277_6650.n1 a_11277_6650.t6 160.666
R6330 a_11277_6650.n2 a_11277_6650.n1 91.507
R6331 a_11277_6650.t3 a_11277_6650.n4 28.568
R6332 a_11277_6650.n0 a_11277_6650.t2 28.565
R6333 a_11277_6650.n0 a_11277_6650.t1 28.565
R6334 a_11277_6650.n3 a_11277_6650.t0 19.061
R6335 a_11277_6650.n4 a_11277_6650.n3 1.005
R6336 a_12470_24163.n4 a_12470_24163.t9 214.335
R6337 a_12470_24163.t7 a_12470_24163.n4 214.335
R6338 a_12470_24163.n5 a_12470_24163.t7 143.851
R6339 a_12470_24163.n5 a_12470_24163.t10 135.658
R6340 a_12470_24163.n4 a_12470_24163.t8 80.333
R6341 a_12470_24163.n0 a_12470_24163.t5 28.565
R6342 a_12470_24163.n0 a_12470_24163.t3 28.565
R6343 a_12470_24163.n2 a_12470_24163.t1 28.565
R6344 a_12470_24163.n2 a_12470_24163.t6 28.565
R6345 a_12470_24163.t0 a_12470_24163.n7 28.565
R6346 a_12470_24163.n7 a_12470_24163.t2 28.565
R6347 a_12470_24163.n1 a_12470_24163.t4 9.714
R6348 a_12470_24163.n1 a_12470_24163.n0 1.003
R6349 a_12470_24163.n6 a_12470_24163.n3 0.833
R6350 a_12470_24163.n3 a_12470_24163.n2 0.653
R6351 a_12470_24163.n7 a_12470_24163.n6 0.653
R6352 a_12470_24163.n3 a_12470_24163.n1 0.341
R6353 a_12470_24163.n6 a_12470_24163.n5 0.032
R6354 a_13060_23726.t5 a_13060_23726.t4 574.43
R6355 a_13060_23726.n0 a_13060_23726.t7 285.109
R6356 a_13060_23726.n2 a_13060_23726.n1 197.217
R6357 a_13060_23726.n4 a_13060_23726.n3 192.754
R6358 a_13060_23726.n0 a_13060_23726.t6 160.666
R6359 a_13060_23726.n1 a_13060_23726.t5 160.666
R6360 a_13060_23726.n1 a_13060_23726.n0 114.829
R6361 a_13060_23726.n3 a_13060_23726.t1 28.568
R6362 a_13060_23726.n4 a_13060_23726.t2 28.565
R6363 a_13060_23726.t3 a_13060_23726.n4 28.565
R6364 a_13060_23726.n2 a_13060_23726.t0 18.838
R6365 a_13060_23726.n3 a_13060_23726.n2 1.129
R6366 a_7308_25153.n2 a_7308_25153.t5 318.922
R6367 a_7308_25153.n1 a_7308_25153.t4 273.935
R6368 a_7308_25153.n1 a_7308_25153.t6 273.935
R6369 a_7308_25153.n2 a_7308_25153.t7 269.116
R6370 a_7308_25153.n4 a_7308_25153.n0 193.227
R6371 a_7308_25153.t5 a_7308_25153.n1 179.142
R6372 a_7308_25153.n3 a_7308_25153.n2 106.999
R6373 a_7308_25153.t3 a_7308_25153.n4 28.568
R6374 a_7308_25153.n0 a_7308_25153.t1 28.565
R6375 a_7308_25153.n0 a_7308_25153.t2 28.565
R6376 a_7308_25153.n3 a_7308_25153.t0 18.149
R6377 a_7308_25153.n4 a_7308_25153.n3 3.726
R6378 a_7853_24460.n0 a_7853_24460.t1 14.282
R6379 a_7853_24460.t5 a_7853_24460.n0 14.282
R6380 a_7853_24460.n0 a_7853_24460.n12 90.416
R6381 a_7853_24460.n12 a_7853_24460.n11 50.575
R6382 a_7853_24460.n12 a_7853_24460.n8 74.302
R6383 a_7853_24460.n11 a_7853_24460.n10 157.665
R6384 a_7853_24460.n10 a_7853_24460.t4 8.7
R6385 a_7853_24460.n10 a_7853_24460.t0 8.7
R6386 a_7853_24460.n11 a_7853_24460.n9 122.999
R6387 a_7853_24460.n9 a_7853_24460.t3 14.282
R6388 a_7853_24460.n9 a_7853_24460.t2 14.282
R6389 a_7853_24460.n8 a_7853_24460.n7 90.436
R6390 a_7853_24460.n7 a_7853_24460.t6 14.282
R6391 a_7853_24460.n7 a_7853_24460.t7 14.282
R6392 a_7853_24460.n8 a_7853_24460.n1 342.688
R6393 a_7853_24460.n1 a_7853_24460.n6 126.566
R6394 a_7853_24460.n6 a_7853_24460.t12 294.653
R6395 a_7853_24460.n6 a_7853_24460.t10 111.663
R6396 a_7853_24460.n1 a_7853_24460.n5 552.333
R6397 a_7853_24460.n5 a_7853_24460.n4 6.615
R6398 a_7853_24460.n4 a_7853_24460.t9 93.989
R6399 a_7853_24460.n5 a_7853_24460.n3 97.816
R6400 a_7853_24460.n3 a_7853_24460.t11 80.333
R6401 a_7853_24460.n3 a_7853_24460.t13 394.151
R6402 a_7853_24460.t13 a_7853_24460.n2 269.523
R6403 a_7853_24460.n2 a_7853_24460.t14 160.666
R6404 a_7853_24460.n2 a_7853_24460.t15 269.523
R6405 a_7853_24460.n4 a_7853_24460.t8 198.043
R6406 a_7395_21658.t6 a_7395_21658.t7 574.43
R6407 a_7395_21658.n0 a_7395_21658.t4 285.109
R6408 a_7395_21658.n2 a_7395_21658.n1 197.215
R6409 a_7395_21658.n4 a_7395_21658.n3 192.754
R6410 a_7395_21658.n0 a_7395_21658.t5 160.666
R6411 a_7395_21658.n1 a_7395_21658.t6 160.666
R6412 a_7395_21658.n1 a_7395_21658.n0 114.829
R6413 a_7395_21658.n3 a_7395_21658.t3 28.568
R6414 a_7395_21658.n4 a_7395_21658.t2 28.565
R6415 a_7395_21658.t0 a_7395_21658.n4 28.565
R6416 a_7395_21658.n2 a_7395_21658.t1 18.838
R6417 a_7395_21658.n3 a_7395_21658.n2 1.129
R6418 a_7101_21684.n0 a_7101_21684.t1 14.282
R6419 a_7101_21684.n0 a_7101_21684.t2 14.282
R6420 a_7101_21684.n1 a_7101_21684.t4 14.282
R6421 a_7101_21684.n1 a_7101_21684.t5 14.282
R6422 a_7101_21684.n3 a_7101_21684.t3 14.282
R6423 a_7101_21684.t0 a_7101_21684.n3 14.282
R6424 a_7101_21684.n2 a_7101_21684.n0 2.546
R6425 a_7101_21684.n2 a_7101_21684.n1 2.367
R6426 a_7101_21684.n3 a_7101_21684.n2 0.001
R6427 a_6966_21028.t6 a_6966_21028.n2 404.877
R6428 a_6966_21028.n1 a_6966_21028.t8 210.902
R6429 a_6966_21028.n3 a_6966_21028.t6 136.949
R6430 a_6966_21028.n2 a_6966_21028.n1 107.801
R6431 a_6966_21028.n1 a_6966_21028.t7 80.333
R6432 a_6966_21028.n2 a_6966_21028.t5 80.333
R6433 a_6966_21028.n0 a_6966_21028.t0 17.4
R6434 a_6966_21028.n0 a_6966_21028.t4 17.4
R6435 a_6966_21028.n4 a_6966_21028.t1 15.032
R6436 a_6966_21028.n5 a_6966_21028.t2 14.282
R6437 a_6966_21028.t3 a_6966_21028.n5 14.282
R6438 a_6966_21028.n5 a_6966_21028.n4 1.65
R6439 a_6966_21028.n3 a_6966_21028.n0 0.657
R6440 a_6966_21028.n4 a_6966_21028.n3 0.614
R6441 a_4150_5439.n0 a_4150_5439.t9 214.335
R6442 a_4150_5439.t7 a_4150_5439.n0 214.335
R6443 a_4150_5439.n1 a_4150_5439.t7 143.851
R6444 a_4150_5439.n1 a_4150_5439.t10 135.658
R6445 a_4150_5439.n0 a_4150_5439.t8 80.333
R6446 a_4150_5439.n2 a_4150_5439.t5 28.565
R6447 a_4150_5439.n2 a_4150_5439.t6 28.565
R6448 a_4150_5439.n4 a_4150_5439.t4 28.565
R6449 a_4150_5439.n4 a_4150_5439.t2 28.565
R6450 a_4150_5439.t1 a_4150_5439.n7 28.565
R6451 a_4150_5439.n7 a_4150_5439.t3 28.565
R6452 a_4150_5439.n6 a_4150_5439.t0 9.714
R6453 a_4150_5439.n7 a_4150_5439.n6 1.003
R6454 a_4150_5439.n5 a_4150_5439.n3 0.833
R6455 a_4150_5439.n3 a_4150_5439.n2 0.653
R6456 a_4150_5439.n5 a_4150_5439.n4 0.653
R6457 a_4150_5439.n6 a_4150_5439.n5 0.341
R6458 a_4150_5439.n3 a_4150_5439.n1 0.032
R6459 a_4740_5002.t4 a_4740_5002.t6 574.43
R6460 a_4740_5002.n0 a_4740_5002.t5 285.109
R6461 a_4740_5002.n2 a_4740_5002.n1 211.136
R6462 a_4740_5002.n4 a_4740_5002.n3 192.754
R6463 a_4740_5002.n0 a_4740_5002.t7 160.666
R6464 a_4740_5002.n1 a_4740_5002.t4 160.666
R6465 a_4740_5002.n1 a_4740_5002.n0 114.829
R6466 a_4740_5002.n3 a_4740_5002.t1 28.568
R6467 a_4740_5002.n4 a_4740_5002.t2 28.565
R6468 a_4740_5002.t3 a_4740_5002.n4 28.565
R6469 a_4740_5002.n2 a_4740_5002.t0 19.084
R6470 a_4740_5002.n3 a_4740_5002.n2 1.051
R6471 a_6041_4129.t0 a_6041_4129.n0 14.282
R6472 a_6041_4129.n0 a_6041_4129.t2 14.282
R6473 a_6041_4129.n0 a_6041_4129.n12 90.436
R6474 a_6041_4129.n8 a_6041_4129.n11 50.575
R6475 a_6041_4129.n12 a_6041_4129.n8 74.302
R6476 a_6041_4129.n11 a_6041_4129.n10 157.665
R6477 a_6041_4129.n10 a_6041_4129.t3 8.7
R6478 a_6041_4129.n10 a_6041_4129.t7 8.7
R6479 a_6041_4129.n11 a_6041_4129.n9 122.999
R6480 a_6041_4129.n9 a_6041_4129.t5 14.282
R6481 a_6041_4129.n9 a_6041_4129.t4 14.282
R6482 a_6041_4129.n8 a_6041_4129.n7 90.416
R6483 a_6041_4129.n7 a_6041_4129.t6 14.282
R6484 a_6041_4129.n7 a_6041_4129.t1 14.282
R6485 a_6041_4129.n12 a_6041_4129.n1 342.688
R6486 a_6041_4129.n1 a_6041_4129.n6 126.566
R6487 a_6041_4129.n6 a_6041_4129.t11 294.653
R6488 a_6041_4129.n6 a_6041_4129.t12 111.663
R6489 a_6041_4129.n1 a_6041_4129.n5 552.333
R6490 a_6041_4129.n5 a_6041_4129.n4 6.615
R6491 a_6041_4129.n4 a_6041_4129.t13 93.989
R6492 a_6041_4129.n5 a_6041_4129.n3 97.816
R6493 a_6041_4129.n3 a_6041_4129.t8 80.333
R6494 a_6041_4129.n3 a_6041_4129.t9 394.151
R6495 a_6041_4129.t9 a_6041_4129.n2 269.523
R6496 a_6041_4129.n2 a_6041_4129.t10 160.666
R6497 a_6041_4129.n2 a_6041_4129.t15 269.523
R6498 a_6041_4129.n4 a_6041_4129.t14 198.043
R6499 a_7394_4822.n1 a_7394_4822.t7 318.922
R6500 a_7394_4822.n0 a_7394_4822.t4 273.935
R6501 a_7394_4822.n0 a_7394_4822.t5 273.935
R6502 a_7394_4822.n1 a_7394_4822.t6 269.116
R6503 a_7394_4822.n4 a_7394_4822.n3 193.227
R6504 a_7394_4822.t7 a_7394_4822.n0 179.142
R6505 a_7394_4822.n2 a_7394_4822.n1 106.999
R6506 a_7394_4822.n3 a_7394_4822.t1 28.568
R6507 a_7394_4822.t3 a_7394_4822.n4 28.565
R6508 a_7394_4822.n4 a_7394_4822.t2 28.565
R6509 a_7394_4822.n2 a_7394_4822.t0 18.149
R6510 a_7394_4822.n3 a_7394_4822.n2 3.726
R6511 a_5962_25770.n0 a_5962_25770.t10 214.335
R6512 a_5962_25770.t8 a_5962_25770.n0 214.335
R6513 a_5962_25770.n1 a_5962_25770.t8 143.851
R6514 a_5962_25770.n1 a_5962_25770.t7 135.658
R6515 a_5962_25770.n0 a_5962_25770.t9 80.333
R6516 a_5962_25770.n2 a_5962_25770.t0 28.565
R6517 a_5962_25770.n2 a_5962_25770.t1 28.565
R6518 a_5962_25770.n4 a_5962_25770.t2 28.565
R6519 a_5962_25770.n4 a_5962_25770.t5 28.565
R6520 a_5962_25770.n7 a_5962_25770.t6 28.565
R6521 a_5962_25770.t3 a_5962_25770.n7 28.565
R6522 a_5962_25770.n6 a_5962_25770.t4 9.714
R6523 a_5962_25770.n7 a_5962_25770.n6 1.003
R6524 a_5962_25770.n5 a_5962_25770.n3 0.833
R6525 a_5962_25770.n3 a_5962_25770.n2 0.653
R6526 a_5962_25770.n5 a_5962_25770.n4 0.653
R6527 a_5962_25770.n6 a_5962_25770.n5 0.341
R6528 a_5962_25770.n3 a_5962_25770.n1 0.032
R6529 a_6552_25333.t5 a_6552_25333.t4 574.43
R6530 a_6552_25333.n0 a_6552_25333.t7 285.109
R6531 a_6552_25333.n2 a_6552_25333.n1 211.136
R6532 a_6552_25333.n4 a_6552_25333.n3 192.754
R6533 a_6552_25333.n0 a_6552_25333.t6 160.666
R6534 a_6552_25333.n1 a_6552_25333.t5 160.666
R6535 a_6552_25333.n1 a_6552_25333.n0 114.829
R6536 a_6552_25333.n3 a_6552_25333.t1 28.568
R6537 a_6552_25333.n4 a_6552_25333.t2 28.565
R6538 a_6552_25333.t3 a_6552_25333.n4 28.565
R6539 a_6552_25333.n2 a_6552_25333.t0 19.084
R6540 a_6552_25333.n3 a_6552_25333.n2 1.051
R6541 a_17361_11239.n4 a_17361_11239.t9 214.335
R6542 a_17361_11239.t7 a_17361_11239.n4 214.335
R6543 a_17361_11239.n5 a_17361_11239.t7 143.851
R6544 a_17361_11239.n5 a_17361_11239.t10 135.658
R6545 a_17361_11239.n4 a_17361_11239.t8 80.333
R6546 a_17361_11239.n0 a_17361_11239.t5 28.565
R6547 a_17361_11239.n0 a_17361_11239.t6 28.565
R6548 a_17361_11239.n2 a_17361_11239.t1 28.565
R6549 a_17361_11239.n2 a_17361_11239.t4 28.565
R6550 a_17361_11239.t2 a_17361_11239.n7 28.565
R6551 a_17361_11239.n7 a_17361_11239.t0 28.565
R6552 a_17361_11239.n1 a_17361_11239.t3 9.714
R6553 a_17361_11239.n1 a_17361_11239.n0 1.003
R6554 a_17361_11239.n6 a_17361_11239.n3 0.833
R6555 a_17361_11239.n3 a_17361_11239.n2 0.653
R6556 a_17361_11239.n7 a_17361_11239.n6 0.653
R6557 a_17361_11239.n3 a_17361_11239.n1 0.341
R6558 a_17361_11239.n6 a_17361_11239.n5 0.032
R6559 a_4145_3835.n0 a_4145_3835.t10 214.335
R6560 a_4145_3835.t9 a_4145_3835.n0 214.335
R6561 a_4145_3835.n1 a_4145_3835.t9 143.851
R6562 a_4145_3835.n1 a_4145_3835.t7 135.658
R6563 a_4145_3835.n0 a_4145_3835.t8 80.333
R6564 a_4145_3835.n2 a_4145_3835.t1 28.565
R6565 a_4145_3835.n2 a_4145_3835.t2 28.565
R6566 a_4145_3835.n4 a_4145_3835.t3 28.565
R6567 a_4145_3835.n4 a_4145_3835.t5 28.565
R6568 a_4145_3835.t0 a_4145_3835.n7 28.565
R6569 a_4145_3835.n7 a_4145_3835.t4 28.565
R6570 a_4145_3835.n6 a_4145_3835.t6 9.714
R6571 a_4145_3835.n7 a_4145_3835.n6 1.003
R6572 a_4145_3835.n5 a_4145_3835.n3 0.833
R6573 a_4145_3835.n3 a_4145_3835.n2 0.653
R6574 a_4145_3835.n5 a_4145_3835.n4 0.653
R6575 a_4145_3835.n6 a_4145_3835.n5 0.341
R6576 a_4145_3835.n3 a_4145_3835.n1 0.032
R6577 a_4735_3398.t5 a_4735_3398.t6 574.43
R6578 a_4735_3398.n0 a_4735_3398.t7 285.109
R6579 a_4735_3398.n2 a_4735_3398.n1 197.217
R6580 a_4735_3398.n4 a_4735_3398.n3 192.754
R6581 a_4735_3398.n0 a_4735_3398.t4 160.666
R6582 a_4735_3398.n1 a_4735_3398.t5 160.666
R6583 a_4735_3398.n1 a_4735_3398.n0 114.829
R6584 a_4735_3398.n3 a_4735_3398.t1 28.568
R6585 a_4735_3398.t3 a_4735_3398.n4 28.565
R6586 a_4735_3398.n4 a_4735_3398.t2 28.565
R6587 a_4735_3398.n2 a_4735_3398.t0 18.838
R6588 a_4735_3398.n3 a_4735_3398.n2 1.129
R6589 a_23918_5413.n5 a_23918_5413.n4 501.28
R6590 a_23918_5413.t14 a_23918_5413.t10 437.233
R6591 a_23918_5413.t4 a_23918_5413.t11 415.315
R6592 a_23918_5413.t19 a_23918_5413.n2 313.873
R6593 a_23918_5413.n4 a_23918_5413.t18 294.986
R6594 a_23918_5413.n1 a_23918_5413.t6 272.288
R6595 a_23918_5413.n5 a_23918_5413.t7 236.01
R6596 a_23918_5413.n9 a_23918_5413.t14 216.627
R6597 a_23918_5413.n7 a_23918_5413.t4 216.069
R6598 a_23918_5413.n8 a_23918_5413.t15 214.686
R6599 a_23918_5413.t10 a_23918_5413.n8 214.686
R6600 a_23918_5413.n6 a_23918_5413.t13 214.335
R6601 a_23918_5413.t11 a_23918_5413.n6 214.335
R6602 a_23918_5413.n11 a_23918_5413.n0 192.754
R6603 a_23918_5413.n3 a_23918_5413.t19 190.152
R6604 a_23918_5413.n3 a_23918_5413.t5 190.152
R6605 a_23918_5413.n1 a_23918_5413.t12 160.666
R6606 a_23918_5413.n2 a_23918_5413.t9 160.666
R6607 a_23918_5413.n7 a_23918_5413.n5 148.384
R6608 a_23918_5413.n4 a_23918_5413.t17 110.859
R6609 a_23918_5413.n2 a_23918_5413.n1 96.129
R6610 a_23918_5413.n8 a_23918_5413.t16 80.333
R6611 a_23918_5413.n6 a_23918_5413.t8 80.333
R6612 a_23918_5413.t7 a_23918_5413.n3 80.333
R6613 a_23918_5413.n10 a_23918_5413.n9 47.31
R6614 a_23918_5413.t0 a_23918_5413.n11 28.568
R6615 a_23918_5413.n0 a_23918_5413.t2 28.565
R6616 a_23918_5413.n0 a_23918_5413.t3 28.565
R6617 a_23918_5413.n10 a_23918_5413.t1 18.466
R6618 a_23918_5413.n9 a_23918_5413.n7 2.697
R6619 a_23918_5413.n11 a_23918_5413.n10 1.161
R6620 a_24210_3198.t0 a_24210_3198.t1 17.4
R6621 a_n3604_15973.n1 a_n3604_15973.t4 318.119
R6622 a_n3604_15973.n1 a_n3604_15973.t5 269.919
R6623 a_n3604_15973.n0 a_n3604_15973.t6 267.256
R6624 a_n3604_15973.n0 a_n3604_15973.t7 267.256
R6625 a_n3604_15973.n4 a_n3604_15973.n3 193.227
R6626 a_n3604_15973.t4 a_n3604_15973.n0 160.666
R6627 a_n3604_15973.n2 a_n3604_15973.n1 106.999
R6628 a_n3604_15973.n3 a_n3604_15973.t3 28.568
R6629 a_n3604_15973.n4 a_n3604_15973.t2 28.565
R6630 a_n3604_15973.t0 a_n3604_15973.n4 28.565
R6631 a_n3604_15973.n2 a_n3604_15973.t1 18.149
R6632 a_n3604_15973.n3 a_n3604_15973.n2 3.726
R6633 a_n3804_15135.t3 a_n3804_15135.n0 14.282
R6634 a_n3804_15135.n0 a_n3804_15135.t4 14.282
R6635 a_n3804_15135.n0 a_n3804_15135.n9 0.999
R6636 a_n3804_15135.n9 a_n3804_15135.n6 0.2
R6637 a_n3804_15135.n6 a_n3804_15135.n8 0.575
R6638 a_n3804_15135.n9 a_n3804_15135.t5 16.058
R6639 a_n3804_15135.n8 a_n3804_15135.n7 0.999
R6640 a_n3804_15135.n7 a_n3804_15135.t0 14.282
R6641 a_n3804_15135.n7 a_n3804_15135.t2 14.282
R6642 a_n3804_15135.n8 a_n3804_15135.t1 16.058
R6643 a_n3804_15135.n6 a_n3804_15135.n4 0.227
R6644 a_n3804_15135.n4 a_n3804_15135.n5 1.511
R6645 a_n3804_15135.n5 a_n3804_15135.t11 14.282
R6646 a_n3804_15135.n5 a_n3804_15135.t9 14.282
R6647 a_n3804_15135.n4 a_n3804_15135.n1 0.669
R6648 a_n3804_15135.n1 a_n3804_15135.n2 0.001
R6649 a_n3804_15135.n1 a_n3804_15135.n3 267.767
R6650 a_n3804_15135.n3 a_n3804_15135.t8 14.282
R6651 a_n3804_15135.n3 a_n3804_15135.t6 14.282
R6652 a_n3804_15135.n2 a_n3804_15135.t7 14.282
R6653 a_n3804_15135.n2 a_n3804_15135.t10 14.282
R6654 a_18055_19249.n6 a_18055_19249.n5 501.28
R6655 a_18055_19249.t18 a_18055_19249.t17 437.233
R6656 a_18055_19249.t8 a_18055_19249.t12 415.315
R6657 a_18055_19249.t16 a_18055_19249.n3 313.873
R6658 a_18055_19249.n5 a_18055_19249.t13 294.986
R6659 a_18055_19249.n2 a_18055_19249.t4 272.288
R6660 a_18055_19249.n6 a_18055_19249.t15 236.009
R6661 a_18055_19249.n9 a_18055_19249.t18 216.627
R6662 a_18055_19249.n7 a_18055_19249.t8 216.111
R6663 a_18055_19249.n8 a_18055_19249.t5 214.686
R6664 a_18055_19249.t17 a_18055_19249.n8 214.686
R6665 a_18055_19249.n1 a_18055_19249.t10 214.335
R6666 a_18055_19249.t12 a_18055_19249.n1 214.335
R6667 a_18055_19249.n4 a_18055_19249.t14 190.152
R6668 a_18055_19249.n4 a_18055_19249.t16 190.152
R6669 a_18055_19249.n2 a_18055_19249.t19 160.666
R6670 a_18055_19249.n3 a_18055_19249.t9 160.666
R6671 a_18055_19249.n7 a_18055_19249.n6 148.428
R6672 a_18055_19249.n5 a_18055_19249.t7 110.859
R6673 a_18055_19249.n3 a_18055_19249.n2 96.129
R6674 a_18055_19249.n8 a_18055_19249.t6 80.333
R6675 a_18055_19249.n1 a_18055_19249.t11 80.333
R6676 a_18055_19249.t15 a_18055_19249.n4 80.333
R6677 a_18055_19249.n0 a_18055_19249.t2 28.57
R6678 a_18055_19249.n11 a_18055_19249.t1 28.565
R6679 a_18055_19249.t0 a_18055_19249.n11 28.565
R6680 a_18055_19249.n0 a_18055_19249.t3 17.638
R6681 a_18055_19249.n10 a_18055_19249.n9 5.55
R6682 a_18055_19249.n9 a_18055_19249.n7 2.923
R6683 a_18055_19249.n11 a_18055_19249.n10 0.693
R6684 a_18055_19249.n10 a_18055_19249.n0 0.597
R6685 a_18597_18853.n0 a_18597_18853.t2 14.282
R6686 a_18597_18853.t0 a_18597_18853.n0 14.282
R6687 a_18597_18853.n0 a_18597_18853.n9 0.999
R6688 a_18597_18853.n9 a_18597_18853.n6 0.2
R6689 a_18597_18853.n6 a_18597_18853.n8 0.575
R6690 a_18597_18853.n8 a_18597_18853.t1 16.058
R6691 a_18597_18853.n8 a_18597_18853.n7 0.999
R6692 a_18597_18853.n7 a_18597_18853.t11 14.282
R6693 a_18597_18853.n7 a_18597_18853.t3 14.282
R6694 a_18597_18853.n9 a_18597_18853.t7 16.058
R6695 a_18597_18853.n6 a_18597_18853.n4 0.227
R6696 a_18597_18853.n4 a_18597_18853.n5 1.511
R6697 a_18597_18853.n5 a_18597_18853.t10 14.282
R6698 a_18597_18853.n5 a_18597_18853.t9 14.282
R6699 a_18597_18853.n4 a_18597_18853.n1 0.669
R6700 a_18597_18853.n1 a_18597_18853.n2 0.001
R6701 a_18597_18853.n1 a_18597_18853.n3 267.767
R6702 a_18597_18853.n3 a_18597_18853.t5 14.282
R6703 a_18597_18853.n3 a_18597_18853.t4 14.282
R6704 a_18597_18853.n2 a_18597_18853.t6 14.282
R6705 a_18597_18853.n2 a_18597_18853.t8 14.282
R6706 A[5].n6 A[5].t9 3756.03
R6707 A[5].n16 A[5].n6 2196.31
R6708 A[5].n11 A[5].n10 535.449
R6709 A[5].t11 A[5].t12 437.233
R6710 A[5].t9 A[5].t31 437.233
R6711 A[5].t19 A[5].t22 437.233
R6712 A[5].t28 A[5].t5 437.233
R6713 A[5].t14 A[5].t20 415.315
R6714 A[5].t30 A[5].t15 415.315
R6715 A[5].t10 A[5].n8 313.873
R6716 A[5].n10 A[5].t7 294.986
R6717 A[5].n7 A[5].t4 272.288
R6718 A[5].n5 A[5].t30 256.298
R6719 A[5].n11 A[5].t25 245.184
R6720 A[5].n3 A[5].t11 219.994
R6721 A[5].n13 A[5].t28 218.627
R6722 A[5].n3 A[5].t14 217.552
R6723 A[5].n15 A[5].t19 217.023
R6724 A[5].n1 A[5].t8 214.686
R6725 A[5].t12 A[5].n1 214.686
R6726 A[5].n0 A[5].t27 214.686
R6727 A[5].t31 A[5].n0 214.686
R6728 A[5].n14 A[5].t2 214.686
R6729 A[5].t22 A[5].n14 214.686
R6730 A[5].n12 A[5].t13 214.686
R6731 A[5].t5 A[5].n12 214.686
R6732 A[5].n2 A[5].t1 214.335
R6733 A[5].t20 A[5].n2 214.335
R6734 A[5].n4 A[5].t16 214.335
R6735 A[5].t15 A[5].n4 214.335
R6736 A[5].n9 A[5].t24 190.152
R6737 A[5].n9 A[5].t10 190.152
R6738 A[5].n7 A[5].t3 160.666
R6739 A[5].n8 A[5].t18 160.666
R6740 A[5].n10 A[5].t17 110.859
R6741 A[5].n8 A[5].n7 96.129
R6742 A[5].n2 A[5].t0 80.333
R6743 A[5].n1 A[5].t21 80.333
R6744 A[5].n4 A[5].t26 80.333
R6745 A[5].n0 A[5].t29 80.333
R6746 A[5].n14 A[5].t23 80.333
R6747 A[5].t25 A[5].n9 80.333
R6748 A[5].n12 A[5].t6 80.333
R6749 A[5].n16 A[5].n15 45.674
R6750 A[5].n13 A[5].n11 14.9
R6751 A[5] A[5].n16 2.638
R6752 A[5].n15 A[5].n13 2.599
R6753 A[5].n5 A[5].n3 0.426
R6754 A[5].n6 A[5].n5 0.09
R6755 a_1246_10551.n2 a_1246_10551.t9 214.335
R6756 a_1246_10551.t7 a_1246_10551.n2 214.335
R6757 a_1246_10551.n3 a_1246_10551.t7 143.851
R6758 a_1246_10551.n3 a_1246_10551.t10 135.658
R6759 a_1246_10551.n2 a_1246_10551.t8 80.333
R6760 a_1246_10551.n4 a_1246_10551.t3 28.565
R6761 a_1246_10551.n4 a_1246_10551.t4 28.565
R6762 a_1246_10551.n0 a_1246_10551.t5 28.565
R6763 a_1246_10551.n0 a_1246_10551.t6 28.565
R6764 a_1246_10551.n7 a_1246_10551.t2 28.565
R6765 a_1246_10551.t0 a_1246_10551.n7 28.565
R6766 a_1246_10551.n1 a_1246_10551.t1 9.714
R6767 a_1246_10551.n1 a_1246_10551.n0 1.003
R6768 a_1246_10551.n6 a_1246_10551.n5 0.833
R6769 a_1246_10551.n5 a_1246_10551.n4 0.653
R6770 a_1246_10551.n7 a_1246_10551.n6 0.653
R6771 a_1246_10551.n6 a_1246_10551.n1 0.341
R6772 a_1246_10551.n5 a_1246_10551.n3 0.032
R6773 a_4965_19545.n1 a_4965_19545.t6 318.922
R6774 a_4965_19545.n0 a_4965_19545.t5 274.739
R6775 a_4965_19545.n0 a_4965_19545.t7 274.739
R6776 a_4965_19545.n1 a_4965_19545.t4 269.116
R6777 a_4965_19545.t6 a_4965_19545.n0 179.946
R6778 a_4965_19545.n2 a_4965_19545.n1 105.178
R6779 a_4965_19545.t3 a_4965_19545.n4 29.444
R6780 a_4965_19545.n3 a_4965_19545.t1 28.565
R6781 a_4965_19545.n3 a_4965_19545.t2 28.565
R6782 a_4965_19545.n2 a_4965_19545.t0 18.145
R6783 a_4965_19545.n4 a_4965_19545.n2 2.878
R6784 a_4965_19545.n4 a_4965_19545.n3 0.764
R6785 a_5623_18120.t0 a_5623_18120.t1 380.209
R6786 a_14507_1337.n0 a_14507_1337.t9 214.335
R6787 a_14507_1337.t7 a_14507_1337.n0 214.335
R6788 a_14507_1337.n1 a_14507_1337.t7 143.85
R6789 a_14507_1337.n1 a_14507_1337.t8 135.66
R6790 a_14507_1337.n0 a_14507_1337.t10 80.333
R6791 a_14507_1337.n2 a_14507_1337.t1 28.565
R6792 a_14507_1337.n2 a_14507_1337.t2 28.565
R6793 a_14507_1337.n4 a_14507_1337.t0 28.565
R6794 a_14507_1337.n4 a_14507_1337.t4 28.565
R6795 a_14507_1337.n7 a_14507_1337.t5 28.565
R6796 a_14507_1337.t3 a_14507_1337.n7 28.565
R6797 a_14507_1337.n6 a_14507_1337.t6 9.714
R6798 a_14507_1337.n7 a_14507_1337.n6 1.003
R6799 a_14507_1337.n5 a_14507_1337.n3 0.836
R6800 a_14507_1337.n5 a_14507_1337.n4 0.653
R6801 a_14507_1337.n3 a_14507_1337.n2 0.65
R6802 a_14507_1337.n6 a_14507_1337.n5 0.341
R6803 a_14507_1337.n3 a_14507_1337.n1 0.032
R6804 a_15097_1774.n7 a_15097_1774.n6 861.987
R6805 a_15097_1774.n6 a_15097_1774.n5 560.726
R6806 a_15097_1774.t13 a_15097_1774.t11 415.315
R6807 a_15097_1774.t4 a_15097_1774.t14 415.315
R6808 a_15097_1774.n2 a_15097_1774.t12 394.151
R6809 a_15097_1774.n5 a_15097_1774.t8 294.653
R6810 a_15097_1774.n1 a_15097_1774.t18 269.523
R6811 a_15097_1774.t12 a_15097_1774.n1 269.523
R6812 a_15097_1774.n9 a_15097_1774.t13 217.716
R6813 a_15097_1774.n8 a_15097_1774.t15 214.335
R6814 a_15097_1774.t11 a_15097_1774.n8 214.335
R6815 a_15097_1774.n0 a_15097_1774.t16 214.335
R6816 a_15097_1774.t14 a_15097_1774.n0 214.335
R6817 a_15097_1774.n7 a_15097_1774.t4 198.921
R6818 a_15097_1774.n3 a_15097_1774.t17 198.043
R6819 a_15097_1774.n12 a_15097_1774.n11 192.754
R6820 a_15097_1774.n1 a_15097_1774.t7 160.666
R6821 a_15097_1774.n5 a_15097_1774.t10 111.663
R6822 a_15097_1774.n4 a_15097_1774.n2 97.816
R6823 a_15097_1774.n3 a_15097_1774.t9 93.989
R6824 a_15097_1774.n8 a_15097_1774.t5 80.333
R6825 a_15097_1774.n2 a_15097_1774.t19 80.333
R6826 a_15097_1774.n0 a_15097_1774.t6 80.333
R6827 a_15097_1774.n6 a_15097_1774.n4 65.07
R6828 a_15097_1774.n11 a_15097_1774.t2 28.568
R6829 a_15097_1774.n12 a_15097_1774.t1 28.565
R6830 a_15097_1774.t3 a_15097_1774.n12 28.565
R6831 a_15097_1774.n10 a_15097_1774.t0 18.826
R6832 a_15097_1774.n9 a_15097_1774.n7 16.411
R6833 a_15097_1774.n4 a_15097_1774.n3 6.615
R6834 a_15097_1774.n10 a_15097_1774.n9 5.027
R6835 a_15097_1774.n11 a_15097_1774.n10 1.101
R6836 a_7947_9909.n0 a_7947_9909.t5 14.282
R6837 a_7947_9909.t0 a_7947_9909.n0 14.282
R6838 a_7947_9909.n0 a_7947_9909.n14 90.416
R6839 a_7947_9909.n14 a_7947_9909.n13 50.575
R6840 a_7947_9909.n14 a_7947_9909.n10 74.302
R6841 a_7947_9909.n13 a_7947_9909.n12 157.665
R6842 a_7947_9909.n12 a_7947_9909.t6 8.7
R6843 a_7947_9909.n12 a_7947_9909.t7 8.7
R6844 a_7947_9909.n13 a_7947_9909.n11 122.999
R6845 a_7947_9909.n11 a_7947_9909.t4 14.282
R6846 a_7947_9909.n11 a_7947_9909.t3 14.282
R6847 a_7947_9909.n10 a_7947_9909.n9 90.436
R6848 a_7947_9909.n9 a_7947_9909.t2 14.282
R6849 a_7947_9909.n9 a_7947_9909.t1 14.282
R6850 a_7947_9909.n1 a_7947_9909.t18 220.285
R6851 a_7947_9909.n10 a_7947_9909.n1 3509.5
R6852 a_7947_9909.n1 a_7947_9909.n8 61.538
R6853 a_7947_9909.n8 a_7947_9909.n3 465.933
R6854 a_7947_9909.n8 a_7947_9909.n7 163.88
R6855 a_7947_9909.n7 a_7947_9909.n6 6.615
R6856 a_7947_9909.n6 a_7947_9909.t13 93.989
R6857 a_7947_9909.n7 a_7947_9909.n5 97.816
R6858 a_7947_9909.n5 a_7947_9909.t16 80.333
R6859 a_7947_9909.n5 a_7947_9909.t19 394.151
R6860 a_7947_9909.t19 a_7947_9909.n4 269.523
R6861 a_7947_9909.n4 a_7947_9909.t8 160.666
R6862 a_7947_9909.n4 a_7947_9909.t9 269.523
R6863 a_7947_9909.n6 a_7947_9909.t12 198.043
R6864 a_7947_9909.n3 a_7947_9909.t14 294.653
R6865 a_7947_9909.n3 a_7947_9909.t17 111.663
R6866 a_7947_9909.t18 a_7947_9909.t10 415.315
R6867 a_7947_9909.t10 a_7947_9909.n2 214.335
R6868 a_7947_9909.n2 a_7947_9909.t11 80.333
R6869 a_7947_9909.n2 a_7947_9909.t15 214.335
R6870 a_31891_13791.n5 a_31891_13791.n7 0.575
R6871 a_31891_13791.n9 a_31891_13791.n5 0.2
R6872 a_31891_13791.t0 a_31891_13791.n9 16.058
R6873 a_31891_13791.n9 a_31891_13791.n8 0.999
R6874 a_31891_13791.n8 a_31891_13791.t2 14.282
R6875 a_31891_13791.n8 a_31891_13791.t1 14.282
R6876 a_31891_13791.n7 a_31891_13791.n6 0.999
R6877 a_31891_13791.n6 a_31891_13791.t6 14.282
R6878 a_31891_13791.n6 a_31891_13791.t8 14.282
R6879 a_31891_13791.n7 a_31891_13791.t7 16.058
R6880 a_31891_13791.n5 a_31891_13791.n3 0.227
R6881 a_31891_13791.n3 a_31891_13791.n4 1.511
R6882 a_31891_13791.n4 a_31891_13791.t3 14.282
R6883 a_31891_13791.n4 a_31891_13791.t5 14.282
R6884 a_31891_13791.n3 a_31891_13791.n0 0.669
R6885 a_31891_13791.n0 a_31891_13791.n1 0.001
R6886 a_31891_13791.n0 a_31891_13791.n2 267.767
R6887 a_31891_13791.n2 a_31891_13791.t10 14.282
R6888 a_31891_13791.n2 a_31891_13791.t11 14.282
R6889 a_31891_13791.n1 a_31891_13791.t4 14.282
R6890 a_31891_13791.n1 a_31891_13791.t9 14.282
R6891 A[1].n4 A[1].n3 535.449
R6892 A[1].t11 A[1].t6 437.233
R6893 A[1].t7 A[1].t9 437.233
R6894 A[1].t12 A[1].n1 313.873
R6895 A[1].n3 A[1].t15 294.986
R6896 A[1].n0 A[1].t14 272.288
R6897 A[1].n4 A[1].t1 245.184
R6898 A[1].n6 A[1].t7 218.628
R6899 A[1].n8 A[1].t11 217.024
R6900 A[1].n7 A[1].t13 214.686
R6901 A[1].t6 A[1].n7 214.686
R6902 A[1].n5 A[1].t4 214.686
R6903 A[1].t9 A[1].n5 214.686
R6904 A[1].n2 A[1].t12 190.152
R6905 A[1].n2 A[1].t3 190.152
R6906 A[1].n0 A[1].t0 160.666
R6907 A[1].n1 A[1].t2 160.666
R6908 A[1].n3 A[1].t10 110.859
R6909 A[1].n1 A[1].n0 96.129
R6910 A[1].n7 A[1].t5 80.333
R6911 A[1].t1 A[1].n2 80.333
R6912 A[1].n5 A[1].t8 80.333
R6913 A[1] A[1].n8 24.959
R6914 A[1].n6 A[1].n4 14.9
R6915 A[1].n8 A[1].n6 2.599
R6916 a_14248_24457.n0 a_14248_24457.n9 1.511
R6917 a_14248_24457.t3 a_14248_24457.n0 14.282
R6918 a_14248_24457.n0 a_14248_24457.t4 14.282
R6919 a_14248_24457.n9 a_14248_24457.n5 0.227
R6920 a_14248_24457.n9 a_14248_24457.n6 0.669
R6921 a_14248_24457.n6 a_14248_24457.n7 0.001
R6922 a_14248_24457.n6 a_14248_24457.n8 267.767
R6923 a_14248_24457.n8 a_14248_24457.t2 14.282
R6924 a_14248_24457.n8 a_14248_24457.t1 14.282
R6925 a_14248_24457.n7 a_14248_24457.t5 14.282
R6926 a_14248_24457.n7 a_14248_24457.t0 14.282
R6927 a_14248_24457.n5 a_14248_24457.n2 0.575
R6928 a_14248_24457.n5 a_14248_24457.n4 0.2
R6929 a_14248_24457.n4 a_14248_24457.t9 16.058
R6930 a_14248_24457.n4 a_14248_24457.n3 0.999
R6931 a_14248_24457.n3 a_14248_24457.t7 14.282
R6932 a_14248_24457.n3 a_14248_24457.t8 14.282
R6933 a_14248_24457.n2 a_14248_24457.n1 0.999
R6934 a_14248_24457.n1 a_14248_24457.t10 14.282
R6935 a_14248_24457.n1 a_14248_24457.t11 14.282
R6936 a_14248_24457.n2 a_14248_24457.t6 16.058
R6937 a_14490_4127.n0 a_14490_4127.n13 122.999
R6938 a_14490_4127.t1 a_14490_4127.n0 14.282
R6939 a_14490_4127.n0 a_14490_4127.t4 14.282
R6940 a_14490_4127.n13 a_14490_4127.n11 50.575
R6941 a_14490_4127.n11 a_14490_4127.n9 74.302
R6942 a_14490_4127.n13 a_14490_4127.n12 157.665
R6943 a_14490_4127.n12 a_14490_4127.t3 8.7
R6944 a_14490_4127.n12 a_14490_4127.t0 8.7
R6945 a_14490_4127.n11 a_14490_4127.n10 90.416
R6946 a_14490_4127.n10 a_14490_4127.t2 14.282
R6947 a_14490_4127.n10 a_14490_4127.t7 14.282
R6948 a_14490_4127.n9 a_14490_4127.n8 90.436
R6949 a_14490_4127.n8 a_14490_4127.t5 14.282
R6950 a_14490_4127.n8 a_14490_4127.t6 14.282
R6951 a_14490_4127.n9 a_14490_4127.n1 1712.43
R6952 a_14490_4127.n1 a_14490_4127.t8 217.826
R6953 a_14490_4127.n1 a_14490_4127.n6 133.839
R6954 a_14490_4127.t8 a_14490_4127.t16 437.233
R6955 a_14490_4127.t16 a_14490_4127.n7 214.686
R6956 a_14490_4127.n7 a_14490_4127.t9 80.333
R6957 a_14490_4127.n7 a_14490_4127.t12 214.686
R6958 a_14490_4127.n6 a_14490_4127.n2 563.136
R6959 a_14490_4127.n6 a_14490_4127.t17 178.973
R6960 a_14490_4127.t17 a_14490_4127.n5 80.333
R6961 a_14490_4127.n5 a_14490_4127.t18 190.152
R6962 a_14490_4127.n5 a_14490_4127.t10 190.152
R6963 a_14490_4127.t10 a_14490_4127.n4 313.873
R6964 a_14490_4127.n4 a_14490_4127.t14 160.666
R6965 a_14490_4127.n4 a_14490_4127.n3 96.129
R6966 a_14490_4127.n3 a_14490_4127.t11 160.666
R6967 a_14490_4127.n3 a_14490_4127.t13 272.288
R6968 a_14490_4127.n2 a_14490_4127.t15 294.986
R6969 a_14490_4127.n2 a_14490_4127.t19 110.859
R6970 a_33377_2547.n4 a_33377_2547.t9 214.335
R6971 a_33377_2547.t8 a_33377_2547.n4 214.335
R6972 a_33377_2547.n5 a_33377_2547.t8 143.851
R6973 a_33377_2547.n5 a_33377_2547.t7 135.658
R6974 a_33377_2547.n4 a_33377_2547.t10 80.333
R6975 a_33377_2547.n0 a_33377_2547.t2 28.565
R6976 a_33377_2547.n0 a_33377_2547.t1 28.565
R6977 a_33377_2547.n2 a_33377_2547.t6 28.565
R6978 a_33377_2547.n2 a_33377_2547.t0 28.565
R6979 a_33377_2547.t4 a_33377_2547.n7 28.565
R6980 a_33377_2547.n7 a_33377_2547.t5 28.565
R6981 a_33377_2547.n1 a_33377_2547.t3 9.714
R6982 a_33377_2547.n1 a_33377_2547.n0 1.003
R6983 a_33377_2547.n6 a_33377_2547.n3 0.833
R6984 a_33377_2547.n3 a_33377_2547.n2 0.653
R6985 a_33377_2547.n7 a_33377_2547.n6 0.653
R6986 a_33377_2547.n3 a_33377_2547.n1 0.341
R6987 a_33377_2547.n6 a_33377_2547.n5 0.032
R6988 a_33614_1910.t0 a_33614_1910.t1 17.4
R6989 B[5].n12 B[5].n6 973.987
R6990 B[5].n11 B[5].n7 592.056
R6991 B[5].t13 B[5].t1 437.233
R6992 B[5].t23 B[5].t14 437.233
R6993 B[5].t3 B[5].t0 415.315
R6994 B[5].t20 B[5].t9 415.315
R6995 B[5].t18 B[5].n9 313.069
R6996 B[5].n7 B[5].t17 294.986
R6997 B[5].n8 B[5].t11 271.484
R6998 B[5].n2 B[5].t20 240.379
R6999 B[5].n5 B[5].t23 227.856
R7000 B[5].n2 B[5].t3 218.339
R7001 B[5].n5 B[5].t13 218.225
R7002 B[5].n3 B[5].t21 214.686
R7003 B[5].t1 B[5].n3 214.686
R7004 B[5].n4 B[5].t2 214.686
R7005 B[5].t14 B[5].n4 214.686
R7006 B[5].n1 B[5].t8 214.335
R7007 B[5].t0 B[5].n1 214.335
R7008 B[5].n0 B[5].t16 214.335
R7009 B[5].t9 B[5].n0 214.335
R7010 B[5].n11 B[5].t10 204.672
R7011 B[5].n10 B[5].t18 190.955
R7012 B[5].n10 B[5].t4 190.955
R7013 B[5].n9 B[5].t22 160.666
R7014 B[5].n8 B[5].t5 160.666
R7015 B[5].n7 B[5].t7 110.859
R7016 B[5].n9 B[5].n8 96.129
R7017 B[5].n1 B[5].t6 80.333
R7018 B[5].n0 B[5].t12 80.333
R7019 B[5].n3 B[5].t15 80.333
R7020 B[5].n4 B[5].t19 80.333
R7021 B[5].t10 B[5].n10 80.333
R7022 B[5].n12 B[5].n11 46.001
R7023 B[5].n6 B[5].n2 28.897
R7024 B[5] B[5].n12 27.064
R7025 B[5].n6 B[5].n5 7.414
R7026 a_14467_15035.n2 a_14467_15035.t10 214.335
R7027 a_14467_15035.t8 a_14467_15035.n2 214.335
R7028 a_14467_15035.n3 a_14467_15035.t8 143.851
R7029 a_14467_15035.n3 a_14467_15035.t7 135.658
R7030 a_14467_15035.n2 a_14467_15035.t9 80.333
R7031 a_14467_15035.n4 a_14467_15035.t0 28.565
R7032 a_14467_15035.n4 a_14467_15035.t1 28.565
R7033 a_14467_15035.n0 a_14467_15035.t5 28.565
R7034 a_14467_15035.n0 a_14467_15035.t6 28.565
R7035 a_14467_15035.t2 a_14467_15035.n7 28.565
R7036 a_14467_15035.n7 a_14467_15035.t4 28.565
R7037 a_14467_15035.n1 a_14467_15035.t3 9.714
R7038 a_14467_15035.n1 a_14467_15035.n0 1.003
R7039 a_14467_15035.n6 a_14467_15035.n5 0.833
R7040 a_14467_15035.n5 a_14467_15035.n4 0.653
R7041 a_14467_15035.n7 a_14467_15035.n6 0.653
R7042 a_14467_15035.n6 a_14467_15035.n1 0.341
R7043 a_14467_15035.n5 a_14467_15035.n3 0.032
R7044 a_8508_14599.n4 a_8508_14599.n3 535.449
R7045 a_8508_14599.t6 a_8508_14599.t4 437.233
R7046 a_8508_14599.t14 a_8508_14599.t9 437.233
R7047 a_8508_14599.t10 a_8508_14599.n1 313.873
R7048 a_8508_14599.n3 a_8508_14599.t18 294.986
R7049 a_8508_14599.n0 a_8508_14599.t17 272.288
R7050 a_8508_14599.n4 a_8508_14599.t11 245.184
R7051 a_8508_14599.n6 a_8508_14599.t14 218.628
R7052 a_8508_14599.n8 a_8508_14599.t6 217.024
R7053 a_8508_14599.n7 a_8508_14599.t15 214.686
R7054 a_8508_14599.t4 a_8508_14599.n7 214.686
R7055 a_8508_14599.n5 a_8508_14599.t8 214.686
R7056 a_8508_14599.t9 a_8508_14599.n5 214.686
R7057 a_8508_14599.n11 a_8508_14599.n10 192.754
R7058 a_8508_14599.n2 a_8508_14599.t10 190.152
R7059 a_8508_14599.n2 a_8508_14599.t19 190.152
R7060 a_8508_14599.n0 a_8508_14599.t12 160.666
R7061 a_8508_14599.n1 a_8508_14599.t13 160.666
R7062 a_8508_14599.n3 a_8508_14599.t7 110.859
R7063 a_8508_14599.n1 a_8508_14599.n0 96.129
R7064 a_8508_14599.n7 a_8508_14599.t16 80.333
R7065 a_8508_14599.t11 a_8508_14599.n2 80.333
R7066 a_8508_14599.n5 a_8508_14599.t5 80.333
R7067 a_8508_14599.n10 a_8508_14599.t1 28.568
R7068 a_8508_14599.t0 a_8508_14599.n11 28.565
R7069 a_8508_14599.n11 a_8508_14599.t2 28.565
R7070 a_8508_14599.n9 a_8508_14599.t3 18.819
R7071 a_8508_14599.n6 a_8508_14599.n4 14.9
R7072 a_8508_14599.n9 a_8508_14599.n8 2.96
R7073 a_8508_14599.n8 a_8508_14599.n6 2.599
R7074 a_8508_14599.n10 a_8508_14599.n9 1.098
R7075 a_10693_12957.n2 a_10693_12957.t10 214.335
R7076 a_10693_12957.t8 a_10693_12957.n2 214.335
R7077 a_10693_12957.n3 a_10693_12957.t8 143.851
R7078 a_10693_12957.n3 a_10693_12957.t7 135.658
R7079 a_10693_12957.n2 a_10693_12957.t9 80.333
R7080 a_10693_12957.n4 a_10693_12957.t6 28.565
R7081 a_10693_12957.n4 a_10693_12957.t5 28.565
R7082 a_10693_12957.n0 a_10693_12957.t1 28.565
R7083 a_10693_12957.n0 a_10693_12957.t2 28.565
R7084 a_10693_12957.t4 a_10693_12957.n7 28.565
R7085 a_10693_12957.n7 a_10693_12957.t3 28.565
R7086 a_10693_12957.n1 a_10693_12957.t0 9.714
R7087 a_10693_12957.n1 a_10693_12957.n0 1.003
R7088 a_10693_12957.n6 a_10693_12957.n5 0.833
R7089 a_10693_12957.n5 a_10693_12957.n4 0.653
R7090 a_10693_12957.n7 a_10693_12957.n6 0.653
R7091 a_10693_12957.n6 a_10693_12957.n1 0.341
R7092 a_10693_12957.n5 a_10693_12957.n3 0.032
R7093 a_28608_18536.n0 a_28608_18536.t10 214.335
R7094 a_28608_18536.t8 a_28608_18536.n0 214.335
R7095 a_28608_18536.n1 a_28608_18536.t8 143.851
R7096 a_28608_18536.n1 a_28608_18536.t9 135.658
R7097 a_28608_18536.n0 a_28608_18536.t7 80.333
R7098 a_28608_18536.n2 a_28608_18536.t6 28.565
R7099 a_28608_18536.n2 a_28608_18536.t5 28.565
R7100 a_28608_18536.n4 a_28608_18536.t4 28.565
R7101 a_28608_18536.n4 a_28608_18536.t1 28.565
R7102 a_28608_18536.n7 a_28608_18536.t2 28.565
R7103 a_28608_18536.t0 a_28608_18536.n7 28.565
R7104 a_28608_18536.n3 a_28608_18536.t3 9.714
R7105 a_28608_18536.n3 a_28608_18536.n2 1.003
R7106 a_28608_18536.n6 a_28608_18536.n5 0.833
R7107 a_28608_18536.n5 a_28608_18536.n4 0.653
R7108 a_28608_18536.n7 a_28608_18536.n6 0.653
R7109 a_28608_18536.n5 a_28608_18536.n3 0.341
R7110 a_28608_18536.n6 a_28608_18536.n1 0.032
R7111 a_27000_21662.t7 a_27000_21662.t4 574.43
R7112 a_27000_21662.n0 a_27000_21662.t5 285.109
R7113 a_27000_21662.n2 a_27000_21662.n1 197.215
R7114 a_27000_21662.n4 a_27000_21662.n3 192.754
R7115 a_27000_21662.n0 a_27000_21662.t6 160.666
R7116 a_27000_21662.n1 a_27000_21662.t7 160.666
R7117 a_27000_21662.n1 a_27000_21662.n0 114.829
R7118 a_27000_21662.n3 a_27000_21662.t1 28.568
R7119 a_27000_21662.n4 a_27000_21662.t2 28.565
R7120 a_27000_21662.t3 a_27000_21662.n4 28.565
R7121 a_27000_21662.n2 a_27000_21662.t0 18.838
R7122 a_27000_21662.n3 a_27000_21662.n2 1.129
R7123 a_7953_1332.n0 a_7953_1332.t9 214.335
R7124 a_7953_1332.t8 a_7953_1332.n0 214.335
R7125 a_7953_1332.n1 a_7953_1332.t8 143.85
R7126 a_7953_1332.n1 a_7953_1332.t7 135.66
R7127 a_7953_1332.n0 a_7953_1332.t10 80.333
R7128 a_7953_1332.n2 a_7953_1332.t2 28.565
R7129 a_7953_1332.n2 a_7953_1332.t1 28.565
R7130 a_7953_1332.n4 a_7953_1332.t6 28.565
R7131 a_7953_1332.n4 a_7953_1332.t3 28.565
R7132 a_7953_1332.t4 a_7953_1332.n7 28.565
R7133 a_7953_1332.n7 a_7953_1332.t5 28.565
R7134 a_7953_1332.n3 a_7953_1332.t0 9.714
R7135 a_7953_1332.n3 a_7953_1332.n2 1.003
R7136 a_7953_1332.n6 a_7953_1332.n5 0.836
R7137 a_7953_1332.n5 a_7953_1332.n4 0.653
R7138 a_7953_1332.n7 a_7953_1332.n6 0.65
R7139 a_7953_1332.n5 a_7953_1332.n3 0.341
R7140 a_7953_1332.n6 a_7953_1332.n1 0.032
R7141 B[4].n5 B[4].t15 1361.95
R7142 B[4].n4 B[4].t21 1211.76
R7143 B[4].n10 B[4].n6 592.056
R7144 B[4].n5 B[4].t11 561.041
R7145 B[4].t15 B[4].t18 437.233
R7146 B[4].t11 B[4].t4 437.233
R7147 B[4].t21 B[4].t22 415.315
R7148 B[4].t23 B[4].t16 415.315
R7149 B[4].t1 B[4].n8 313.069
R7150 B[4].n6 B[4].t5 294.986
R7151 B[4].n7 B[4].t17 271.484
R7152 B[4].n4 B[4].t23 219.359
R7153 B[4].n0 B[4].t13 214.686
R7154 B[4].t18 B[4].n0 214.686
R7155 B[4].n1 B[4].t9 214.686
R7156 B[4].t4 B[4].n1 214.686
R7157 B[4].n2 B[4].t0 214.335
R7158 B[4].t22 B[4].n2 214.335
R7159 B[4].n3 B[4].t20 214.335
R7160 B[4].t16 B[4].n3 214.335
R7161 B[4].n10 B[4].t14 204.672
R7162 B[4].n9 B[4].t1 190.955
R7163 B[4].n9 B[4].t6 190.955
R7164 B[4].n8 B[4].t3 160.666
R7165 B[4].n7 B[4].t7 160.666
R7166 B[4].n6 B[4].t12 110.859
R7167 B[4].n8 B[4].n7 96.129
R7168 B[4].n0 B[4].t2 80.333
R7169 B[4].n1 B[4].t10 80.333
R7170 B[4].n2 B[4].t8 80.333
R7171 B[4].n3 B[4].t19 80.333
R7172 B[4].t14 B[4].n9 80.333
R7173 B[4].n11 B[4].n10 52.607
R7174 B[4] B[4].n11 16.139
R7175 B[4].n11 B[4].n5 1.607
R7176 B[4].n5 B[4].n4 1.018
R7177 a_1227_7273.n4 a_1227_7273.t7 214.335
R7178 a_1227_7273.t10 a_1227_7273.n4 214.335
R7179 a_1227_7273.n5 a_1227_7273.t10 143.851
R7180 a_1227_7273.n5 a_1227_7273.t9 135.658
R7181 a_1227_7273.n4 a_1227_7273.t8 80.333
R7182 a_1227_7273.n0 a_1227_7273.t4 28.565
R7183 a_1227_7273.n0 a_1227_7273.t6 28.565
R7184 a_1227_7273.n2 a_1227_7273.t0 28.565
R7185 a_1227_7273.n2 a_1227_7273.t5 28.565
R7186 a_1227_7273.t2 a_1227_7273.n7 28.565
R7187 a_1227_7273.n7 a_1227_7273.t1 28.565
R7188 a_1227_7273.n1 a_1227_7273.t3 9.714
R7189 a_1227_7273.n1 a_1227_7273.n0 1.003
R7190 a_1227_7273.n6 a_1227_7273.n3 0.833
R7191 a_1227_7273.n3 a_1227_7273.n2 0.653
R7192 a_1227_7273.n7 a_1227_7273.n6 0.653
R7193 a_1227_7273.n3 a_1227_7273.n1 0.341
R7194 a_1227_7273.n6 a_1227_7273.n5 0.032
R7195 a_15810_27293.t5 a_15810_27293.n2 404.877
R7196 a_15810_27293.n1 a_15810_27293.t7 210.902
R7197 a_15810_27293.n3 a_15810_27293.t5 136.943
R7198 a_15810_27293.n2 a_15810_27293.n1 107.801
R7199 a_15810_27293.n1 a_15810_27293.t6 80.333
R7200 a_15810_27293.n2 a_15810_27293.t8 80.333
R7201 a_15810_27293.n0 a_15810_27293.t0 17.4
R7202 a_15810_27293.n0 a_15810_27293.t2 17.4
R7203 a_15810_27293.n4 a_15810_27293.t3 15.032
R7204 a_15810_27293.t1 a_15810_27293.n5 14.282
R7205 a_15810_27293.n5 a_15810_27293.t4 14.282
R7206 a_15810_27293.n5 a_15810_27293.n4 1.65
R7207 a_15810_27293.n3 a_15810_27293.n0 0.672
R7208 a_15810_27293.n4 a_15810_27293.n3 0.665
R7209 a_16074_26710.n6 a_16074_26710.n5 501.28
R7210 a_16074_26710.t16 a_16074_26710.t18 437.233
R7211 a_16074_26710.t4 a_16074_26710.t17 415.315
R7212 a_16074_26710.t7 a_16074_26710.n3 313.873
R7213 a_16074_26710.n5 a_16074_26710.t14 294.986
R7214 a_16074_26710.n2 a_16074_26710.t10 272.288
R7215 a_16074_26710.n6 a_16074_26710.t8 236.01
R7216 a_16074_26710.n9 a_16074_26710.t16 216.627
R7217 a_16074_26710.n7 a_16074_26710.t4 216.111
R7218 a_16074_26710.n8 a_16074_26710.t19 214.686
R7219 a_16074_26710.t18 a_16074_26710.n8 214.686
R7220 a_16074_26710.n1 a_16074_26710.t6 214.335
R7221 a_16074_26710.t17 a_16074_26710.n1 214.335
R7222 a_16074_26710.n4 a_16074_26710.t7 190.152
R7223 a_16074_26710.n4 a_16074_26710.t13 190.152
R7224 a_16074_26710.n2 a_16074_26710.t11 160.666
R7225 a_16074_26710.n3 a_16074_26710.t12 160.666
R7226 a_16074_26710.n7 a_16074_26710.n6 148.428
R7227 a_16074_26710.n5 a_16074_26710.t9 110.859
R7228 a_16074_26710.n3 a_16074_26710.n2 96.129
R7229 a_16074_26710.n8 a_16074_26710.t15 80.333
R7230 a_16074_26710.n1 a_16074_26710.t5 80.333
R7231 a_16074_26710.t8 a_16074_26710.n4 80.333
R7232 a_16074_26710.n0 a_16074_26710.t1 28.57
R7233 a_16074_26710.n11 a_16074_26710.t2 28.565
R7234 a_16074_26710.t3 a_16074_26710.n11 28.565
R7235 a_16074_26710.n0 a_16074_26710.t0 17.638
R7236 a_16074_26710.n10 a_16074_26710.n9 5.6
R7237 a_16074_26710.n9 a_16074_26710.n7 2.923
R7238 a_16074_26710.n11 a_16074_26710.n10 0.69
R7239 a_16074_26710.n10 a_16074_26710.n0 0.6
R7240 a_36755_23013.t0 a_36755_23013.n0 14.282
R7241 a_36755_23013.n0 a_36755_23013.t2 14.282
R7242 a_36755_23013.n0 a_36755_23013.n1 258.161
R7243 a_36755_23013.n1 a_36755_23013.n7 4.366
R7244 a_36755_23013.n7 a_36755_23013.n5 0.852
R7245 a_36755_23013.n5 a_36755_23013.n6 258.161
R7246 a_36755_23013.n6 a_36755_23013.t5 14.282
R7247 a_36755_23013.n6 a_36755_23013.t6 14.282
R7248 a_36755_23013.n5 a_36755_23013.t4 14.283
R7249 a_36755_23013.n7 a_36755_23013.n4 73.514
R7250 a_36755_23013.n4 a_36755_23013.t8 1551.5
R7251 a_36755_23013.t8 a_36755_23013.n3 656.576
R7252 a_36755_23013.n3 a_36755_23013.t1 8.7
R7253 a_36755_23013.n3 a_36755_23013.t7 8.7
R7254 a_36755_23013.n4 a_36755_23013.t9 224.129
R7255 a_36755_23013.t9 a_36755_23013.n2 207.225
R7256 a_36755_23013.n2 a_36755_23013.t11 207.225
R7257 a_36755_23013.n2 a_36755_23013.t10 80.333
R7258 a_36755_23013.n1 a_36755_23013.t3 14.283
R7259 Y[0].n1 Y[0].n0 185.55
R7260 Y[0].n1 Y[0].t3 28.568
R7261 Y[0].n0 Y[0].t1 28.565
R7262 Y[0].n0 Y[0].t2 28.565
R7263 Y[0].n2 Y[0].t0 20.393
R7264 Y[0].n2 Y[0].n1 1.831
R7265 Y[0].n3 Y[0].n2 1.048
R7266 Y[0] Y[0].n3 0.052
R7267 Y[0].n3 Y[0] 0.046
R7268 a_30359_11881.n4 a_30359_11881.n3 563.136
R7269 a_30359_11881.t11 a_30359_11881.t14 437.233
R7270 a_30359_11881.t5 a_30359_11881.n1 313.873
R7271 a_30359_11881.n3 a_30359_11881.t10 294.986
R7272 a_30359_11881.n0 a_30359_11881.t4 272.288
R7273 a_30359_11881.n6 a_30359_11881.t11 217.824
R7274 a_30359_11881.n5 a_30359_11881.t12 214.686
R7275 a_30359_11881.t14 a_30359_11881.n5 214.686
R7276 a_30359_11881.n9 a_30359_11881.n8 192.754
R7277 a_30359_11881.n2 a_30359_11881.t5 190.152
R7278 a_30359_11881.n2 a_30359_11881.t9 190.152
R7279 a_30359_11881.n4 a_30359_11881.t6 178.973
R7280 a_30359_11881.n0 a_30359_11881.t7 160.666
R7281 a_30359_11881.n1 a_30359_11881.t8 160.666
R7282 a_30359_11881.n6 a_30359_11881.n4 133.838
R7283 a_30359_11881.n3 a_30359_11881.t15 110.859
R7284 a_30359_11881.n1 a_30359_11881.n0 96.129
R7285 a_30359_11881.t6 a_30359_11881.n2 80.333
R7286 a_30359_11881.n5 a_30359_11881.t13 80.333
R7287 a_30359_11881.n8 a_30359_11881.t1 28.568
R7288 a_30359_11881.n9 a_30359_11881.t2 28.565
R7289 a_30359_11881.t3 a_30359_11881.n9 28.565
R7290 a_30359_11881.n7 a_30359_11881.t0 18.822
R7291 a_30359_11881.n7 a_30359_11881.n6 5.647
R7292 a_30359_11881.n8 a_30359_11881.n7 1.105
R7293 a_n3608_55.n1 a_n3608_55.t6 318.119
R7294 a_n3608_55.n1 a_n3608_55.t5 269.919
R7295 a_n3608_55.n0 a_n3608_55.t7 267.853
R7296 a_n3608_55.n0 a_n3608_55.t4 267.853
R7297 a_n3608_55.t6 a_n3608_55.n0 160.666
R7298 a_n3608_55.n2 a_n3608_55.n1 107.263
R7299 a_n3608_55.t0 a_n3608_55.n4 29.444
R7300 a_n3608_55.n3 a_n3608_55.t2 28.565
R7301 a_n3608_55.n3 a_n3608_55.t1 28.565
R7302 a_n3608_55.n2 a_n3608_55.t3 18.145
R7303 a_n3608_55.n4 a_n3608_55.n2 2.878
R7304 a_n3608_55.n4 a_n3608_55.n3 0.764
R7305 a_n3808_656.n0 a_n3808_656.t1 14.282
R7306 a_n3808_656.t0 a_n3808_656.n0 14.282
R7307 a_n3808_656.n0 a_n3808_656.n9 0.999
R7308 a_n3808_656.n9 a_n3808_656.n6 0.2
R7309 a_n3808_656.n6 a_n3808_656.n8 0.575
R7310 a_n3808_656.n9 a_n3808_656.t2 16.058
R7311 a_n3808_656.n8 a_n3808_656.n7 0.999
R7312 a_n3808_656.n7 a_n3808_656.t4 14.282
R7313 a_n3808_656.n7 a_n3808_656.t5 14.282
R7314 a_n3808_656.n8 a_n3808_656.t3 16.058
R7315 a_n3808_656.n6 a_n3808_656.n4 0.227
R7316 a_n3808_656.n4 a_n3808_656.n5 1.511
R7317 a_n3808_656.n5 a_n3808_656.t11 14.282
R7318 a_n3808_656.n5 a_n3808_656.t9 14.282
R7319 a_n3808_656.n4 a_n3808_656.n1 0.669
R7320 a_n3808_656.n1 a_n3808_656.n2 0.001
R7321 a_n3808_656.n1 a_n3808_656.n3 267.767
R7322 a_n3808_656.n3 a_n3808_656.t7 14.282
R7323 a_n3808_656.n3 a_n3808_656.t8 14.282
R7324 a_n3808_656.n2 a_n3808_656.t6 14.282
R7325 a_n3808_656.n2 a_n3808_656.t10 14.282
R7326 a_n3115_713.n0 a_n3115_713.t6 14.282
R7327 a_n3115_713.t4 a_n3115_713.n0 14.282
R7328 a_n3115_713.n4 a_n3115_713.n2 74.302
R7329 a_n3115_713.n6 a_n3115_713.n4 50.575
R7330 a_n3115_713.n0 a_n3115_713.n6 110.084
R7331 a_n3115_713.n2 a_n3115_713.n7 664.97
R7332 a_n3115_713.n7 a_n3115_713.n9 16.411
R7333 a_n3115_713.n9 a_n3115_713.t21 198.921
R7334 a_n3115_713.t21 a_n3115_713.t20 415.315
R7335 a_n3115_713.t20 a_n3115_713.n16 214.335
R7336 a_n3115_713.n16 a_n3115_713.t15 80.333
R7337 a_n3115_713.n16 a_n3115_713.t14 214.335
R7338 a_n3115_713.n9 a_n3115_713.n15 861.987
R7339 a_n3115_713.n15 a_n3115_713.n10 560.726
R7340 a_n3115_713.n15 a_n3115_713.n14 65.07
R7341 a_n3115_713.n14 a_n3115_713.n13 6.615
R7342 a_n3115_713.n13 a_n3115_713.t18 93.989
R7343 a_n3115_713.n13 a_n3115_713.t23 198.043
R7344 a_n3115_713.n14 a_n3115_713.n12 97.816
R7345 a_n3115_713.n12 a_n3115_713.t17 80.333
R7346 a_n3115_713.n12 a_n3115_713.t10 394.151
R7347 a_n3115_713.t10 a_n3115_713.n11 269.523
R7348 a_n3115_713.n11 a_n3115_713.t9 160.666
R7349 a_n3115_713.n11 a_n3115_713.t8 269.523
R7350 a_n3115_713.n10 a_n3115_713.t13 294.653
R7351 a_n3115_713.n10 a_n3115_713.t22 111.663
R7352 a_n3115_713.n7 a_n3115_713.t16 217.716
R7353 a_n3115_713.t16 a_n3115_713.t19 415.315
R7354 a_n3115_713.t19 a_n3115_713.n8 214.335
R7355 a_n3115_713.n8 a_n3115_713.t12 80.333
R7356 a_n3115_713.n8 a_n3115_713.t11 214.335
R7357 a_n3115_713.n6 a_n3115_713.n5 157.665
R7358 a_n3115_713.n5 a_n3115_713.t7 8.7
R7359 a_n3115_713.n5 a_n3115_713.t3 8.7
R7360 a_n3115_713.n4 a_n3115_713.n3 90.416
R7361 a_n3115_713.n3 a_n3115_713.t0 14.282
R7362 a_n3115_713.n3 a_n3115_713.t5 14.282
R7363 a_n3115_713.n2 a_n3115_713.n1 90.436
R7364 a_n3115_713.n1 a_n3115_713.t2 14.282
R7365 a_n3115_713.n1 a_n3115_713.t1 14.282
R7366 a_25465_19523.n0 a_25465_19523.n12 90.436
R7367 a_25465_19523.t0 a_25465_19523.n0 14.282
R7368 a_25465_19523.n0 a_25465_19523.t1 14.282
R7369 a_25465_19523.n12 a_25465_19523.n9 74.302
R7370 a_25465_19523.n9 a_25465_19523.n11 50.575
R7371 a_25465_19523.n11 a_25465_19523.n10 157.665
R7372 a_25465_19523.n10 a_25465_19523.t7 8.7
R7373 a_25465_19523.n10 a_25465_19523.t5 8.7
R7374 a_25465_19523.n9 a_25465_19523.n8 90.416
R7375 a_25465_19523.n8 a_25465_19523.t2 14.282
R7376 a_25465_19523.n8 a_25465_19523.t6 14.282
R7377 a_25465_19523.n11 a_25465_19523.n7 122.746
R7378 a_25465_19523.n7 a_25465_19523.t3 14.282
R7379 a_25465_19523.n7 a_25465_19523.t4 14.282
R7380 a_25465_19523.n12 a_25465_19523.n1 342.688
R7381 a_25465_19523.n1 a_25465_19523.n6 126.566
R7382 a_25465_19523.n6 a_25465_19523.t15 294.653
R7383 a_25465_19523.n6 a_25465_19523.t9 111.663
R7384 a_25465_19523.n1 a_25465_19523.n5 552.333
R7385 a_25465_19523.n5 a_25465_19523.n4 6.615
R7386 a_25465_19523.n4 a_25465_19523.t10 93.989
R7387 a_25465_19523.n4 a_25465_19523.t11 198.043
R7388 a_25465_19523.n5 a_25465_19523.n3 97.816
R7389 a_25465_19523.n3 a_25465_19523.t12 80.333
R7390 a_25465_19523.n3 a_25465_19523.t8 394.151
R7391 a_25465_19523.t8 a_25465_19523.n2 269.523
R7392 a_25465_19523.n2 a_25465_19523.t14 160.666
R7393 a_25465_19523.n2 a_25465_19523.t13 269.523
R7394 a_25110_18856.t0 a_25110_18856.n0 14.282
R7395 a_25110_18856.n0 a_25110_18856.t5 14.282
R7396 a_25110_18856.n0 a_25110_18856.n9 0.999
R7397 a_25110_18856.n6 a_25110_18856.n8 0.2
R7398 a_25110_18856.n9 a_25110_18856.n6 0.575
R7399 a_25110_18856.n9 a_25110_18856.t4 16.058
R7400 a_25110_18856.n8 a_25110_18856.n7 0.999
R7401 a_25110_18856.n7 a_25110_18856.t11 14.282
R7402 a_25110_18856.n7 a_25110_18856.t9 14.282
R7403 a_25110_18856.n8 a_25110_18856.t10 16.058
R7404 a_25110_18856.n6 a_25110_18856.n4 0.227
R7405 a_25110_18856.n4 a_25110_18856.n5 1.511
R7406 a_25110_18856.n5 a_25110_18856.t1 14.282
R7407 a_25110_18856.n5 a_25110_18856.t3 14.282
R7408 a_25110_18856.n4 a_25110_18856.n1 0.669
R7409 a_25110_18856.n1 a_25110_18856.n2 0.001
R7410 a_25110_18856.n1 a_25110_18856.n3 267.767
R7411 a_25110_18856.n3 a_25110_18856.t6 14.282
R7412 a_25110_18856.n3 a_25110_18856.t7 14.282
R7413 a_25110_18856.n2 a_25110_18856.t8 14.282
R7414 a_25110_18856.n2 a_25110_18856.t2 14.282
R7415 a_n3606_9768.n2 a_n3606_9768.t6 318.119
R7416 a_n3606_9768.n2 a_n3606_9768.t4 269.919
R7417 a_n3606_9768.n1 a_n3606_9768.t7 267.256
R7418 a_n3606_9768.n1 a_n3606_9768.t5 267.256
R7419 a_n3606_9768.n4 a_n3606_9768.n0 193.227
R7420 a_n3606_9768.t6 a_n3606_9768.n1 160.666
R7421 a_n3606_9768.n3 a_n3606_9768.n2 106.999
R7422 a_n3606_9768.t0 a_n3606_9768.n4 28.568
R7423 a_n3606_9768.n0 a_n3606_9768.t2 28.565
R7424 a_n3606_9768.n0 a_n3606_9768.t1 28.565
R7425 a_n3606_9768.n3 a_n3606_9768.t3 18.149
R7426 a_n3606_9768.n4 a_n3606_9768.n3 3.726
R7427 a_n3113_8987.n0 a_n3113_8987.t6 14.282
R7428 a_n3113_8987.t0 a_n3113_8987.n0 14.282
R7429 a_n3113_8987.n0 a_n3113_8987.n16 90.436
R7430 a_n3113_8987.n16 a_n3113_8987.n2 74.302
R7431 a_n3113_8987.n2 a_n3113_8987.n4 50.575
R7432 a_n3113_8987.n4 a_n3113_8987.n5 110.084
R7433 a_n3113_8987.n16 a_n3113_8987.n6 214.569
R7434 a_n3113_8987.n6 a_n3113_8987.n8 16.411
R7435 a_n3113_8987.n8 a_n3113_8987.t14 198.921
R7436 a_n3113_8987.t14 a_n3113_8987.t15 415.315
R7437 a_n3113_8987.t15 a_n3113_8987.n15 214.335
R7438 a_n3113_8987.n15 a_n3113_8987.t22 80.333
R7439 a_n3113_8987.n15 a_n3113_8987.t20 214.335
R7440 a_n3113_8987.n8 a_n3113_8987.n14 861.987
R7441 a_n3113_8987.n14 a_n3113_8987.n9 560.726
R7442 a_n3113_8987.n14 a_n3113_8987.n13 65.07
R7443 a_n3113_8987.n13 a_n3113_8987.n12 6.615
R7444 a_n3113_8987.n12 a_n3113_8987.t23 93.989
R7445 a_n3113_8987.n13 a_n3113_8987.n11 97.816
R7446 a_n3113_8987.n11 a_n3113_8987.t8 80.333
R7447 a_n3113_8987.n11 a_n3113_8987.t11 394.151
R7448 a_n3113_8987.t11 a_n3113_8987.n10 269.523
R7449 a_n3113_8987.n10 a_n3113_8987.t12 160.666
R7450 a_n3113_8987.n10 a_n3113_8987.t13 269.523
R7451 a_n3113_8987.n12 a_n3113_8987.t19 198.043
R7452 a_n3113_8987.n9 a_n3113_8987.t10 294.653
R7453 a_n3113_8987.n9 a_n3113_8987.t9 111.663
R7454 a_n3113_8987.n6 a_n3113_8987.t21 217.716
R7455 a_n3113_8987.t21 a_n3113_8987.t17 415.315
R7456 a_n3113_8987.t17 a_n3113_8987.n7 214.335
R7457 a_n3113_8987.n7 a_n3113_8987.t18 80.333
R7458 a_n3113_8987.n7 a_n3113_8987.t16 214.335
R7459 a_n3113_8987.n5 a_n3113_8987.t2 14.282
R7460 a_n3113_8987.n5 a_n3113_8987.t3 14.282
R7461 a_n3113_8987.n4 a_n3113_8987.n3 157.665
R7462 a_n3113_8987.n3 a_n3113_8987.t7 8.7
R7463 a_n3113_8987.n3 a_n3113_8987.t4 8.7
R7464 a_n3113_8987.n2 a_n3113_8987.n1 90.416
R7465 a_n3113_8987.n1 a_n3113_8987.t5 14.282
R7466 a_n3113_8987.n1 a_n3113_8987.t1 14.282
R7467 a_n2381_8987.t0 a_n2381_8987.t1 379.845
R7468 a_19554_12761.t8 a_19554_12761.n2 404.877
R7469 a_19554_12761.n1 a_19554_12761.t7 210.902
R7470 a_19554_12761.n3 a_19554_12761.t8 136.943
R7471 a_19554_12761.n2 a_19554_12761.n1 107.801
R7472 a_19554_12761.n1 a_19554_12761.t6 80.333
R7473 a_19554_12761.n2 a_19554_12761.t5 80.333
R7474 a_19554_12761.n0 a_19554_12761.t0 17.4
R7475 a_19554_12761.n0 a_19554_12761.t3 17.4
R7476 a_19554_12761.n4 a_19554_12761.t4 15.032
R7477 a_19554_12761.n5 a_19554_12761.t2 14.282
R7478 a_19554_12761.t1 a_19554_12761.n5 14.282
R7479 a_19554_12761.n5 a_19554_12761.n4 1.65
R7480 a_19554_12761.n3 a_19554_12761.n0 0.672
R7481 a_19554_12761.n4 a_19554_12761.n3 0.665
R7482 a_19818_12178.t4 a_19818_12178.t7 800.071
R7483 a_19818_12178.n3 a_19818_12178.n2 672.951
R7484 a_19818_12178.n1 a_19818_12178.t6 285.109
R7485 a_19818_12178.n2 a_19818_12178.t4 193.602
R7486 a_19818_12178.n1 a_19818_12178.t5 160.666
R7487 a_19818_12178.n2 a_19818_12178.n1 91.507
R7488 a_19818_12178.t3 a_19818_12178.n4 28.57
R7489 a_19818_12178.n0 a_19818_12178.t1 28.565
R7490 a_19818_12178.n0 a_19818_12178.t2 28.565
R7491 a_19818_12178.n4 a_19818_12178.t0 17.638
R7492 a_19818_12178.n3 a_19818_12178.n0 0.69
R7493 a_19818_12178.n4 a_19818_12178.n3 0.6
R7494 a_31464_14484.n2 a_31464_14484.t4 318.922
R7495 a_31464_14484.n1 a_31464_14484.t6 273.935
R7496 a_31464_14484.n1 a_31464_14484.t5 273.935
R7497 a_31464_14484.n2 a_31464_14484.t7 269.116
R7498 a_31464_14484.n4 a_31464_14484.n0 193.227
R7499 a_31464_14484.t4 a_31464_14484.n1 179.142
R7500 a_31464_14484.n3 a_31464_14484.n2 106.999
R7501 a_31464_14484.t3 a_31464_14484.n4 28.568
R7502 a_31464_14484.n0 a_31464_14484.t1 28.565
R7503 a_31464_14484.n0 a_31464_14484.t2 28.565
R7504 a_31464_14484.n3 a_31464_14484.t0 18.149
R7505 a_31464_14484.n4 a_31464_14484.n3 3.726
R7506 a_32009_13791.n0 a_32009_13791.t1 14.282
R7507 a_32009_13791.t0 a_32009_13791.n0 14.282
R7508 a_32009_13791.n0 a_32009_13791.n8 90.436
R7509 a_32009_13791.n4 a_32009_13791.n7 50.575
R7510 a_32009_13791.n8 a_32009_13791.n4 74.302
R7511 a_32009_13791.n7 a_32009_13791.n6 157.665
R7512 a_32009_13791.n6 a_32009_13791.t6 8.7
R7513 a_32009_13791.n6 a_32009_13791.t7 8.7
R7514 a_32009_13791.n7 a_32009_13791.n5 122.999
R7515 a_32009_13791.n5 a_32009_13791.t3 14.282
R7516 a_32009_13791.n5 a_32009_13791.t5 14.282
R7517 a_32009_13791.n4 a_32009_13791.n3 90.416
R7518 a_32009_13791.n3 a_32009_13791.t4 14.282
R7519 a_32009_13791.n3 a_32009_13791.t2 14.282
R7520 a_32009_13791.n8 a_32009_13791.n1 1216.25
R7521 a_32009_13791.n1 a_32009_13791.t10 408.806
R7522 a_32009_13791.t9 a_32009_13791.n2 160.666
R7523 a_32009_13791.n1 a_32009_13791.t9 989.744
R7524 a_32009_13791.n2 a_32009_13791.t8 287.241
R7525 a_32009_13791.n2 a_32009_13791.t11 287.241
R7526 opcode[0].n5 opcode[0].n4 501.28
R7527 opcode[0].t17 opcode[0].t20 437.233
R7528 opcode[0].n56 opcode[0].n51 436.21
R7529 opcode[0].n50 opcode[0].n45 436.21
R7530 opcode[0].n44 opcode[0].n39 436.21
R7531 opcode[0].n38 opcode[0].n33 436.21
R7532 opcode[0].n32 opcode[0].n27 436.21
R7533 opcode[0].n26 opcode[0].n21 436.21
R7534 opcode[0].n20 opcode[0].n15 436.21
R7535 opcode[0].n14 opcode[0].n9 436.21
R7536 opcode[0].t76 opcode[0].t0 415.315
R7537 opcode[0].n54 opcode[0].t26 393.348
R7538 opcode[0].n48 opcode[0].t52 393.348
R7539 opcode[0].n42 opcode[0].t31 393.348
R7540 opcode[0].n36 opcode[0].t78 393.348
R7541 opcode[0].n30 opcode[0].t13 393.348
R7542 opcode[0].n24 opcode[0].t73 393.348
R7543 opcode[0].n18 opcode[0].t58 393.348
R7544 opcode[0].n12 opcode[0].t15 393.348
R7545 opcode[0].t12 opcode[0].n2 313.873
R7546 opcode[0].n4 opcode[0].t47 294.986
R7547 opcode[0].n51 opcode[0].t62 294.653
R7548 opcode[0].n45 opcode[0].t36 294.653
R7549 opcode[0].n39 opcode[0].t7 294.653
R7550 opcode[0].n33 opcode[0].t38 294.653
R7551 opcode[0].n27 opcode[0].t74 294.653
R7552 opcode[0].n21 opcode[0].t57 294.653
R7553 opcode[0].n15 opcode[0].t4 294.653
R7554 opcode[0].n9 opcode[0].t3 294.653
R7555 opcode[0].n1 opcode[0].t32 272.288
R7556 opcode[0].n53 opcode[0].t59 270.326
R7557 opcode[0].t26 opcode[0].n53 270.326
R7558 opcode[0].n47 opcode[0].t69 270.326
R7559 opcode[0].t52 opcode[0].n47 270.326
R7560 opcode[0].n41 opcode[0].t64 270.326
R7561 opcode[0].t31 opcode[0].n41 270.326
R7562 opcode[0].n35 opcode[0].t14 270.326
R7563 opcode[0].t78 opcode[0].n35 270.326
R7564 opcode[0].n29 opcode[0].t33 270.326
R7565 opcode[0].t13 opcode[0].n29 270.326
R7566 opcode[0].n23 opcode[0].t49 270.326
R7567 opcode[0].t73 opcode[0].n23 270.326
R7568 opcode[0].n17 opcode[0].t16 270.326
R7569 opcode[0].t58 opcode[0].n17 270.326
R7570 opcode[0].n11 opcode[0].t37 270.326
R7571 opcode[0].t15 opcode[0].n11 270.326
R7572 opcode[0].n56 opcode[0].n55 248.23
R7573 opcode[0].n50 opcode[0].n49 248.23
R7574 opcode[0].n44 opcode[0].n43 248.23
R7575 opcode[0].n38 opcode[0].n37 248.23
R7576 opcode[0].n32 opcode[0].n31 248.23
R7577 opcode[0].n26 opcode[0].n25 248.23
R7578 opcode[0].n20 opcode[0].n19 248.23
R7579 opcode[0].n14 opcode[0].n13 248.23
R7580 opcode[0].n5 opcode[0].t42 236.01
R7581 opcode[0].n8 opcode[0].t17 216.627
R7582 opcode[0].n6 opcode[0].t76 216.111
R7583 opcode[0].n7 opcode[0].t5 214.686
R7584 opcode[0].t20 opcode[0].n7 214.686
R7585 opcode[0].n0 opcode[0].t27 214.335
R7586 opcode[0].t0 opcode[0].n0 214.335
R7587 opcode[0].n52 opcode[0].t41 197.241
R7588 opcode[0].n46 opcode[0].t45 197.241
R7589 opcode[0].n40 opcode[0].t23 197.241
R7590 opcode[0].n34 opcode[0].t70 197.241
R7591 opcode[0].n28 opcode[0].t8 197.241
R7592 opcode[0].n22 opcode[0].t67 197.241
R7593 opcode[0].n16 opcode[0].t54 197.241
R7594 opcode[0].n10 opcode[0].t68 197.241
R7595 opcode[0].n3 opcode[0].t12 190.152
R7596 opcode[0].n3 opcode[0].t43 190.152
R7597 opcode[0].n1 opcode[0].t35 160.666
R7598 opcode[0].n2 opcode[0].t51 160.666
R7599 opcode[0].n53 opcode[0].t72 160.666
R7600 opcode[0].n47 opcode[0].t22 160.666
R7601 opcode[0].n41 opcode[0].t77 160.666
R7602 opcode[0].n35 opcode[0].t44 160.666
R7603 opcode[0].n29 opcode[0].t61 160.666
R7604 opcode[0].n23 opcode[0].t63 160.666
R7605 opcode[0].n17 opcode[0].t30 160.666
R7606 opcode[0].n11 opcode[0].t65 160.666
R7607 opcode[0].n6 opcode[0].n5 148.428
R7608 opcode[0].n57 opcode[0].n56 121.522
R7609 opcode[0].n63 opcode[0].n14 119.477
R7610 opcode[0].n62 opcode[0].n20 118.483
R7611 opcode[0].n59 opcode[0].n38 118.277
R7612 opcode[0].n60 opcode[0].n32 118.275
R7613 opcode[0].n61 opcode[0].n26 118.132
R7614 opcode[0].n57 opcode[0].n50 118.08
R7615 opcode[0].n58 opcode[0].n44 118.08
R7616 opcode[0].n51 opcode[0].t29 111.663
R7617 opcode[0].n45 opcode[0].t55 111.663
R7618 opcode[0].n39 opcode[0].t48 111.663
R7619 opcode[0].n33 opcode[0].t1 111.663
R7620 opcode[0].n27 opcode[0].t75 111.663
R7621 opcode[0].n21 opcode[0].t21 111.663
R7622 opcode[0].n15 opcode[0].t46 111.663
R7623 opcode[0].n9 opcode[0].t34 111.663
R7624 opcode[0].n4 opcode[0].t71 110.859
R7625 opcode[0].n55 opcode[0].n54 97.816
R7626 opcode[0].n49 opcode[0].n48 97.816
R7627 opcode[0].n43 opcode[0].n42 97.816
R7628 opcode[0].n37 opcode[0].n36 97.816
R7629 opcode[0].n31 opcode[0].n30 97.816
R7630 opcode[0].n25 opcode[0].n24 97.816
R7631 opcode[0].n19 opcode[0].n18 97.816
R7632 opcode[0].n13 opcode[0].n12 97.816
R7633 opcode[0].n2 opcode[0].n1 96.129
R7634 opcode[0].n52 opcode[0].t10 93.989
R7635 opcode[0].n46 opcode[0].t39 93.989
R7636 opcode[0].n40 opcode[0].t11 93.989
R7637 opcode[0].n34 opcode[0].t40 93.989
R7638 opcode[0].n28 opcode[0].t53 93.989
R7639 opcode[0].n22 opcode[0].t50 93.989
R7640 opcode[0].n16 opcode[0].t19 93.989
R7641 opcode[0].n10 opcode[0].t60 93.989
R7642 opcode[0].n7 opcode[0].t79 80.333
R7643 opcode[0].n0 opcode[0].t24 80.333
R7644 opcode[0].t42 opcode[0].n3 80.333
R7645 opcode[0].n54 opcode[0].t56 80.333
R7646 opcode[0].n48 opcode[0].t6 80.333
R7647 opcode[0].n42 opcode[0].t2 80.333
R7648 opcode[0].n36 opcode[0].t9 80.333
R7649 opcode[0].n30 opcode[0].t25 80.333
R7650 opcode[0].n24 opcode[0].t18 80.333
R7651 opcode[0].n18 opcode[0].t66 80.333
R7652 opcode[0].n12 opcode[0].t28 80.333
R7653 opcode[0].n64 opcode[0].n63 11.636
R7654 opcode[0].n55 opcode[0].n52 6.615
R7655 opcode[0].n49 opcode[0].n46 6.615
R7656 opcode[0].n43 opcode[0].n40 6.615
R7657 opcode[0].n37 opcode[0].n34 6.615
R7658 opcode[0].n31 opcode[0].n28 6.615
R7659 opcode[0].n25 opcode[0].n22 6.615
R7660 opcode[0].n19 opcode[0].n16 6.615
R7661 opcode[0].n13 opcode[0].n10 6.615
R7662 opcode[0].n63 opcode[0].n62 3.481
R7663 opcode[0].n60 opcode[0].n59 3.446
R7664 opcode[0].n58 opcode[0].n57 3.446
R7665 opcode[0].n59 opcode[0].n58 3.445
R7666 opcode[0].n61 opcode[0].n60 3.44
R7667 opcode[0].n62 opcode[0].n61 3.433
R7668 opcode[0].n64 opcode[0].n8 3.293
R7669 opcode[0].n8 opcode[0].n6 2.923
R7670 opcode[0] opcode[0].n64 2.149
R7671 a_5957_24166.n0 a_5957_24166.t9 214.335
R7672 a_5957_24166.t7 a_5957_24166.n0 214.335
R7673 a_5957_24166.n1 a_5957_24166.t7 143.851
R7674 a_5957_24166.n1 a_5957_24166.t10 135.658
R7675 a_5957_24166.n0 a_5957_24166.t8 80.333
R7676 a_5957_24166.n2 a_5957_24166.t0 28.565
R7677 a_5957_24166.n2 a_5957_24166.t1 28.565
R7678 a_5957_24166.n4 a_5957_24166.t2 28.565
R7679 a_5957_24166.n4 a_5957_24166.t6 28.565
R7680 a_5957_24166.n7 a_5957_24166.t5 28.565
R7681 a_5957_24166.t3 a_5957_24166.n7 28.565
R7682 a_5957_24166.n6 a_5957_24166.t4 9.714
R7683 a_5957_24166.n7 a_5957_24166.n6 1.003
R7684 a_5957_24166.n5 a_5957_24166.n3 0.833
R7685 a_5957_24166.n3 a_5957_24166.n2 0.653
R7686 a_5957_24166.n5 a_5957_24166.n4 0.653
R7687 a_5957_24166.n6 a_5957_24166.n5 0.341
R7688 a_5957_24166.n3 a_5957_24166.n1 0.032
R7689 a_36751_13711.t0 a_36751_13711.n9 104.259
R7690 a_36751_13711.n9 a_36751_13711.n2 77.784
R7691 a_36751_13711.n2 a_36751_13711.n4 77.456
R7692 a_36751_13711.n4 a_36751_13711.n6 77.456
R7693 a_36751_13711.n6 a_36751_13711.n7 75.815
R7694 a_36751_13711.n7 a_36751_13711.n8 167.433
R7695 a_36751_13711.n8 a_36751_13711.t5 14.282
R7696 a_36751_13711.n8 a_36751_13711.t4 14.282
R7697 a_36751_13711.n7 a_36751_13711.t3 104.259
R7698 a_36751_13711.n6 a_36751_13711.n5 89.977
R7699 a_36751_13711.n5 a_36751_13711.t8 14.282
R7700 a_36751_13711.n5 a_36751_13711.t6 14.282
R7701 a_36751_13711.n4 a_36751_13711.n3 89.977
R7702 a_36751_13711.n3 a_36751_13711.t9 14.282
R7703 a_36751_13711.n3 a_36751_13711.t7 14.282
R7704 a_36751_13711.n2 a_36751_13711.n1 89.977
R7705 a_36751_13711.n1 a_36751_13711.t10 14.282
R7706 a_36751_13711.n1 a_36751_13711.t11 14.282
R7707 a_36751_13711.n9 a_36751_13711.n0 167.433
R7708 a_36751_13711.n0 a_36751_13711.t1 14.282
R7709 a_36751_13711.n0 a_36751_13711.t2 14.282
R7710 a_20955_6381.n8 a_20955_6381.n7 861.987
R7711 a_20955_6381.n7 a_20955_6381.n6 560.726
R7712 a_20955_6381.t16 a_20955_6381.t10 415.315
R7713 a_20955_6381.t15 a_20955_6381.t7 415.315
R7714 a_20955_6381.n3 a_20955_6381.t13 394.151
R7715 a_20955_6381.n6 a_20955_6381.t6 294.653
R7716 a_20955_6381.n2 a_20955_6381.t4 269.523
R7717 a_20955_6381.t13 a_20955_6381.n2 269.523
R7718 a_20955_6381.n10 a_20955_6381.t16 217.716
R7719 a_20955_6381.n9 a_20955_6381.t19 214.335
R7720 a_20955_6381.t10 a_20955_6381.n9 214.335
R7721 a_20955_6381.n1 a_20955_6381.t18 214.335
R7722 a_20955_6381.t7 a_20955_6381.n1 214.335
R7723 a_20955_6381.n8 a_20955_6381.t15 198.921
R7724 a_20955_6381.n4 a_20955_6381.t17 198.043
R7725 a_20955_6381.n2 a_20955_6381.t14 160.666
R7726 a_20955_6381.n6 a_20955_6381.t5 111.663
R7727 a_20955_6381.n5 a_20955_6381.n3 97.816
R7728 a_20955_6381.n4 a_20955_6381.t8 93.989
R7729 a_20955_6381.n9 a_20955_6381.t12 80.333
R7730 a_20955_6381.n3 a_20955_6381.t9 80.333
R7731 a_20955_6381.n1 a_20955_6381.t11 80.333
R7732 a_20955_6381.n7 a_20955_6381.n5 65.07
R7733 a_20955_6381.n0 a_20955_6381.t3 28.57
R7734 a_20955_6381.t0 a_20955_6381.n12 28.565
R7735 a_20955_6381.n12 a_20955_6381.t1 28.565
R7736 a_20955_6381.n0 a_20955_6381.t2 17.638
R7737 a_20955_6381.n10 a_20955_6381.n8 16.411
R7738 a_20955_6381.n11 a_20955_6381.n10 7.315
R7739 a_20955_6381.n5 a_20955_6381.n4 6.615
R7740 a_20955_6381.n12 a_20955_6381.n11 0.69
R7741 a_20955_6381.n11 a_20955_6381.n0 0.6
R7742 a_25759_9997.t0 a_25759_9997.n7 16.058
R7743 a_25759_9997.n7 a_25759_9997.n5 0.575
R7744 a_25759_9997.n5 a_25759_9997.n9 0.2
R7745 a_25759_9997.n9 a_25759_9997.t10 16.058
R7746 a_25759_9997.n9 a_25759_9997.n8 0.999
R7747 a_25759_9997.n8 a_25759_9997.t9 14.282
R7748 a_25759_9997.n8 a_25759_9997.t4 14.282
R7749 a_25759_9997.n7 a_25759_9997.n6 0.999
R7750 a_25759_9997.n6 a_25759_9997.t2 14.282
R7751 a_25759_9997.n6 a_25759_9997.t1 14.282
R7752 a_25759_9997.n5 a_25759_9997.n3 0.227
R7753 a_25759_9997.n3 a_25759_9997.n4 1.511
R7754 a_25759_9997.n4 a_25759_9997.t7 14.282
R7755 a_25759_9997.n4 a_25759_9997.t6 14.282
R7756 a_25759_9997.n3 a_25759_9997.n0 0.669
R7757 a_25759_9997.n0 a_25759_9997.n1 0.001
R7758 a_25759_9997.n0 a_25759_9997.n2 267.767
R7759 a_25759_9997.n2 a_25759_9997.t3 14.282
R7760 a_25759_9997.n2 a_25759_9997.t11 14.282
R7761 a_25759_9997.n1 a_25759_9997.t8 14.282
R7762 a_25759_9997.n1 a_25759_9997.t5 14.282
R7763 a_13599_21654.t6 a_13599_21654.t7 800.071
R7764 a_13599_21654.n3 a_13599_21654.n2 659.095
R7765 a_13599_21654.n1 a_13599_21654.t4 285.109
R7766 a_13599_21654.n2 a_13599_21654.t6 193.602
R7767 a_13599_21654.n4 a_13599_21654.n0 192.754
R7768 a_13599_21654.n1 a_13599_21654.t5 160.666
R7769 a_13599_21654.n2 a_13599_21654.n1 91.507
R7770 a_13599_21654.t3 a_13599_21654.n4 28.568
R7771 a_13599_21654.n0 a_13599_21654.t1 28.565
R7772 a_13599_21654.n0 a_13599_21654.t2 28.565
R7773 a_13599_21654.n3 a_13599_21654.t0 19.063
R7774 a_13599_21654.n4 a_13599_21654.n3 1.005
R7775 a_17296_5412.n6 a_17296_5412.n5 501.28
R7776 a_17296_5412.t9 a_17296_5412.t5 437.233
R7777 a_17296_5412.t13 a_17296_5412.t8 415.315
R7778 a_17296_5412.t10 a_17296_5412.n3 313.873
R7779 a_17296_5412.n5 a_17296_5412.t6 294.986
R7780 a_17296_5412.n2 a_17296_5412.t15 272.288
R7781 a_17296_5412.n6 a_17296_5412.t11 236.01
R7782 a_17296_5412.n9 a_17296_5412.t9 216.627
R7783 a_17296_5412.n7 a_17296_5412.t13 216.111
R7784 a_17296_5412.n8 a_17296_5412.t4 214.686
R7785 a_17296_5412.t5 a_17296_5412.n8 214.686
R7786 a_17296_5412.n1 a_17296_5412.t14 214.335
R7787 a_17296_5412.t8 a_17296_5412.n1 214.335
R7788 a_17296_5412.n4 a_17296_5412.t10 190.152
R7789 a_17296_5412.n4 a_17296_5412.t16 190.152
R7790 a_17296_5412.n2 a_17296_5412.t7 160.666
R7791 a_17296_5412.n3 a_17296_5412.t17 160.666
R7792 a_17296_5412.n7 a_17296_5412.n6 148.428
R7793 a_17296_5412.n5 a_17296_5412.t19 110.859
R7794 a_17296_5412.n3 a_17296_5412.n2 96.129
R7795 a_17296_5412.n8 a_17296_5412.t12 80.333
R7796 a_17296_5412.n1 a_17296_5412.t18 80.333
R7797 a_17296_5412.t11 a_17296_5412.n4 80.333
R7798 a_17296_5412.n0 a_17296_5412.t1 28.57
R7799 a_17296_5412.n11 a_17296_5412.t3 28.565
R7800 a_17296_5412.t0 a_17296_5412.n11 28.565
R7801 a_17296_5412.n0 a_17296_5412.t2 17.638
R7802 a_17296_5412.n10 a_17296_5412.n9 6.64
R7803 a_17296_5412.n9 a_17296_5412.n7 2.923
R7804 a_17296_5412.n11 a_17296_5412.n10 0.69
R7805 a_17296_5412.n10 a_17296_5412.n0 0.6
R7806 a_17356_5438.n4 a_17356_5438.t10 214.335
R7807 a_17356_5438.t8 a_17356_5438.n4 214.335
R7808 a_17356_5438.n5 a_17356_5438.t8 143.851
R7809 a_17356_5438.n5 a_17356_5438.t9 135.658
R7810 a_17356_5438.n4 a_17356_5438.t7 80.333
R7811 a_17356_5438.n0 a_17356_5438.t4 28.565
R7812 a_17356_5438.n0 a_17356_5438.t6 28.565
R7813 a_17356_5438.n2 a_17356_5438.t1 28.565
R7814 a_17356_5438.n2 a_17356_5438.t5 28.565
R7815 a_17356_5438.n7 a_17356_5438.t0 28.565
R7816 a_17356_5438.t2 a_17356_5438.n7 28.565
R7817 a_17356_5438.n1 a_17356_5438.t3 9.714
R7818 a_17356_5438.n1 a_17356_5438.n0 1.003
R7819 a_17356_5438.n6 a_17356_5438.n3 0.833
R7820 a_17356_5438.n3 a_17356_5438.n2 0.653
R7821 a_17356_5438.n7 a_17356_5438.n6 0.653
R7822 a_17356_5438.n3 a_17356_5438.n1 0.341
R7823 a_17356_5438.n6 a_17356_5438.n5 0.032
R7824 a_1833_4076.n7 a_1833_4076.n6 861.987
R7825 a_1833_4076.n6 a_1833_4076.n5 560.726
R7826 a_1833_4076.t11 a_1833_4076.t6 415.315
R7827 a_1833_4076.t12 a_1833_4076.t7 415.315
R7828 a_1833_4076.n2 a_1833_4076.t5 394.151
R7829 a_1833_4076.n5 a_1833_4076.t17 294.653
R7830 a_1833_4076.n1 a_1833_4076.t10 269.523
R7831 a_1833_4076.t5 a_1833_4076.n1 269.523
R7832 a_1833_4076.n9 a_1833_4076.t11 217.716
R7833 a_1833_4076.n8 a_1833_4076.t8 214.335
R7834 a_1833_4076.t6 a_1833_4076.n8 214.335
R7835 a_1833_4076.n0 a_1833_4076.t13 214.335
R7836 a_1833_4076.t7 a_1833_4076.n0 214.335
R7837 a_1833_4076.n7 a_1833_4076.t12 198.921
R7838 a_1833_4076.n3 a_1833_4076.t9 198.043
R7839 a_1833_4076.n12 a_1833_4076.n11 192.754
R7840 a_1833_4076.n1 a_1833_4076.t16 160.666
R7841 a_1833_4076.n5 a_1833_4076.t19 111.663
R7842 a_1833_4076.n4 a_1833_4076.n2 97.816
R7843 a_1833_4076.n3 a_1833_4076.t4 93.989
R7844 a_1833_4076.n8 a_1833_4076.t14 80.333
R7845 a_1833_4076.n2 a_1833_4076.t15 80.333
R7846 a_1833_4076.n0 a_1833_4076.t18 80.333
R7847 a_1833_4076.n6 a_1833_4076.n4 65.07
R7848 a_1833_4076.n11 a_1833_4076.t2 28.568
R7849 a_1833_4076.t0 a_1833_4076.n12 28.565
R7850 a_1833_4076.n12 a_1833_4076.t1 28.565
R7851 a_1833_4076.n10 a_1833_4076.t3 18.825
R7852 a_1833_4076.n9 a_1833_4076.n7 16.411
R7853 a_1833_4076.n4 a_1833_4076.n3 6.615
R7854 a_1833_4076.n10 a_1833_4076.n9 2.988
R7855 a_1833_4076.n11 a_1833_4076.n10 1.105
R7856 a_5496_4822.n1 a_5496_4822.t5 318.922
R7857 a_5496_4822.n0 a_5496_4822.t6 273.935
R7858 a_5496_4822.n0 a_5496_4822.t7 273.935
R7859 a_5496_4822.n1 a_5496_4822.t4 269.116
R7860 a_5496_4822.n4 a_5496_4822.n3 193.227
R7861 a_5496_4822.t5 a_5496_4822.n0 179.142
R7862 a_5496_4822.n2 a_5496_4822.n1 106.999
R7863 a_5496_4822.n3 a_5496_4822.t2 28.568
R7864 a_5496_4822.n4 a_5496_4822.t1 28.565
R7865 a_5496_4822.t3 a_5496_4822.n4 28.565
R7866 a_5496_4822.n2 a_5496_4822.t0 18.149
R7867 a_5496_4822.n3 a_5496_4822.n2 3.726
R7868 a_1836_10114.n7 a_1836_10114.n6 861.987
R7869 a_1836_10114.n6 a_1836_10114.n5 560.726
R7870 a_1836_10114.t12 a_1836_10114.t4 415.315
R7871 a_1836_10114.t11 a_1836_10114.t14 415.315
R7872 a_1836_10114.n2 a_1836_10114.t16 394.151
R7873 a_1836_10114.n5 a_1836_10114.t19 294.653
R7874 a_1836_10114.n1 a_1836_10114.t18 269.523
R7875 a_1836_10114.t16 a_1836_10114.n1 269.523
R7876 a_1836_10114.n9 a_1836_10114.t12 217.716
R7877 a_1836_10114.n8 a_1836_10114.t7 214.335
R7878 a_1836_10114.t4 a_1836_10114.n8 214.335
R7879 a_1836_10114.n0 a_1836_10114.t6 214.335
R7880 a_1836_10114.t14 a_1836_10114.n0 214.335
R7881 a_1836_10114.n7 a_1836_10114.t11 198.921
R7882 a_1836_10114.n3 a_1836_10114.t8 198.043
R7883 a_1836_10114.n12 a_1836_10114.n11 192.754
R7884 a_1836_10114.n1 a_1836_10114.t17 160.666
R7885 a_1836_10114.n5 a_1836_10114.t10 111.663
R7886 a_1836_10114.n4 a_1836_10114.n2 97.816
R7887 a_1836_10114.n3 a_1836_10114.t9 93.989
R7888 a_1836_10114.n8 a_1836_10114.t5 80.333
R7889 a_1836_10114.n2 a_1836_10114.t13 80.333
R7890 a_1836_10114.n0 a_1836_10114.t15 80.333
R7891 a_1836_10114.n6 a_1836_10114.n4 65.07
R7892 a_1836_10114.n11 a_1836_10114.t1 28.568
R7893 a_1836_10114.n12 a_1836_10114.t2 28.565
R7894 a_1836_10114.t3 a_1836_10114.n12 28.565
R7895 a_1836_10114.n10 a_1836_10114.t0 18.825
R7896 a_1836_10114.n9 a_1836_10114.n7 16.411
R7897 a_1836_10114.n4 a_1836_10114.n3 6.615
R7898 a_1836_10114.n10 a_1836_10114.n9 2.757
R7899 a_1836_10114.n11 a_1836_10114.n10 1.105
R7900 a_4144_12869.n0 a_4144_12869.t10 214.335
R7901 a_4144_12869.t8 a_4144_12869.n0 214.335
R7902 a_4144_12869.n1 a_4144_12869.t8 143.851
R7903 a_4144_12869.n1 a_4144_12869.t7 135.658
R7904 a_4144_12869.n0 a_4144_12869.t9 80.333
R7905 a_4144_12869.n2 a_4144_12869.t0 28.565
R7906 a_4144_12869.n2 a_4144_12869.t1 28.565
R7907 a_4144_12869.n4 a_4144_12869.t2 28.565
R7908 a_4144_12869.n4 a_4144_12869.t6 28.565
R7909 a_4144_12869.n7 a_4144_12869.t5 28.565
R7910 a_4144_12869.t4 a_4144_12869.n7 28.565
R7911 a_4144_12869.n6 a_4144_12869.t3 9.714
R7912 a_4144_12869.n7 a_4144_12869.n6 1.003
R7913 a_4144_12869.n5 a_4144_12869.n3 0.833
R7914 a_4144_12869.n3 a_4144_12869.n2 0.653
R7915 a_4144_12869.n5 a_4144_12869.n4 0.653
R7916 a_4144_12869.n6 a_4144_12869.n5 0.341
R7917 a_4144_12869.n3 a_4144_12869.n1 0.032
R7918 a_12475_25767.n0 a_12475_25767.t7 214.335
R7919 a_12475_25767.t9 a_12475_25767.n0 214.335
R7920 a_12475_25767.n1 a_12475_25767.t9 143.851
R7921 a_12475_25767.n1 a_12475_25767.t8 135.658
R7922 a_12475_25767.n0 a_12475_25767.t10 80.333
R7923 a_12475_25767.n2 a_12475_25767.t5 28.565
R7924 a_12475_25767.n2 a_12475_25767.t4 28.565
R7925 a_12475_25767.n4 a_12475_25767.t3 28.565
R7926 a_12475_25767.n4 a_12475_25767.t2 28.565
R7927 a_12475_25767.n7 a_12475_25767.t1 28.565
R7928 a_12475_25767.t0 a_12475_25767.n7 28.565
R7929 a_12475_25767.n6 a_12475_25767.t6 9.714
R7930 a_12475_25767.n7 a_12475_25767.n6 1.003
R7931 a_12475_25767.n5 a_12475_25767.n3 0.833
R7932 a_12475_25767.n3 a_12475_25767.n2 0.653
R7933 a_12475_25767.n5 a_12475_25767.n4 0.653
R7934 a_12475_25767.n6 a_12475_25767.n5 0.341
R7935 a_12475_25767.n3 a_12475_25767.n1 0.032
R7936 a_13065_25330.t6 a_13065_25330.t5 574.43
R7937 a_13065_25330.n1 a_13065_25330.t4 285.109
R7938 a_13065_25330.n3 a_13065_25330.n2 211.136
R7939 a_13065_25330.n4 a_13065_25330.n0 192.754
R7940 a_13065_25330.n1 a_13065_25330.t7 160.666
R7941 a_13065_25330.n2 a_13065_25330.t6 160.666
R7942 a_13065_25330.n2 a_13065_25330.n1 114.829
R7943 a_13065_25330.t3 a_13065_25330.n4 28.568
R7944 a_13065_25330.n0 a_13065_25330.t1 28.565
R7945 a_13065_25330.n0 a_13065_25330.t2 28.565
R7946 a_13065_25330.n3 a_13065_25330.t0 19.084
R7947 a_13065_25330.n4 a_13065_25330.n3 1.051
R7948 a_14784_4101.n1 a_14784_4101.t5 318.922
R7949 a_14784_4101.n0 a_14784_4101.t7 274.739
R7950 a_14784_4101.n0 a_14784_4101.t6 274.739
R7951 a_14784_4101.n1 a_14784_4101.t4 269.116
R7952 a_14784_4101.t5 a_14784_4101.n0 179.946
R7953 a_14784_4101.n2 a_14784_4101.n1 105.178
R7954 a_14784_4101.t3 a_14784_4101.n4 29.444
R7955 a_14784_4101.n3 a_14784_4101.t2 28.565
R7956 a_14784_4101.n3 a_14784_4101.t1 28.565
R7957 a_14784_4101.n2 a_14784_4101.t0 18.145
R7958 a_14784_4101.n4 a_14784_4101.n2 2.878
R7959 a_14784_4101.n4 a_14784_4101.n3 0.764
R7960 a_14490_3395.t0 a_14490_3395.t1 380.209
R7961 A[4].n16 A[4].n6 1956.22
R7962 A[4].n6 A[4].n4 1494.07
R7963 A[4].n11 A[4].n10 535.449
R7964 A[4].t1 A[4].t3 437.233
R7965 A[4].t28 A[4].t29 437.233
R7966 A[4].t26 A[4].t20 437.233
R7967 A[4].t31 A[4].t2 437.233
R7968 A[4].t8 A[4].t21 437.233
R7969 A[4].t30 A[4].t24 415.315
R7970 A[4].t13 A[4].n8 313.873
R7971 A[4].n10 A[4].t17 294.986
R7972 A[4].n7 A[4].t14 272.288
R7973 A[4].n11 A[4].t11 245.184
R7974 A[4].n3 A[4].t28 224.833
R7975 A[4].n4 A[4].t30 219.944
R7976 A[4].n13 A[4].t8 218.627
R7977 A[4].n6 A[4].t26 217.054
R7978 A[4].n15 A[4].t31 217.023
R7979 A[4].n3 A[4].t1 216.198
R7980 A[4].n2 A[4].t27 214.686
R7981 A[4].t3 A[4].n2 214.686
R7982 A[4].n1 A[4].t18 214.686
R7983 A[4].t29 A[4].n1 214.686
R7984 A[4].n5 A[4].t7 214.686
R7985 A[4].t20 A[4].n5 214.686
R7986 A[4].n14 A[4].t5 214.686
R7987 A[4].t2 A[4].n14 214.686
R7988 A[4].n12 A[4].t23 214.686
R7989 A[4].t21 A[4].n12 214.686
R7990 A[4].n0 A[4].t0 214.335
R7991 A[4].t24 A[4].n0 214.335
R7992 A[4].n9 A[4].t9 190.152
R7993 A[4].n9 A[4].t13 190.152
R7994 A[4].n7 A[4].t12 160.666
R7995 A[4].n8 A[4].t10 160.666
R7996 A[4].n10 A[4].t25 110.859
R7997 A[4].n8 A[4].n7 96.129
R7998 A[4].n0 A[4].t15 80.333
R7999 A[4].n2 A[4].t16 80.333
R8000 A[4].n1 A[4].t6 80.333
R8001 A[4].n5 A[4].t19 80.333
R8002 A[4].n14 A[4].t4 80.333
R8003 A[4].t11 A[4].n9 80.333
R8004 A[4].n12 A[4].t22 80.333
R8005 A[4].n16 A[4].n15 53.076
R8006 A[4].n4 A[4].n3 34.046
R8007 A[4].n13 A[4].n11 14.9
R8008 A[4] A[4].n16 2.676
R8009 A[4].n15 A[4].n13 2.599
R8010 a_16264_24457.n0 a_16264_24457.n8 122.999
R8011 a_16264_24457.t1 a_16264_24457.n0 14.282
R8012 a_16264_24457.n0 a_16264_24457.t2 14.282
R8013 a_16264_24457.n8 a_16264_24457.n6 50.575
R8014 a_16264_24457.n6 a_16264_24457.n4 74.302
R8015 a_16264_24457.n8 a_16264_24457.n7 157.665
R8016 a_16264_24457.n7 a_16264_24457.t4 8.7
R8017 a_16264_24457.n7 a_16264_24457.t0 8.7
R8018 a_16264_24457.n6 a_16264_24457.n5 90.416
R8019 a_16264_24457.n5 a_16264_24457.t3 14.282
R8020 a_16264_24457.n5 a_16264_24457.t5 14.282
R8021 a_16264_24457.n4 a_16264_24457.n3 90.436
R8022 a_16264_24457.n3 a_16264_24457.t6 14.282
R8023 a_16264_24457.n3 a_16264_24457.t7 14.282
R8024 a_16264_24457.n4 a_16264_24457.n1 2011.09
R8025 a_16264_24457.t9 a_16264_24457.n2 160.666
R8026 a_16264_24457.n1 a_16264_24457.t9 867.393
R8027 a_16264_24457.n2 a_16264_24457.t10 287.241
R8028 a_16264_24457.n2 a_16264_24457.t11 287.241
R8029 a_16264_24457.n1 a_16264_24457.t8 545.094
R8030 a_38088_20578.t0 a_38088_20578.t1 17.4
R8031 a_n3606_7699.n1 a_n3606_7699.t5 318.119
R8032 a_n3606_7699.n1 a_n3606_7699.t7 269.919
R8033 a_n3606_7699.n0 a_n3606_7699.t6 267.256
R8034 a_n3606_7699.n0 a_n3606_7699.t4 267.256
R8035 a_n3606_7699.n4 a_n3606_7699.n3 193.227
R8036 a_n3606_7699.t5 a_n3606_7699.n0 160.666
R8037 a_n3606_7699.n2 a_n3606_7699.n1 106.999
R8038 a_n3606_7699.n3 a_n3606_7699.t1 28.568
R8039 a_n3606_7699.n4 a_n3606_7699.t2 28.565
R8040 a_n3606_7699.t3 a_n3606_7699.n4 28.565
R8041 a_n3606_7699.n2 a_n3606_7699.t0 18.149
R8042 a_n3606_7699.n3 a_n3606_7699.n2 3.726
R8043 a_13051_26980.t6 a_13051_26980.t7 800.071
R8044 a_13051_26980.n3 a_13051_26980.n2 659.097
R8045 a_13051_26980.n1 a_13051_26980.t5 285.109
R8046 a_13051_26980.n2 a_13051_26980.t6 193.602
R8047 a_13051_26980.n4 a_13051_26980.n0 192.754
R8048 a_13051_26980.n1 a_13051_26980.t4 160.666
R8049 a_13051_26980.n2 a_13051_26980.n1 91.507
R8050 a_13051_26980.t0 a_13051_26980.n4 28.568
R8051 a_13051_26980.n0 a_13051_26980.t3 28.565
R8052 a_13051_26980.n0 a_13051_26980.t1 28.565
R8053 a_13051_26980.n3 a_13051_26980.t2 19.061
R8054 a_13051_26980.n4 a_13051_26980.n3 1.005
R8055 a_14786_27289.n0 a_14786_27289.t0 14.282
R8056 a_14786_27289.n0 a_14786_27289.t4 14.282
R8057 a_14786_27289.n1 a_14786_27289.t1 14.282
R8058 a_14786_27289.n1 a_14786_27289.t2 14.282
R8059 a_14786_27289.n3 a_14786_27289.t5 14.282
R8060 a_14786_27289.t3 a_14786_27289.n3 14.282
R8061 a_14786_27289.n3 a_14786_27289.n2 2.546
R8062 a_14786_27289.n2 a_14786_27289.n1 2.367
R8063 a_14786_27289.n2 a_14786_27289.n0 0.001
R8064 a_21439_4102.n1 a_21439_4102.t4 318.922
R8065 a_21439_4102.n0 a_21439_4102.t5 274.739
R8066 a_21439_4102.n0 a_21439_4102.t6 274.739
R8067 a_21439_4102.n1 a_21439_4102.t7 269.116
R8068 a_21439_4102.t4 a_21439_4102.n0 179.946
R8069 a_21439_4102.n2 a_21439_4102.n1 105.178
R8070 a_21439_4102.n3 a_21439_4102.t1 29.444
R8071 a_21439_4102.n4 a_21439_4102.t2 28.565
R8072 a_21439_4102.t3 a_21439_4102.n4 28.565
R8073 a_21439_4102.n2 a_21439_4102.t0 18.145
R8074 a_21439_4102.n3 a_21439_4102.n2 2.878
R8075 a_21439_4102.n4 a_21439_4102.n3 0.764
R8076 a_21027_4128.t0 a_21027_4128.n0 14.282
R8077 a_21027_4128.n0 a_21027_4128.t5 14.282
R8078 a_21027_4128.n0 a_21027_4128.n9 0.999
R8079 a_21027_4128.n9 a_21027_4128.n6 0.575
R8080 a_21027_4128.n6 a_21027_4128.n8 0.2
R8081 a_21027_4128.n8 a_21027_4128.t9 16.058
R8082 a_21027_4128.n8 a_21027_4128.n7 0.999
R8083 a_21027_4128.n7 a_21027_4128.t10 14.282
R8084 a_21027_4128.n7 a_21027_4128.t11 14.282
R8085 a_21027_4128.n9 a_21027_4128.t4 16.058
R8086 a_21027_4128.n6 a_21027_4128.n4 0.227
R8087 a_21027_4128.n4 a_21027_4128.n5 1.511
R8088 a_21027_4128.n5 a_21027_4128.t6 14.282
R8089 a_21027_4128.n5 a_21027_4128.t8 14.282
R8090 a_21027_4128.n4 a_21027_4128.n1 0.669
R8091 a_21027_4128.n1 a_21027_4128.n2 0.001
R8092 a_21027_4128.n1 a_21027_4128.n3 267.767
R8093 a_21027_4128.n3 a_21027_4128.t3 14.282
R8094 a_21027_4128.n3 a_21027_4128.t1 14.282
R8095 a_21027_4128.n2 a_21027_4128.t7 14.282
R8096 a_21027_4128.n2 a_21027_4128.t2 14.282
R8097 a_21145_4128.n0 a_21145_4128.t2 14.282
R8098 a_21145_4128.t1 a_21145_4128.n0 14.282
R8099 a_21145_4128.n0 a_21145_4128.n15 122.999
R8100 a_21145_4128.n15 a_21145_4128.n13 50.575
R8101 a_21145_4128.n13 a_21145_4128.n11 74.302
R8102 a_21145_4128.n15 a_21145_4128.n14 157.665
R8103 a_21145_4128.n14 a_21145_4128.t0 8.7
R8104 a_21145_4128.n14 a_21145_4128.t4 8.7
R8105 a_21145_4128.n13 a_21145_4128.n12 90.416
R8106 a_21145_4128.n12 a_21145_4128.t3 14.282
R8107 a_21145_4128.n12 a_21145_4128.t6 14.282
R8108 a_21145_4128.n11 a_21145_4128.n10 90.436
R8109 a_21145_4128.n10 a_21145_4128.t7 14.282
R8110 a_21145_4128.n10 a_21145_4128.t5 14.282
R8111 a_21145_4128.n11 a_21145_4128.n9 220.49
R8112 a_21145_4128.n9 a_21145_4128.n2 2.599
R8113 a_21145_4128.n2 a_21145_4128.t16 218.628
R8114 a_21145_4128.t16 a_21145_4128.t8 437.233
R8115 a_21145_4128.t8 a_21145_4128.n8 214.686
R8116 a_21145_4128.n8 a_21145_4128.t18 80.333
R8117 a_21145_4128.n8 a_21145_4128.t17 214.686
R8118 a_21145_4128.n2 a_21145_4128.n3 14.9
R8119 a_21145_4128.n3 a_21145_4128.n7 535.449
R8120 a_21145_4128.n7 a_21145_4128.t12 294.986
R8121 a_21145_4128.n7 a_21145_4128.t11 110.859
R8122 a_21145_4128.n3 a_21145_4128.t9 245.184
R8123 a_21145_4128.t9 a_21145_4128.n6 80.333
R8124 a_21145_4128.n6 a_21145_4128.t14 190.152
R8125 a_21145_4128.n6 a_21145_4128.t13 190.152
R8126 a_21145_4128.t13 a_21145_4128.n5 313.873
R8127 a_21145_4128.n5 a_21145_4128.t23 160.666
R8128 a_21145_4128.n5 a_21145_4128.n4 96.129
R8129 a_21145_4128.n4 a_21145_4128.t10 160.666
R8130 a_21145_4128.n4 a_21145_4128.t19 272.288
R8131 a_21145_4128.n9 a_21145_4128.t20 217.024
R8132 a_21145_4128.t20 a_21145_4128.t15 437.233
R8133 a_21145_4128.t15 a_21145_4128.n1 214.686
R8134 a_21145_4128.n1 a_21145_4128.t22 80.333
R8135 a_21145_4128.n1 a_21145_4128.t21 214.686
R8136 a_n3113_6918.t1 a_n3113_6918.n0 14.282
R8137 a_n3113_6918.n0 a_n3113_6918.t6 14.282
R8138 a_n3113_6918.n0 a_n3113_6918.n16 90.416
R8139 a_n3113_6918.n16 a_n3113_6918.n2 74.302
R8140 a_n3113_6918.n16 a_n3113_6918.n4 50.575
R8141 a_n3113_6918.n4 a_n3113_6918.n5 110.084
R8142 a_n3113_6918.n2 a_n3113_6918.n6 213.889
R8143 a_n3113_6918.n6 a_n3113_6918.n8 16.411
R8144 a_n3113_6918.n8 a_n3113_6918.t21 198.921
R8145 a_n3113_6918.t21 a_n3113_6918.t20 415.315
R8146 a_n3113_6918.t20 a_n3113_6918.n15 214.335
R8147 a_n3113_6918.n15 a_n3113_6918.t19 80.333
R8148 a_n3113_6918.n15 a_n3113_6918.t23 214.335
R8149 a_n3113_6918.n8 a_n3113_6918.n14 861.987
R8150 a_n3113_6918.n14 a_n3113_6918.n9 560.726
R8151 a_n3113_6918.n14 a_n3113_6918.n13 65.07
R8152 a_n3113_6918.n13 a_n3113_6918.n12 6.615
R8153 a_n3113_6918.n12 a_n3113_6918.t11 93.989
R8154 a_n3113_6918.n12 a_n3113_6918.t9 198.043
R8155 a_n3113_6918.n13 a_n3113_6918.n11 97.816
R8156 a_n3113_6918.n11 a_n3113_6918.t10 80.333
R8157 a_n3113_6918.n11 a_n3113_6918.t17 394.151
R8158 a_n3113_6918.t17 a_n3113_6918.n10 269.523
R8159 a_n3113_6918.n10 a_n3113_6918.t14 160.666
R8160 a_n3113_6918.n10 a_n3113_6918.t13 269.523
R8161 a_n3113_6918.n9 a_n3113_6918.t15 294.653
R8162 a_n3113_6918.n9 a_n3113_6918.t12 111.663
R8163 a_n3113_6918.n6 a_n3113_6918.t22 217.716
R8164 a_n3113_6918.t22 a_n3113_6918.t8 415.315
R8165 a_n3113_6918.t8 a_n3113_6918.n7 214.335
R8166 a_n3113_6918.n7 a_n3113_6918.t18 80.333
R8167 a_n3113_6918.n7 a_n3113_6918.t16 214.335
R8168 a_n3113_6918.n5 a_n3113_6918.t5 14.282
R8169 a_n3113_6918.n5 a_n3113_6918.t4 14.282
R8170 a_n3113_6918.n4 a_n3113_6918.n3 157.665
R8171 a_n3113_6918.n3 a_n3113_6918.t0 8.7
R8172 a_n3113_6918.n3 a_n3113_6918.t7 8.7
R8173 a_n3113_6918.n2 a_n3113_6918.n1 90.436
R8174 a_n3113_6918.n1 a_n3113_6918.t2 14.282
R8175 a_n3113_6918.n1 a_n3113_6918.t3 14.282
R8176 a_28617_21790.n0 a_28617_21790.t8 214.335
R8177 a_28617_21790.t10 a_28617_21790.n0 214.335
R8178 a_28617_21790.n1 a_28617_21790.t10 143.851
R8179 a_28617_21790.n1 a_28617_21790.t7 135.658
R8180 a_28617_21790.n0 a_28617_21790.t9 80.333
R8181 a_28617_21790.n4 a_28617_21790.t1 28.565
R8182 a_28617_21790.n4 a_28617_21790.t2 28.565
R8183 a_28617_21790.n2 a_28617_21790.t4 28.565
R8184 a_28617_21790.n2 a_28617_21790.t5 28.565
R8185 a_28617_21790.t3 a_28617_21790.n7 28.565
R8186 a_28617_21790.n7 a_28617_21790.t6 28.565
R8187 a_28617_21790.n5 a_28617_21790.t0 9.714
R8188 a_28617_21790.n5 a_28617_21790.n4 1.003
R8189 a_28617_21790.n6 a_28617_21790.n3 0.833
R8190 a_28617_21790.n3 a_28617_21790.n2 0.653
R8191 a_28617_21790.n7 a_28617_21790.n6 0.653
R8192 a_28617_21790.n6 a_28617_21790.n5 0.341
R8193 a_28617_21790.n3 a_28617_21790.n1 0.032
R8194 a_12475_18822.n1 a_12475_18822.t5 318.922
R8195 a_12475_18822.n0 a_12475_18822.t4 273.935
R8196 a_12475_18822.n0 a_12475_18822.t6 273.935
R8197 a_12475_18822.n1 a_12475_18822.t7 269.116
R8198 a_12475_18822.n4 a_12475_18822.n3 193.227
R8199 a_12475_18822.t5 a_12475_18822.n0 179.142
R8200 a_12475_18822.n2 a_12475_18822.n1 106.999
R8201 a_12475_18822.n3 a_12475_18822.t2 28.568
R8202 a_12475_18822.t0 a_12475_18822.n4 28.565
R8203 a_12475_18822.n4 a_12475_18822.t1 28.565
R8204 a_12475_18822.n2 a_12475_18822.t3 18.149
R8205 a_12475_18822.n3 a_12475_18822.n2 3.726
R8206 opcode[1].n11 opcode[1].t8 1374.48
R8207 opcode[1].n6 opcode[1].t41 1374.48
R8208 opcode[1].n1 opcode[1].t60 1374.48
R8209 opcode[1].n23 opcode[1].t10 1374.48
R8210 opcode[1].n28 opcode[1].t61 1374.48
R8211 opcode[1].n33 opcode[1].t59 1374.48
R8212 opcode[1].n42 opcode[1].t38 1374.48
R8213 opcode[1].n48 opcode[1].t52 1374.48
R8214 opcode[1].n14 opcode[1].t57 622.488
R8215 opcode[1].n8 opcode[1].t55 622.488
R8216 opcode[1].n3 opcode[1].t29 622.488
R8217 opcode[1].n25 opcode[1].t46 622.488
R8218 opcode[1].n30 opcode[1].t36 622.488
R8219 opcode[1].n35 opcode[1].t33 622.488
R8220 opcode[1].n38 opcode[1].t13 622.488
R8221 opcode[1].n50 opcode[1].t30 622.488
R8222 opcode[1].n14 opcode[1].t34 610.283
R8223 opcode[1].n8 opcode[1].t54 610.283
R8224 opcode[1].n3 opcode[1].t11 610.283
R8225 opcode[1].n25 opcode[1].t27 610.283
R8226 opcode[1].n30 opcode[1].t17 610.283
R8227 opcode[1].n35 opcode[1].t9 610.283
R8228 opcode[1].n38 opcode[1].t53 610.283
R8229 opcode[1].n50 opcode[1].t63 610.283
R8230 opcode[1].n11 opcode[1].t5 325.68
R8231 opcode[1].n6 opcode[1].t21 325.68
R8232 opcode[1].n1 opcode[1].t40 325.68
R8233 opcode[1].n23 opcode[1].t56 325.68
R8234 opcode[1].n28 opcode[1].t47 325.68
R8235 opcode[1].n33 opcode[1].t28 325.68
R8236 opcode[1].n42 opcode[1].t2 325.68
R8237 opcode[1].n48 opcode[1].t26 325.68
R8238 opcode[1].n13 opcode[1].t22 287.241
R8239 opcode[1].n13 opcode[1].t32 287.241
R8240 opcode[1].n7 opcode[1].t20 287.241
R8241 opcode[1].n7 opcode[1].t50 287.241
R8242 opcode[1].n2 opcode[1].t39 287.241
R8243 opcode[1].n2 opcode[1].t0 287.241
R8244 opcode[1].n24 opcode[1].t6 287.241
R8245 opcode[1].n24 opcode[1].t23 287.241
R8246 opcode[1].n29 opcode[1].t43 287.241
R8247 opcode[1].n29 opcode[1].t7 287.241
R8248 opcode[1].n34 opcode[1].t45 287.241
R8249 opcode[1].n34 opcode[1].t3 287.241
R8250 opcode[1].n37 opcode[1].t37 287.241
R8251 opcode[1].n37 opcode[1].t49 287.241
R8252 opcode[1].n49 opcode[1].t35 287.241
R8253 opcode[1].n49 opcode[1].t1 287.241
R8254 opcode[1].n10 opcode[1].t19 207.225
R8255 opcode[1].t5 opcode[1].n10 207.225
R8256 opcode[1].n5 opcode[1].t51 207.225
R8257 opcode[1].t21 opcode[1].n5 207.225
R8258 opcode[1].n0 opcode[1].t4 207.225
R8259 opcode[1].t40 opcode[1].n0 207.225
R8260 opcode[1].n22 opcode[1].t24 207.225
R8261 opcode[1].t56 opcode[1].n22 207.225
R8262 opcode[1].n27 opcode[1].t14 207.225
R8263 opcode[1].t47 opcode[1].n27 207.225
R8264 opcode[1].n32 opcode[1].t58 207.225
R8265 opcode[1].t28 opcode[1].n32 207.225
R8266 opcode[1].n41 opcode[1].t18 207.225
R8267 opcode[1].t2 opcode[1].n41 207.225
R8268 opcode[1].n47 opcode[1].t48 207.225
R8269 opcode[1].t26 opcode[1].n47 207.225
R8270 opcode[1].t57 opcode[1].n13 160.666
R8271 opcode[1].t55 opcode[1].n7 160.666
R8272 opcode[1].t29 opcode[1].n2 160.666
R8273 opcode[1].t46 opcode[1].n24 160.666
R8274 opcode[1].t36 opcode[1].n29 160.666
R8275 opcode[1].t33 opcode[1].n34 160.666
R8276 opcode[1].t13 opcode[1].n37 160.666
R8277 opcode[1].t30 opcode[1].n49 160.666
R8278 opcode[1].n10 opcode[1].t42 80.333
R8279 opcode[1].n5 opcode[1].t15 80.333
R8280 opcode[1].n0 opcode[1].t16 80.333
R8281 opcode[1].n22 opcode[1].t31 80.333
R8282 opcode[1].n27 opcode[1].t25 80.333
R8283 opcode[1].n32 opcode[1].t62 80.333
R8284 opcode[1].n41 opcode[1].t44 80.333
R8285 opcode[1].n47 opcode[1].t12 80.333
R8286 opcode[1] opcode[1].n56 56.443
R8287 opcode[1].n52 opcode[1].n51 7.802
R8288 opcode[1].n20 opcode[1].n19 7.174
R8289 opcode[1].n54 opcode[1].n31 4.102
R8290 opcode[1].n53 opcode[1].n36 4.1
R8291 opcode[1].n20 opcode[1].n9 4.052
R8292 opcode[1].n21 opcode[1].n4 4.046
R8293 opcode[1].n55 opcode[1].n26 3.999
R8294 opcode[1].n52 opcode[1].n46 3.828
R8295 opcode[1].n55 opcode[1].n54 3.777
R8296 opcode[1].n54 opcode[1].n53 3.707
R8297 opcode[1].n21 opcode[1].n20 3.693
R8298 opcode[1].n53 opcode[1].n52 3.693
R8299 opcode[1].n56 opcode[1].n21 3.625
R8300 opcode[1].n15 opcode[1].n14 2.07
R8301 opcode[1].n39 opcode[1].n38 1.715
R8302 opcode[1].n9 opcode[1].n8 1.614
R8303 opcode[1].n4 opcode[1].n3 1.614
R8304 opcode[1].n26 opcode[1].n25 1.614
R8305 opcode[1].n31 opcode[1].n30 1.614
R8306 opcode[1].n36 opcode[1].n35 1.614
R8307 opcode[1].n51 opcode[1].n50 1.614
R8308 opcode[1].n46 opcode[1].n45 0.243
R8309 opcode[1].n19 opcode[1].n18 0.236
R8310 opcode[1].n18 opcode[1].n17 0.086
R8311 opcode[1].n56 opcode[1].n55 0.08
R8312 opcode[1].n45 opcode[1].n44 0.056
R8313 opcode[1].n9 opcode[1].n6 0.003
R8314 opcode[1].n4 opcode[1].n1 0.003
R8315 opcode[1].n26 opcode[1].n23 0.003
R8316 opcode[1].n31 opcode[1].n28 0.003
R8317 opcode[1].n36 opcode[1].n33 0.003
R8318 opcode[1].n51 opcode[1].n48 0.003
R8319 opcode[1].n17 opcode[1].n16 0.002
R8320 opcode[1].n44 opcode[1].n40 0.002
R8321 opcode[1].n12 opcode[1].n11 0.001
R8322 opcode[1].n43 opcode[1].n42 0.001
R8323 opcode[1].n40 opcode[1].n39 0.001
R8324 opcode[1].n16 opcode[1].n15 0.001
R8325 opcode[1].n17 opcode[1].n12 0.001
R8326 opcode[1].n44 opcode[1].n43 0.001
R8327 a_36751_16855.t0 a_36751_16855.n9 104.259
R8328 a_36751_16855.n9 a_36751_16855.n2 77.784
R8329 a_36751_16855.n2 a_36751_16855.n4 77.456
R8330 a_36751_16855.n4 a_36751_16855.n6 77.456
R8331 a_36751_16855.n6 a_36751_16855.n7 75.815
R8332 a_36751_16855.n7 a_36751_16855.n8 167.433
R8333 a_36751_16855.n8 a_36751_16855.t3 14.282
R8334 a_36751_16855.n8 a_36751_16855.t2 14.282
R8335 a_36751_16855.n7 a_36751_16855.t4 104.259
R8336 a_36751_16855.n6 a_36751_16855.n5 89.977
R8337 a_36751_16855.n5 a_36751_16855.t9 14.282
R8338 a_36751_16855.n5 a_36751_16855.t10 14.282
R8339 a_36751_16855.n4 a_36751_16855.n3 89.977
R8340 a_36751_16855.n3 a_36751_16855.t5 14.282
R8341 a_36751_16855.n3 a_36751_16855.t11 14.282
R8342 a_36751_16855.n2 a_36751_16855.n1 89.977
R8343 a_36751_16855.n1 a_36751_16855.t7 14.282
R8344 a_36751_16855.n1 a_36751_16855.t6 14.282
R8345 a_36751_16855.n9 a_36751_16855.n0 167.433
R8346 a_36751_16855.n0 a_36751_16855.t8 14.282
R8347 a_36751_16855.n0 a_36751_16855.t1 14.282
R8348 a_15719_25150.n2 a_15719_25150.t5 318.922
R8349 a_15719_25150.n1 a_15719_25150.t4 273.935
R8350 a_15719_25150.n1 a_15719_25150.t6 273.935
R8351 a_15719_25150.n2 a_15719_25150.t7 269.116
R8352 a_15719_25150.n4 a_15719_25150.n0 193.227
R8353 a_15719_25150.t5 a_15719_25150.n1 179.142
R8354 a_15719_25150.n3 a_15719_25150.n2 106.999
R8355 a_15719_25150.t0 a_15719_25150.n4 28.568
R8356 a_15719_25150.n0 a_15719_25150.t1 28.565
R8357 a_15719_25150.n0 a_15719_25150.t3 28.565
R8358 a_15719_25150.n3 a_15719_25150.t2 18.149
R8359 a_15719_25150.n4 a_15719_25150.n3 3.726
R8360 a_16146_24457.n0 a_16146_24457.n1 0.001
R8361 a_16146_24457.t0 a_16146_24457.n0 14.282
R8362 a_16146_24457.n0 a_16146_24457.t6 14.282
R8363 a_16146_24457.n1 a_16146_24457.n9 267.767
R8364 a_16146_24457.n9 a_16146_24457.t7 14.282
R8365 a_16146_24457.n9 a_16146_24457.t8 14.282
R8366 a_16146_24457.n1 a_16146_24457.n7 0.669
R8367 a_16146_24457.n7 a_16146_24457.n8 1.511
R8368 a_16146_24457.n8 a_16146_24457.t2 14.282
R8369 a_16146_24457.n8 a_16146_24457.t1 14.282
R8370 a_16146_24457.n7 a_16146_24457.n6 0.227
R8371 a_16146_24457.n6 a_16146_24457.n3 0.575
R8372 a_16146_24457.n6 a_16146_24457.n5 0.2
R8373 a_16146_24457.n5 a_16146_24457.t11 16.058
R8374 a_16146_24457.n5 a_16146_24457.n4 0.999
R8375 a_16146_24457.n4 a_16146_24457.t9 14.282
R8376 a_16146_24457.n4 a_16146_24457.t10 14.282
R8377 a_16146_24457.n3 a_16146_24457.n2 0.999
R8378 a_16146_24457.n2 a_16146_24457.t4 14.282
R8379 a_16146_24457.n2 a_16146_24457.t3 14.282
R8380 a_16146_24457.n3 a_16146_24457.t5 16.058
R8381 a_n3608_5631.n1 a_n3608_5631.t4 318.119
R8382 a_n3608_5631.n1 a_n3608_5631.t5 269.919
R8383 a_n3608_5631.n0 a_n3608_5631.t6 267.256
R8384 a_n3608_5631.n0 a_n3608_5631.t7 267.256
R8385 a_n3608_5631.n4 a_n3608_5631.n3 193.227
R8386 a_n3608_5631.t4 a_n3608_5631.n0 160.666
R8387 a_n3608_5631.n2 a_n3608_5631.n1 106.999
R8388 a_n3608_5631.n3 a_n3608_5631.t1 28.568
R8389 a_n3608_5631.n4 a_n3608_5631.t2 28.565
R8390 a_n3608_5631.t3 a_n3608_5631.n4 28.565
R8391 a_n3608_5631.n2 a_n3608_5631.t0 18.149
R8392 a_n3608_5631.n3 a_n3608_5631.n2 3.726
R8393 a_30359_8848.n4 a_30359_8848.n3 563.136
R8394 a_30359_8848.t5 a_30359_8848.t15 437.233
R8395 a_30359_8848.t9 a_30359_8848.n1 313.873
R8396 a_30359_8848.n3 a_30359_8848.t12 294.986
R8397 a_30359_8848.n0 a_30359_8848.t6 272.288
R8398 a_30359_8848.n6 a_30359_8848.t5 217.824
R8399 a_30359_8848.n5 a_30359_8848.t13 214.686
R8400 a_30359_8848.t15 a_30359_8848.n5 214.686
R8401 a_30359_8848.n9 a_30359_8848.n8 192.754
R8402 a_30359_8848.n2 a_30359_8848.t9 190.152
R8403 a_30359_8848.n2 a_30359_8848.t8 190.152
R8404 a_30359_8848.n4 a_30359_8848.t10 178.973
R8405 a_30359_8848.n0 a_30359_8848.t7 160.666
R8406 a_30359_8848.n1 a_30359_8848.t11 160.666
R8407 a_30359_8848.n6 a_30359_8848.n4 133.838
R8408 a_30359_8848.n3 a_30359_8848.t4 110.859
R8409 a_30359_8848.n1 a_30359_8848.n0 96.129
R8410 a_30359_8848.t10 a_30359_8848.n2 80.333
R8411 a_30359_8848.n5 a_30359_8848.t14 80.333
R8412 a_30359_8848.n8 a_30359_8848.t2 28.568
R8413 a_30359_8848.n9 a_30359_8848.t3 28.565
R8414 a_30359_8848.t0 a_30359_8848.n9 28.565
R8415 a_30359_8848.n7 a_30359_8848.t1 18.824
R8416 a_30359_8848.n7 a_30359_8848.n6 5.567
R8417 a_30359_8848.n8 a_30359_8848.n7 1.105
R8418 a_32305_9674.n1 a_32305_9674.t7 318.922
R8419 a_32305_9674.n0 a_32305_9674.t4 274.739
R8420 a_32305_9674.n0 a_32305_9674.t6 274.739
R8421 a_32305_9674.n1 a_32305_9674.t5 269.116
R8422 a_32305_9674.t7 a_32305_9674.n0 179.946
R8423 a_32305_9674.n2 a_32305_9674.n1 107.263
R8424 a_32305_9674.t3 a_32305_9674.n4 29.444
R8425 a_32305_9674.n3 a_32305_9674.t1 28.565
R8426 a_32305_9674.n3 a_32305_9674.t2 28.565
R8427 a_32305_9674.n2 a_32305_9674.t0 18.145
R8428 a_32305_9674.n4 a_32305_9674.n2 2.878
R8429 a_32305_9674.n4 a_32305_9674.n3 0.764
R8430 a_21444_9903.n1 a_21444_9903.t7 318.922
R8431 a_21444_9903.n0 a_21444_9903.t4 274.739
R8432 a_21444_9903.n0 a_21444_9903.t5 274.739
R8433 a_21444_9903.n1 a_21444_9903.t6 269.116
R8434 a_21444_9903.t7 a_21444_9903.n0 179.946
R8435 a_21444_9903.n2 a_21444_9903.n1 105.178
R8436 a_21444_9903.n3 a_21444_9903.t1 29.444
R8437 a_21444_9903.n4 a_21444_9903.t2 28.565
R8438 a_21444_9903.t3 a_21444_9903.n4 28.565
R8439 a_21444_9903.n2 a_21444_9903.t0 18.145
R8440 a_21444_9903.n3 a_21444_9903.n2 2.878
R8441 a_21444_9903.n4 a_21444_9903.n3 0.764
R8442 a_21032_9929.t0 a_21032_9929.n7 16.058
R8443 a_21032_9929.n7 a_21032_9929.n5 0.575
R8444 a_21032_9929.n5 a_21032_9929.n9 0.2
R8445 a_21032_9929.n9 a_21032_9929.t6 16.058
R8446 a_21032_9929.n9 a_21032_9929.n8 0.999
R8447 a_21032_9929.n8 a_21032_9929.t7 14.282
R8448 a_21032_9929.n8 a_21032_9929.t5 14.282
R8449 a_21032_9929.n7 a_21032_9929.n6 0.999
R8450 a_21032_9929.n6 a_21032_9929.t11 14.282
R8451 a_21032_9929.n6 a_21032_9929.t4 14.282
R8452 a_21032_9929.n5 a_21032_9929.n3 0.227
R8453 a_21032_9929.n3 a_21032_9929.n4 1.511
R8454 a_21032_9929.n4 a_21032_9929.t1 14.282
R8455 a_21032_9929.n4 a_21032_9929.t2 14.282
R8456 a_21032_9929.n3 a_21032_9929.n0 0.669
R8457 a_21032_9929.n0 a_21032_9929.n1 0.001
R8458 a_21032_9929.n0 a_21032_9929.n2 267.767
R8459 a_21032_9929.n2 a_21032_9929.t9 14.282
R8460 a_21032_9929.n2 a_21032_9929.t8 14.282
R8461 a_21032_9929.n1 a_21032_9929.t3 14.282
R8462 a_21032_9929.n1 a_21032_9929.t10 14.282
R8463 a_21156_1325.n2 a_21156_1325.t10 214.335
R8464 a_21156_1325.t7 a_21156_1325.n2 214.335
R8465 a_21156_1325.n3 a_21156_1325.t7 143.85
R8466 a_21156_1325.n3 a_21156_1325.t8 135.66
R8467 a_21156_1325.n2 a_21156_1325.t9 80.333
R8468 a_21156_1325.n4 a_21156_1325.t5 28.565
R8469 a_21156_1325.n4 a_21156_1325.t4 28.565
R8470 a_21156_1325.n0 a_21156_1325.t3 28.565
R8471 a_21156_1325.n0 a_21156_1325.t1 28.565
R8472 a_21156_1325.n7 a_21156_1325.t6 28.565
R8473 a_21156_1325.t0 a_21156_1325.n7 28.565
R8474 a_21156_1325.n1 a_21156_1325.t2 9.714
R8475 a_21156_1325.n1 a_21156_1325.n0 1.003
R8476 a_21156_1325.n6 a_21156_1325.n5 0.836
R8477 a_21156_1325.n7 a_21156_1325.n6 0.653
R8478 a_21156_1325.n5 a_21156_1325.n4 0.65
R8479 a_21156_1325.n6 a_21156_1325.n1 0.341
R8480 a_21156_1325.n5 a_21156_1325.n3 0.032
R8481 a_21746_1762.n7 a_21746_1762.n6 861.987
R8482 a_21746_1762.n6 a_21746_1762.n5 560.726
R8483 a_21746_1762.t7 a_21746_1762.t19 415.315
R8484 a_21746_1762.t12 a_21746_1762.t8 415.315
R8485 a_21746_1762.n2 a_21746_1762.t15 394.151
R8486 a_21746_1762.n5 a_21746_1762.t16 294.653
R8487 a_21746_1762.n1 a_21746_1762.t5 269.523
R8488 a_21746_1762.t15 a_21746_1762.n1 269.523
R8489 a_21746_1762.n9 a_21746_1762.t7 217.716
R8490 a_21746_1762.n8 a_21746_1762.t9 214.335
R8491 a_21746_1762.t19 a_21746_1762.n8 214.335
R8492 a_21746_1762.n0 a_21746_1762.t4 214.335
R8493 a_21746_1762.t8 a_21746_1762.n0 214.335
R8494 a_21746_1762.n7 a_21746_1762.t12 198.921
R8495 a_21746_1762.n3 a_21746_1762.t10 198.043
R8496 a_21746_1762.n12 a_21746_1762.n11 192.754
R8497 a_21746_1762.n1 a_21746_1762.t11 160.666
R8498 a_21746_1762.n5 a_21746_1762.t14 111.663
R8499 a_21746_1762.n4 a_21746_1762.n2 97.816
R8500 a_21746_1762.n3 a_21746_1762.t17 93.989
R8501 a_21746_1762.n8 a_21746_1762.t13 80.333
R8502 a_21746_1762.n2 a_21746_1762.t6 80.333
R8503 a_21746_1762.n0 a_21746_1762.t18 80.333
R8504 a_21746_1762.n6 a_21746_1762.n4 65.07
R8505 a_21746_1762.n11 a_21746_1762.t1 28.568
R8506 a_21746_1762.n12 a_21746_1762.t2 28.565
R8507 a_21746_1762.t3 a_21746_1762.n12 28.565
R8508 a_21746_1762.n10 a_21746_1762.t0 18.827
R8509 a_21746_1762.n9 a_21746_1762.n7 16.411
R8510 a_21746_1762.n4 a_21746_1762.n3 6.615
R8511 a_21746_1762.n10 a_21746_1762.n9 4.58
R8512 a_21746_1762.n11 a_21746_1762.n10 1.105
R8513 a_18952_19520.n0 a_18952_19520.t6 14.282
R8514 a_18952_19520.t0 a_18952_19520.n0 14.282
R8515 a_18952_19520.n0 a_18952_19520.n12 90.416
R8516 a_18952_19520.n12 a_18952_19520.n9 74.302
R8517 a_18952_19520.n12 a_18952_19520.n11 50.575
R8518 a_18952_19520.n11 a_18952_19520.n10 157.665
R8519 a_18952_19520.n10 a_18952_19520.t7 8.7
R8520 a_18952_19520.n10 a_18952_19520.t2 8.7
R8521 a_18952_19520.n9 a_18952_19520.n8 90.436
R8522 a_18952_19520.n8 a_18952_19520.t5 14.282
R8523 a_18952_19520.n8 a_18952_19520.t4 14.282
R8524 a_18952_19520.n11 a_18952_19520.n7 122.746
R8525 a_18952_19520.n7 a_18952_19520.t1 14.282
R8526 a_18952_19520.n7 a_18952_19520.t3 14.282
R8527 a_18952_19520.n9 a_18952_19520.n1 342.688
R8528 a_18952_19520.n1 a_18952_19520.n6 126.566
R8529 a_18952_19520.n6 a_18952_19520.t10 294.653
R8530 a_18952_19520.n6 a_18952_19520.t14 111.663
R8531 a_18952_19520.n1 a_18952_19520.n5 552.333
R8532 a_18952_19520.n5 a_18952_19520.n4 6.615
R8533 a_18952_19520.n4 a_18952_19520.t12 93.989
R8534 a_18952_19520.n4 a_18952_19520.t13 198.043
R8535 a_18952_19520.n5 a_18952_19520.n3 97.816
R8536 a_18952_19520.n3 a_18952_19520.t11 80.333
R8537 a_18952_19520.n3 a_18952_19520.t9 394.151
R8538 a_18952_19520.t9 a_18952_19520.n2 269.523
R8539 a_18952_19520.n2 a_18952_19520.t15 160.666
R8540 a_18952_19520.n2 a_18952_19520.t8 269.523
R8541 a_10702_9703.n4 a_10702_9703.t8 214.335
R8542 a_10702_9703.t7 a_10702_9703.n4 214.335
R8543 a_10702_9703.n5 a_10702_9703.t7 143.851
R8544 a_10702_9703.n5 a_10702_9703.t9 135.658
R8545 a_10702_9703.n4 a_10702_9703.t10 80.333
R8546 a_10702_9703.n0 a_10702_9703.t4 28.565
R8547 a_10702_9703.n0 a_10702_9703.t3 28.565
R8548 a_10702_9703.n2 a_10702_9703.t5 28.565
R8549 a_10702_9703.n2 a_10702_9703.t2 28.565
R8550 a_10702_9703.t0 a_10702_9703.n7 28.565
R8551 a_10702_9703.n7 a_10702_9703.t6 28.565
R8552 a_10702_9703.n1 a_10702_9703.t1 9.714
R8553 a_10702_9703.n1 a_10702_9703.n0 1.003
R8554 a_10702_9703.n6 a_10702_9703.n3 0.833
R8555 a_10702_9703.n3 a_10702_9703.n2 0.653
R8556 a_10702_9703.n7 a_10702_9703.n6 0.653
R8557 a_10702_9703.n3 a_10702_9703.n1 0.341
R8558 a_10702_9703.n6 a_10702_9703.n5 0.032
R8559 a_14660_24431.n1 a_14660_24431.t6 318.922
R8560 a_14660_24431.n0 a_14660_24431.t5 274.739
R8561 a_14660_24431.n0 a_14660_24431.t7 274.739
R8562 a_14660_24431.n1 a_14660_24431.t4 269.116
R8563 a_14660_24431.t6 a_14660_24431.n0 179.946
R8564 a_14660_24431.n2 a_14660_24431.n1 107.263
R8565 a_14660_24431.n3 a_14660_24431.t2 29.444
R8566 a_14660_24431.t3 a_14660_24431.n4 28.565
R8567 a_14660_24431.n4 a_14660_24431.t1 28.565
R8568 a_14660_24431.n2 a_14660_24431.t0 18.145
R8569 a_14660_24431.n3 a_14660_24431.n2 2.878
R8570 a_14660_24431.n4 a_14660_24431.n3 0.764
R8571 a_27458_24456.n0 a_27458_24456.n12 122.999
R8572 a_27458_24456.n0 a_27458_24456.t2 14.282
R8573 a_27458_24456.t1 a_27458_24456.n0 14.282
R8574 a_27458_24456.n12 a_27458_24456.n10 50.575
R8575 a_27458_24456.n10 a_27458_24456.n8 74.302
R8576 a_27458_24456.n12 a_27458_24456.n11 157.665
R8577 a_27458_24456.n11 a_27458_24456.t0 8.7
R8578 a_27458_24456.n11 a_27458_24456.t4 8.7
R8579 a_27458_24456.n10 a_27458_24456.n9 90.416
R8580 a_27458_24456.n9 a_27458_24456.t5 14.282
R8581 a_27458_24456.n9 a_27458_24456.t6 14.282
R8582 a_27458_24456.n8 a_27458_24456.n7 90.436
R8583 a_27458_24456.n7 a_27458_24456.t7 14.282
R8584 a_27458_24456.n7 a_27458_24456.t3 14.282
R8585 a_27458_24456.n8 a_27458_24456.n1 342.688
R8586 a_27458_24456.n1 a_27458_24456.n6 126.566
R8587 a_27458_24456.n6 a_27458_24456.t15 294.653
R8588 a_27458_24456.n6 a_27458_24456.t14 111.663
R8589 a_27458_24456.n1 a_27458_24456.n5 552.333
R8590 a_27458_24456.n5 a_27458_24456.n4 6.615
R8591 a_27458_24456.n4 a_27458_24456.t12 93.989
R8592 a_27458_24456.n5 a_27458_24456.n3 97.816
R8593 a_27458_24456.n3 a_27458_24456.t13 80.333
R8594 a_27458_24456.n3 a_27458_24456.t8 394.151
R8595 a_27458_24456.t8 a_27458_24456.n2 269.523
R8596 a_27458_24456.n2 a_27458_24456.t9 160.666
R8597 a_27458_24456.n2 a_27458_24456.t10 269.523
R8598 a_27458_24456.n4 a_27458_24456.t11 198.043
R8599 a_29238_24456.t0 a_29238_24456.n0 14.282
R8600 a_29238_24456.n0 a_29238_24456.t1 14.282
R8601 a_29238_24456.n0 a_29238_24456.n9 0.999
R8602 a_29238_24456.n6 a_29238_24456.n8 0.575
R8603 a_29238_24456.n9 a_29238_24456.n6 0.2
R8604 a_29238_24456.n9 a_29238_24456.t2 16.058
R8605 a_29238_24456.n8 a_29238_24456.n7 0.999
R8606 a_29238_24456.n7 a_29238_24456.t7 14.282
R8607 a_29238_24456.n7 a_29238_24456.t8 14.282
R8608 a_29238_24456.n8 a_29238_24456.t6 16.058
R8609 a_29238_24456.n6 a_29238_24456.n4 0.227
R8610 a_29238_24456.n4 a_29238_24456.n5 1.511
R8611 a_29238_24456.n5 a_29238_24456.t11 14.282
R8612 a_29238_24456.n5 a_29238_24456.t10 14.282
R8613 a_29238_24456.n4 a_29238_24456.n1 0.669
R8614 a_29238_24456.n1 a_29238_24456.n2 0.001
R8615 a_29238_24456.n1 a_29238_24456.n3 267.767
R8616 a_29238_24456.n3 a_29238_24456.t4 14.282
R8617 a_29238_24456.n3 a_29238_24456.t5 14.282
R8618 a_29238_24456.n2 a_29238_24456.t9 14.282
R8619 a_29238_24456.n2 a_29238_24456.t3 14.282
R8620 a_17351_3834.n0 a_17351_3834.t8 214.335
R8621 a_17351_3834.t7 a_17351_3834.n0 214.335
R8622 a_17351_3834.n1 a_17351_3834.t7 143.851
R8623 a_17351_3834.n1 a_17351_3834.t9 135.658
R8624 a_17351_3834.n0 a_17351_3834.t10 80.333
R8625 a_17351_3834.n2 a_17351_3834.t3 28.565
R8626 a_17351_3834.n2 a_17351_3834.t2 28.565
R8627 a_17351_3834.n4 a_17351_3834.t4 28.565
R8628 a_17351_3834.n4 a_17351_3834.t5 28.565
R8629 a_17351_3834.t1 a_17351_3834.n7 28.565
R8630 a_17351_3834.n7 a_17351_3834.t6 28.565
R8631 a_17351_3834.n6 a_17351_3834.t0 9.714
R8632 a_17351_3834.n7 a_17351_3834.n6 1.003
R8633 a_17351_3834.n5 a_17351_3834.n3 0.833
R8634 a_17351_3834.n3 a_17351_3834.n2 0.653
R8635 a_17351_3834.n5 a_17351_3834.n4 0.653
R8636 a_17351_3834.n6 a_17351_3834.n5 0.341
R8637 a_17351_3834.n3 a_17351_3834.n1 0.032
R8638 a_17941_3397.t4 a_17941_3397.t5 574.43
R8639 a_17941_3397.n0 a_17941_3397.t6 285.109
R8640 a_17941_3397.n2 a_17941_3397.n1 197.217
R8641 a_17941_3397.n4 a_17941_3397.n3 192.754
R8642 a_17941_3397.n0 a_17941_3397.t7 160.666
R8643 a_17941_3397.n1 a_17941_3397.t4 160.666
R8644 a_17941_3397.n1 a_17941_3397.n0 114.829
R8645 a_17941_3397.n3 a_17941_3397.t2 28.568
R8646 a_17941_3397.n4 a_17941_3397.t1 28.565
R8647 a_17941_3397.t3 a_17941_3397.n4 28.565
R8648 a_17941_3397.n2 a_17941_3397.t0 18.838
R8649 a_17941_3397.n3 a_17941_3397.n2 1.129
R8650 a_7939_4129.n0 a_7939_4129.t3 14.282
R8651 a_7939_4129.t0 a_7939_4129.n0 14.282
R8652 a_7939_4129.n0 a_7939_4129.n15 90.416
R8653 a_7939_4129.n15 a_7939_4129.n14 50.575
R8654 a_7939_4129.n15 a_7939_4129.n11 74.302
R8655 a_7939_4129.n14 a_7939_4129.n13 157.665
R8656 a_7939_4129.n13 a_7939_4129.t5 8.7
R8657 a_7939_4129.n13 a_7939_4129.t7 8.7
R8658 a_7939_4129.n14 a_7939_4129.n12 122.999
R8659 a_7939_4129.n12 a_7939_4129.t4 14.282
R8660 a_7939_4129.n12 a_7939_4129.t2 14.282
R8661 a_7939_4129.n11 a_7939_4129.n10 90.436
R8662 a_7939_4129.n10 a_7939_4129.t1 14.282
R8663 a_7939_4129.n10 a_7939_4129.t6 14.282
R8664 a_7939_4129.n11 a_7939_4129.n9 220.358
R8665 a_7939_4129.n9 a_7939_4129.n2 2.596
R8666 a_7939_4129.n2 a_7939_4129.t11 218.628
R8667 a_7939_4129.t11 a_7939_4129.t23 437.233
R8668 a_7939_4129.t23 a_7939_4129.n8 214.686
R8669 a_7939_4129.n8 a_7939_4129.t12 80.333
R8670 a_7939_4129.n8 a_7939_4129.t19 214.686
R8671 a_7939_4129.n2 a_7939_4129.n3 14.9
R8672 a_7939_4129.n3 a_7939_4129.n7 535.449
R8673 a_7939_4129.n7 a_7939_4129.t8 294.986
R8674 a_7939_4129.n7 a_7939_4129.t13 110.859
R8675 a_7939_4129.n3 a_7939_4129.t9 245.184
R8676 a_7939_4129.t9 a_7939_4129.n6 80.333
R8677 a_7939_4129.n6 a_7939_4129.t20 190.152
R8678 a_7939_4129.n6 a_7939_4129.t14 190.152
R8679 a_7939_4129.t14 a_7939_4129.n5 313.873
R8680 a_7939_4129.n5 a_7939_4129.t22 160.666
R8681 a_7939_4129.n5 a_7939_4129.n4 96.129
R8682 a_7939_4129.n4 a_7939_4129.t17 160.666
R8683 a_7939_4129.n4 a_7939_4129.t15 272.288
R8684 a_7939_4129.n9 a_7939_4129.t16 217.023
R8685 a_7939_4129.t16 a_7939_4129.t10 437.233
R8686 a_7939_4129.t10 a_7939_4129.n1 214.686
R8687 a_7939_4129.n1 a_7939_4129.t18 80.333
R8688 a_7939_4129.n1 a_7939_4129.t21 214.686
R8689 a_12828_3395.t0 a_12828_3395.t1 17.4
R8690 a_26157_25329.t7 a_26157_25329.t6 574.43
R8691 a_26157_25329.n0 a_26157_25329.t5 285.109
R8692 a_26157_25329.n2 a_26157_25329.n1 211.136
R8693 a_26157_25329.n4 a_26157_25329.n3 192.754
R8694 a_26157_25329.n0 a_26157_25329.t4 160.666
R8695 a_26157_25329.n1 a_26157_25329.t7 160.666
R8696 a_26157_25329.n1 a_26157_25329.n0 114.829
R8697 a_26157_25329.n3 a_26157_25329.t3 28.568
R8698 a_26157_25329.n4 a_26157_25329.t2 28.565
R8699 a_26157_25329.t1 a_26157_25329.n4 28.565
R8700 a_26157_25329.n2 a_26157_25329.t0 19.084
R8701 a_26157_25329.n3 a_26157_25329.n2 1.051
R8702 a_29020_27292.n0 a_29020_27292.t5 14.282
R8703 a_29020_27292.n0 a_29020_27292.t3 14.282
R8704 a_29020_27292.n1 a_29020_27292.t2 14.282
R8705 a_29020_27292.n1 a_29020_27292.t1 14.282
R8706 a_29020_27292.t0 a_29020_27292.n3 14.282
R8707 a_29020_27292.n3 a_29020_27292.t4 14.282
R8708 a_29020_27292.n2 a_29020_27292.n0 2.546
R8709 a_29020_27292.n2 a_29020_27292.n1 2.367
R8710 a_29020_27292.n3 a_29020_27292.n2 0.001
R8711 a_28902_27292.t5 a_28902_27292.n2 404.877
R8712 a_28902_27292.n1 a_28902_27292.t7 210.902
R8713 a_28902_27292.n3 a_28902_27292.t5 136.943
R8714 a_28902_27292.n2 a_28902_27292.n1 107.801
R8715 a_28902_27292.n1 a_28902_27292.t6 80.333
R8716 a_28902_27292.n2 a_28902_27292.t8 80.333
R8717 a_28902_27292.n0 a_28902_27292.t0 17.4
R8718 a_28902_27292.n0 a_28902_27292.t4 17.4
R8719 a_28902_27292.n4 a_28902_27292.t1 15.032
R8720 a_28902_27292.n5 a_28902_27292.t2 14.282
R8721 a_28902_27292.t3 a_28902_27292.n5 14.282
R8722 a_28902_27292.n5 a_28902_27292.n4 1.65
R8723 a_28902_27292.n3 a_28902_27292.n0 0.672
R8724 a_28902_27292.n4 a_28902_27292.n3 0.665
R8725 a_7749_6382.n8 a_7749_6382.n7 861.987
R8726 a_7749_6382.n7 a_7749_6382.n6 560.726
R8727 a_7749_6382.t11 a_7749_6382.t4 415.315
R8728 a_7749_6382.t14 a_7749_6382.t19 415.315
R8729 a_7749_6382.n3 a_7749_6382.t5 394.151
R8730 a_7749_6382.n6 a_7749_6382.t6 294.653
R8731 a_7749_6382.n2 a_7749_6382.t15 269.523
R8732 a_7749_6382.t5 a_7749_6382.n2 269.523
R8733 a_7749_6382.n10 a_7749_6382.t11 217.716
R8734 a_7749_6382.n9 a_7749_6382.t10 214.335
R8735 a_7749_6382.t4 a_7749_6382.n9 214.335
R8736 a_7749_6382.n1 a_7749_6382.t9 214.335
R8737 a_7749_6382.t19 a_7749_6382.n1 214.335
R8738 a_7749_6382.n8 a_7749_6382.t14 198.921
R8739 a_7749_6382.n4 a_7749_6382.t16 198.043
R8740 a_7749_6382.n2 a_7749_6382.t13 160.666
R8741 a_7749_6382.n6 a_7749_6382.t12 111.663
R8742 a_7749_6382.n5 a_7749_6382.n3 97.816
R8743 a_7749_6382.n4 a_7749_6382.t17 93.989
R8744 a_7749_6382.n9 a_7749_6382.t8 80.333
R8745 a_7749_6382.n3 a_7749_6382.t18 80.333
R8746 a_7749_6382.n1 a_7749_6382.t7 80.333
R8747 a_7749_6382.n7 a_7749_6382.n5 65.07
R8748 a_7749_6382.n0 a_7749_6382.t2 28.57
R8749 a_7749_6382.t0 a_7749_6382.n12 28.565
R8750 a_7749_6382.n12 a_7749_6382.t3 28.565
R8751 a_7749_6382.n0 a_7749_6382.t1 17.638
R8752 a_7749_6382.n10 a_7749_6382.n8 16.411
R8753 a_7749_6382.n11 a_7749_6382.n10 8.712
R8754 a_7749_6382.n5 a_7749_6382.n4 6.615
R8755 a_7749_6382.n12 a_7749_6382.n11 0.69
R8756 a_7749_6382.n11 a_7749_6382.n0 0.6
R8757 a_n2379_15428.t0 a_n2379_15428.t1 17.4
R8758 a_23978_5439.n2 a_23978_5439.t8 214.335
R8759 a_23978_5439.t10 a_23978_5439.n2 214.335
R8760 a_23978_5439.n3 a_23978_5439.t10 143.851
R8761 a_23978_5439.n3 a_23978_5439.t7 135.658
R8762 a_23978_5439.n2 a_23978_5439.t9 80.333
R8763 a_23978_5439.n4 a_23978_5439.t6 28.565
R8764 a_23978_5439.n4 a_23978_5439.t4 28.565
R8765 a_23978_5439.n0 a_23978_5439.t1 28.565
R8766 a_23978_5439.n0 a_23978_5439.t2 28.565
R8767 a_23978_5439.n7 a_23978_5439.t5 28.565
R8768 a_23978_5439.t3 a_23978_5439.n7 28.565
R8769 a_23978_5439.n1 a_23978_5439.t0 9.714
R8770 a_23978_5439.n1 a_23978_5439.n0 1.003
R8771 a_23978_5439.n6 a_23978_5439.n5 0.833
R8772 a_23978_5439.n5 a_23978_5439.n4 0.653
R8773 a_23978_5439.n7 a_23978_5439.n6 0.653
R8774 a_23978_5439.n6 a_23978_5439.n1 0.341
R8775 a_23978_5439.n5 a_23978_5439.n3 0.032
R8776 a_24568_5002.t4 a_24568_5002.t5 574.43
R8777 a_24568_5002.n1 a_24568_5002.t7 285.109
R8778 a_24568_5002.n3 a_24568_5002.n2 211.136
R8779 a_24568_5002.n4 a_24568_5002.n0 192.754
R8780 a_24568_5002.n1 a_24568_5002.t6 160.666
R8781 a_24568_5002.n2 a_24568_5002.t4 160.666
R8782 a_24568_5002.n2 a_24568_5002.n1 114.829
R8783 a_24568_5002.t3 a_24568_5002.n4 28.568
R8784 a_24568_5002.n0 a_24568_5002.t2 28.565
R8785 a_24568_5002.n0 a_24568_5002.t1 28.565
R8786 a_24568_5002.n3 a_24568_5002.t0 19.084
R8787 a_24568_5002.n4 a_24568_5002.n3 1.051
R8788 a_n3608_4192.n1 a_n3608_4192.t4 318.119
R8789 a_n3608_4192.n1 a_n3608_4192.t6 269.919
R8790 a_n3608_4192.n0 a_n3608_4192.t7 267.853
R8791 a_n3608_4192.n0 a_n3608_4192.t5 267.853
R8792 a_n3608_4192.t4 a_n3608_4192.n0 160.666
R8793 a_n3608_4192.n2 a_n3608_4192.n1 107.263
R8794 a_n3608_4192.t3 a_n3608_4192.n4 29.444
R8795 a_n3608_4192.n3 a_n3608_4192.t1 28.565
R8796 a_n3608_4192.n3 a_n3608_4192.t2 28.565
R8797 a_n3608_4192.n2 a_n3608_4192.t0 18.145
R8798 a_n3608_4192.n4 a_n3608_4192.n2 2.878
R8799 a_n3608_4192.n4 a_n3608_4192.n3 0.764
R8800 a_n3115_4850.t0 a_n3115_4850.n0 14.282
R8801 a_n3115_4850.n0 a_n3115_4850.t5 14.282
R8802 a_n3115_4850.n0 a_n3115_4850.n16 90.416
R8803 a_n3115_4850.n16 a_n3115_4850.n2 74.302
R8804 a_n3115_4850.n16 a_n3115_4850.n4 50.575
R8805 a_n3115_4850.n4 a_n3115_4850.n5 110.084
R8806 a_n3115_4850.n2 a_n3115_4850.n6 670.431
R8807 a_n3115_4850.n6 a_n3115_4850.n8 16.411
R8808 a_n3115_4850.n8 a_n3115_4850.t22 198.921
R8809 a_n3115_4850.t22 a_n3115_4850.t18 415.315
R8810 a_n3115_4850.t18 a_n3115_4850.n15 214.335
R8811 a_n3115_4850.n15 a_n3115_4850.t17 80.333
R8812 a_n3115_4850.n15 a_n3115_4850.t16 214.335
R8813 a_n3115_4850.n8 a_n3115_4850.n14 861.987
R8814 a_n3115_4850.n14 a_n3115_4850.n9 560.726
R8815 a_n3115_4850.n14 a_n3115_4850.n13 65.07
R8816 a_n3115_4850.n13 a_n3115_4850.n12 6.615
R8817 a_n3115_4850.n12 a_n3115_4850.t20 93.989
R8818 a_n3115_4850.n12 a_n3115_4850.t21 198.043
R8819 a_n3115_4850.n13 a_n3115_4850.n11 97.816
R8820 a_n3115_4850.n11 a_n3115_4850.t19 80.333
R8821 a_n3115_4850.n11 a_n3115_4850.t9 394.151
R8822 a_n3115_4850.t9 a_n3115_4850.n10 269.523
R8823 a_n3115_4850.n10 a_n3115_4850.t11 160.666
R8824 a_n3115_4850.n10 a_n3115_4850.t8 269.523
R8825 a_n3115_4850.n9 a_n3115_4850.t15 294.653
R8826 a_n3115_4850.n9 a_n3115_4850.t23 111.663
R8827 a_n3115_4850.n6 a_n3115_4850.t10 217.716
R8828 a_n3115_4850.t10 a_n3115_4850.t14 415.315
R8829 a_n3115_4850.t14 a_n3115_4850.n7 214.335
R8830 a_n3115_4850.n7 a_n3115_4850.t13 80.333
R8831 a_n3115_4850.n7 a_n3115_4850.t12 214.335
R8832 a_n3115_4850.n5 a_n3115_4850.t7 14.282
R8833 a_n3115_4850.n5 a_n3115_4850.t6 14.282
R8834 a_n3115_4850.n4 a_n3115_4850.n3 157.665
R8835 a_n3115_4850.n3 a_n3115_4850.t3 8.7
R8836 a_n3115_4850.n3 a_n3115_4850.t4 8.7
R8837 a_n3115_4850.n2 a_n3115_4850.n1 90.436
R8838 a_n3115_4850.n1 a_n3115_4850.t1 14.282
R8839 a_n3115_4850.n1 a_n3115_4850.t2 14.282
R8840 a_n3808_4793.n9 a_n3808_4793.n8 267.767
R8841 a_n3808_4793.n1 a_n3808_4793.t10 16.058
R8842 a_n3808_4793.n3 a_n3808_4793.t4 16.058
R8843 a_n3808_4793.n0 a_n3808_4793.t11 14.282
R8844 a_n3808_4793.n0 a_n3808_4793.t9 14.282
R8845 a_n3808_4793.n2 a_n3808_4793.t3 14.282
R8846 a_n3808_4793.n2 a_n3808_4793.t5 14.282
R8847 a_n3808_4793.n5 a_n3808_4793.t8 14.282
R8848 a_n3808_4793.n5 a_n3808_4793.t6 14.282
R8849 a_n3808_4793.n7 a_n3808_4793.t7 14.282
R8850 a_n3808_4793.n7 a_n3808_4793.t1 14.282
R8851 a_n3808_4793.t2 a_n3808_4793.n9 14.282
R8852 a_n3808_4793.n9 a_n3808_4793.t0 14.282
R8853 a_n3808_4793.n6 a_n3808_4793.n5 1.511
R8854 a_n3808_4793.n1 a_n3808_4793.n0 0.999
R8855 a_n3808_4793.n3 a_n3808_4793.n2 0.999
R8856 a_n3808_4793.n8 a_n3808_4793.n6 0.669
R8857 a_n3808_4793.n4 a_n3808_4793.n1 0.575
R8858 a_n3808_4793.n6 a_n3808_4793.n4 0.227
R8859 a_n3808_4793.n4 a_n3808_4793.n3 0.2
R8860 a_n3808_4793.n8 a_n3808_4793.n7 0.001
R8861 a_4748_10782.t4 a_4748_10782.t5 574.43
R8862 a_4748_10782.n1 a_4748_10782.t7 285.109
R8863 a_4748_10782.n3 a_4748_10782.n2 211.136
R8864 a_4748_10782.n4 a_4748_10782.n0 192.754
R8865 a_4748_10782.n1 a_4748_10782.t6 160.666
R8866 a_4748_10782.n2 a_4748_10782.t4 160.666
R8867 a_4748_10782.n2 a_4748_10782.n1 114.829
R8868 a_4748_10782.t1 a_4748_10782.n4 28.568
R8869 a_4748_10782.n0 a_4748_10782.t3 28.565
R8870 a_4748_10782.n0 a_4748_10782.t2 28.565
R8871 a_4748_10782.n3 a_4748_10782.t0 19.084
R8872 a_4748_10782.n4 a_4748_10782.n3 1.051
R8873 a_7493_12745.t6 a_7493_12745.n2 404.877
R8874 a_7493_12745.n1 a_7493_12745.t8 210.902
R8875 a_7493_12745.n3 a_7493_12745.t6 136.943
R8876 a_7493_12745.n2 a_7493_12745.n1 107.801
R8877 a_7493_12745.n1 a_7493_12745.t7 80.333
R8878 a_7493_12745.n2 a_7493_12745.t5 80.333
R8879 a_7493_12745.n0 a_7493_12745.t0 17.4
R8880 a_7493_12745.n0 a_7493_12745.t1 17.4
R8881 a_7493_12745.n4 a_7493_12745.t4 15.032
R8882 a_7493_12745.t2 a_7493_12745.n5 14.282
R8883 a_7493_12745.n5 a_7493_12745.t3 14.282
R8884 a_7493_12745.n5 a_7493_12745.n4 1.65
R8885 a_7493_12745.n3 a_7493_12745.n0 0.672
R8886 a_7493_12745.n4 a_7493_12745.n3 0.665
R8887 a_7611_12745.n1 a_7611_12745.t1 14.282
R8888 a_7611_12745.n1 a_7611_12745.t2 14.282
R8889 a_7611_12745.n0 a_7611_12745.t3 14.282
R8890 a_7611_12745.n0 a_7611_12745.t4 14.282
R8891 a_7611_12745.t0 a_7611_12745.n3 14.282
R8892 a_7611_12745.n3 a_7611_12745.t5 14.282
R8893 a_7611_12745.n2 a_7611_12745.n0 2.546
R8894 a_7611_12745.n3 a_7611_12745.n2 2.367
R8895 a_7611_12745.n2 a_7611_12745.n1 0.001
R8896 a_6863_19545.n1 a_6863_19545.t5 318.922
R8897 a_6863_19545.n0 a_6863_19545.t4 274.739
R8898 a_6863_19545.n0 a_6863_19545.t6 274.739
R8899 a_6863_19545.n1 a_6863_19545.t7 269.116
R8900 a_6863_19545.t5 a_6863_19545.n0 179.946
R8901 a_6863_19545.n2 a_6863_19545.n1 107.263
R8902 a_6863_19545.n3 a_6863_19545.t2 29.444
R8903 a_6863_19545.n4 a_6863_19545.t3 28.565
R8904 a_6863_19545.t0 a_6863_19545.n4 28.565
R8905 a_6863_19545.n2 a_6863_19545.t1 18.145
R8906 a_6863_19545.n3 a_6863_19545.n2 2.878
R8907 a_6863_19545.n4 a_6863_19545.n3 0.764
R8908 a_7403_18852.n5 a_7403_18852.n7 0.2
R8909 a_7403_18852.n9 a_7403_18852.n5 0.575
R8910 a_7403_18852.t0 a_7403_18852.n9 16.058
R8911 a_7403_18852.n9 a_7403_18852.n8 0.999
R8912 a_7403_18852.n8 a_7403_18852.t4 14.282
R8913 a_7403_18852.n8 a_7403_18852.t5 14.282
R8914 a_7403_18852.n7 a_7403_18852.n6 0.999
R8915 a_7403_18852.n6 a_7403_18852.t10 14.282
R8916 a_7403_18852.n6 a_7403_18852.t9 14.282
R8917 a_7403_18852.n7 a_7403_18852.t11 16.058
R8918 a_7403_18852.n5 a_7403_18852.n3 0.227
R8919 a_7403_18852.n3 a_7403_18852.n4 1.511
R8920 a_7403_18852.n4 a_7403_18852.t2 14.282
R8921 a_7403_18852.n4 a_7403_18852.t1 14.282
R8922 a_7403_18852.n3 a_7403_18852.n0 0.669
R8923 a_7403_18852.n0 a_7403_18852.n1 0.001
R8924 a_7403_18852.n0 a_7403_18852.n2 267.767
R8925 a_7403_18852.n2 a_7403_18852.t8 14.282
R8926 a_7403_18852.n2 a_7403_18852.t7 14.282
R8927 a_7403_18852.n1 a_7403_18852.t6 14.282
R8928 a_7403_18852.n1 a_7403_18852.t3 14.282
R8929 a_28811_25149.n2 a_28811_25149.t5 318.922
R8930 a_28811_25149.n1 a_28811_25149.t4 273.935
R8931 a_28811_25149.n1 a_28811_25149.t6 273.935
R8932 a_28811_25149.n2 a_28811_25149.t7 269.116
R8933 a_28811_25149.n4 a_28811_25149.n0 193.227
R8934 a_28811_25149.t5 a_28811_25149.n1 179.142
R8935 a_28811_25149.n3 a_28811_25149.n2 106.999
R8936 a_28811_25149.t3 a_28811_25149.n4 28.568
R8937 a_28811_25149.n0 a_28811_25149.t1 28.565
R8938 a_28811_25149.n0 a_28811_25149.t2 28.565
R8939 a_28811_25149.n3 a_28811_25149.t0 18.149
R8940 a_28811_25149.n4 a_28811_25149.n3 3.726
R8941 a_29356_24456.n0 a_29356_24456.t4 14.282
R8942 a_29356_24456.t0 a_29356_24456.n0 14.282
R8943 a_29356_24456.n0 a_29356_24456.n8 90.416
R8944 a_29356_24456.n8 a_29356_24456.n7 50.575
R8945 a_29356_24456.n8 a_29356_24456.n4 74.302
R8946 a_29356_24456.n7 a_29356_24456.n6 157.665
R8947 a_29356_24456.n6 a_29356_24456.t3 8.7
R8948 a_29356_24456.n6 a_29356_24456.t7 8.7
R8949 a_29356_24456.n7 a_29356_24456.n5 122.999
R8950 a_29356_24456.n5 a_29356_24456.t6 14.282
R8951 a_29356_24456.n5 a_29356_24456.t5 14.282
R8952 a_29356_24456.n4 a_29356_24456.n3 90.436
R8953 a_29356_24456.n3 a_29356_24456.t1 14.282
R8954 a_29356_24456.n3 a_29356_24456.t2 14.282
R8955 a_29356_24456.n4 a_29356_24456.n1 449.112
R8956 a_29356_24456.t11 a_29356_24456.n2 160.666
R8957 a_29356_24456.n1 a_29356_24456.t11 867.393
R8958 a_29356_24456.n2 a_29356_24456.t9 287.241
R8959 a_29356_24456.n2 a_29356_24456.t8 287.241
R8960 a_29356_24456.n1 a_29356_24456.t10 545.094
R8961 a_9751_24460.t0 a_9751_24460.n0 14.282
R8962 a_9751_24460.n0 a_9751_24460.t2 14.282
R8963 a_9751_24460.n0 a_9751_24460.n8 90.436
R8964 a_9751_24460.n4 a_9751_24460.n7 50.575
R8965 a_9751_24460.n8 a_9751_24460.n4 74.302
R8966 a_9751_24460.n7 a_9751_24460.n6 157.665
R8967 a_9751_24460.n6 a_9751_24460.t5 8.7
R8968 a_9751_24460.n6 a_9751_24460.t7 8.7
R8969 a_9751_24460.n7 a_9751_24460.n5 122.999
R8970 a_9751_24460.n5 a_9751_24460.t6 14.282
R8971 a_9751_24460.n5 a_9751_24460.t3 14.282
R8972 a_9751_24460.n4 a_9751_24460.n3 90.416
R8973 a_9751_24460.n3 a_9751_24460.t4 14.282
R8974 a_9751_24460.n3 a_9751_24460.t1 14.282
R8975 a_9751_24460.n8 a_9751_24460.n1 3155.65
R8976 a_9751_24460.t10 a_9751_24460.n2 160.666
R8977 a_9751_24460.n1 a_9751_24460.t10 867.393
R8978 a_9751_24460.n2 a_9751_24460.t9 287.241
R8979 a_9751_24460.n2 a_9751_24460.t11 287.241
R8980 a_9751_24460.n1 a_9751_24460.t8 545.094
R8981 a_38088_23722.t0 a_38088_23722.t1 17.4
R8982 B[3].n11 B[3].n7 592.056
R8983 B[3].t1 B[3].t19 437.233
R8984 B[3].t21 B[3].t5 437.233
R8985 B[3].t16 B[3].t12 437.233
R8986 B[3].t8 B[3].t10 415.315
R8987 B[3].t3 B[3].n9 313.069
R8988 B[3].n7 B[3].t6 294.986
R8989 B[3].n8 B[3].t23 271.484
R8990 B[3].n2 B[3].t8 225.375
R8991 B[3].n5 B[3].t16 223.992
R8992 B[3].n5 B[3].t21 217.885
R8993 B[3].n2 B[3].t1 216.848
R8994 B[3].n1 B[3].t17 214.686
R8995 B[3].t19 B[3].n1 214.686
R8996 B[3].n3 B[3].t7 214.686
R8997 B[3].t5 B[3].n3 214.686
R8998 B[3].n4 B[3].t2 214.686
R8999 B[3].t12 B[3].n4 214.686
R9000 B[3].n0 B[3].t13 214.335
R9001 B[3].t10 B[3].n0 214.335
R9002 B[3].n11 B[3].t22 204.672
R9003 B[3].n10 B[3].t3 190.955
R9004 B[3].n10 B[3].t14 190.955
R9005 B[3].n9 B[3].t9 160.666
R9006 B[3].n8 B[3].t15 160.666
R9007 B[3].n7 B[3].t20 110.859
R9008 B[3].n9 B[3].n8 96.129
R9009 B[3].n1 B[3].t18 80.333
R9010 B[3].n0 B[3].t4 80.333
R9011 B[3].n3 B[3].t0 80.333
R9012 B[3].n4 B[3].t11 80.333
R9013 B[3].t22 B[3].n10 80.333
R9014 B[3].n6 B[3].n2 62.925
R9015 B[3].n12 B[3].n11 45.981
R9016 B[3] B[3].n12 19.531
R9017 B[3].n12 B[3].n6 13.481
R9018 B[3].n6 B[3].n5 0.469
R9019 a_1243_4513.n2 a_1243_4513.t8 214.335
R9020 a_1243_4513.t7 a_1243_4513.n2 214.335
R9021 a_1243_4513.n3 a_1243_4513.t7 143.851
R9022 a_1243_4513.n3 a_1243_4513.t9 135.658
R9023 a_1243_4513.n2 a_1243_4513.t10 80.333
R9024 a_1243_4513.n4 a_1243_4513.t1 28.565
R9025 a_1243_4513.n4 a_1243_4513.t0 28.565
R9026 a_1243_4513.n0 a_1243_4513.t6 28.565
R9027 a_1243_4513.n0 a_1243_4513.t4 28.565
R9028 a_1243_4513.t2 a_1243_4513.n7 28.565
R9029 a_1243_4513.n7 a_1243_4513.t5 28.565
R9030 a_1243_4513.n1 a_1243_4513.t3 9.714
R9031 a_1243_4513.n1 a_1243_4513.n0 1.003
R9032 a_1243_4513.n6 a_1243_4513.n5 0.833
R9033 a_1243_4513.n5 a_1243_4513.n4 0.653
R9034 a_1243_4513.n7 a_1243_4513.n6 0.653
R9035 a_1243_4513.n6 a_1243_4513.n1 0.341
R9036 a_1243_4513.n5 a_1243_4513.n3 0.032
R9037 a_4734_12432.t5 a_4734_12432.t4 800.071
R9038 a_4734_12432.n2 a_4734_12432.n1 659.097
R9039 a_4734_12432.n0 a_4734_12432.t7 285.109
R9040 a_4734_12432.n1 a_4734_12432.t5 193.602
R9041 a_4734_12432.n4 a_4734_12432.n3 192.754
R9042 a_4734_12432.n0 a_4734_12432.t6 160.666
R9043 a_4734_12432.n1 a_4734_12432.n0 91.507
R9044 a_4734_12432.n3 a_4734_12432.t1 28.568
R9045 a_4734_12432.n4 a_4734_12432.t2 28.565
R9046 a_4734_12432.t3 a_4734_12432.n4 28.565
R9047 a_4734_12432.n2 a_4734_12432.t0 19.061
R9048 a_4734_12432.n3 a_4734_12432.n2 1.005
R9049 a_21202_27284.t6 a_21202_27284.n2 404.877
R9050 a_21202_27284.n1 a_21202_27284.t8 210.902
R9051 a_21202_27284.n3 a_21202_27284.t6 136.943
R9052 a_21202_27284.n2 a_21202_27284.n1 107.801
R9053 a_21202_27284.n1 a_21202_27284.t7 80.333
R9054 a_21202_27284.n2 a_21202_27284.t5 80.333
R9055 a_21202_27284.n0 a_21202_27284.t0 17.4
R9056 a_21202_27284.n0 a_21202_27284.t1 17.4
R9057 a_21202_27284.n4 a_21202_27284.t3 15.032
R9058 a_21202_27284.t2 a_21202_27284.n5 14.282
R9059 a_21202_27284.n5 a_21202_27284.t4 14.282
R9060 a_21202_27284.n5 a_21202_27284.n4 1.65
R9061 a_21202_27284.n3 a_21202_27284.n0 0.672
R9062 a_21202_27284.n4 a_21202_27284.n3 0.665
R9063 a_19247_4128.n0 a_19247_4128.t7 14.282
R9064 a_19247_4128.t0 a_19247_4128.n0 14.282
R9065 a_19247_4128.n0 a_19247_4128.n12 90.436
R9066 a_19247_4128.n8 a_19247_4128.n11 50.575
R9067 a_19247_4128.n12 a_19247_4128.n8 74.302
R9068 a_19247_4128.n11 a_19247_4128.n10 157.665
R9069 a_19247_4128.n10 a_19247_4128.t4 8.7
R9070 a_19247_4128.n10 a_19247_4128.t1 8.7
R9071 a_19247_4128.n11 a_19247_4128.n9 122.999
R9072 a_19247_4128.n9 a_19247_4128.t6 14.282
R9073 a_19247_4128.n9 a_19247_4128.t5 14.282
R9074 a_19247_4128.n8 a_19247_4128.n7 90.416
R9075 a_19247_4128.n7 a_19247_4128.t2 14.282
R9076 a_19247_4128.n7 a_19247_4128.t3 14.282
R9077 a_19247_4128.n12 a_19247_4128.n1 342.688
R9078 a_19247_4128.n1 a_19247_4128.n6 126.566
R9079 a_19247_4128.n6 a_19247_4128.t13 294.653
R9080 a_19247_4128.n6 a_19247_4128.t15 111.663
R9081 a_19247_4128.n1 a_19247_4128.n5 552.333
R9082 a_19247_4128.n5 a_19247_4128.n4 6.615
R9083 a_19247_4128.n4 a_19247_4128.t14 93.989
R9084 a_19247_4128.n5 a_19247_4128.n3 97.816
R9085 a_19247_4128.n3 a_19247_4128.t11 80.333
R9086 a_19247_4128.n3 a_19247_4128.t8 394.151
R9087 a_19247_4128.t8 a_19247_4128.n2 269.523
R9088 a_19247_4128.n2 a_19247_4128.t12 160.666
R9089 a_19247_4128.n2 a_19247_4128.t10 269.523
R9090 a_19247_4128.n4 a_19247_4128.t9 198.043
R9091 a_7402_10602.n1 a_7402_10602.t4 318.922
R9092 a_7402_10602.n0 a_7402_10602.t5 273.935
R9093 a_7402_10602.n0 a_7402_10602.t6 273.935
R9094 a_7402_10602.n1 a_7402_10602.t7 269.116
R9095 a_7402_10602.n4 a_7402_10602.n3 193.227
R9096 a_7402_10602.t4 a_7402_10602.n0 179.142
R9097 a_7402_10602.n2 a_7402_10602.n1 106.999
R9098 a_7402_10602.n3 a_7402_10602.t3 28.568
R9099 a_7402_10602.n4 a_7402_10602.t1 28.565
R9100 a_7402_10602.t0 a_7402_10602.n4 28.565
R9101 a_7402_10602.n2 a_7402_10602.t2 18.149
R9102 a_7402_10602.n3 a_7402_10602.n2 3.726
R9103 a_7829_9909.n0 a_7829_9909.t8 14.282
R9104 a_7829_9909.t0 a_7829_9909.n0 14.282
R9105 a_7829_9909.n1 a_7829_9909.n9 0.001
R9106 a_7829_9909.n0 a_7829_9909.n1 267.767
R9107 a_7829_9909.n9 a_7829_9909.t10 14.282
R9108 a_7829_9909.n9 a_7829_9909.t4 14.282
R9109 a_7829_9909.n1 a_7829_9909.n7 0.669
R9110 a_7829_9909.n7 a_7829_9909.n8 1.511
R9111 a_7829_9909.n8 a_7829_9909.t11 14.282
R9112 a_7829_9909.n8 a_7829_9909.t9 14.282
R9113 a_7829_9909.n7 a_7829_9909.n6 0.227
R9114 a_7829_9909.n6 a_7829_9909.n3 0.575
R9115 a_7829_9909.n6 a_7829_9909.n5 0.2
R9116 a_7829_9909.n5 a_7829_9909.t2 16.058
R9117 a_7829_9909.n5 a_7829_9909.n4 0.999
R9118 a_7829_9909.n4 a_7829_9909.t1 14.282
R9119 a_7829_9909.n4 a_7829_9909.t3 14.282
R9120 a_7829_9909.n3 a_7829_9909.n2 0.999
R9121 a_7829_9909.n2 a_7829_9909.t7 14.282
R9122 a_7829_9909.n2 a_7829_9909.t5 14.282
R9123 a_7829_9909.n3 a_7829_9909.t6 16.058
R9124 a_29837_4295.n4 a_29837_4295.t9 214.335
R9125 a_29837_4295.t8 a_29837_4295.n4 214.335
R9126 a_29837_4295.n5 a_29837_4295.t8 143.851
R9127 a_29837_4295.n5 a_29837_4295.t7 135.658
R9128 a_29837_4295.n4 a_29837_4295.t10 80.333
R9129 a_29837_4295.n0 a_29837_4295.t3 28.565
R9130 a_29837_4295.n0 a_29837_4295.t2 28.565
R9131 a_29837_4295.n2 a_29837_4295.t5 28.565
R9132 a_29837_4295.n2 a_29837_4295.t4 28.565
R9133 a_29837_4295.t0 a_29837_4295.n7 28.565
R9134 a_29837_4295.n7 a_29837_4295.t6 28.565
R9135 a_29837_4295.n1 a_29837_4295.t1 9.714
R9136 a_29837_4295.n1 a_29837_4295.n0 1.003
R9137 a_29837_4295.n6 a_29837_4295.n3 0.833
R9138 a_29837_4295.n3 a_29837_4295.n2 0.653
R9139 a_29837_4295.n7 a_29837_4295.n6 0.653
R9140 a_29837_4295.n3 a_29837_4295.n1 0.341
R9141 a_29837_4295.n6 a_29837_4295.n5 0.032
R9142 a_30074_3658.t0 a_30074_3658.t1 17.4
R9143 a_1844_12699.n4 a_1844_12699.n3 535.449
R9144 a_1844_12699.t4 a_1844_12699.t16 437.233
R9145 a_1844_12699.t17 a_1844_12699.t8 437.233
R9146 a_1844_12699.t5 a_1844_12699.n1 313.873
R9147 a_1844_12699.n3 a_1844_12699.t14 294.986
R9148 a_1844_12699.n0 a_1844_12699.t6 272.288
R9149 a_1844_12699.n4 a_1844_12699.t7 245.184
R9150 a_1844_12699.n6 a_1844_12699.t17 218.628
R9151 a_1844_12699.n8 a_1844_12699.t4 217.024
R9152 a_1844_12699.n7 a_1844_12699.t9 214.686
R9153 a_1844_12699.t16 a_1844_12699.n7 214.686
R9154 a_1844_12699.n5 a_1844_12699.t10 214.686
R9155 a_1844_12699.t8 a_1844_12699.n5 214.686
R9156 a_1844_12699.n11 a_1844_12699.n10 192.754
R9157 a_1844_12699.n2 a_1844_12699.t5 190.152
R9158 a_1844_12699.n2 a_1844_12699.t13 190.152
R9159 a_1844_12699.n0 a_1844_12699.t11 160.666
R9160 a_1844_12699.n1 a_1844_12699.t12 160.666
R9161 a_1844_12699.n3 a_1844_12699.t18 110.859
R9162 a_1844_12699.n1 a_1844_12699.n0 96.129
R9163 a_1844_12699.n7 a_1844_12699.t15 80.333
R9164 a_1844_12699.t7 a_1844_12699.n2 80.333
R9165 a_1844_12699.n5 a_1844_12699.t19 80.333
R9166 a_1844_12699.n10 a_1844_12699.t2 28.568
R9167 a_1844_12699.t0 a_1844_12699.n11 28.565
R9168 a_1844_12699.n11 a_1844_12699.t1 28.565
R9169 a_1844_12699.n9 a_1844_12699.t3 18.726
R9170 a_1844_12699.n6 a_1844_12699.n4 14.9
R9171 a_1844_12699.n8 a_1844_12699.n6 2.599
R9172 a_1844_12699.n9 a_1844_12699.n8 2.514
R9173 a_1844_12699.n10 a_1844_12699.n9 1.123
R9174 a_4381_12232.t0 a_4381_12232.t1 17.4
R9175 a_20900_24452.n0 a_20900_24452.t6 14.282
R9176 a_20900_24452.t0 a_20900_24452.n0 14.282
R9177 a_20900_24452.n0 a_20900_24452.n12 90.416
R9178 a_20900_24452.n12 a_20900_24452.n11 50.575
R9179 a_20900_24452.n12 a_20900_24452.n8 74.302
R9180 a_20900_24452.n11 a_20900_24452.n10 157.665
R9181 a_20900_24452.n10 a_20900_24452.t4 8.7
R9182 a_20900_24452.n10 a_20900_24452.t3 8.7
R9183 a_20900_24452.n11 a_20900_24452.n9 122.999
R9184 a_20900_24452.n9 a_20900_24452.t5 14.282
R9185 a_20900_24452.n9 a_20900_24452.t7 14.282
R9186 a_20900_24452.n8 a_20900_24452.n7 90.436
R9187 a_20900_24452.n7 a_20900_24452.t1 14.282
R9188 a_20900_24452.n7 a_20900_24452.t2 14.282
R9189 a_20900_24452.n8 a_20900_24452.n1 342.688
R9190 a_20900_24452.n1 a_20900_24452.n6 126.566
R9191 a_20900_24452.n6 a_20900_24452.t14 294.653
R9192 a_20900_24452.n6 a_20900_24452.t8 111.663
R9193 a_20900_24452.n1 a_20900_24452.n5 552.333
R9194 a_20900_24452.n5 a_20900_24452.n4 6.615
R9195 a_20900_24452.n4 a_20900_24452.t12 93.989
R9196 a_20900_24452.n5 a_20900_24452.n3 97.816
R9197 a_20900_24452.n3 a_20900_24452.t13 80.333
R9198 a_20900_24452.n3 a_20900_24452.t15 394.151
R9199 a_20900_24452.t15 a_20900_24452.n2 269.523
R9200 a_20900_24452.n2 a_20900_24452.t10 160.666
R9201 a_20900_24452.n2 a_20900_24452.t9 269.523
R9202 a_20900_24452.n4 a_20900_24452.t11 198.043
R9203 a_22253_25145.n2 a_22253_25145.t5 318.922
R9204 a_22253_25145.n1 a_22253_25145.t4 273.935
R9205 a_22253_25145.n1 a_22253_25145.t6 273.935
R9206 a_22253_25145.n2 a_22253_25145.t7 269.116
R9207 a_22253_25145.n4 a_22253_25145.n0 193.227
R9208 a_22253_25145.t5 a_22253_25145.n1 179.142
R9209 a_22253_25145.n3 a_22253_25145.n2 106.999
R9210 a_22253_25145.t3 a_22253_25145.n4 28.568
R9211 a_22253_25145.n0 a_22253_25145.t1 28.565
R9212 a_22253_25145.n0 a_22253_25145.t2 28.565
R9213 a_22253_25145.n3 a_22253_25145.t0 18.149
R9214 a_22253_25145.n4 a_22253_25145.n3 3.726
R9215 a_26571_21032.t7 a_26571_21032.n2 404.877
R9216 a_26571_21032.n1 a_26571_21032.t5 210.902
R9217 a_26571_21032.n3 a_26571_21032.t7 136.949
R9218 a_26571_21032.n2 a_26571_21032.n1 107.801
R9219 a_26571_21032.n1 a_26571_21032.t6 80.333
R9220 a_26571_21032.n2 a_26571_21032.t8 80.333
R9221 a_26571_21032.n0 a_26571_21032.t3 17.4
R9222 a_26571_21032.n0 a_26571_21032.t0 17.4
R9223 a_26571_21032.n4 a_26571_21032.t2 15.032
R9224 a_26571_21032.t1 a_26571_21032.n5 14.282
R9225 a_26571_21032.n5 a_26571_21032.t4 14.282
R9226 a_26571_21032.n5 a_26571_21032.n4 1.65
R9227 a_26571_21032.n3 a_26571_21032.n0 0.657
R9228 a_26571_21032.n4 a_26571_21032.n3 0.614
R9229 a_25504_21666.t6 a_25504_21666.t7 800.071
R9230 a_25504_21666.n3 a_25504_21666.n2 672.95
R9231 a_25504_21666.n1 a_25504_21666.t4 285.109
R9232 a_25504_21666.n2 a_25504_21666.t6 193.602
R9233 a_25504_21666.n1 a_25504_21666.t5 160.666
R9234 a_25504_21666.n2 a_25504_21666.n1 91.507
R9235 a_25504_21666.n0 a_25504_21666.t1 28.57
R9236 a_25504_21666.n4 a_25504_21666.t2 28.565
R9237 a_25504_21666.t3 a_25504_21666.n4 28.565
R9238 a_25504_21666.n0 a_25504_21666.t0 17.638
R9239 a_25504_21666.n4 a_25504_21666.n3 0.693
R9240 a_25504_21666.n3 a_25504_21666.n0 0.597
R9241 a_27340_24456.t3 a_27340_24456.n0 14.282
R9242 a_27340_24456.n0 a_27340_24456.t9 14.282
R9243 a_27340_24456.n0 a_27340_24456.n9 0.999
R9244 a_27340_24456.n9 a_27340_24456.n6 0.575
R9245 a_27340_24456.n6 a_27340_24456.n8 0.2
R9246 a_27340_24456.n8 a_27340_24456.t5 16.058
R9247 a_27340_24456.n8 a_27340_24456.n7 0.999
R9248 a_27340_24456.n7 a_27340_24456.t10 14.282
R9249 a_27340_24456.n7 a_27340_24456.t11 14.282
R9250 a_27340_24456.n9 a_27340_24456.t4 16.058
R9251 a_27340_24456.n6 a_27340_24456.n4 0.227
R9252 a_27340_24456.n4 a_27340_24456.n5 1.511
R9253 a_27340_24456.n5 a_27340_24456.t8 14.282
R9254 a_27340_24456.n5 a_27340_24456.t7 14.282
R9255 a_27340_24456.n4 a_27340_24456.n1 0.669
R9256 a_27340_24456.n1 a_27340_24456.n2 0.001
R9257 a_27340_24456.n1 a_27340_24456.n3 267.767
R9258 a_27340_24456.n3 a_27340_24456.t1 14.282
R9259 a_27340_24456.n3 a_27340_24456.t0 14.282
R9260 a_27340_24456.n2 a_27340_24456.t6 14.282
R9261 a_27340_24456.n2 a_27340_24456.t2 14.282
R9262 a_15928_27293.n0 a_15928_27293.t3 14.282
R9263 a_15928_27293.n0 a_15928_27293.t4 14.282
R9264 a_15928_27293.n1 a_15928_27293.t2 14.282
R9265 a_15928_27293.n1 a_15928_27293.t1 14.282
R9266 a_15928_27293.t0 a_15928_27293.n3 14.282
R9267 a_15928_27293.n3 a_15928_27293.t5 14.282
R9268 a_15928_27293.n2 a_15928_27293.n0 2.546
R9269 a_15928_27293.n2 a_15928_27293.n1 2.367
R9270 a_15928_27293.n3 a_15928_27293.n2 0.001
R9271 a_27420_18830.n2 a_27420_18830.t4 318.922
R9272 a_27420_18830.n1 a_27420_18830.t7 273.935
R9273 a_27420_18830.n1 a_27420_18830.t5 273.935
R9274 a_27420_18830.n2 a_27420_18830.t6 269.116
R9275 a_27420_18830.n4 a_27420_18830.n0 193.227
R9276 a_27420_18830.t4 a_27420_18830.n1 179.142
R9277 a_27420_18830.n3 a_27420_18830.n2 106.999
R9278 a_27420_18830.t3 a_27420_18830.n4 28.568
R9279 a_27420_18830.n0 a_27420_18830.t1 28.565
R9280 a_27420_18830.n0 a_27420_18830.t2 28.565
R9281 a_27420_18830.n3 a_27420_18830.t0 18.149
R9282 a_27420_18830.n4 a_27420_18830.n3 3.726
R9283 a_24568_19252.n6 a_24568_19252.n5 501.28
R9284 a_24568_19252.t7 a_24568_19252.t6 437.233
R9285 a_24568_19252.t18 a_24568_19252.t8 415.315
R9286 a_24568_19252.t15 a_24568_19252.n3 313.873
R9287 a_24568_19252.n5 a_24568_19252.t17 294.986
R9288 a_24568_19252.n2 a_24568_19252.t16 272.288
R9289 a_24568_19252.n6 a_24568_19252.t13 236.009
R9290 a_24568_19252.n9 a_24568_19252.t7 216.627
R9291 a_24568_19252.n7 a_24568_19252.t18 216.111
R9292 a_24568_19252.n8 a_24568_19252.t11 214.686
R9293 a_24568_19252.t6 a_24568_19252.n8 214.686
R9294 a_24568_19252.n1 a_24568_19252.t5 214.335
R9295 a_24568_19252.t8 a_24568_19252.n1 214.335
R9296 a_24568_19252.n4 a_24568_19252.t12 190.152
R9297 a_24568_19252.n4 a_24568_19252.t15 190.152
R9298 a_24568_19252.n2 a_24568_19252.t14 160.666
R9299 a_24568_19252.n3 a_24568_19252.t9 160.666
R9300 a_24568_19252.n7 a_24568_19252.n6 148.428
R9301 a_24568_19252.n5 a_24568_19252.t4 110.859
R9302 a_24568_19252.n3 a_24568_19252.n2 96.129
R9303 a_24568_19252.n8 a_24568_19252.t10 80.333
R9304 a_24568_19252.n1 a_24568_19252.t19 80.333
R9305 a_24568_19252.t13 a_24568_19252.n4 80.333
R9306 a_24568_19252.n0 a_24568_19252.t1 28.57
R9307 a_24568_19252.n11 a_24568_19252.t2 28.565
R9308 a_24568_19252.t3 a_24568_19252.n11 28.565
R9309 a_24568_19252.n0 a_24568_19252.t0 17.638
R9310 a_24568_19252.n10 a_24568_19252.n9 10.943
R9311 a_24568_19252.n9 a_24568_19252.n7 2.923
R9312 a_24568_19252.n11 a_24568_19252.n10 0.69
R9313 a_24568_19252.n10 a_24568_19252.n0 0.6
R9314 a_24570_19549.n1 a_24570_19549.t7 318.922
R9315 a_24570_19549.n0 a_24570_19549.t6 274.739
R9316 a_24570_19549.n0 a_24570_19549.t4 274.739
R9317 a_24570_19549.n1 a_24570_19549.t5 269.116
R9318 a_24570_19549.t7 a_24570_19549.n0 179.946
R9319 a_24570_19549.n2 a_24570_19549.n1 105.178
R9320 a_24570_19549.t3 a_24570_19549.n4 29.444
R9321 a_24570_19549.n3 a_24570_19549.t1 28.565
R9322 a_24570_19549.n3 a_24570_19549.t2 28.565
R9323 a_24570_19549.n2 a_24570_19549.t0 18.145
R9324 a_24570_19549.n4 a_24570_19549.n2 2.878
R9325 a_24570_19549.n4 a_24570_19549.n3 0.764
R9326 a_6049_9909.n0 a_6049_9909.n12 122.999
R9327 a_6049_9909.t0 a_6049_9909.n0 14.282
R9328 a_6049_9909.n0 a_6049_9909.t7 14.282
R9329 a_6049_9909.n12 a_6049_9909.n10 50.575
R9330 a_6049_9909.n10 a_6049_9909.n8 74.302
R9331 a_6049_9909.n12 a_6049_9909.n11 157.665
R9332 a_6049_9909.n11 a_6049_9909.t6 8.7
R9333 a_6049_9909.n11 a_6049_9909.t1 8.7
R9334 a_6049_9909.n10 a_6049_9909.n9 90.416
R9335 a_6049_9909.n9 a_6049_9909.t5 14.282
R9336 a_6049_9909.n9 a_6049_9909.t3 14.282
R9337 a_6049_9909.n8 a_6049_9909.n7 90.436
R9338 a_6049_9909.n7 a_6049_9909.t2 14.282
R9339 a_6049_9909.n7 a_6049_9909.t4 14.282
R9340 a_6049_9909.n8 a_6049_9909.n1 342.688
R9341 a_6049_9909.n1 a_6049_9909.n6 126.566
R9342 a_6049_9909.n6 a_6049_9909.t12 294.653
R9343 a_6049_9909.n6 a_6049_9909.t14 111.663
R9344 a_6049_9909.n1 a_6049_9909.n5 552.333
R9345 a_6049_9909.n5 a_6049_9909.n4 6.615
R9346 a_6049_9909.n4 a_6049_9909.t8 93.989
R9347 a_6049_9909.n5 a_6049_9909.n3 97.816
R9348 a_6049_9909.n3 a_6049_9909.t9 80.333
R9349 a_6049_9909.n3 a_6049_9909.t13 394.151
R9350 a_6049_9909.t13 a_6049_9909.n2 269.523
R9351 a_6049_9909.n2 a_6049_9909.t10 160.666
R9352 a_6049_9909.n2 a_6049_9909.t11 269.523
R9353 a_6049_9909.n4 a_6049_9909.t15 198.043
R9354 a_36751_1089.t0 a_36751_1089.n0 14.282
R9355 a_36751_1089.n0 a_36751_1089.t2 14.282
R9356 a_36751_1089.n0 a_36751_1089.n9 89.977
R9357 a_36751_1089.n4 a_36751_1089.n2 77.784
R9358 a_36751_1089.n6 a_36751_1089.n4 77.456
R9359 a_36751_1089.n9 a_36751_1089.n6 77.456
R9360 a_36751_1089.n9 a_36751_1089.n7 75.815
R9361 a_36751_1089.n7 a_36751_1089.n8 167.433
R9362 a_36751_1089.n8 a_36751_1089.t4 14.282
R9363 a_36751_1089.n8 a_36751_1089.t1 14.282
R9364 a_36751_1089.n7 a_36751_1089.t5 104.259
R9365 a_36751_1089.n6 a_36751_1089.n5 89.977
R9366 a_36751_1089.n5 a_36751_1089.t9 14.282
R9367 a_36751_1089.n5 a_36751_1089.t3 14.282
R9368 a_36751_1089.n4 a_36751_1089.n3 89.977
R9369 a_36751_1089.n3 a_36751_1089.t11 14.282
R9370 a_36751_1089.n3 a_36751_1089.t10 14.282
R9371 a_36751_1089.n2 a_36751_1089.t6 104.259
R9372 a_36751_1089.n2 a_36751_1089.n1 167.433
R9373 a_36751_1089.n1 a_36751_1089.t7 14.282
R9374 a_36751_1089.n1 a_36751_1089.t8 14.282
R9375 a_33375_14481.n0 a_33375_14481.t10 214.335
R9376 a_33375_14481.t8 a_33375_14481.n0 214.335
R9377 a_33375_14481.n1 a_33375_14481.t8 143.851
R9378 a_33375_14481.n1 a_33375_14481.t7 135.658
R9379 a_33375_14481.n0 a_33375_14481.t9 80.333
R9380 a_33375_14481.n2 a_33375_14481.t4 28.565
R9381 a_33375_14481.n2 a_33375_14481.t5 28.565
R9382 a_33375_14481.n4 a_33375_14481.t6 28.565
R9383 a_33375_14481.n4 a_33375_14481.t1 28.565
R9384 a_33375_14481.n7 a_33375_14481.t2 28.565
R9385 a_33375_14481.t3 a_33375_14481.n7 28.565
R9386 a_33375_14481.n6 a_33375_14481.t0 9.714
R9387 a_33375_14481.n7 a_33375_14481.n6 1.003
R9388 a_33375_14481.n5 a_33375_14481.n3 0.833
R9389 a_33375_14481.n3 a_33375_14481.n2 0.653
R9390 a_33375_14481.n5 a_33375_14481.n4 0.653
R9391 a_33375_14481.n6 a_33375_14481.n5 0.341
R9392 a_33375_14481.n3 a_33375_14481.n1 0.032
R9393 a_5623_18852.t0 a_5623_18852.n0 14.282
R9394 a_5623_18852.n0 a_5623_18852.t6 14.282
R9395 a_5623_18852.n0 a_5623_18852.n8 90.416
R9396 a_5623_18852.n8 a_5623_18852.n5 74.302
R9397 a_5623_18852.n8 a_5623_18852.n7 50.575
R9398 a_5623_18852.n7 a_5623_18852.n6 157.665
R9399 a_5623_18852.n6 a_5623_18852.t7 8.7
R9400 a_5623_18852.n6 a_5623_18852.t3 8.7
R9401 a_5623_18852.n5 a_5623_18852.n4 90.436
R9402 a_5623_18852.n4 a_5623_18852.t2 14.282
R9403 a_5623_18852.n4 a_5623_18852.t1 14.282
R9404 a_5623_18852.n7 a_5623_18852.n3 122.746
R9405 a_5623_18852.n3 a_5623_18852.t5 14.282
R9406 a_5623_18852.n3 a_5623_18852.t4 14.282
R9407 a_5623_18852.n5 a_5623_18852.n1 293.294
R9408 a_5623_18852.t11 a_5623_18852.n2 160.666
R9409 a_5623_18852.n1 a_5623_18852.t11 867.393
R9410 a_5623_18852.n2 a_5623_18852.t9 287.241
R9411 a_5623_18852.n2 a_5623_18852.t8 287.241
R9412 a_5623_18852.n1 a_5623_18852.t10 545.094
R9413 a_5505_18852.n3 a_5505_18852.n1 267.767
R9414 a_5505_18852.n7 a_5505_18852.t3 16.058
R9415 a_5505_18852.t2 a_5505_18852.n9 16.058
R9416 a_5505_18852.n2 a_5505_18852.t8 14.282
R9417 a_5505_18852.n2 a_5505_18852.t9 14.282
R9418 a_5505_18852.n1 a_5505_18852.t10 14.282
R9419 a_5505_18852.n1 a_5505_18852.t11 14.282
R9420 a_5505_18852.n4 a_5505_18852.t7 14.282
R9421 a_5505_18852.n4 a_5505_18852.t6 14.282
R9422 a_5505_18852.n0 a_5505_18852.t0 14.282
R9423 a_5505_18852.n0 a_5505_18852.t1 14.282
R9424 a_5505_18852.n6 a_5505_18852.t4 14.282
R9425 a_5505_18852.n6 a_5505_18852.t5 14.282
R9426 a_5505_18852.n5 a_5505_18852.n4 1.511
R9427 a_5505_18852.n9 a_5505_18852.n0 0.999
R9428 a_5505_18852.n7 a_5505_18852.n6 0.999
R9429 a_5505_18852.n5 a_5505_18852.n3 0.669
R9430 a_5505_18852.n8 a_5505_18852.n7 0.575
R9431 a_5505_18852.n8 a_5505_18852.n5 0.227
R9432 a_5505_18852.n9 a_5505_18852.n8 0.2
R9433 a_5505_18852.n3 a_5505_18852.n2 0.001
R9434 a_4158_11219.n0 a_4158_11219.t8 214.335
R9435 a_4158_11219.t9 a_4158_11219.n0 214.335
R9436 a_4158_11219.n1 a_4158_11219.t9 143.851
R9437 a_4158_11219.n1 a_4158_11219.t7 135.658
R9438 a_4158_11219.n0 a_4158_11219.t10 80.333
R9439 a_4158_11219.n2 a_4158_11219.t3 28.565
R9440 a_4158_11219.n2 a_4158_11219.t1 28.565
R9441 a_4158_11219.n4 a_4158_11219.t2 28.565
R9442 a_4158_11219.n4 a_4158_11219.t4 28.565
R9443 a_4158_11219.n7 a_4158_11219.t6 28.565
R9444 a_4158_11219.t0 a_4158_11219.n7 28.565
R9445 a_4158_11219.n6 a_4158_11219.t5 9.714
R9446 a_4158_11219.n7 a_4158_11219.n6 1.003
R9447 a_4158_11219.n5 a_4158_11219.n3 0.833
R9448 a_4158_11219.n3 a_4158_11219.n2 0.653
R9449 a_4158_11219.n5 a_4158_11219.n4 0.653
R9450 a_4158_11219.n6 a_4158_11219.n5 0.341
R9451 a_4158_11219.n3 a_4158_11219.n1 0.032
R9452 a_6253_21662.t6 a_6253_21662.t7 574.43
R9453 a_6253_21662.n1 a_6253_21662.t4 285.109
R9454 a_6253_21662.n3 a_6253_21662.n2 211.134
R9455 a_6253_21662.n4 a_6253_21662.n0 192.754
R9456 a_6253_21662.n1 a_6253_21662.t5 160.666
R9457 a_6253_21662.n2 a_6253_21662.t6 160.666
R9458 a_6253_21662.n2 a_6253_21662.n1 114.829
R9459 a_6253_21662.t3 a_6253_21662.n4 28.568
R9460 a_6253_21662.n0 a_6253_21662.t1 28.565
R9461 a_6253_21662.n0 a_6253_21662.t2 28.565
R9462 a_6253_21662.n3 a_6253_21662.t0 19.087
R9463 a_6253_21662.n4 a_6253_21662.n3 1.051
R9464 a_5824_21032.t5 a_5824_21032.n2 404.877
R9465 a_5824_21032.n1 a_5824_21032.t7 210.902
R9466 a_5824_21032.n3 a_5824_21032.t5 136.949
R9467 a_5824_21032.n2 a_5824_21032.n1 107.801
R9468 a_5824_21032.n1 a_5824_21032.t8 80.333
R9469 a_5824_21032.n2 a_5824_21032.t6 80.333
R9470 a_5824_21032.n0 a_5824_21032.t1 17.4
R9471 a_5824_21032.n0 a_5824_21032.t0 17.4
R9472 a_5824_21032.n4 a_5824_21032.t2 15.032
R9473 a_5824_21032.n5 a_5824_21032.t3 14.282
R9474 a_5824_21032.t4 a_5824_21032.n5 14.282
R9475 a_5824_21032.n5 a_5824_21032.n4 1.65
R9476 a_5824_21032.n3 a_5824_21032.n0 0.657
R9477 a_5824_21032.n4 a_5824_21032.n3 0.614
R9478 a_6343_9883.n1 a_6343_9883.t5 318.922
R9479 a_6343_9883.n0 a_6343_9883.t6 274.739
R9480 a_6343_9883.n0 a_6343_9883.t7 274.739
R9481 a_6343_9883.n1 a_6343_9883.t4 269.116
R9482 a_6343_9883.t5 a_6343_9883.n0 179.946
R9483 a_6343_9883.n2 a_6343_9883.n1 107.263
R9484 a_6343_9883.n3 a_6343_9883.t1 29.444
R9485 a_6343_9883.n4 a_6343_9883.t2 28.565
R9486 a_6343_9883.t3 a_6343_9883.n4 28.565
R9487 a_6343_9883.n2 a_6343_9883.t0 18.145
R9488 a_6343_9883.n3 a_6343_9883.n2 2.878
R9489 a_6343_9883.n4 a_6343_9883.n3 0.764
R9490 a_n3604_10397.n1 a_n3604_10397.t4 318.119
R9491 a_n3604_10397.n1 a_n3604_10397.t5 269.919
R9492 a_n3604_10397.n0 a_n3604_10397.t6 267.853
R9493 a_n3604_10397.n0 a_n3604_10397.t7 267.853
R9494 a_n3604_10397.t4 a_n3604_10397.n0 160.666
R9495 a_n3604_10397.n2 a_n3604_10397.n1 107.263
R9496 a_n3604_10397.n3 a_n3604_10397.t3 29.444
R9497 a_n3604_10397.t0 a_n3604_10397.n4 28.565
R9498 a_n3604_10397.n4 a_n3604_10397.t1 28.565
R9499 a_n3604_10397.n2 a_n3604_10397.t2 18.145
R9500 a_n3604_10397.n3 a_n3604_10397.n2 2.878
R9501 a_n3604_10397.n4 a_n3604_10397.n3 0.764
R9502 a_n3111_11055.t0 a_n3111_11055.n0 14.282
R9503 a_n3111_11055.n0 a_n3111_11055.t2 14.282
R9504 a_n3111_11055.n0 a_n3111_11055.n16 90.436
R9505 a_n3111_11055.n16 a_n3111_11055.n2 74.302
R9506 a_n3111_11055.n2 a_n3111_11055.n4 50.575
R9507 a_n3111_11055.n4 a_n3111_11055.n5 110.084
R9508 a_n3111_11055.n16 a_n3111_11055.n6 210.799
R9509 a_n3111_11055.n6 a_n3111_11055.n8 16.411
R9510 a_n3111_11055.n8 a_n3111_11055.t10 198.921
R9511 a_n3111_11055.t10 a_n3111_11055.t11 415.315
R9512 a_n3111_11055.t11 a_n3111_11055.n15 214.335
R9513 a_n3111_11055.n15 a_n3111_11055.t12 80.333
R9514 a_n3111_11055.n15 a_n3111_11055.t17 214.335
R9515 a_n3111_11055.n8 a_n3111_11055.n14 861.987
R9516 a_n3111_11055.n14 a_n3111_11055.n9 560.726
R9517 a_n3111_11055.n14 a_n3111_11055.n13 65.07
R9518 a_n3111_11055.n13 a_n3111_11055.n12 6.615
R9519 a_n3111_11055.n12 a_n3111_11055.t21 93.989
R9520 a_n3111_11055.n13 a_n3111_11055.n11 97.816
R9521 a_n3111_11055.n11 a_n3111_11055.t8 80.333
R9522 a_n3111_11055.n11 a_n3111_11055.t13 394.151
R9523 a_n3111_11055.t13 a_n3111_11055.n10 269.523
R9524 a_n3111_11055.n10 a_n3111_11055.t18 160.666
R9525 a_n3111_11055.n10 a_n3111_11055.t19 269.523
R9526 a_n3111_11055.n12 a_n3111_11055.t20 198.043
R9527 a_n3111_11055.n9 a_n3111_11055.t9 294.653
R9528 a_n3111_11055.n9 a_n3111_11055.t16 111.663
R9529 a_n3111_11055.n6 a_n3111_11055.t22 217.716
R9530 a_n3111_11055.t22 a_n3111_11055.t23 415.315
R9531 a_n3111_11055.t23 a_n3111_11055.n7 214.335
R9532 a_n3111_11055.n7 a_n3111_11055.t14 80.333
R9533 a_n3111_11055.n7 a_n3111_11055.t15 214.335
R9534 a_n3111_11055.n5 a_n3111_11055.t7 14.282
R9535 a_n3111_11055.n5 a_n3111_11055.t5 14.282
R9536 a_n3111_11055.n4 a_n3111_11055.n3 157.665
R9537 a_n3111_11055.n3 a_n3111_11055.t3 8.7
R9538 a_n3111_11055.n3 a_n3111_11055.t4 8.7
R9539 a_n3111_11055.n2 a_n3111_11055.n1 90.416
R9540 a_n3111_11055.n1 a_n3111_11055.t1 14.282
R9541 a_n3111_11055.n1 a_n3111_11055.t6 14.282
R9542 a_n3804_10998.t3 a_n3804_10998.n0 14.282
R9543 a_n3804_10998.n0 a_n3804_10998.t7 14.282
R9544 a_n3804_10998.n1 a_n3804_10998.n9 0.001
R9545 a_n3804_10998.n0 a_n3804_10998.n1 267.767
R9546 a_n3804_10998.n9 a_n3804_10998.t8 14.282
R9547 a_n3804_10998.n9 a_n3804_10998.t6 14.282
R9548 a_n3804_10998.n1 a_n3804_10998.n7 0.669
R9549 a_n3804_10998.n7 a_n3804_10998.n8 1.511
R9550 a_n3804_10998.n8 a_n3804_10998.t5 14.282
R9551 a_n3804_10998.n8 a_n3804_10998.t4 14.282
R9552 a_n3804_10998.n7 a_n3804_10998.n6 0.227
R9553 a_n3804_10998.n6 a_n3804_10998.n5 0.2
R9554 a_n3804_10998.n6 a_n3804_10998.n3 0.575
R9555 a_n3804_10998.n5 a_n3804_10998.t0 16.058
R9556 a_n3804_10998.n5 a_n3804_10998.n4 0.999
R9557 a_n3804_10998.n4 a_n3804_10998.t2 14.282
R9558 a_n3804_10998.n4 a_n3804_10998.t1 14.282
R9559 a_n3804_10998.n3 a_n3804_10998.n2 0.999
R9560 a_n3804_10998.n2 a_n3804_10998.t10 14.282
R9561 a_n3804_10998.n2 a_n3804_10998.t11 14.282
R9562 a_n3804_10998.n3 a_n3804_10998.t9 16.058
R9563 a_12811_21658.t7 a_12811_21658.t5 574.43
R9564 a_12811_21658.n1 a_12811_21658.t6 285.109
R9565 a_12811_21658.n3 a_12811_21658.n2 211.134
R9566 a_12811_21658.n4 a_12811_21658.n0 192.754
R9567 a_12811_21658.n1 a_12811_21658.t4 160.666
R9568 a_12811_21658.n2 a_12811_21658.t7 160.666
R9569 a_12811_21658.n2 a_12811_21658.n1 114.829
R9570 a_12811_21658.t3 a_12811_21658.n4 28.568
R9571 a_12811_21658.n0 a_12811_21658.t1 28.565
R9572 a_12811_21658.n0 a_12811_21658.t2 28.565
R9573 a_12811_21658.n3 a_12811_21658.t0 19.087
R9574 a_12811_21658.n4 a_12811_21658.n3 1.051
R9575 a_12382_21028.t5 a_12382_21028.n3 404.877
R9576 a_12382_21028.n2 a_12382_21028.t6 210.902
R9577 a_12382_21028.n4 a_12382_21028.t5 136.949
R9578 a_12382_21028.n3 a_12382_21028.n2 107.801
R9579 a_12382_21028.n2 a_12382_21028.t7 80.333
R9580 a_12382_21028.n3 a_12382_21028.t8 80.333
R9581 a_12382_21028.n1 a_12382_21028.t1 17.4
R9582 a_12382_21028.n1 a_12382_21028.t0 17.4
R9583 a_12382_21028.t2 a_12382_21028.n5 15.032
R9584 a_12382_21028.n0 a_12382_21028.t4 14.282
R9585 a_12382_21028.n0 a_12382_21028.t3 14.282
R9586 a_12382_21028.n5 a_12382_21028.n0 1.65
R9587 a_12382_21028.n4 a_12382_21028.n1 0.657
R9588 a_12382_21028.n5 a_12382_21028.n4 0.614
R9589 a_12517_21684.n1 a_12517_21684.t4 14.282
R9590 a_12517_21684.n1 a_12517_21684.t1 14.282
R9591 a_12517_21684.n0 a_12517_21684.t3 14.282
R9592 a_12517_21684.n0 a_12517_21684.t5 14.282
R9593 a_12517_21684.n3 a_12517_21684.t2 14.282
R9594 a_12517_21684.t0 a_12517_21684.n3 14.282
R9595 a_12517_21684.n2 a_12517_21684.n0 2.546
R9596 a_12517_21684.n3 a_12517_21684.n2 2.367
R9597 a_12517_21684.n2 a_12517_21684.n1 0.001
R9598 a_n3606_12466.n1 a_n3606_12466.t7 318.119
R9599 a_n3606_12466.n1 a_n3606_12466.t6 269.919
R9600 a_n3606_12466.n0 a_n3606_12466.t4 267.853
R9601 a_n3606_12466.n0 a_n3606_12466.t5 267.853
R9602 a_n3606_12466.t7 a_n3606_12466.n0 160.666
R9603 a_n3606_12466.n2 a_n3606_12466.n1 107.263
R9604 a_n3606_12466.t0 a_n3606_12466.n4 29.444
R9605 a_n3606_12466.n3 a_n3606_12466.t3 28.565
R9606 a_n3606_12466.n3 a_n3606_12466.t2 28.565
R9607 a_n3606_12466.n2 a_n3606_12466.t1 18.145
R9608 a_n3606_12466.n4 a_n3606_12466.n2 2.878
R9609 a_n3606_12466.n4 a_n3606_12466.n3 0.764
R9610 a_n3806_13067.t0 a_n3806_13067.n7 16.058
R9611 a_n3806_13067.n5 a_n3806_13067.n9 0.2
R9612 a_n3806_13067.n7 a_n3806_13067.n5 0.575
R9613 a_n3806_13067.n9 a_n3806_13067.t4 16.058
R9614 a_n3806_13067.n9 a_n3806_13067.n8 0.999
R9615 a_n3806_13067.n8 a_n3806_13067.t6 14.282
R9616 a_n3806_13067.n8 a_n3806_13067.t5 14.282
R9617 a_n3806_13067.n7 a_n3806_13067.n6 0.999
R9618 a_n3806_13067.n6 a_n3806_13067.t11 14.282
R9619 a_n3806_13067.n6 a_n3806_13067.t10 14.282
R9620 a_n3806_13067.n5 a_n3806_13067.n3 0.227
R9621 a_n3806_13067.n3 a_n3806_13067.n4 1.511
R9622 a_n3806_13067.n4 a_n3806_13067.t2 14.282
R9623 a_n3806_13067.n4 a_n3806_13067.t1 14.282
R9624 a_n3806_13067.n3 a_n3806_13067.n0 0.669
R9625 a_n3806_13067.n0 a_n3806_13067.n1 0.001
R9626 a_n3806_13067.n0 a_n3806_13067.n2 267.767
R9627 a_n3806_13067.n2 a_n3806_13067.t7 14.282
R9628 a_n3806_13067.n2 a_n3806_13067.t8 14.282
R9629 a_n3806_13067.n1 a_n3806_13067.t9 14.282
R9630 a_n3806_13067.n1 a_n3806_13067.t3 14.282
R9631 a_n3113_13124.n0 a_n3113_13124.t6 14.282
R9632 a_n3113_13124.t0 a_n3113_13124.n0 14.282
R9633 a_n3113_13124.n4 a_n3113_13124.n2 74.302
R9634 a_n3113_13124.n6 a_n3113_13124.n4 50.575
R9635 a_n3113_13124.n0 a_n3113_13124.n6 110.084
R9636 a_n3113_13124.n2 a_n3113_13124.n7 206.242
R9637 a_n3113_13124.n7 a_n3113_13124.n9 16.411
R9638 a_n3113_13124.n9 a_n3113_13124.t17 198.921
R9639 a_n3113_13124.t17 a_n3113_13124.t15 415.315
R9640 a_n3113_13124.t15 a_n3113_13124.n16 214.335
R9641 a_n3113_13124.n16 a_n3113_13124.t16 80.333
R9642 a_n3113_13124.n16 a_n3113_13124.t19 214.335
R9643 a_n3113_13124.n9 a_n3113_13124.n15 861.987
R9644 a_n3113_13124.n15 a_n3113_13124.n10 560.726
R9645 a_n3113_13124.n15 a_n3113_13124.n14 65.07
R9646 a_n3113_13124.n14 a_n3113_13124.n13 6.615
R9647 a_n3113_13124.n13 a_n3113_13124.t22 93.989
R9648 a_n3113_13124.n14 a_n3113_13124.n12 97.816
R9649 a_n3113_13124.n12 a_n3113_13124.t8 80.333
R9650 a_n3113_13124.n12 a_n3113_13124.t13 394.151
R9651 a_n3113_13124.t13 a_n3113_13124.n11 269.523
R9652 a_n3113_13124.n11 a_n3113_13124.t14 160.666
R9653 a_n3113_13124.n11 a_n3113_13124.t18 269.523
R9654 a_n3113_13124.n13 a_n3113_13124.t21 198.043
R9655 a_n3113_13124.n10 a_n3113_13124.t23 294.653
R9656 a_n3113_13124.n10 a_n3113_13124.t9 111.663
R9657 a_n3113_13124.n7 a_n3113_13124.t20 217.716
R9658 a_n3113_13124.t20 a_n3113_13124.t10 415.315
R9659 a_n3113_13124.t10 a_n3113_13124.n8 214.335
R9660 a_n3113_13124.n8 a_n3113_13124.t11 80.333
R9661 a_n3113_13124.n8 a_n3113_13124.t12 214.335
R9662 a_n3113_13124.n6 a_n3113_13124.n5 157.665
R9663 a_n3113_13124.n5 a_n3113_13124.t1 8.7
R9664 a_n3113_13124.n5 a_n3113_13124.t5 8.7
R9665 a_n3113_13124.n4 a_n3113_13124.n3 90.416
R9666 a_n3113_13124.n3 a_n3113_13124.t4 14.282
R9667 a_n3113_13124.n3 a_n3113_13124.t7 14.282
R9668 a_n3113_13124.n2 a_n3113_13124.n1 90.436
R9669 a_n3113_13124.n1 a_n3113_13124.t3 14.282
R9670 a_n3113_13124.n1 a_n3113_13124.t2 14.282
R9671 a_20355_25145.n1 a_20355_25145.t7 318.922
R9672 a_20355_25145.n0 a_20355_25145.t5 273.935
R9673 a_20355_25145.n0 a_20355_25145.t6 273.935
R9674 a_20355_25145.n1 a_20355_25145.t4 269.116
R9675 a_20355_25145.n4 a_20355_25145.n3 193.227
R9676 a_20355_25145.t7 a_20355_25145.n0 179.142
R9677 a_20355_25145.n2 a_20355_25145.n1 106.999
R9678 a_20355_25145.n3 a_20355_25145.t2 28.568
R9679 a_20355_25145.t3 a_20355_25145.n4 28.565
R9680 a_20355_25145.n4 a_20355_25145.t1 28.565
R9681 a_20355_25145.n2 a_20355_25145.t0 18.149
R9682 a_20355_25145.n3 a_20355_25145.n2 3.726
R9683 a_10930_12320.t0 a_10930_12320.t1 17.4
R9684 a_5923_4129.n0 a_5923_4129.t11 14.282
R9685 a_5923_4129.t0 a_5923_4129.n0 14.282
R9686 a_5923_4129.n1 a_5923_4129.n9 0.001
R9687 a_5923_4129.n0 a_5923_4129.n1 267.767
R9688 a_5923_4129.n9 a_5923_4129.t8 14.282
R9689 a_5923_4129.n9 a_5923_4129.t10 14.282
R9690 a_5923_4129.n1 a_5923_4129.n7 0.669
R9691 a_5923_4129.n7 a_5923_4129.n8 1.511
R9692 a_5923_4129.n8 a_5923_4129.t9 14.282
R9693 a_5923_4129.n8 a_5923_4129.t7 14.282
R9694 a_5923_4129.n7 a_5923_4129.n6 0.227
R9695 a_5923_4129.n6 a_5923_4129.n3 0.575
R9696 a_5923_4129.n6 a_5923_4129.n5 0.2
R9697 a_5923_4129.n5 a_5923_4129.t3 16.058
R9698 a_5923_4129.n5 a_5923_4129.n4 0.999
R9699 a_5923_4129.n4 a_5923_4129.t2 14.282
R9700 a_5923_4129.n4 a_5923_4129.t1 14.282
R9701 a_5923_4129.n3 a_5923_4129.n2 0.999
R9702 a_5923_4129.n2 a_5923_4129.t6 14.282
R9703 a_5923_4129.n2 a_5923_4129.t4 14.282
R9704 a_5923_4129.n3 a_5923_4129.t5 16.058
R9705 a_22104_21787.n0 a_22104_21787.t7 214.335
R9706 a_22104_21787.t9 a_22104_21787.n0 214.335
R9707 a_22104_21787.n1 a_22104_21787.t9 143.851
R9708 a_22104_21787.n1 a_22104_21787.t10 135.658
R9709 a_22104_21787.n0 a_22104_21787.t8 80.333
R9710 a_22104_21787.n2 a_22104_21787.t6 28.565
R9711 a_22104_21787.n2 a_22104_21787.t4 28.565
R9712 a_22104_21787.n4 a_22104_21787.t5 28.565
R9713 a_22104_21787.n4 a_22104_21787.t0 28.565
R9714 a_22104_21787.n7 a_22104_21787.t1 28.565
R9715 a_22104_21787.t2 a_22104_21787.n7 28.565
R9716 a_22104_21787.n3 a_22104_21787.t3 9.714
R9717 a_22104_21787.n3 a_22104_21787.n2 1.003
R9718 a_22104_21787.n6 a_22104_21787.n5 0.833
R9719 a_22104_21787.n5 a_22104_21787.n4 0.653
R9720 a_22104_21787.n7 a_22104_21787.n6 0.653
R9721 a_22104_21787.n5 a_22104_21787.n3 0.341
R9722 a_22104_21787.n6 a_22104_21787.n1 0.032
R9723 a_10701_5437.n4 a_10701_5437.t7 214.335
R9724 a_10701_5437.t10 a_10701_5437.n4 214.335
R9725 a_10701_5437.n5 a_10701_5437.t10 143.851
R9726 a_10701_5437.n5 a_10701_5437.t8 135.658
R9727 a_10701_5437.n4 a_10701_5437.t9 80.333
R9728 a_10701_5437.n0 a_10701_5437.t1 28.565
R9729 a_10701_5437.n0 a_10701_5437.t3 28.565
R9730 a_10701_5437.n2 a_10701_5437.t6 28.565
R9731 a_10701_5437.n2 a_10701_5437.t2 28.565
R9732 a_10701_5437.t4 a_10701_5437.n7 28.565
R9733 a_10701_5437.n7 a_10701_5437.t5 28.565
R9734 a_10701_5437.n1 a_10701_5437.t0 9.714
R9735 a_10701_5437.n1 a_10701_5437.n0 1.003
R9736 a_10701_5437.n6 a_10701_5437.n3 0.833
R9737 a_10701_5437.n3 a_10701_5437.n2 0.653
R9738 a_10701_5437.n7 a_10701_5437.n6 0.653
R9739 a_10701_5437.n3 a_10701_5437.n1 0.341
R9740 a_10701_5437.n6 a_10701_5437.n5 0.032
R9741 a_11291_5000.t4 a_11291_5000.t6 574.43
R9742 a_11291_5000.n1 a_11291_5000.t5 285.109
R9743 a_11291_5000.n3 a_11291_5000.n2 211.136
R9744 a_11291_5000.n4 a_11291_5000.n0 192.754
R9745 a_11291_5000.n1 a_11291_5000.t7 160.666
R9746 a_11291_5000.n2 a_11291_5000.t4 160.666
R9747 a_11291_5000.n2 a_11291_5000.n1 114.829
R9748 a_11291_5000.t3 a_11291_5000.n4 28.568
R9749 a_11291_5000.n0 a_11291_5000.t2 28.565
R9750 a_11291_5000.n0 a_11291_5000.t1 28.565
R9751 a_11291_5000.n3 a_11291_5000.t0 19.084
R9752 a_11291_5000.n4 a_11291_5000.n3 1.051
R9753 a_26468_19549.n1 a_26468_19549.t6 318.922
R9754 a_26468_19549.n0 a_26468_19549.t5 274.739
R9755 a_26468_19549.n0 a_26468_19549.t7 274.739
R9756 a_26468_19549.n1 a_26468_19549.t4 269.116
R9757 a_26468_19549.t6 a_26468_19549.n0 179.946
R9758 a_26468_19549.n2 a_26468_19549.n1 107.263
R9759 a_26468_19549.t3 a_26468_19549.n4 29.444
R9760 a_26468_19549.n3 a_26468_19549.t1 28.565
R9761 a_26468_19549.n3 a_26468_19549.t2 28.565
R9762 a_26468_19549.n2 a_26468_19549.t0 18.145
R9763 a_26468_19549.n4 a_26468_19549.n2 2.878
R9764 a_26468_19549.n4 a_26468_19549.n3 0.764
R9765 a_27126_18124.t0 a_27126_18124.t1 380.209
R9766 a_36701_11276.n2 a_36701_11276.t5 448.381
R9767 a_36701_11276.n1 a_36701_11276.t6 287.241
R9768 a_36701_11276.n1 a_36701_11276.t4 287.241
R9769 a_36701_11276.n0 a_36701_11276.t7 247.733
R9770 a_36701_11276.n4 a_36701_11276.n3 182.117
R9771 a_36701_11276.t5 a_36701_11276.n1 160.666
R9772 a_36701_11276.n3 a_36701_11276.t1 28.568
R9773 a_36701_11276.n4 a_36701_11276.t2 28.565
R9774 a_36701_11276.t3 a_36701_11276.n4 28.565
R9775 a_36701_11276.n0 a_36701_11276.t0 18.127
R9776 a_36701_11276.n2 a_36701_11276.n0 4.036
R9777 a_36701_11276.n3 a_36701_11276.n2 0.937
R9778 a_36755_10509.n0 a_36755_10509.t11 14.282
R9779 a_36755_10509.t0 a_36755_10509.n0 14.282
R9780 a_36755_10509.n0 a_36755_10509.n1 167.433
R9781 a_36755_10509.n1 a_36755_10509.n3 77.784
R9782 a_36755_10509.n3 a_36755_10509.n5 77.456
R9783 a_36755_10509.n5 a_36755_10509.n7 77.456
R9784 a_36755_10509.n7 a_36755_10509.n8 75.815
R9785 a_36755_10509.n8 a_36755_10509.n9 167.433
R9786 a_36755_10509.n9 a_36755_10509.t1 14.282
R9787 a_36755_10509.n9 a_36755_10509.t3 14.282
R9788 a_36755_10509.n8 a_36755_10509.t2 104.259
R9789 a_36755_10509.n7 a_36755_10509.n6 89.977
R9790 a_36755_10509.n6 a_36755_10509.t8 14.282
R9791 a_36755_10509.n6 a_36755_10509.t7 14.282
R9792 a_36755_10509.n5 a_36755_10509.n4 89.977
R9793 a_36755_10509.n4 a_36755_10509.t4 14.282
R9794 a_36755_10509.n4 a_36755_10509.t9 14.282
R9795 a_36755_10509.n3 a_36755_10509.n2 89.977
R9796 a_36755_10509.n2 a_36755_10509.t6 14.282
R9797 a_36755_10509.n2 a_36755_10509.t5 14.282
R9798 a_36755_10509.n1 a_36755_10509.t10 104.259
R9799 a_36755_10391.t0 a_36755_10391.n0 14.282
R9800 a_36755_10391.n0 a_36755_10391.t6 14.282
R9801 a_36755_10391.n0 a_36755_10391.n1 258.161
R9802 a_36755_10391.n1 a_36755_10391.t7 14.283
R9803 a_36755_10391.n1 a_36755_10391.n5 0.852
R9804 a_36755_10391.n5 a_36755_10391.n6 4.366
R9805 a_36755_10391.n6 a_36755_10391.n7 258.161
R9806 a_36755_10391.n7 a_36755_10391.t5 14.282
R9807 a_36755_10391.n7 a_36755_10391.t4 14.282
R9808 a_36755_10391.n6 a_36755_10391.t3 14.283
R9809 a_36755_10391.n5 a_36755_10391.n4 73.514
R9810 a_36755_10391.n4 a_36755_10391.t11 1551.5
R9811 a_36755_10391.t11 a_36755_10391.n3 656.576
R9812 a_36755_10391.n3 a_36755_10391.t2 8.7
R9813 a_36755_10391.n3 a_36755_10391.t1 8.7
R9814 a_36755_10391.n4 a_36755_10391.t8 224.129
R9815 a_36755_10391.t8 a_36755_10391.n2 207.225
R9816 a_36755_10391.n2 a_36755_10391.t10 207.225
R9817 a_36755_10391.n2 a_36755_10391.t9 80.333
R9818 a_20600_4821.n2 a_20600_4821.t5 318.922
R9819 a_20600_4821.n1 a_20600_4821.t6 273.935
R9820 a_20600_4821.n1 a_20600_4821.t7 273.935
R9821 a_20600_4821.n2 a_20600_4821.t4 269.116
R9822 a_20600_4821.n4 a_20600_4821.n0 193.227
R9823 a_20600_4821.t5 a_20600_4821.n1 179.142
R9824 a_20600_4821.n3 a_20600_4821.n2 106.999
R9825 a_20600_4821.t3 a_20600_4821.n4 28.568
R9826 a_20600_4821.n0 a_20600_4821.t2 28.565
R9827 a_20600_4821.n0 a_20600_4821.t1 28.565
R9828 a_20600_4821.n3 a_20600_4821.t0 18.149
R9829 a_20600_4821.n4 a_20600_4821.n3 3.726
R9830 a_21145_3396.t0 a_21145_3396.t1 380.209
R9831 a_8543_1769.n7 a_8543_1769.n6 861.987
R9832 a_8543_1769.n6 a_8543_1769.n5 560.726
R9833 a_8543_1769.t6 a_8543_1769.t16 415.315
R9834 a_8543_1769.t7 a_8543_1769.t17 415.315
R9835 a_8543_1769.n2 a_8543_1769.t13 394.151
R9836 a_8543_1769.n5 a_8543_1769.t9 294.653
R9837 a_8543_1769.n1 a_8543_1769.t15 269.523
R9838 a_8543_1769.t13 a_8543_1769.n1 269.523
R9839 a_8543_1769.n9 a_8543_1769.t6 217.716
R9840 a_8543_1769.n8 a_8543_1769.t19 214.335
R9841 a_8543_1769.t16 a_8543_1769.n8 214.335
R9842 a_8543_1769.n0 a_8543_1769.t8 214.335
R9843 a_8543_1769.t17 a_8543_1769.n0 214.335
R9844 a_8543_1769.n7 a_8543_1769.t7 198.921
R9845 a_8543_1769.n3 a_8543_1769.t4 198.043
R9846 a_8543_1769.n12 a_8543_1769.n11 192.754
R9847 a_8543_1769.n1 a_8543_1769.t5 160.666
R9848 a_8543_1769.n5 a_8543_1769.t18 111.663
R9849 a_8543_1769.n4 a_8543_1769.n2 97.816
R9850 a_8543_1769.n3 a_8543_1769.t14 93.989
R9851 a_8543_1769.n8 a_8543_1769.t11 80.333
R9852 a_8543_1769.n2 a_8543_1769.t10 80.333
R9853 a_8543_1769.n0 a_8543_1769.t12 80.333
R9854 a_8543_1769.n6 a_8543_1769.n4 65.07
R9855 a_8543_1769.n11 a_8543_1769.t2 28.568
R9856 a_8543_1769.n12 a_8543_1769.t1 28.565
R9857 a_8543_1769.t3 a_8543_1769.n12 28.565
R9858 a_8543_1769.n10 a_8543_1769.t0 18.827
R9859 a_8543_1769.n9 a_8543_1769.n7 16.411
R9860 a_8543_1769.n4 a_8543_1769.n3 6.615
R9861 a_8543_1769.n10 a_8543_1769.n9 4.997
R9862 a_8543_1769.n11 a_8543_1769.n10 1.105
R9863 a_12047_4820.n2 a_12047_4820.t4 318.922
R9864 a_12047_4820.n1 a_12047_4820.t5 273.935
R9865 a_12047_4820.n1 a_12047_4820.t6 273.935
R9866 a_12047_4820.n2 a_12047_4820.t7 269.116
R9867 a_12047_4820.n4 a_12047_4820.n0 193.227
R9868 a_12047_4820.t4 a_12047_4820.n1 179.142
R9869 a_12047_4820.n3 a_12047_4820.n2 106.999
R9870 a_12047_4820.t3 a_12047_4820.n4 28.568
R9871 a_12047_4820.n0 a_12047_4820.t2 28.565
R9872 a_12047_4820.n0 a_12047_4820.t1 28.565
R9873 a_12047_4820.n3 a_12047_4820.t0 18.149
R9874 a_12047_4820.n4 a_12047_4820.n3 3.726
R9875 a_20495_18853.t0 a_20495_18853.n0 14.282
R9876 a_20495_18853.n0 a_20495_18853.t1 14.282
R9877 a_20495_18853.n0 a_20495_18853.n9 0.999
R9878 a_20495_18853.n6 a_20495_18853.n8 0.2
R9879 a_20495_18853.n9 a_20495_18853.n6 0.575
R9880 a_20495_18853.n9 a_20495_18853.t2 16.058
R9881 a_20495_18853.n8 a_20495_18853.n7 0.999
R9882 a_20495_18853.n7 a_20495_18853.t3 14.282
R9883 a_20495_18853.n7 a_20495_18853.t5 14.282
R9884 a_20495_18853.n8 a_20495_18853.t4 16.058
R9885 a_20495_18853.n6 a_20495_18853.n4 0.227
R9886 a_20495_18853.n4 a_20495_18853.n5 1.511
R9887 a_20495_18853.n5 a_20495_18853.t6 14.282
R9888 a_20495_18853.n5 a_20495_18853.t7 14.282
R9889 a_20495_18853.n4 a_20495_18853.n1 0.669
R9890 a_20495_18853.n1 a_20495_18853.n2 0.001
R9891 a_20495_18853.n1 a_20495_18853.n3 267.767
R9892 a_20495_18853.n3 a_20495_18853.t9 14.282
R9893 a_20495_18853.n3 a_20495_18853.t11 14.282
R9894 a_20495_18853.n2 a_20495_18853.t10 14.282
R9895 a_20495_18853.n2 a_20495_18853.t8 14.282
R9896 B[1].n4 B[1].n0 592.056
R9897 B[1].t6 B[1].n2 313.069
R9898 B[1].n0 B[1].t7 294.986
R9899 B[1].n1 B[1].t5 271.484
R9900 B[1].n4 B[1].t4 204.672
R9901 B[1].n3 B[1].t6 190.955
R9902 B[1].n3 B[1].t1 190.955
R9903 B[1].n2 B[1].t0 160.666
R9904 B[1].n1 B[1].t3 160.666
R9905 B[1].n0 B[1].t2 110.859
R9906 B[1].n2 B[1].n1 96.129
R9907 B[1].t4 B[1].n3 80.333
R9908 B[1] B[1].n4 55.108
R9909 a_28061_4103.n1 a_28061_4103.t7 318.922
R9910 a_28061_4103.n0 a_28061_4103.t4 274.739
R9911 a_28061_4103.n0 a_28061_4103.t5 274.739
R9912 a_28061_4103.n1 a_28061_4103.t6 269.116
R9913 a_28061_4103.t7 a_28061_4103.n0 179.946
R9914 a_28061_4103.n2 a_28061_4103.n1 105.178
R9915 a_28061_4103.t3 a_28061_4103.n4 29.444
R9916 a_28061_4103.n3 a_28061_4103.t2 28.565
R9917 a_28061_4103.n3 a_28061_4103.t1 28.565
R9918 a_28061_4103.n2 a_28061_4103.t0 18.145
R9919 a_28061_4103.n4 a_28061_4103.n2 2.878
R9920 a_28061_4103.n4 a_28061_4103.n3 0.764
R9921 a_19134_9929.t3 a_19134_9929.n0 14.282
R9922 a_19134_9929.n0 a_19134_9929.t5 14.282
R9923 a_19134_9929.n1 a_19134_9929.n9 0.001
R9924 a_19134_9929.n0 a_19134_9929.n1 267.767
R9925 a_19134_9929.n9 a_19134_9929.t0 14.282
R9926 a_19134_9929.n9 a_19134_9929.t4 14.282
R9927 a_19134_9929.n1 a_19134_9929.n7 0.669
R9928 a_19134_9929.n7 a_19134_9929.n8 1.511
R9929 a_19134_9929.n8 a_19134_9929.t2 14.282
R9930 a_19134_9929.n8 a_19134_9929.t1 14.282
R9931 a_19134_9929.n7 a_19134_9929.n6 0.227
R9932 a_19134_9929.n6 a_19134_9929.n3 0.575
R9933 a_19134_9929.n6 a_19134_9929.n5 0.2
R9934 a_19134_9929.n5 a_19134_9929.t9 16.058
R9935 a_19134_9929.n5 a_19134_9929.n4 0.999
R9936 a_19134_9929.n4 a_19134_9929.t8 14.282
R9937 a_19134_9929.n4 a_19134_9929.t7 14.282
R9938 a_19134_9929.n3 a_19134_9929.n2 0.999
R9939 a_19134_9929.n2 a_19134_9929.t10 14.282
R9940 a_19134_9929.n2 a_19134_9929.t11 14.282
R9941 a_19134_9929.n3 a_19134_9929.t6 16.058
R9942 a_36701_20754.n2 a_36701_20754.t4 448.381
R9943 a_36701_20754.n1 a_36701_20754.t6 287.241
R9944 a_36701_20754.n1 a_36701_20754.t7 287.241
R9945 a_36701_20754.n0 a_36701_20754.t5 247.733
R9946 a_36701_20754.n4 a_36701_20754.n3 182.117
R9947 a_36701_20754.t4 a_36701_20754.n1 160.666
R9948 a_36701_20754.n3 a_36701_20754.t2 28.568
R9949 a_36701_20754.t3 a_36701_20754.n4 28.565
R9950 a_36701_20754.n4 a_36701_20754.t1 28.565
R9951 a_36701_20754.n0 a_36701_20754.t0 18.127
R9952 a_36701_20754.n2 a_36701_20754.n0 4.036
R9953 a_36701_20754.n3 a_36701_20754.n2 0.937
R9954 a_36755_19869.n0 a_36755_19869.t2 14.282
R9955 a_36755_19869.t0 a_36755_19869.n0 14.282
R9956 a_36755_19869.n0 a_36755_19869.n1 258.161
R9957 a_36755_19869.n1 a_36755_19869.t1 14.283
R9958 a_36755_19869.n1 a_36755_19869.n5 0.852
R9959 a_36755_19869.n5 a_36755_19869.n6 4.366
R9960 a_36755_19869.n6 a_36755_19869.n7 258.161
R9961 a_36755_19869.n7 a_36755_19869.t3 14.282
R9962 a_36755_19869.n7 a_36755_19869.t5 14.282
R9963 a_36755_19869.n6 a_36755_19869.t4 14.283
R9964 a_36755_19869.n5 a_36755_19869.n4 73.514
R9965 a_36755_19869.n4 a_36755_19869.t8 1551.5
R9966 a_36755_19869.t8 a_36755_19869.n3 656.576
R9967 a_36755_19869.n3 a_36755_19869.t6 8.7
R9968 a_36755_19869.n3 a_36755_19869.t7 8.7
R9969 a_36755_19869.n4 a_36755_19869.t11 224.129
R9970 a_36755_19869.t11 a_36755_19869.n2 207.225
R9971 a_36755_19869.n2 a_36755_19869.t10 207.225
R9972 a_36755_19869.n2 a_36755_19869.t9 80.333
R9973 a_36755_19987.t6 a_36755_19987.n9 104.259
R9974 a_36755_19987.n3 a_36755_19987.n1 77.784
R9975 a_36755_19987.n5 a_36755_19987.n3 77.456
R9976 a_36755_19987.n7 a_36755_19987.n5 77.456
R9977 a_36755_19987.n9 a_36755_19987.n7 75.815
R9978 a_36755_19987.n9 a_36755_19987.n8 167.433
R9979 a_36755_19987.n8 a_36755_19987.t7 14.282
R9980 a_36755_19987.n8 a_36755_19987.t8 14.282
R9981 a_36755_19987.n7 a_36755_19987.n6 89.977
R9982 a_36755_19987.n6 a_36755_19987.t5 14.282
R9983 a_36755_19987.n6 a_36755_19987.t4 14.282
R9984 a_36755_19987.n5 a_36755_19987.n4 89.977
R9985 a_36755_19987.n4 a_36755_19987.t11 14.282
R9986 a_36755_19987.n4 a_36755_19987.t3 14.282
R9987 a_36755_19987.n3 a_36755_19987.n2 89.977
R9988 a_36755_19987.n2 a_36755_19987.t10 14.282
R9989 a_36755_19987.n2 a_36755_19987.t9 14.282
R9990 a_36755_19987.n1 a_36755_19987.t0 104.259
R9991 a_36755_19987.n1 a_36755_19987.n0 167.433
R9992 a_36755_19987.n0 a_36755_19987.t1 14.282
R9993 a_36755_19987.n0 a_36755_19987.t2 14.282
R9994 a_9206_25153.n2 a_9206_25153.t4 318.922
R9995 a_9206_25153.n1 a_9206_25153.t7 273.935
R9996 a_9206_25153.n1 a_9206_25153.t5 273.935
R9997 a_9206_25153.n2 a_9206_25153.t6 269.116
R9998 a_9206_25153.n4 a_9206_25153.n0 193.227
R9999 a_9206_25153.t4 a_9206_25153.n1 179.142
R10000 a_9206_25153.n3 a_9206_25153.n2 106.999
R10001 a_9206_25153.t3 a_9206_25153.n4 28.568
R10002 a_9206_25153.n0 a_9206_25153.t1 28.565
R10003 a_9206_25153.n0 a_9206_25153.t2 28.565
R10004 a_9206_25153.n3 a_9206_25153.t0 18.149
R10005 a_9206_25153.n4 a_9206_25153.n3 3.726
R10006 a_23973_3835.n4 a_23973_3835.t8 214.335
R10007 a_23973_3835.t7 a_23973_3835.n4 214.335
R10008 a_23973_3835.n5 a_23973_3835.t7 143.851
R10009 a_23973_3835.n5 a_23973_3835.t9 135.658
R10010 a_23973_3835.n4 a_23973_3835.t10 80.333
R10011 a_23973_3835.n0 a_23973_3835.t4 28.565
R10012 a_23973_3835.n0 a_23973_3835.t5 28.565
R10013 a_23973_3835.n2 a_23973_3835.t1 28.565
R10014 a_23973_3835.n2 a_23973_3835.t6 28.565
R10015 a_23973_3835.n7 a_23973_3835.t0 28.565
R10016 a_23973_3835.t2 a_23973_3835.n7 28.565
R10017 a_23973_3835.n1 a_23973_3835.t3 9.714
R10018 a_23973_3835.n1 a_23973_3835.n0 1.003
R10019 a_23973_3835.n6 a_23973_3835.n3 0.833
R10020 a_23973_3835.n3 a_23973_3835.n2 0.653
R10021 a_23973_3835.n7 a_23973_3835.n6 0.653
R10022 a_23973_3835.n3 a_23973_3835.n1 0.341
R10023 a_23973_3835.n6 a_23973_3835.n5 0.032
R10024 a_26163_4103.n1 a_26163_4103.t5 318.922
R10025 a_26163_4103.n0 a_26163_4103.t6 274.739
R10026 a_26163_4103.n0 a_26163_4103.t7 274.739
R10027 a_26163_4103.n1 a_26163_4103.t4 269.116
R10028 a_26163_4103.t5 a_26163_4103.n0 179.946
R10029 a_26163_4103.n2 a_26163_4103.n1 107.263
R10030 a_26163_4103.n3 a_26163_4103.t1 29.444
R10031 a_26163_4103.t3 a_26163_4103.n4 28.565
R10032 a_26163_4103.n4 a_26163_4103.t2 28.565
R10033 a_26163_4103.n2 a_26163_4103.t0 18.145
R10034 a_26163_4103.n3 a_26163_4103.n2 2.878
R10035 a_26163_4103.n4 a_26163_4103.n3 0.764
R10036 a_25869_3397.t0 a_25869_3397.t1 380.209
R10037 a_36755_7247.n0 a_36755_7247.t3 14.282
R10038 a_36755_7247.t0 a_36755_7247.n0 14.282
R10039 a_36755_7247.n0 a_36755_7247.n1 258.161
R10040 a_36755_7247.n1 a_36755_7247.t1 14.283
R10041 a_36755_7247.n1 a_36755_7247.n5 0.852
R10042 a_36755_7247.n5 a_36755_7247.n6 4.366
R10043 a_36755_7247.n6 a_36755_7247.n7 258.161
R10044 a_36755_7247.n7 a_36755_7247.t4 14.282
R10045 a_36755_7247.n7 a_36755_7247.t5 14.282
R10046 a_36755_7247.n6 a_36755_7247.t6 14.283
R10047 a_36755_7247.n5 a_36755_7247.n4 73.514
R10048 a_36755_7247.n4 a_36755_7247.t10 1551.5
R10049 a_36755_7247.t10 a_36755_7247.n3 656.576
R10050 a_36755_7247.n3 a_36755_7247.t7 8.7
R10051 a_36755_7247.n3 a_36755_7247.t2 8.7
R10052 a_36755_7247.n4 a_36755_7247.t9 224.129
R10053 a_36755_7247.t9 a_36755_7247.n2 207.225
R10054 a_36755_7247.n2 a_36755_7247.t8 207.225
R10055 a_36755_7247.n2 a_36755_7247.t11 80.333
R10056 Y[5].n1 Y[5].n0 185.55
R10057 Y[5].n1 Y[5].t2 28.568
R10058 Y[5].n0 Y[5].t3 28.565
R10059 Y[5].n0 Y[5].t1 28.565
R10060 Y[5].n2 Y[5].t0 20.393
R10061 Y[5].n2 Y[5].n1 1.834
R10062 Y[5].n3 Y[5].n2 1.047
R10063 Y[5] Y[5].n3 0.052
R10064 Y[5].n3 Y[5] 0.046
R10065 a_19813_6377.t6 a_19813_6377.t5 800.071
R10066 a_19813_6377.n3 a_19813_6377.n2 672.951
R10067 a_19813_6377.n1 a_19813_6377.t7 285.109
R10068 a_19813_6377.n2 a_19813_6377.t6 193.602
R10069 a_19813_6377.n1 a_19813_6377.t4 160.666
R10070 a_19813_6377.n2 a_19813_6377.n1 91.507
R10071 a_19813_6377.n0 a_19813_6377.t2 28.57
R10072 a_19813_6377.n4 a_19813_6377.t3 28.565
R10073 a_19813_6377.t0 a_19813_6377.n4 28.565
R10074 a_19813_6377.n0 a_19813_6377.t1 17.638
R10075 a_19813_6377.n4 a_19813_6377.n3 0.69
R10076 a_19813_6377.n3 a_19813_6377.n0 0.6
R10077 a_20809_6964.n0 a_20809_6964.t2 14.282
R10078 a_20809_6964.n0 a_20809_6964.t1 14.282
R10079 a_20809_6964.n1 a_20809_6964.t3 14.282
R10080 a_20809_6964.n1 a_20809_6964.t5 14.282
R10081 a_20809_6964.n3 a_20809_6964.t4 14.282
R10082 a_20809_6964.t0 a_20809_6964.n3 14.282
R10083 a_20809_6964.n2 a_20809_6964.n0 2.546
R10084 a_20809_6964.n2 a_20809_6964.n1 2.367
R10085 a_20809_6964.n3 a_20809_6964.n2 0.001
R10086 A[0].n4 A[0].n3 535.449
R10087 A[0].t3 A[0].t2 437.233
R10088 A[0].t13 A[0].t15 437.233
R10089 A[0].t4 A[0].n1 313.873
R10090 A[0].n3 A[0].t11 294.986
R10091 A[0].n0 A[0].t5 272.288
R10092 A[0].n4 A[0].t8 245.184
R10093 A[0].n6 A[0].t13 218.628
R10094 A[0].n8 A[0].t3 217.024
R10095 A[0].n7 A[0].t12 214.686
R10096 A[0].t2 A[0].n7 214.686
R10097 A[0].n5 A[0].t10 214.686
R10098 A[0].t15 A[0].n5 214.686
R10099 A[0].n2 A[0].t4 190.152
R10100 A[0].n2 A[0].t9 190.152
R10101 A[0].n0 A[0].t6 160.666
R10102 A[0].n1 A[0].t7 160.666
R10103 A[0].n3 A[0].t0 110.859
R10104 A[0].n1 A[0].n0 96.129
R10105 A[0].n7 A[0].t1 80.333
R10106 A[0].t8 A[0].n2 80.333
R10107 A[0].n5 A[0].t14 80.333
R10108 A[0].n6 A[0].n4 14.9
R10109 A[0] A[0].n8 7.849
R10110 A[0].n8 A[0].n6 2.599
R10111 a_8147_24434.n1 a_8147_24434.t5 318.922
R10112 a_8147_24434.n0 a_8147_24434.t4 274.739
R10113 a_8147_24434.n0 a_8147_24434.t6 274.739
R10114 a_8147_24434.n1 a_8147_24434.t7 269.116
R10115 a_8147_24434.t5 a_8147_24434.n0 179.946
R10116 a_8147_24434.n2 a_8147_24434.n1 107.263
R10117 a_8147_24434.n3 a_8147_24434.t1 29.444
R10118 a_8147_24434.n4 a_8147_24434.t2 28.565
R10119 a_8147_24434.t3 a_8147_24434.n4 28.565
R10120 a_8147_24434.n2 a_8147_24434.t0 18.145
R10121 a_8147_24434.n3 a_8147_24434.n2 2.878
R10122 a_8147_24434.n4 a_8147_24434.n3 0.764
R10123 a_1817_6836.n5 a_1817_6836.n4 535.449
R10124 a_1817_6836.t18 a_1817_6836.t13 437.233
R10125 a_1817_6836.t14 a_1817_6836.t8 437.233
R10126 a_1817_6836.t17 a_1817_6836.n2 313.873
R10127 a_1817_6836.n4 a_1817_6836.t10 294.986
R10128 a_1817_6836.n1 a_1817_6836.t4 272.288
R10129 a_1817_6836.n5 a_1817_6836.t9 245.184
R10130 a_1817_6836.n7 a_1817_6836.t14 218.628
R10131 a_1817_6836.n9 a_1817_6836.t18 217.026
R10132 a_1817_6836.n8 a_1817_6836.t11 214.686
R10133 a_1817_6836.t13 a_1817_6836.n8 214.686
R10134 a_1817_6836.n6 a_1817_6836.t7 214.686
R10135 a_1817_6836.t8 a_1817_6836.n6 214.686
R10136 a_1817_6836.n11 a_1817_6836.n0 192.754
R10137 a_1817_6836.n3 a_1817_6836.t17 190.152
R10138 a_1817_6836.n3 a_1817_6836.t5 190.152
R10139 a_1817_6836.n1 a_1817_6836.t12 160.666
R10140 a_1817_6836.n2 a_1817_6836.t19 160.666
R10141 a_1817_6836.n4 a_1817_6836.t15 110.859
R10142 a_1817_6836.n2 a_1817_6836.n1 96.129
R10143 a_1817_6836.n8 a_1817_6836.t6 80.333
R10144 a_1817_6836.t9 a_1817_6836.n3 80.333
R10145 a_1817_6836.n6 a_1817_6836.t16 80.333
R10146 a_1817_6836.t3 a_1817_6836.n11 28.568
R10147 a_1817_6836.n0 a_1817_6836.t2 28.565
R10148 a_1817_6836.n0 a_1817_6836.t1 28.565
R10149 a_1817_6836.n10 a_1817_6836.t0 18.722
R10150 a_1817_6836.n7 a_1817_6836.n5 14.9
R10151 a_1817_6836.n9 a_1817_6836.n7 2.603
R10152 a_1817_6836.n10 a_1817_6836.n9 2.382
R10153 a_1817_6836.n11 a_1817_6836.n10 1.281
R10154 B[0].n4 B[0].n0 592.056
R10155 B[0].t0 B[0].n2 313.069
R10156 B[0].n0 B[0].t3 294.986
R10157 B[0].n1 B[0].t2 271.484
R10158 B[0].n4 B[0].t6 204.672
R10159 B[0].n3 B[0].t0 190.955
R10160 B[0].n3 B[0].t5 190.955
R10161 B[0].n2 B[0].t4 160.666
R10162 B[0].n1 B[0].t1 160.666
R10163 B[0].n0 B[0].t7 110.859
R10164 B[0].n2 B[0].n1 96.129
R10165 B[0].t6 B[0].n3 80.333
R10166 B[0] B[0].n4 46.892
R10167 a_n3604_14534.n1 a_n3604_14534.t4 318.119
R10168 a_n3604_14534.n1 a_n3604_14534.t6 269.919
R10169 a_n3604_14534.n0 a_n3604_14534.t5 267.853
R10170 a_n3604_14534.n0 a_n3604_14534.t7 267.853
R10171 a_n3604_14534.t4 a_n3604_14534.n0 160.666
R10172 a_n3604_14534.n2 a_n3604_14534.n1 107.263
R10173 a_n3604_14534.n3 a_n3604_14534.t2 29.444
R10174 a_n3604_14534.t3 a_n3604_14534.n4 28.565
R10175 a_n3604_14534.n4 a_n3604_14534.t1 28.565
R10176 a_n3604_14534.n2 a_n3604_14534.t0 18.145
R10177 a_n3604_14534.n3 a_n3604_14534.n2 2.878
R10178 a_n3604_14534.n4 a_n3604_14534.n3 0.764
R10179 a_14932_26706.t4 a_14932_26706.t7 800.071
R10180 a_14932_26706.n3 a_14932_26706.n2 672.951
R10181 a_14932_26706.n1 a_14932_26706.t6 285.109
R10182 a_14932_26706.n2 a_14932_26706.t4 193.602
R10183 a_14932_26706.n1 a_14932_26706.t5 160.666
R10184 a_14932_26706.n2 a_14932_26706.n1 91.507
R10185 a_14932_26706.n0 a_14932_26706.t3 28.57
R10186 a_14932_26706.t0 a_14932_26706.n4 28.565
R10187 a_14932_26706.n4 a_14932_26706.t1 28.565
R10188 a_14932_26706.n0 a_14932_26706.t2 17.638
R10189 a_14932_26706.n4 a_14932_26706.n3 0.69
R10190 a_14932_26706.n3 a_14932_26706.n0 0.6
R10191 a_17593_4801.t0 a_17593_4801.t1 17.4
R10192 a_22095_18533.n0 a_22095_18533.t7 214.335
R10193 a_22095_18533.t9 a_22095_18533.n0 214.335
R10194 a_22095_18533.n1 a_22095_18533.t9 143.851
R10195 a_22095_18533.n1 a_22095_18533.t10 135.658
R10196 a_22095_18533.n0 a_22095_18533.t8 80.333
R10197 a_22095_18533.n2 a_22095_18533.t4 28.565
R10198 a_22095_18533.n2 a_22095_18533.t5 28.565
R10199 a_22095_18533.n4 a_22095_18533.t6 28.565
R10200 a_22095_18533.n4 a_22095_18533.t0 28.565
R10201 a_22095_18533.n7 a_22095_18533.t1 28.565
R10202 a_22095_18533.t2 a_22095_18533.n7 28.565
R10203 a_22095_18533.n3 a_22095_18533.t3 9.714
R10204 a_22095_18533.n3 a_22095_18533.n2 1.003
R10205 a_22095_18533.n6 a_22095_18533.n5 0.833
R10206 a_22095_18533.n5 a_22095_18533.n4 0.653
R10207 a_22095_18533.n7 a_22095_18533.n6 0.653
R10208 a_22095_18533.n5 a_22095_18533.n3 0.341
R10209 a_22095_18533.n6 a_22095_18533.n1 0.032
R10210 a_20487_21659.t6 a_20487_21659.t7 574.43
R10211 a_20487_21659.n1 a_20487_21659.t4 285.109
R10212 a_20487_21659.n3 a_20487_21659.n2 197.215
R10213 a_20487_21659.n4 a_20487_21659.n0 192.754
R10214 a_20487_21659.n1 a_20487_21659.t5 160.666
R10215 a_20487_21659.n2 a_20487_21659.t6 160.666
R10216 a_20487_21659.n2 a_20487_21659.n1 114.829
R10217 a_20487_21659.t3 a_20487_21659.n4 28.568
R10218 a_20487_21659.n0 a_20487_21659.t1 28.565
R10219 a_20487_21659.n0 a_20487_21659.t2 28.565
R10220 a_20487_21659.n3 a_20487_21659.t0 18.838
R10221 a_20487_21659.n4 a_20487_21659.n3 1.129
R10222 a_13945_4820.n1 a_13945_4820.t7 318.922
R10223 a_13945_4820.n0 a_13945_4820.t4 273.935
R10224 a_13945_4820.n0 a_13945_4820.t5 273.935
R10225 a_13945_4820.n1 a_13945_4820.t6 269.116
R10226 a_13945_4820.n4 a_13945_4820.n3 193.227
R10227 a_13945_4820.t7 a_13945_4820.n0 179.142
R10228 a_13945_4820.n2 a_13945_4820.n1 106.999
R10229 a_13945_4820.n3 a_13945_4820.t2 28.568
R10230 a_13945_4820.n4 a_13945_4820.t1 28.565
R10231 a_13945_4820.t3 a_13945_4820.n4 28.565
R10232 a_13945_4820.n2 a_13945_4820.t0 18.149
R10233 a_13945_4820.n3 a_13945_4820.n2 3.726
R10234 a_18707_10622.n2 a_18707_10622.t6 318.922
R10235 a_18707_10622.n1 a_18707_10622.t4 273.935
R10236 a_18707_10622.n1 a_18707_10622.t7 273.935
R10237 a_18707_10622.n2 a_18707_10622.t5 269.116
R10238 a_18707_10622.n4 a_18707_10622.n0 193.227
R10239 a_18707_10622.t6 a_18707_10622.n1 179.142
R10240 a_18707_10622.n3 a_18707_10622.n2 106.999
R10241 a_18707_10622.t3 a_18707_10622.n4 28.568
R10242 a_18707_10622.n0 a_18707_10622.t1 28.565
R10243 a_18707_10622.n0 a_18707_10622.t2 28.565
R10244 a_18707_10622.n3 a_18707_10622.t0 18.149
R10245 a_18707_10622.n4 a_18707_10622.n3 3.726
R10246 a_19252_9929.t5 a_19252_9929.n0 14.282
R10247 a_19252_9929.n0 a_19252_9929.t7 14.282
R10248 a_19252_9929.n0 a_19252_9929.n12 90.436
R10249 a_19252_9929.n8 a_19252_9929.n11 50.575
R10250 a_19252_9929.n12 a_19252_9929.n8 74.302
R10251 a_19252_9929.n11 a_19252_9929.n10 157.665
R10252 a_19252_9929.n10 a_19252_9929.t4 8.7
R10253 a_19252_9929.n10 a_19252_9929.t0 8.7
R10254 a_19252_9929.n11 a_19252_9929.n9 122.999
R10255 a_19252_9929.n9 a_19252_9929.t3 14.282
R10256 a_19252_9929.n9 a_19252_9929.t2 14.282
R10257 a_19252_9929.n8 a_19252_9929.n7 90.416
R10258 a_19252_9929.n7 a_19252_9929.t1 14.282
R10259 a_19252_9929.n7 a_19252_9929.t6 14.282
R10260 a_19252_9929.n12 a_19252_9929.n1 342.688
R10261 a_19252_9929.n1 a_19252_9929.n6 126.566
R10262 a_19252_9929.n6 a_19252_9929.t11 294.653
R10263 a_19252_9929.n6 a_19252_9929.t12 111.663
R10264 a_19252_9929.n1 a_19252_9929.n5 552.333
R10265 a_19252_9929.n5 a_19252_9929.n4 6.615
R10266 a_19252_9929.n4 a_19252_9929.t14 93.989
R10267 a_19252_9929.n5 a_19252_9929.n3 97.816
R10268 a_19252_9929.n3 a_19252_9929.t15 80.333
R10269 a_19252_9929.n3 a_19252_9929.t8 394.151
R10270 a_19252_9929.t8 a_19252_9929.n2 269.523
R10271 a_19252_9929.n2 a_19252_9929.t9 160.666
R10272 a_19252_9929.n2 a_19252_9929.t10 269.523
R10273 a_19252_9929.n4 a_19252_9929.t13 198.043
R10274 a_36697_5000.n3 a_36697_5000.t7 448.381
R10275 a_36697_5000.n2 a_36697_5000.t4 287.241
R10276 a_36697_5000.n2 a_36697_5000.t6 287.241
R10277 a_36697_5000.n1 a_36697_5000.t5 247.733
R10278 a_36697_5000.n4 a_36697_5000.n0 182.117
R10279 a_36697_5000.t7 a_36697_5000.n2 160.666
R10280 a_36697_5000.t3 a_36697_5000.n4 28.568
R10281 a_36697_5000.n0 a_36697_5000.t1 28.565
R10282 a_36697_5000.n0 a_36697_5000.t2 28.565
R10283 a_36697_5000.n1 a_36697_5000.t0 18.127
R10284 a_36697_5000.n3 a_36697_5000.n1 4.036
R10285 a_36697_5000.n4 a_36697_5000.n3 0.937
R10286 a_23926_11281.n6 a_23926_11281.n5 501.28
R10287 a_23926_11281.t15 a_23926_11281.t9 437.233
R10288 a_23926_11281.t14 a_23926_11281.t10 415.315
R10289 a_23926_11281.t4 a_23926_11281.n3 313.873
R10290 a_23926_11281.n5 a_23926_11281.t7 294.986
R10291 a_23926_11281.n2 a_23926_11281.t16 272.288
R10292 a_23926_11281.n6 a_23926_11281.t5 236.01
R10293 a_23926_11281.n9 a_23926_11281.t15 216.627
R10294 a_23926_11281.n7 a_23926_11281.t14 216.111
R10295 a_23926_11281.n8 a_23926_11281.t11 214.686
R10296 a_23926_11281.t9 a_23926_11281.n8 214.686
R10297 a_23926_11281.n1 a_23926_11281.t12 214.335
R10298 a_23926_11281.t10 a_23926_11281.n1 214.335
R10299 a_23926_11281.n4 a_23926_11281.t4 190.152
R10300 a_23926_11281.n4 a_23926_11281.t6 190.152
R10301 a_23926_11281.n2 a_23926_11281.t18 160.666
R10302 a_23926_11281.n3 a_23926_11281.t19 160.666
R10303 a_23926_11281.n7 a_23926_11281.n6 148.428
R10304 a_23926_11281.n5 a_23926_11281.t13 110.859
R10305 a_23926_11281.n3 a_23926_11281.n2 96.129
R10306 a_23926_11281.n8 a_23926_11281.t8 80.333
R10307 a_23926_11281.n1 a_23926_11281.t17 80.333
R10308 a_23926_11281.t5 a_23926_11281.n4 80.333
R10309 a_23926_11281.t1 a_23926_11281.n11 28.57
R10310 a_23926_11281.n0 a_23926_11281.t3 28.565
R10311 a_23926_11281.n0 a_23926_11281.t2 28.565
R10312 a_23926_11281.n11 a_23926_11281.t0 17.638
R10313 a_23926_11281.n10 a_23926_11281.n9 11.942
R10314 a_23926_11281.n9 a_23926_11281.n7 2.923
R10315 a_23926_11281.n10 a_23926_11281.n0 0.69
R10316 a_23926_11281.n11 a_23926_11281.n10 0.6
R10317 a_28069_9971.n1 a_28069_9971.t4 318.922
R10318 a_28069_9971.n0 a_28069_9971.t5 274.739
R10319 a_28069_9971.n0 a_28069_9971.t6 274.739
R10320 a_28069_9971.n1 a_28069_9971.t7 269.116
R10321 a_28069_9971.t4 a_28069_9971.n0 179.946
R10322 a_28069_9971.n2 a_28069_9971.n1 105.178
R10323 a_28069_9971.n3 a_28069_9971.t1 29.444
R10324 a_28069_9971.n4 a_28069_9971.t2 28.565
R10325 a_28069_9971.t3 a_28069_9971.n4 28.565
R10326 a_28069_9971.n2 a_28069_9971.t0 18.145
R10327 a_28069_9971.n3 a_28069_9971.n2 2.878
R10328 a_28069_9971.n4 a_28069_9971.n3 0.764
R10329 a_27775_9997.n0 a_27775_9997.n8 122.999
R10330 a_27775_9997.t2 a_27775_9997.n0 14.282
R10331 a_27775_9997.n0 a_27775_9997.t7 14.282
R10332 a_27775_9997.n8 a_27775_9997.n6 50.575
R10333 a_27775_9997.n6 a_27775_9997.n4 74.302
R10334 a_27775_9997.n8 a_27775_9997.n7 157.665
R10335 a_27775_9997.n7 a_27775_9997.t1 8.7
R10336 a_27775_9997.n7 a_27775_9997.t0 8.7
R10337 a_27775_9997.n6 a_27775_9997.n5 90.416
R10338 a_27775_9997.n5 a_27775_9997.t3 14.282
R10339 a_27775_9997.n5 a_27775_9997.t6 14.282
R10340 a_27775_9997.n4 a_27775_9997.n3 90.436
R10341 a_27775_9997.n3 a_27775_9997.t5 14.282
R10342 a_27775_9997.n3 a_27775_9997.t4 14.282
R10343 a_27775_9997.n4 a_27775_9997.n1 670.272
R10344 a_27775_9997.n1 a_27775_9997.t11 408.806
R10345 a_27775_9997.t9 a_27775_9997.n2 160.666
R10346 a_27775_9997.n1 a_27775_9997.t9 989.744
R10347 a_27775_9997.n2 a_27775_9997.t8 287.241
R10348 a_27775_9997.n2 a_27775_9997.t10 287.241
R10349 a_36751_4233.t0 a_36751_4233.n9 104.259
R10350 a_36751_4233.n9 a_36751_4233.n2 77.784
R10351 a_36751_4233.n2 a_36751_4233.n4 77.456
R10352 a_36751_4233.n4 a_36751_4233.n6 77.456
R10353 a_36751_4233.n6 a_36751_4233.n7 75.815
R10354 a_36751_4233.n7 a_36751_4233.n8 167.433
R10355 a_36751_4233.n8 a_36751_4233.t10 14.282
R10356 a_36751_4233.n8 a_36751_4233.t9 14.282
R10357 a_36751_4233.n7 a_36751_4233.t11 104.259
R10358 a_36751_4233.n6 a_36751_4233.n5 89.977
R10359 a_36751_4233.n5 a_36751_4233.t4 14.282
R10360 a_36751_4233.n5 a_36751_4233.t5 14.282
R10361 a_36751_4233.n4 a_36751_4233.n3 89.977
R10362 a_36751_4233.n3 a_36751_4233.t7 14.282
R10363 a_36751_4233.n3 a_36751_4233.t3 14.282
R10364 a_36751_4233.n2 a_36751_4233.n1 89.977
R10365 a_36751_4233.n1 a_36751_4233.t6 14.282
R10366 a_36751_4233.n1 a_36751_4233.t8 14.282
R10367 a_36751_4233.n9 a_36751_4233.n0 167.433
R10368 a_36751_4233.n0 a_36751_4233.t2 14.282
R10369 a_36751_4233.n0 a_36751_4233.t1 14.282
R10370 a_32011_9700.t1 a_32011_9700.n0 14.282
R10371 a_32011_9700.n0 a_32011_9700.t2 14.282
R10372 a_32011_9700.n0 a_32011_9700.n8 122.999
R10373 a_32011_9700.n8 a_32011_9700.n6 50.575
R10374 a_32011_9700.n6 a_32011_9700.n4 74.302
R10375 a_32011_9700.n8 a_32011_9700.n7 157.665
R10376 a_32011_9700.n7 a_32011_9700.t0 8.7
R10377 a_32011_9700.n7 a_32011_9700.t7 8.7
R10378 a_32011_9700.n6 a_32011_9700.n5 90.416
R10379 a_32011_9700.n5 a_32011_9700.t3 14.282
R10380 a_32011_9700.n5 a_32011_9700.t4 14.282
R10381 a_32011_9700.n4 a_32011_9700.n3 90.436
R10382 a_32011_9700.n3 a_32011_9700.t6 14.282
R10383 a_32011_9700.n3 a_32011_9700.t5 14.282
R10384 a_32011_9700.n4 a_32011_9700.n1 653.122
R10385 a_32011_9700.n1 a_32011_9700.t10 408.806
R10386 a_32011_9700.t9 a_32011_9700.n2 160.666
R10387 a_32011_9700.n1 a_32011_9700.t9 989.744
R10388 a_32011_9700.n2 a_32011_9700.t8 287.241
R10389 a_32011_9700.n2 a_32011_9700.t11 287.241
R10390 a_21136_23720.t0 a_21136_23720.t1 17.4
R10391 a_22344_27288.t7 a_22344_27288.n2 404.877
R10392 a_22344_27288.n1 a_22344_27288.t8 210.902
R10393 a_22344_27288.n3 a_22344_27288.t7 136.943
R10394 a_22344_27288.n2 a_22344_27288.n1 107.801
R10395 a_22344_27288.n1 a_22344_27288.t5 80.333
R10396 a_22344_27288.n2 a_22344_27288.t6 80.333
R10397 a_22344_27288.n0 a_22344_27288.t4 17.4
R10398 a_22344_27288.n0 a_22344_27288.t0 17.4
R10399 a_22344_27288.n4 a_22344_27288.t3 15.032
R10400 a_22344_27288.t1 a_22344_27288.n5 14.282
R10401 a_22344_27288.n5 a_22344_27288.t2 14.282
R10402 a_22344_27288.n5 a_22344_27288.n4 1.65
R10403 a_22344_27288.n3 a_22344_27288.n0 0.672
R10404 a_22344_27288.n4 a_22344_27288.n3 0.665
R10405 a_22608_26705.n6 a_22608_26705.n5 501.28
R10406 a_22608_26705.t8 a_22608_26705.t9 437.233
R10407 a_22608_26705.t16 a_22608_26705.t17 415.315
R10408 a_22608_26705.t10 a_22608_26705.n3 313.873
R10409 a_22608_26705.n5 a_22608_26705.t19 294.986
R10410 a_22608_26705.n2 a_22608_26705.t12 272.288
R10411 a_22608_26705.n6 a_22608_26705.t4 236.01
R10412 a_22608_26705.n9 a_22608_26705.t8 216.627
R10413 a_22608_26705.n7 a_22608_26705.t16 216.111
R10414 a_22608_26705.n8 a_22608_26705.t6 214.686
R10415 a_22608_26705.t9 a_22608_26705.n8 214.686
R10416 a_22608_26705.n1 a_22608_26705.t15 214.335
R10417 a_22608_26705.t17 a_22608_26705.n1 214.335
R10418 a_22608_26705.n4 a_22608_26705.t10 190.152
R10419 a_22608_26705.n4 a_22608_26705.t5 190.152
R10420 a_22608_26705.n2 a_22608_26705.t13 160.666
R10421 a_22608_26705.n3 a_22608_26705.t14 160.666
R10422 a_22608_26705.n7 a_22608_26705.n6 148.428
R10423 a_22608_26705.n5 a_22608_26705.t11 110.859
R10424 a_22608_26705.n3 a_22608_26705.n2 96.129
R10425 a_22608_26705.n8 a_22608_26705.t7 80.333
R10426 a_22608_26705.n1 a_22608_26705.t18 80.333
R10427 a_22608_26705.t4 a_22608_26705.n4 80.333
R10428 a_22608_26705.n0 a_22608_26705.t2 28.57
R10429 a_22608_26705.n11 a_22608_26705.t1 28.565
R10430 a_22608_26705.t3 a_22608_26705.n11 28.565
R10431 a_22608_26705.n0 a_22608_26705.t0 17.638
R10432 a_22608_26705.n10 a_22608_26705.n9 5.767
R10433 a_22608_26705.n9 a_22608_26705.n7 2.923
R10434 a_22608_26705.n11 a_22608_26705.n10 0.69
R10435 a_22608_26705.n10 a_22608_26705.n0 0.6
R10436 a_19546_9903.n1 a_19546_9903.t5 318.922
R10437 a_19546_9903.n0 a_19546_9903.t6 274.739
R10438 a_19546_9903.n0 a_19546_9903.t7 274.739
R10439 a_19546_9903.n1 a_19546_9903.t4 269.116
R10440 a_19546_9903.t5 a_19546_9903.n0 179.946
R10441 a_19546_9903.n2 a_19546_9903.n1 107.263
R10442 a_19546_9903.n3 a_19546_9903.t2 29.444
R10443 a_19546_9903.n4 a_19546_9903.t1 28.565
R10444 a_19546_9903.t0 a_19546_9903.n4 28.565
R10445 a_19546_9903.n2 a_19546_9903.t3 18.145
R10446 a_19546_9903.n3 a_19546_9903.n2 2.878
R10447 a_19546_9903.n4 a_19546_9903.n3 0.764
R10448 a_19252_9197.t0 a_19252_9197.t1 380.209
R10449 a_5948_27420.n2 a_5948_27420.t10 214.335
R10450 a_5948_27420.t8 a_5948_27420.n2 214.335
R10451 a_5948_27420.n3 a_5948_27420.t8 143.851
R10452 a_5948_27420.n3 a_5948_27420.t7 135.658
R10453 a_5948_27420.n2 a_5948_27420.t9 80.333
R10454 a_5948_27420.n4 a_5948_27420.t0 28.565
R10455 a_5948_27420.n4 a_5948_27420.t1 28.565
R10456 a_5948_27420.n0 a_5948_27420.t6 28.565
R10457 a_5948_27420.n0 a_5948_27420.t4 28.565
R10458 a_5948_27420.t2 a_5948_27420.n7 28.565
R10459 a_5948_27420.n7 a_5948_27420.t5 28.565
R10460 a_5948_27420.n1 a_5948_27420.t3 9.714
R10461 a_5948_27420.n1 a_5948_27420.n0 1.003
R10462 a_5948_27420.n6 a_5948_27420.n5 0.833
R10463 a_5948_27420.n5 a_5948_27420.n4 0.653
R10464 a_5948_27420.n7 a_5948_27420.n6 0.653
R10465 a_5948_27420.n6 a_5948_27420.n1 0.341
R10466 a_5948_27420.n5 a_5948_27420.n3 0.032
R10467 a_12892_9971.n1 a_12892_9971.t7 318.922
R10468 a_12892_9971.n0 a_12892_9971.t4 274.739
R10469 a_12892_9971.n0 a_12892_9971.t5 274.739
R10470 a_12892_9971.n1 a_12892_9971.t6 269.116
R10471 a_12892_9971.t7 a_12892_9971.n0 179.946
R10472 a_12892_9971.n2 a_12892_9971.n1 107.263
R10473 a_12892_9971.n3 a_12892_9971.t1 29.444
R10474 a_12892_9971.n4 a_12892_9971.t2 28.565
R10475 a_12892_9971.t3 a_12892_9971.n4 28.565
R10476 a_12892_9971.n2 a_12892_9971.t0 18.145
R10477 a_12892_9971.n3 a_12892_9971.n2 2.878
R10478 a_12892_9971.n4 a_12892_9971.n3 0.764
R10479 a_32305_6179.n1 a_32305_6179.t5 318.922
R10480 a_32305_6179.n0 a_32305_6179.t6 274.739
R10481 a_32305_6179.n0 a_32305_6179.t7 274.739
R10482 a_32305_6179.n1 a_32305_6179.t4 269.116
R10483 a_32305_6179.t5 a_32305_6179.n0 179.946
R10484 a_32305_6179.n2 a_32305_6179.n1 107.263
R10485 a_32305_6179.n3 a_32305_6179.t2 29.444
R10486 a_32305_6179.t3 a_32305_6179.n4 28.565
R10487 a_32305_6179.n4 a_32305_6179.t1 28.565
R10488 a_32305_6179.n2 a_32305_6179.t0 18.145
R10489 a_32305_6179.n3 a_32305_6179.n2 2.878
R10490 a_32305_6179.n4 a_32305_6179.n3 0.764
R10491 a_32011_5473.t0 a_32011_5473.t1 380.209
R10492 a_14378_9997.n0 a_14378_9997.n9 1.511
R10493 a_14378_9997.n0 a_14378_9997.t11 14.282
R10494 a_14378_9997.t0 a_14378_9997.n0 14.282
R10495 a_14378_9997.n9 a_14378_9997.n5 0.227
R10496 a_14378_9997.n9 a_14378_9997.n6 0.669
R10497 a_14378_9997.n6 a_14378_9997.n7 0.001
R10498 a_14378_9997.n6 a_14378_9997.n8 267.767
R10499 a_14378_9997.n8 a_14378_9997.t3 14.282
R10500 a_14378_9997.n8 a_14378_9997.t4 14.282
R10501 a_14378_9997.n7 a_14378_9997.t10 14.282
R10502 a_14378_9997.n7 a_14378_9997.t5 14.282
R10503 a_14378_9997.n5 a_14378_9997.n2 0.575
R10504 a_14378_9997.n5 a_14378_9997.n4 0.2
R10505 a_14378_9997.n4 a_14378_9997.t2 16.058
R10506 a_14378_9997.n4 a_14378_9997.n3 0.999
R10507 a_14378_9997.n3 a_14378_9997.t6 14.282
R10508 a_14378_9997.n3 a_14378_9997.t1 14.282
R10509 a_14378_9997.n2 a_14378_9997.n1 0.999
R10510 a_14378_9997.n1 a_14378_9997.t8 14.282
R10511 a_14378_9997.n1 a_14378_9997.t9 14.282
R10512 a_14378_9997.n2 a_14378_9997.t7 16.058
R10513 a_25567_25766.n2 a_25567_25766.t9 214.335
R10514 a_25567_25766.t7 a_25567_25766.n2 214.335
R10515 a_25567_25766.n3 a_25567_25766.t7 143.851
R10516 a_25567_25766.n3 a_25567_25766.t10 135.658
R10517 a_25567_25766.n2 a_25567_25766.t8 80.333
R10518 a_25567_25766.n4 a_25567_25766.t1 28.565
R10519 a_25567_25766.n4 a_25567_25766.t0 28.565
R10520 a_25567_25766.n0 a_25567_25766.t5 28.565
R10521 a_25567_25766.n0 a_25567_25766.t6 28.565
R10522 a_25567_25766.t2 a_25567_25766.n7 28.565
R10523 a_25567_25766.n7 a_25567_25766.t4 28.565
R10524 a_25567_25766.n1 a_25567_25766.t3 9.714
R10525 a_25567_25766.n1 a_25567_25766.n0 1.003
R10526 a_25567_25766.n6 a_25567_25766.n5 0.833
R10527 a_25567_25766.n5 a_25567_25766.n4 0.653
R10528 a_25567_25766.n7 a_25567_25766.n6 0.653
R10529 a_25567_25766.n6 a_25567_25766.n1 0.341
R10530 a_25567_25766.n5 a_25567_25766.n3 0.032
R10531 a_19241_23521.t0 a_19241_23521.t1 17.4
R10532 B[7].n4 B[7].n0 592.056
R10533 B[7].t4 B[7].n2 313.069
R10534 B[7].n0 B[7].t1 294.986
R10535 B[7].n1 B[7].t2 271.484
R10536 B[7].n4 B[7].t3 204.672
R10537 B[7].n3 B[7].t4 190.955
R10538 B[7].n3 B[7].t0 190.955
R10539 B[7].n2 B[7].t6 160.666
R10540 B[7].n1 B[7].t7 160.666
R10541 B[7].n0 B[7].t5 110.859
R10542 B[7].n2 B[7].n1 96.129
R10543 B[7] B[7].n4 84.444
R10544 B[7].t3 B[7].n3 80.333
R10545 a_36755_7365.t0 a_36755_7365.n0 14.282
R10546 a_36755_7365.n0 a_36755_7365.t1 14.282
R10547 a_36755_7365.n4 a_36755_7365.n2 77.784
R10548 a_36755_7365.n6 a_36755_7365.n4 77.456
R10549 a_36755_7365.n8 a_36755_7365.n6 77.456
R10550 a_36755_7365.n9 a_36755_7365.n8 75.815
R10551 a_36755_7365.n0 a_36755_7365.n9 167.433
R10552 a_36755_7365.n9 a_36755_7365.t2 104.259
R10553 a_36755_7365.n8 a_36755_7365.n7 89.977
R10554 a_36755_7365.n7 a_36755_7365.t10 14.282
R10555 a_36755_7365.n7 a_36755_7365.t11 14.282
R10556 a_36755_7365.n6 a_36755_7365.n5 89.977
R10557 a_36755_7365.n5 a_36755_7365.t5 14.282
R10558 a_36755_7365.n5 a_36755_7365.t9 14.282
R10559 a_36755_7365.n4 a_36755_7365.n3 89.977
R10560 a_36755_7365.n3 a_36755_7365.t7 14.282
R10561 a_36755_7365.n3 a_36755_7365.t6 14.282
R10562 a_36755_7365.n2 a_36755_7365.t3 104.259
R10563 a_36755_7365.n2 a_36755_7365.n1 167.433
R10564 a_36755_7365.n1 a_36755_7365.t4 14.282
R10565 a_36755_7365.n1 a_36755_7365.t8 14.282
R10566 a_26152_23725.t6 a_26152_23725.t5 574.43
R10567 a_26152_23725.n0 a_26152_23725.t4 285.109
R10568 a_26152_23725.n2 a_26152_23725.n1 197.217
R10569 a_26152_23725.n4 a_26152_23725.n3 192.754
R10570 a_26152_23725.n0 a_26152_23725.t7 160.666
R10571 a_26152_23725.n1 a_26152_23725.t6 160.666
R10572 a_26152_23725.n1 a_26152_23725.n0 114.829
R10573 a_26152_23725.n3 a_26152_23725.t3 28.568
R10574 a_26152_23725.n4 a_26152_23725.t2 28.565
R10575 a_26152_23725.t0 a_26152_23725.n4 28.565
R10576 a_26152_23725.n2 a_26152_23725.t1 18.838
R10577 a_26152_23725.n3 a_26152_23725.n2 1.129
R10578 a_27760_27288.t5 a_27760_27288.n2 404.877
R10579 a_27760_27288.n1 a_27760_27288.t8 210.902
R10580 a_27760_27288.n3 a_27760_27288.t5 136.943
R10581 a_27760_27288.n2 a_27760_27288.n1 107.801
R10582 a_27760_27288.n1 a_27760_27288.t7 80.333
R10583 a_27760_27288.n2 a_27760_27288.t6 80.333
R10584 a_27760_27288.n0 a_27760_27288.t0 17.4
R10585 a_27760_27288.n0 a_27760_27288.t1 17.4
R10586 a_27760_27288.n4 a_27760_27288.t3 15.032
R10587 a_27760_27288.n5 a_27760_27288.t4 14.282
R10588 a_27760_27288.t2 a_27760_27288.n5 14.282
R10589 a_27760_27288.n5 a_27760_27288.n4 1.65
R10590 a_27760_27288.n3 a_27760_27288.n0 0.672
R10591 a_27760_27288.n4 a_27760_27288.n3 0.665
R10592 a_27878_27288.n0 a_27878_27288.t3 14.282
R10593 a_27878_27288.n0 a_27878_27288.t4 14.282
R10594 a_27878_27288.n1 a_27878_27288.t2 14.282
R10595 a_27878_27288.n1 a_27878_27288.t1 14.282
R10596 a_27878_27288.t0 a_27878_27288.n3 14.282
R10597 a_27878_27288.n3 a_27878_27288.t5 14.282
R10598 a_27878_27288.n2 a_27878_27288.n0 2.546
R10599 a_27878_27288.n2 a_27878_27288.n1 2.367
R10600 a_27878_27288.n3 a_27878_27288.n2 0.001
R10601 a_n2381_13360.t0 a_n2381_13360.t1 17.4
R10602 a_6335_4103.n1 a_6335_4103.t5 318.922
R10603 a_6335_4103.n0 a_6335_4103.t6 274.739
R10604 a_6335_4103.n0 a_6335_4103.t7 274.739
R10605 a_6335_4103.n1 a_6335_4103.t4 269.116
R10606 a_6335_4103.t5 a_6335_4103.n0 179.946
R10607 a_6335_4103.n2 a_6335_4103.n1 107.263
R10608 a_6335_4103.t3 a_6335_4103.n4 29.444
R10609 a_6335_4103.n3 a_6335_4103.t2 28.565
R10610 a_6335_4103.n3 a_6335_4103.t1 28.565
R10611 a_6335_4103.n2 a_6335_4103.t0 18.145
R10612 a_6335_4103.n4 a_6335_4103.n2 2.878
R10613 a_6335_4103.n4 a_6335_4103.n3 0.764
R10614 a_6041_3397.t0 a_6041_3397.t1 380.209
R10615 a_36755_23131.t0 a_36755_23131.n0 14.282
R10616 a_36755_23131.n0 a_36755_23131.t7 14.282
R10617 a_36755_23131.n4 a_36755_23131.n2 77.784
R10618 a_36755_23131.n6 a_36755_23131.n4 77.456
R10619 a_36755_23131.n8 a_36755_23131.n6 77.456
R10620 a_36755_23131.n9 a_36755_23131.n8 75.815
R10621 a_36755_23131.n0 a_36755_23131.n9 167.433
R10622 a_36755_23131.n9 a_36755_23131.t8 104.259
R10623 a_36755_23131.n8 a_36755_23131.n7 89.977
R10624 a_36755_23131.n7 a_36755_23131.t5 14.282
R10625 a_36755_23131.n7 a_36755_23131.t6 14.282
R10626 a_36755_23131.n6 a_36755_23131.n5 89.977
R10627 a_36755_23131.n5 a_36755_23131.t11 14.282
R10628 a_36755_23131.n5 a_36755_23131.t4 14.282
R10629 a_36755_23131.n4 a_36755_23131.n3 89.977
R10630 a_36755_23131.n3 a_36755_23131.t10 14.282
R10631 a_36755_23131.n3 a_36755_23131.t9 14.282
R10632 a_36755_23131.n2 a_36755_23131.t1 104.259
R10633 a_36755_23131.n2 a_36755_23131.n1 167.433
R10634 a_36755_23131.n1 a_36755_23131.t3 14.282
R10635 a_36755_23131.n1 a_36755_23131.t2 14.282
R10636 a_14306_12250.n5 a_14306_12250.n4 535.449
R10637 a_14306_12250.t4 a_14306_12250.t14 437.233
R10638 a_14306_12250.t16 a_14306_12250.t11 437.233
R10639 a_14306_12250.t10 a_14306_12250.n2 313.873
R10640 a_14306_12250.n4 a_14306_12250.t18 294.986
R10641 a_14306_12250.n1 a_14306_12250.t6 272.288
R10642 a_14306_12250.n5 a_14306_12250.t15 245.184
R10643 a_14306_12250.n7 a_14306_12250.t16 218.628
R10644 a_14306_12250.n9 a_14306_12250.t4 217.024
R10645 a_14306_12250.n8 a_14306_12250.t19 214.686
R10646 a_14306_12250.t14 a_14306_12250.n8 214.686
R10647 a_14306_12250.n6 a_14306_12250.t13 214.686
R10648 a_14306_12250.t11 a_14306_12250.n6 214.686
R10649 a_14306_12250.n3 a_14306_12250.t10 190.152
R10650 a_14306_12250.n3 a_14306_12250.t5 190.152
R10651 a_14306_12250.n1 a_14306_12250.t12 160.666
R10652 a_14306_12250.n2 a_14306_12250.t9 160.666
R10653 a_14306_12250.n4 a_14306_12250.t7 110.859
R10654 a_14306_12250.n2 a_14306_12250.n1 96.129
R10655 a_14306_12250.n8 a_14306_12250.t8 80.333
R10656 a_14306_12250.t15 a_14306_12250.n3 80.333
R10657 a_14306_12250.n6 a_14306_12250.t17 80.333
R10658 a_14306_12250.n0 a_14306_12250.t1 28.57
R10659 a_14306_12250.n11 a_14306_12250.t3 28.565
R10660 a_14306_12250.t0 a_14306_12250.n11 28.565
R10661 a_14306_12250.n0 a_14306_12250.t2 17.638
R10662 a_14306_12250.n7 a_14306_12250.n5 14.9
R10663 a_14306_12250.n10 a_14306_12250.n9 8.819
R10664 a_14306_12250.n9 a_14306_12250.n7 2.599
R10665 a_14306_12250.n11 a_14306_12250.n10 0.69
R10666 a_14306_12250.n10 a_14306_12250.n0 0.6
R10667 a_17342_7088.n4 a_17342_7088.t8 214.335
R10668 a_17342_7088.t7 a_17342_7088.n4 214.335
R10669 a_17342_7088.n5 a_17342_7088.t7 143.851
R10670 a_17342_7088.n5 a_17342_7088.t9 135.658
R10671 a_17342_7088.n4 a_17342_7088.t10 80.333
R10672 a_17342_7088.n0 a_17342_7088.t6 28.565
R10673 a_17342_7088.n0 a_17342_7088.t4 28.565
R10674 a_17342_7088.n2 a_17342_7088.t1 28.565
R10675 a_17342_7088.n2 a_17342_7088.t5 28.565
R10676 a_17342_7088.n7 a_17342_7088.t0 28.565
R10677 a_17342_7088.t2 a_17342_7088.n7 28.565
R10678 a_17342_7088.n1 a_17342_7088.t3 9.714
R10679 a_17342_7088.n1 a_17342_7088.n0 1.003
R10680 a_17342_7088.n6 a_17342_7088.n3 0.833
R10681 a_17342_7088.n3 a_17342_7088.n2 0.653
R10682 a_17342_7088.n7 a_17342_7088.n6 0.653
R10683 a_17342_7088.n3 a_17342_7088.n1 0.341
R10684 a_17342_7088.n6 a_17342_7088.n5 0.032
R10685 a_17579_6451.t0 a_17579_6451.t1 17.4
R10686 a_36697_17622.n2 a_36697_17622.t4 448.381
R10687 a_36697_17622.n1 a_36697_17622.t5 287.241
R10688 a_36697_17622.n1 a_36697_17622.t7 287.241
R10689 a_36697_17622.n0 a_36697_17622.t6 247.733
R10690 a_36697_17622.n4 a_36697_17622.n3 182.117
R10691 a_36697_17622.t4 a_36697_17622.n1 160.666
R10692 a_36697_17622.n3 a_36697_17622.t1 28.568
R10693 a_36697_17622.n4 a_36697_17622.t2 28.565
R10694 a_36697_17622.t3 a_36697_17622.n4 28.565
R10695 a_36697_17622.n0 a_36697_17622.t0 18.127
R10696 a_36697_17622.n2 a_36697_17622.n0 4.036
R10697 a_36697_17622.n3 a_36697_17622.n2 0.937
R10698 a_36701_8132.n3 a_36701_8132.t5 448.381
R10699 a_36701_8132.n2 a_36701_8132.t6 287.241
R10700 a_36701_8132.n2 a_36701_8132.t4 287.241
R10701 a_36701_8132.n1 a_36701_8132.t7 247.733
R10702 a_36701_8132.n4 a_36701_8132.n0 182.117
R10703 a_36701_8132.t5 a_36701_8132.n2 160.666
R10704 a_36701_8132.t3 a_36701_8132.n4 28.568
R10705 a_36701_8132.n0 a_36701_8132.t1 28.565
R10706 a_36701_8132.n0 a_36701_8132.t2 28.565
R10707 a_36701_8132.n1 a_36701_8132.t0 18.127
R10708 a_36701_8132.n3 a_36701_8132.n1 4.036
R10709 a_36701_8132.n4 a_36701_8132.n3 0.937
R10710 a_12894_6959.t8 a_12894_6959.n3 404.877
R10711 a_12894_6959.n2 a_12894_6959.t7 210.902
R10712 a_12894_6959.n4 a_12894_6959.t8 136.943
R10713 a_12894_6959.n3 a_12894_6959.n2 107.801
R10714 a_12894_6959.n2 a_12894_6959.t6 80.333
R10715 a_12894_6959.n3 a_12894_6959.t5 80.333
R10716 a_12894_6959.n1 a_12894_6959.t4 17.4
R10717 a_12894_6959.n1 a_12894_6959.t2 17.4
R10718 a_12894_6959.t0 a_12894_6959.n5 15.032
R10719 a_12894_6959.n0 a_12894_6959.t3 14.282
R10720 a_12894_6959.n0 a_12894_6959.t1 14.282
R10721 a_12894_6959.n5 a_12894_6959.n0 1.65
R10722 a_12894_6959.n4 a_12894_6959.n1 0.672
R10723 a_12894_6959.n5 a_12894_6959.n4 0.665
R10724 a_13158_6376.t5 a_13158_6376.t6 800.071
R10725 a_13158_6376.n3 a_13158_6376.n2 672.951
R10726 a_13158_6376.n1 a_13158_6376.t7 285.109
R10727 a_13158_6376.n2 a_13158_6376.t5 193.602
R10728 a_13158_6376.n1 a_13158_6376.t4 160.666
R10729 a_13158_6376.n2 a_13158_6376.n1 91.507
R10730 a_13158_6376.t3 a_13158_6376.n4 28.57
R10731 a_13158_6376.n0 a_13158_6376.t1 28.565
R10732 a_13158_6376.n0 a_13158_6376.t2 28.565
R10733 a_13158_6376.n4 a_13158_6376.t0 17.638
R10734 a_13158_6376.n3 a_13158_6376.n0 0.69
R10735 a_13158_6376.n4 a_13158_6376.n3 0.6
R10736 a_19549_6960.t6 a_19549_6960.n2 404.877
R10737 a_19549_6960.n1 a_19549_6960.t8 210.902
R10738 a_19549_6960.n3 a_19549_6960.t6 136.943
R10739 a_19549_6960.n2 a_19549_6960.n1 107.801
R10740 a_19549_6960.n1 a_19549_6960.t5 80.333
R10741 a_19549_6960.n2 a_19549_6960.t7 80.333
R10742 a_19549_6960.n0 a_19549_6960.t0 17.4
R10743 a_19549_6960.n0 a_19549_6960.t1 17.4
R10744 a_19549_6960.n4 a_19549_6960.t4 15.032
R10745 a_19549_6960.n5 a_19549_6960.t3 14.282
R10746 a_19549_6960.t2 a_19549_6960.n5 14.282
R10747 a_19549_6960.n5 a_19549_6960.n4 1.65
R10748 a_19549_6960.n3 a_19549_6960.n0 0.672
R10749 a_19549_6960.n4 a_19549_6960.n3 0.665
R10750 a_19667_6960.n0 a_19667_6960.t3 14.282
R10751 a_19667_6960.n0 a_19667_6960.t5 14.282
R10752 a_19667_6960.n1 a_19667_6960.t1 14.282
R10753 a_19667_6960.n1 a_19667_6960.t2 14.282
R10754 a_19667_6960.t0 a_19667_6960.n3 14.282
R10755 a_19667_6960.n3 a_19667_6960.t4 14.282
R10756 a_19667_6960.n2 a_19667_6960.n0 2.546
R10757 a_19667_6960.n2 a_19667_6960.n1 2.367
R10758 a_19667_6960.n3 a_19667_6960.n2 0.001
R10759 a_27752_24430.n1 a_27752_24430.t7 318.922
R10760 a_27752_24430.n0 a_27752_24430.t6 274.739
R10761 a_27752_24430.n0 a_27752_24430.t4 274.739
R10762 a_27752_24430.n1 a_27752_24430.t5 269.116
R10763 a_27752_24430.t7 a_27752_24430.n0 179.946
R10764 a_27752_24430.n2 a_27752_24430.n1 107.263
R10765 a_27752_24430.t3 a_27752_24430.n4 29.444
R10766 a_27752_24430.n3 a_27752_24430.t1 28.565
R10767 a_27752_24430.n3 a_27752_24430.t2 28.565
R10768 a_27752_24430.n2 a_27752_24430.t0 18.145
R10769 a_27752_24430.n4 a_27752_24430.n2 2.878
R10770 a_27752_24430.n4 a_27752_24430.n3 0.764
R10771 a_36701_23898.n3 a_36701_23898.t6 448.381
R10772 a_36701_23898.n2 a_36701_23898.t7 287.241
R10773 a_36701_23898.n2 a_36701_23898.t4 287.241
R10774 a_36701_23898.n1 a_36701_23898.t5 247.733
R10775 a_36701_23898.n4 a_36701_23898.n0 182.117
R10776 a_36701_23898.t6 a_36701_23898.n2 160.666
R10777 a_36701_23898.t3 a_36701_23898.n4 28.568
R10778 a_36701_23898.n0 a_36701_23898.t1 28.565
R10779 a_36701_23898.n0 a_36701_23898.t2 28.565
R10780 a_36701_23898.n1 a_36701_23898.t0 18.127
R10781 a_36701_23898.n3 a_36701_23898.n1 4.036
R10782 a_36701_23898.n4 a_36701_23898.n3 0.937
R10783 a_32305_1831.n1 a_32305_1831.t7 318.922
R10784 a_32305_1831.n0 a_32305_1831.t4 274.739
R10785 a_32305_1831.n0 a_32305_1831.t6 274.739
R10786 a_32305_1831.n1 a_32305_1831.t5 269.116
R10787 a_32305_1831.t7 a_32305_1831.n0 179.946
R10788 a_32305_1831.n2 a_32305_1831.n1 107.263
R10789 a_32305_1831.n3 a_32305_1831.t1 29.444
R10790 a_32305_1831.n4 a_32305_1831.t2 28.565
R10791 a_32305_1831.t3 a_32305_1831.n4 28.565
R10792 a_32305_1831.n2 a_32305_1831.t0 18.145
R10793 a_32305_1831.n3 a_32305_1831.n2 2.878
R10794 a_32305_1831.n4 a_32305_1831.n3 0.764
R10795 a_26646_21662.t7 a_26646_21662.t4 800.071
R10796 a_26646_21662.n3 a_26646_21662.n2 659.095
R10797 a_26646_21662.n1 a_26646_21662.t5 285.109
R10798 a_26646_21662.n2 a_26646_21662.t7 193.602
R10799 a_26646_21662.n4 a_26646_21662.n0 192.754
R10800 a_26646_21662.n1 a_26646_21662.t6 160.666
R10801 a_26646_21662.n2 a_26646_21662.n1 91.507
R10802 a_26646_21662.t3 a_26646_21662.n4 28.568
R10803 a_26646_21662.n0 a_26646_21662.t1 28.565
R10804 a_26646_21662.n0 a_26646_21662.t2 28.565
R10805 a_26646_21662.n3 a_26646_21662.t0 19.063
R10806 a_26646_21662.n4 a_26646_21662.n3 1.005
R10807 a_4090_5413.n6 a_4090_5413.n5 501.28
R10808 a_4090_5413.t16 a_4090_5413.t11 437.233
R10809 a_4090_5413.t7 a_4090_5413.t13 415.315
R10810 a_4090_5413.t6 a_4090_5413.n3 313.873
R10811 a_4090_5413.n5 a_4090_5413.t19 294.986
R10812 a_4090_5413.n2 a_4090_5413.t12 272.288
R10813 a_4090_5413.n6 a_4090_5413.t18 236.01
R10814 a_4090_5413.n9 a_4090_5413.t16 216.627
R10815 a_4090_5413.n7 a_4090_5413.t7 216.111
R10816 a_4090_5413.n8 a_4090_5413.t14 214.686
R10817 a_4090_5413.t11 a_4090_5413.n8 214.686
R10818 a_4090_5413.n1 a_4090_5413.t4 214.335
R10819 a_4090_5413.t13 a_4090_5413.n1 214.335
R10820 a_4090_5413.n4 a_4090_5413.t6 190.152
R10821 a_4090_5413.n4 a_4090_5413.t8 190.152
R10822 a_4090_5413.n2 a_4090_5413.t15 160.666
R10823 a_4090_5413.n3 a_4090_5413.t10 160.666
R10824 a_4090_5413.n7 a_4090_5413.n6 148.428
R10825 a_4090_5413.n5 a_4090_5413.t5 110.859
R10826 a_4090_5413.n3 a_4090_5413.n2 96.129
R10827 a_4090_5413.n8 a_4090_5413.t17 80.333
R10828 a_4090_5413.n1 a_4090_5413.t9 80.333
R10829 a_4090_5413.t18 a_4090_5413.n4 80.333
R10830 a_4090_5413.t3 a_4090_5413.n11 28.57
R10831 a_4090_5413.n0 a_4090_5413.t1 28.565
R10832 a_4090_5413.n0 a_4090_5413.t2 28.565
R10833 a_4090_5413.n11 a_4090_5413.t0 17.638
R10834 a_4090_5413.n10 a_4090_5413.n9 7.04
R10835 a_4090_5413.n9 a_4090_5413.n7 2.923
R10836 a_4090_5413.n10 a_4090_5413.n0 0.69
R10837 a_4090_5413.n11 a_4090_5413.n10 0.6
R10838 A[2].n4 A[2].n3 535.449
R10839 A[2].t15 A[2].t6 437.233
R10840 A[2].t12 A[2].t3 437.233
R10841 A[2].t7 A[2].n1 313.873
R10842 A[2].n3 A[2].t0 294.986
R10843 A[2].n0 A[2].t1 272.288
R10844 A[2].n4 A[2].t8 245.184
R10845 A[2].n6 A[2].t12 218.628
R10846 A[2].n8 A[2].t15 217.024
R10847 A[2].n7 A[2].t11 214.686
R10848 A[2].t6 A[2].n7 214.686
R10849 A[2].n5 A[2].t4 214.686
R10850 A[2].t3 A[2].n5 214.686
R10851 A[2].n2 A[2].t7 190.152
R10852 A[2].n2 A[2].t10 190.152
R10853 A[2].n0 A[2].t13 160.666
R10854 A[2].n1 A[2].t14 160.666
R10855 A[2].n3 A[2].t9 110.859
R10856 A[2].n1 A[2].n0 96.129
R10857 A[2].n7 A[2].t5 80.333
R10858 A[2].t8 A[2].n2 80.333
R10859 A[2].n5 A[2].t2 80.333
R10860 A[2] A[2].n8 27.013
R10861 A[2].n6 A[2].n4 14.9
R10862 A[2].n8 A[2].n6 2.599
R10863 a_23986_11307.n2 a_23986_11307.t10 214.335
R10864 a_23986_11307.t8 a_23986_11307.n2 214.335
R10865 a_23986_11307.n3 a_23986_11307.t8 143.851
R10866 a_23986_11307.n3 a_23986_11307.t7 135.658
R10867 a_23986_11307.n2 a_23986_11307.t9 80.333
R10868 a_23986_11307.n4 a_23986_11307.t0 28.565
R10869 a_23986_11307.n4 a_23986_11307.t1 28.565
R10870 a_23986_11307.n0 a_23986_11307.t6 28.565
R10871 a_23986_11307.n0 a_23986_11307.t4 28.565
R10872 a_23986_11307.t2 a_23986_11307.n7 28.565
R10873 a_23986_11307.n7 a_23986_11307.t5 28.565
R10874 a_23986_11307.n1 a_23986_11307.t3 9.714
R10875 a_23986_11307.n1 a_23986_11307.n0 1.003
R10876 a_23986_11307.n6 a_23986_11307.n5 0.833
R10877 a_23986_11307.n5 a_23986_11307.n4 0.653
R10878 a_23986_11307.n7 a_23986_11307.n6 0.653
R10879 a_23986_11307.n6 a_23986_11307.n1 0.341
R10880 a_23986_11307.n5 a_23986_11307.n3 0.032
R10881 a_24576_10870.t6 a_24576_10870.t4 574.43
R10882 a_24576_10870.n0 a_24576_10870.t5 285.109
R10883 a_24576_10870.n2 a_24576_10870.n1 211.136
R10884 a_24576_10870.n4 a_24576_10870.n3 192.754
R10885 a_24576_10870.n0 a_24576_10870.t7 160.666
R10886 a_24576_10870.n1 a_24576_10870.t6 160.666
R10887 a_24576_10870.n1 a_24576_10870.n0 114.829
R10888 a_24576_10870.n3 a_24576_10870.t1 28.568
R10889 a_24576_10870.n4 a_24576_10870.t2 28.565
R10890 a_24576_10870.t3 a_24576_10870.n4 28.565
R10891 a_24576_10870.n2 a_24576_10870.t0 19.084
R10892 a_24576_10870.n3 a_24576_10870.n2 1.051
R10893 a_1254_13136.n0 a_1254_13136.t9 214.335
R10894 a_1254_13136.t8 a_1254_13136.n0 214.335
R10895 a_1254_13136.n1 a_1254_13136.t8 143.851
R10896 a_1254_13136.n1 a_1254_13136.t10 135.658
R10897 a_1254_13136.n0 a_1254_13136.t7 80.333
R10898 a_1254_13136.n2 a_1254_13136.t4 28.565
R10899 a_1254_13136.n2 a_1254_13136.t5 28.565
R10900 a_1254_13136.n4 a_1254_13136.t6 28.565
R10901 a_1254_13136.n4 a_1254_13136.t1 28.565
R10902 a_1254_13136.n7 a_1254_13136.t2 28.565
R10903 a_1254_13136.t3 a_1254_13136.n7 28.565
R10904 a_1254_13136.n6 a_1254_13136.t0 9.714
R10905 a_1254_13136.n7 a_1254_13136.n6 1.003
R10906 a_1254_13136.n5 a_1254_13136.n3 0.833
R10907 a_1254_13136.n3 a_1254_13136.n2 0.653
R10908 a_1254_13136.n5 a_1254_13136.n4 0.653
R10909 a_1254_13136.n6 a_1254_13136.n5 0.341
R10910 a_1254_13136.n3 a_1254_13136.n1 0.032
R10911 a_27321_12833.t5 a_27321_12833.n2 404.877
R10912 a_27321_12833.n1 a_27321_12833.t6 210.902
R10913 a_27321_12833.n3 a_27321_12833.t5 136.943
R10914 a_27321_12833.n2 a_27321_12833.n1 107.801
R10915 a_27321_12833.n1 a_27321_12833.t8 80.333
R10916 a_27321_12833.n2 a_27321_12833.t7 80.333
R10917 a_27321_12833.n0 a_27321_12833.t0 17.4
R10918 a_27321_12833.n0 a_27321_12833.t3 17.4
R10919 a_27321_12833.n4 a_27321_12833.t4 15.032
R10920 a_27321_12833.n5 a_27321_12833.t2 14.282
R10921 a_27321_12833.t1 a_27321_12833.n5 14.282
R10922 a_27321_12833.n5 a_27321_12833.n4 1.65
R10923 a_27321_12833.n3 a_27321_12833.n0 0.672
R10924 a_27321_12833.n4 a_27321_12833.n3 0.665
R10925 a_14036_6963.t8 a_14036_6963.n2 404.877
R10926 a_14036_6963.n1 a_14036_6963.t7 210.902
R10927 a_14036_6963.n3 a_14036_6963.t8 136.943
R10928 a_14036_6963.n2 a_14036_6963.n1 107.801
R10929 a_14036_6963.n1 a_14036_6963.t5 80.333
R10930 a_14036_6963.n2 a_14036_6963.t6 80.333
R10931 a_14036_6963.n0 a_14036_6963.t0 17.4
R10932 a_14036_6963.n0 a_14036_6963.t1 17.4
R10933 a_14036_6963.n4 a_14036_6963.t4 15.032
R10934 a_14036_6963.n5 a_14036_6963.t3 14.282
R10935 a_14036_6963.t2 a_14036_6963.n5 14.282
R10936 a_14036_6963.n5 a_14036_6963.n4 1.65
R10937 a_14036_6963.n3 a_14036_6963.n0 0.672
R10938 a_14036_6963.n4 a_14036_6963.n3 0.665
R10939 a_14154_6963.n1 a_14154_6963.t1 14.282
R10940 a_14154_6963.n1 a_14154_6963.t4 14.282
R10941 a_14154_6963.n0 a_14154_6963.t3 14.282
R10942 a_14154_6963.n0 a_14154_6963.t5 14.282
R10943 a_14154_6963.n3 a_14154_6963.t0 14.282
R10944 a_14154_6963.t2 a_14154_6963.n3 14.282
R10945 a_14154_6963.n2 a_14154_6963.n0 2.546
R10946 a_14154_6963.n3 a_14154_6963.n2 2.367
R10947 a_14154_6963.n2 a_14154_6963.n1 0.001
R10948 a_n3606_3562.n1 a_n3606_3562.t5 318.119
R10949 a_n3606_3562.n1 a_n3606_3562.t7 269.919
R10950 a_n3606_3562.n0 a_n3606_3562.t6 267.256
R10951 a_n3606_3562.n0 a_n3606_3562.t4 267.256
R10952 a_n3606_3562.n4 a_n3606_3562.n3 193.227
R10953 a_n3606_3562.t5 a_n3606_3562.n0 160.666
R10954 a_n3606_3562.n2 a_n3606_3562.n1 106.999
R10955 a_n3606_3562.n3 a_n3606_3562.t1 28.568
R10956 a_n3606_3562.n4 a_n3606_3562.t2 28.565
R10957 a_n3606_3562.t3 a_n3606_3562.n4 28.565
R10958 a_n3606_3562.n2 a_n3606_3562.t0 18.149
R10959 a_n3606_3562.n3 a_n3606_3562.n2 3.726
R10960 a_23092_24426.n1 a_23092_24426.t6 318.922
R10961 a_23092_24426.n0 a_23092_24426.t5 274.739
R10962 a_23092_24426.n0 a_23092_24426.t7 274.739
R10963 a_23092_24426.n1 a_23092_24426.t4 269.116
R10964 a_23092_24426.t6 a_23092_24426.n0 179.946
R10965 a_23092_24426.n2 a_23092_24426.n1 105.178
R10966 a_23092_24426.n3 a_23092_24426.t1 29.444
R10967 a_23092_24426.n4 a_23092_24426.t2 28.565
R10968 a_23092_24426.t3 a_23092_24426.n4 28.565
R10969 a_23092_24426.n2 a_23092_24426.t0 18.145
R10970 a_23092_24426.n3 a_23092_24426.n2 2.878
R10971 a_23092_24426.n4 a_23092_24426.n3 0.764
R10972 a_22798_23720.t0 a_22798_23720.t1 380.209
R10973 a_n3606_6260.n1 a_n3606_6260.t6 318.119
R10974 a_n3606_6260.n1 a_n3606_6260.t7 269.919
R10975 a_n3606_6260.n0 a_n3606_6260.t4 267.853
R10976 a_n3606_6260.n0 a_n3606_6260.t5 267.853
R10977 a_n3606_6260.t6 a_n3606_6260.n0 160.666
R10978 a_n3606_6260.n2 a_n3606_6260.n1 107.263
R10979 a_n3606_6260.n3 a_n3606_6260.t2 29.444
R10980 a_n3606_6260.t3 a_n3606_6260.n4 28.565
R10981 a_n3606_6260.n4 a_n3606_6260.t1 28.565
R10982 a_n3606_6260.n2 a_n3606_6260.t0 18.145
R10983 a_n3606_6260.n3 a_n3606_6260.n2 2.878
R10984 a_n3606_6260.n4 a_n3606_6260.n3 0.764
R10985 a_n3806_6861.n8 a_n3806_6861.n7 267.767
R10986 a_n3806_6861.n1 a_n3806_6861.t9 16.058
R10987 a_n3806_6861.n3 a_n3806_6861.t4 16.058
R10988 a_n3806_6861.n0 a_n3806_6861.t10 14.282
R10989 a_n3806_6861.n0 a_n3806_6861.t11 14.282
R10990 a_n3806_6861.n2 a_n3806_6861.t5 14.282
R10991 a_n3806_6861.n2 a_n3806_6861.t3 14.282
R10992 a_n3806_6861.n5 a_n3806_6861.t0 14.282
R10993 a_n3806_6861.n5 a_n3806_6861.t1 14.282
R10994 a_n3806_6861.n7 a_n3806_6861.t7 14.282
R10995 a_n3806_6861.n7 a_n3806_6861.t8 14.282
R10996 a_n3806_6861.t2 a_n3806_6861.n9 14.282
R10997 a_n3806_6861.n9 a_n3806_6861.t6 14.282
R10998 a_n3806_6861.n6 a_n3806_6861.n5 1.511
R10999 a_n3806_6861.n1 a_n3806_6861.n0 0.999
R11000 a_n3806_6861.n3 a_n3806_6861.n2 0.999
R11001 a_n3806_6861.n8 a_n3806_6861.n6 0.669
R11002 a_n3806_6861.n4 a_n3806_6861.n1 0.575
R11003 a_n3806_6861.n6 a_n3806_6861.n4 0.227
R11004 a_n3806_6861.n4 a_n3806_6861.n3 0.2
R11005 a_n3806_6861.n9 a_n3806_6861.n8 0.001
R11006 a_12418_19515.t1 a_12418_19515.n0 14.282
R11007 a_12418_19515.n0 a_12418_19515.t2 14.282
R11008 a_12418_19515.n0 a_12418_19515.n12 122.747
R11009 a_12418_19515.n8 a_12418_19515.n10 74.302
R11010 a_12418_19515.n12 a_12418_19515.n8 50.575
R11011 a_12418_19515.n12 a_12418_19515.n11 157.665
R11012 a_12418_19515.n11 a_12418_19515.t0 8.7
R11013 a_12418_19515.n11 a_12418_19515.t7 8.7
R11014 a_12418_19515.n10 a_12418_19515.n9 90.436
R11015 a_12418_19515.n9 a_12418_19515.t5 14.282
R11016 a_12418_19515.n9 a_12418_19515.t4 14.282
R11017 a_12418_19515.n8 a_12418_19515.n7 90.416
R11018 a_12418_19515.n7 a_12418_19515.t6 14.282
R11019 a_12418_19515.n7 a_12418_19515.t3 14.282
R11020 a_12418_19515.n10 a_12418_19515.n1 342.688
R11021 a_12418_19515.n1 a_12418_19515.n6 126.566
R11022 a_12418_19515.n6 a_12418_19515.t13 294.653
R11023 a_12418_19515.n6 a_12418_19515.t11 111.663
R11024 a_12418_19515.n1 a_12418_19515.n5 552.333
R11025 a_12418_19515.n5 a_12418_19515.n4 6.615
R11026 a_12418_19515.n4 a_12418_19515.t12 93.989
R11027 a_12418_19515.n4 a_12418_19515.t15 198.043
R11028 a_12418_19515.n5 a_12418_19515.n3 97.816
R11029 a_12418_19515.n3 a_12418_19515.t14 80.333
R11030 a_12418_19515.n3 a_12418_19515.t10 394.151
R11031 a_12418_19515.t10 a_12418_19515.n2 269.523
R11032 a_12418_19515.n2 a_12418_19515.t9 160.666
R11033 a_12418_19515.n2 a_12418_19515.t8 269.523
R11034 a_12480_9997.n0 a_12480_9997.t2 14.282
R11035 a_12480_9997.t0 a_12480_9997.n0 14.282
R11036 a_12480_9997.n0 a_12480_9997.n9 0.999
R11037 a_12480_9997.n6 a_12480_9997.n8 0.575
R11038 a_12480_9997.n9 a_12480_9997.n6 0.2
R11039 a_12480_9997.n9 a_12480_9997.t1 16.058
R11040 a_12480_9997.n8 a_12480_9997.n7 0.999
R11041 a_12480_9997.n7 a_12480_9997.t8 14.282
R11042 a_12480_9997.n7 a_12480_9997.t7 14.282
R11043 a_12480_9997.n8 a_12480_9997.t6 16.058
R11044 a_12480_9997.n6 a_12480_9997.n4 0.227
R11045 a_12480_9997.n4 a_12480_9997.n5 1.511
R11046 a_12480_9997.n5 a_12480_9997.t11 14.282
R11047 a_12480_9997.n5 a_12480_9997.t10 14.282
R11048 a_12480_9997.n4 a_12480_9997.n1 0.669
R11049 a_12480_9997.n1 a_12480_9997.n2 0.001
R11050 a_12480_9997.n1 a_12480_9997.n3 267.767
R11051 a_12480_9997.n3 a_12480_9997.t5 14.282
R11052 a_12480_9997.n3 a_12480_9997.t4 14.282
R11053 a_12480_9997.n2 a_12480_9997.t9 14.282
R11054 a_12480_9997.n2 a_12480_9997.t3 14.282
R11055 a_n2383_5086.t0 a_n2383_5086.t1 17.4
R11056 a_17932_6651.t4 a_17932_6651.t7 800.071
R11057 a_17932_6651.n2 a_17932_6651.n1 659.097
R11058 a_17932_6651.n0 a_17932_6651.t5 285.109
R11059 a_17932_6651.n1 a_17932_6651.t4 193.602
R11060 a_17932_6651.n4 a_17932_6651.n3 192.754
R11061 a_17932_6651.n0 a_17932_6651.t6 160.666
R11062 a_17932_6651.n1 a_17932_6651.n0 91.507
R11063 a_17932_6651.n3 a_17932_6651.t2 28.568
R11064 a_17932_6651.n4 a_17932_6651.t1 28.565
R11065 a_17932_6651.t3 a_17932_6651.n4 28.565
R11066 a_17932_6651.n2 a_17932_6651.t0 19.061
R11067 a_17932_6651.n3 a_17932_6651.n2 1.005
R11068 a_7821_4129.t0 a_7821_4129.n0 14.282
R11069 a_7821_4129.n0 a_7821_4129.t1 14.282
R11070 a_7821_4129.n0 a_7821_4129.n9 0.999
R11071 a_7821_4129.n6 a_7821_4129.n8 0.575
R11072 a_7821_4129.n9 a_7821_4129.n6 0.2
R11073 a_7821_4129.n9 a_7821_4129.t8 16.058
R11074 a_7821_4129.n8 a_7821_4129.n7 0.999
R11075 a_7821_4129.n7 a_7821_4129.t2 14.282
R11076 a_7821_4129.n7 a_7821_4129.t3 14.282
R11077 a_7821_4129.n8 a_7821_4129.t4 16.058
R11078 a_7821_4129.n6 a_7821_4129.n4 0.227
R11079 a_7821_4129.n4 a_7821_4129.n5 1.511
R11080 a_7821_4129.n5 a_7821_4129.t11 14.282
R11081 a_7821_4129.n5 a_7821_4129.t10 14.282
R11082 a_7821_4129.n4 a_7821_4129.n1 0.669
R11083 a_7821_4129.n1 a_7821_4129.n2 0.001
R11084 a_7821_4129.n1 a_7821_4129.n3 267.767
R11085 a_7821_4129.n3 a_7821_4129.t5 14.282
R11086 a_7821_4129.n3 a_7821_4129.t7 14.282
R11087 a_7821_4129.n2 a_7821_4129.t9 14.282
R11088 a_7821_4129.n2 a_7821_4129.t6 14.282
R11089 a_12598_9997.n0 a_12598_9997.n12 122.999
R11090 a_12598_9997.t3 a_12598_9997.n0 14.282
R11091 a_12598_9997.n0 a_12598_9997.t6 14.282
R11092 a_12598_9997.n12 a_12598_9997.n10 50.575
R11093 a_12598_9997.n10 a_12598_9997.n8 74.302
R11094 a_12598_9997.n12 a_12598_9997.n11 157.665
R11095 a_12598_9997.n11 a_12598_9997.t4 8.7
R11096 a_12598_9997.n11 a_12598_9997.t7 8.7
R11097 a_12598_9997.n10 a_12598_9997.n9 90.416
R11098 a_12598_9997.n9 a_12598_9997.t5 14.282
R11099 a_12598_9997.n9 a_12598_9997.t2 14.282
R11100 a_12598_9997.n8 a_12598_9997.n7 90.436
R11101 a_12598_9997.n7 a_12598_9997.t0 14.282
R11102 a_12598_9997.n7 a_12598_9997.t1 14.282
R11103 a_12598_9997.n8 a_12598_9997.n1 342.688
R11104 a_12598_9997.n1 a_12598_9997.n6 126.566
R11105 a_12598_9997.n6 a_12598_9997.t13 294.653
R11106 a_12598_9997.n6 a_12598_9997.t15 111.663
R11107 a_12598_9997.n1 a_12598_9997.n5 552.333
R11108 a_12598_9997.n5 a_12598_9997.n4 6.615
R11109 a_12598_9997.n4 a_12598_9997.t11 93.989
R11110 a_12598_9997.n5 a_12598_9997.n3 97.816
R11111 a_12598_9997.n3 a_12598_9997.t12 80.333
R11112 a_12598_9997.n3 a_12598_9997.t14 394.151
R11113 a_12598_9997.t14 a_12598_9997.n2 269.523
R11114 a_12598_9997.n2 a_12598_9997.t8 160.666
R11115 a_12598_9997.n2 a_12598_9997.t9 269.523
R11116 a_12598_9997.n4 a_12598_9997.t10 198.043
R11117 a_12834_9265.t0 a_12834_9265.t1 17.4
R11118 a_26143_26979.t4 a_26143_26979.t6 800.071
R11119 a_26143_26979.n3 a_26143_26979.n2 659.097
R11120 a_26143_26979.n1 a_26143_26979.t7 285.109
R11121 a_26143_26979.n2 a_26143_26979.t4 193.602
R11122 a_26143_26979.n4 a_26143_26979.n0 192.754
R11123 a_26143_26979.n1 a_26143_26979.t5 160.666
R11124 a_26143_26979.n2 a_26143_26979.n1 91.507
R11125 a_26143_26979.t0 a_26143_26979.n4 28.568
R11126 a_26143_26979.n0 a_26143_26979.t1 28.565
R11127 a_26143_26979.n0 a_26143_26979.t3 28.565
R11128 a_26143_26979.n3 a_26143_26979.t2 19.061
R11129 a_26143_26979.n4 a_26143_26979.n3 1.005
R11130 a_27649_4129.n0 a_27649_4129.n1 0.001
R11131 a_27649_4129.t0 a_27649_4129.n0 14.282
R11132 a_27649_4129.n0 a_27649_4129.t11 14.282
R11133 a_27649_4129.n1 a_27649_4129.n9 267.767
R11134 a_27649_4129.n9 a_27649_4129.t9 14.282
R11135 a_27649_4129.n9 a_27649_4129.t10 14.282
R11136 a_27649_4129.n1 a_27649_4129.n7 0.669
R11137 a_27649_4129.n7 a_27649_4129.n8 1.511
R11138 a_27649_4129.n8 a_27649_4129.t7 14.282
R11139 a_27649_4129.n8 a_27649_4129.t8 14.282
R11140 a_27649_4129.n7 a_27649_4129.n6 0.227
R11141 a_27649_4129.n6 a_27649_4129.n3 0.575
R11142 a_27649_4129.n6 a_27649_4129.n5 0.2
R11143 a_27649_4129.n5 a_27649_4129.t5 16.058
R11144 a_27649_4129.n5 a_27649_4129.n4 0.999
R11145 a_27649_4129.n4 a_27649_4129.t6 14.282
R11146 a_27649_4129.n4 a_27649_4129.t4 14.282
R11147 a_27649_4129.n3 a_27649_4129.n2 0.999
R11148 a_27649_4129.n2 a_27649_4129.t1 14.282
R11149 a_27649_4129.n2 a_27649_4129.t2 14.282
R11150 a_27649_4129.n3 a_27649_4129.t3 16.058
R11151 a_25562_24162.n0 a_25562_24162.t10 214.335
R11152 a_25562_24162.t7 a_25562_24162.n0 214.335
R11153 a_25562_24162.n1 a_25562_24162.t7 143.851
R11154 a_25562_24162.n1 a_25562_24162.t8 135.658
R11155 a_25562_24162.n0 a_25562_24162.t9 80.333
R11156 a_25562_24162.n2 a_25562_24162.t6 28.565
R11157 a_25562_24162.n2 a_25562_24162.t4 28.565
R11158 a_25562_24162.n4 a_25562_24162.t5 28.565
R11159 a_25562_24162.n4 a_25562_24162.t1 28.565
R11160 a_25562_24162.n7 a_25562_24162.t2 28.565
R11161 a_25562_24162.t3 a_25562_24162.n7 28.565
R11162 a_25562_24162.n6 a_25562_24162.t0 9.714
R11163 a_25562_24162.n7 a_25562_24162.n6 1.003
R11164 a_25562_24162.n5 a_25562_24162.n3 0.833
R11165 a_25562_24162.n3 a_25562_24162.n2 0.653
R11166 a_25562_24162.n5 a_25562_24162.n4 0.653
R11167 a_25562_24162.n6 a_25562_24162.n5 0.341
R11168 a_25562_24162.n3 a_25562_24162.n1 0.032
R11169 a_n2383_713.t0 a_n2383_713.t1 379.845
R11170 a_33377_6895.n2 a_33377_6895.t7 214.335
R11171 a_33377_6895.t10 a_33377_6895.n2 214.335
R11172 a_33377_6895.n3 a_33377_6895.t10 143.851
R11173 a_33377_6895.n3 a_33377_6895.t8 135.658
R11174 a_33377_6895.n2 a_33377_6895.t9 80.333
R11175 a_33377_6895.n4 a_33377_6895.t5 28.565
R11176 a_33377_6895.n4 a_33377_6895.t6 28.565
R11177 a_33377_6895.n0 a_33377_6895.t1 28.565
R11178 a_33377_6895.n0 a_33377_6895.t3 28.565
R11179 a_33377_6895.t4 a_33377_6895.n7 28.565
R11180 a_33377_6895.n7 a_33377_6895.t2 28.565
R11181 a_33377_6895.n1 a_33377_6895.t0 9.714
R11182 a_33377_6895.n1 a_33377_6895.n0 1.003
R11183 a_33377_6895.n6 a_33377_6895.n5 0.833
R11184 a_33377_6895.n5 a_33377_6895.n4 0.653
R11185 a_33377_6895.n7 a_33377_6895.n6 0.653
R11186 a_33377_6895.n6 a_33377_6895.n1 0.341
R11187 a_33377_6895.n5 a_33377_6895.n3 0.032
R11188 a_10924_6450.t0 a_10924_6450.t1 17.4
R11189 a_13961_18848.n0 a_13961_18848.n1 0.001
R11190 a_13961_18848.n0 a_13961_18848.t2 14.282
R11191 a_13961_18848.t0 a_13961_18848.n0 14.282
R11192 a_13961_18848.n1 a_13961_18848.n9 267.767
R11193 a_13961_18848.n9 a_13961_18848.t3 14.282
R11194 a_13961_18848.n9 a_13961_18848.t4 14.282
R11195 a_13961_18848.n1 a_13961_18848.n7 0.669
R11196 a_13961_18848.n7 a_13961_18848.n8 1.511
R11197 a_13961_18848.n8 a_13961_18848.t1 14.282
R11198 a_13961_18848.n8 a_13961_18848.t11 14.282
R11199 a_13961_18848.n7 a_13961_18848.n6 0.227
R11200 a_13961_18848.n6 a_13961_18848.n3 0.2
R11201 a_13961_18848.n6 a_13961_18848.n5 0.575
R11202 a_13961_18848.n5 a_13961_18848.t6 16.058
R11203 a_13961_18848.n5 a_13961_18848.n4 0.999
R11204 a_13961_18848.n4 a_13961_18848.t7 14.282
R11205 a_13961_18848.n4 a_13961_18848.t5 14.282
R11206 a_13961_18848.n3 a_13961_18848.n2 0.999
R11207 a_13961_18848.n2 a_13961_18848.t8 14.282
R11208 a_13961_18848.n2 a_13961_18848.t10 14.282
R11209 a_13961_18848.n3 a_13961_18848.t9 16.058
R11210 a_10647_11281.n6 a_10647_11281.n5 501.28
R11211 a_10647_11281.t6 a_10647_11281.t18 437.233
R11212 a_10647_11281.t9 a_10647_11281.t4 415.315
R11213 a_10647_11281.t5 a_10647_11281.n3 313.873
R11214 a_10647_11281.n5 a_10647_11281.t8 294.986
R11215 a_10647_11281.n2 a_10647_11281.t10 272.288
R11216 a_10647_11281.n6 a_10647_11281.t12 236.01
R11217 a_10647_11281.n9 a_10647_11281.t6 216.627
R11218 a_10647_11281.n7 a_10647_11281.t9 216.111
R11219 a_10647_11281.n8 a_10647_11281.t16 214.686
R11220 a_10647_11281.t18 a_10647_11281.n8 214.686
R11221 a_10647_11281.n1 a_10647_11281.t14 214.335
R11222 a_10647_11281.t4 a_10647_11281.n1 214.335
R11223 a_10647_11281.n4 a_10647_11281.t5 190.152
R11224 a_10647_11281.n4 a_10647_11281.t13 190.152
R11225 a_10647_11281.n2 a_10647_11281.t11 160.666
R11226 a_10647_11281.n3 a_10647_11281.t7 160.666
R11227 a_10647_11281.n7 a_10647_11281.n6 148.428
R11228 a_10647_11281.n5 a_10647_11281.t15 110.859
R11229 a_10647_11281.n3 a_10647_11281.n2 96.129
R11230 a_10647_11281.n8 a_10647_11281.t17 80.333
R11231 a_10647_11281.n1 a_10647_11281.t19 80.333
R11232 a_10647_11281.t12 a_10647_11281.n4 80.333
R11233 a_10647_11281.n0 a_10647_11281.t2 28.57
R11234 a_10647_11281.n11 a_10647_11281.t1 28.565
R11235 a_10647_11281.t3 a_10647_11281.n11 28.565
R11236 a_10647_11281.n0 a_10647_11281.t0 17.638
R11237 a_10647_11281.n10 a_10647_11281.n9 12.318
R11238 a_10647_11281.n9 a_10647_11281.n7 2.923
R11239 a_10647_11281.n11 a_10647_11281.n10 0.69
R11240 a_10647_11281.n10 a_10647_11281.n0 0.6
R11241 a_27008_18856.n9 a_27008_18856.n8 267.767
R11242 a_27008_18856.n3 a_27008_18856.t5 16.058
R11243 a_27008_18856.n1 a_27008_18856.t10 16.058
R11244 a_27008_18856.n2 a_27008_18856.t3 14.282
R11245 a_27008_18856.n2 a_27008_18856.t4 14.282
R11246 a_27008_18856.n0 a_27008_18856.t11 14.282
R11247 a_27008_18856.n0 a_27008_18856.t9 14.282
R11248 a_27008_18856.n5 a_27008_18856.t6 14.282
R11249 a_27008_18856.n5 a_27008_18856.t7 14.282
R11250 a_27008_18856.n7 a_27008_18856.t8 14.282
R11251 a_27008_18856.n7 a_27008_18856.t0 14.282
R11252 a_27008_18856.n9 a_27008_18856.t1 14.282
R11253 a_27008_18856.t2 a_27008_18856.n9 14.282
R11254 a_27008_18856.n6 a_27008_18856.n5 1.511
R11255 a_27008_18856.n3 a_27008_18856.n2 0.999
R11256 a_27008_18856.n1 a_27008_18856.n0 0.999
R11257 a_27008_18856.n8 a_27008_18856.n6 0.669
R11258 a_27008_18856.n4 a_27008_18856.n1 0.575
R11259 a_27008_18856.n6 a_27008_18856.n4 0.227
R11260 a_27008_18856.n4 a_27008_18856.n3 0.2
R11261 a_27008_18856.n8 a_27008_18856.n7 0.001
R11262 a_36751_971.n0 a_36751_971.t6 14.282
R11263 a_36751_971.t0 a_36751_971.n0 14.282
R11264 a_36751_971.n0 a_36751_971.n1 258.161
R11265 a_36751_971.n1 a_36751_971.n7 4.366
R11266 a_36751_971.n7 a_36751_971.n5 0.852
R11267 a_36751_971.n5 a_36751_971.n6 258.161
R11268 a_36751_971.n6 a_36751_971.t2 14.282
R11269 a_36751_971.n6 a_36751_971.t4 14.282
R11270 a_36751_971.n5 a_36751_971.t3 14.283
R11271 a_36751_971.n7 a_36751_971.n4 73.514
R11272 a_36751_971.n4 a_36751_971.t9 1551.5
R11273 a_36751_971.t9 a_36751_971.n3 656.576
R11274 a_36751_971.n3 a_36751_971.t1 8.7
R11275 a_36751_971.n3 a_36751_971.t7 8.7
R11276 a_36751_971.n4 a_36751_971.t8 224.129
R11277 a_36751_971.t8 a_36751_971.n2 207.225
R11278 a_36751_971.n2 a_36751_971.t11 207.225
R11279 a_36751_971.n2 a_36751_971.t10 80.333
R11280 a_36751_971.n1 a_36751_971.t5 14.283
R11281 Y[7].n1 Y[7].n0 185.55
R11282 Y[7].n1 Y[7].t3 28.568
R11283 Y[7].n0 Y[7].t1 28.565
R11284 Y[7].n0 Y[7].t2 28.565
R11285 Y[7].n2 Y[7].t0 20.393
R11286 Y[7].n2 Y[7].n1 1.886
R11287 Y[7].n3 Y[7].n2 1.307
R11288 Y[7] Y[7].n3 0.05
R11289 Y[7].n3 Y[7] 0.048
R11290 a_4136_7089.n0 a_4136_7089.t9 214.335
R11291 a_4136_7089.t10 a_4136_7089.n0 214.335
R11292 a_4136_7089.n1 a_4136_7089.t10 143.851
R11293 a_4136_7089.n1 a_4136_7089.t7 135.658
R11294 a_4136_7089.n0 a_4136_7089.t8 80.333
R11295 a_4136_7089.n2 a_4136_7089.t5 28.565
R11296 a_4136_7089.n2 a_4136_7089.t4 28.565
R11297 a_4136_7089.n4 a_4136_7089.t6 28.565
R11298 a_4136_7089.n4 a_4136_7089.t1 28.565
R11299 a_4136_7089.t3 a_4136_7089.n7 28.565
R11300 a_4136_7089.n7 a_4136_7089.t2 28.565
R11301 a_4136_7089.n6 a_4136_7089.t0 9.714
R11302 a_4136_7089.n7 a_4136_7089.n6 1.003
R11303 a_4136_7089.n5 a_4136_7089.n3 0.833
R11304 a_4136_7089.n3 a_4136_7089.n2 0.653
R11305 a_4136_7089.n5 a_4136_7089.n4 0.653
R11306 a_4136_7089.n6 a_4136_7089.n5 0.341
R11307 a_4136_7089.n3 a_4136_7089.n1 0.032
R11308 a_27313_6965.t5 a_27313_6965.n2 404.877
R11309 a_27313_6965.n1 a_27313_6965.t8 210.902
R11310 a_27313_6965.n3 a_27313_6965.t5 136.943
R11311 a_27313_6965.n2 a_27313_6965.n1 107.801
R11312 a_27313_6965.n1 a_27313_6965.t7 80.333
R11313 a_27313_6965.n2 a_27313_6965.t6 80.333
R11314 a_27313_6965.n0 a_27313_6965.t4 17.4
R11315 a_27313_6965.n0 a_27313_6965.t2 17.4
R11316 a_27313_6965.n4 a_27313_6965.t3 15.032
R11317 a_27313_6965.n5 a_27313_6965.t1 14.282
R11318 a_27313_6965.t0 a_27313_6965.n5 14.282
R11319 a_27313_6965.n5 a_27313_6965.n4 1.65
R11320 a_27313_6965.n3 a_27313_6965.n0 0.672
R11321 a_27313_6965.n4 a_27313_6965.n3 0.665
R11322 a_27431_6965.n1 a_27431_6965.t5 14.282
R11323 a_27431_6965.n1 a_27431_6965.t1 14.282
R11324 a_27431_6965.n0 a_27431_6965.t2 14.282
R11325 a_27431_6965.n0 a_27431_6965.t3 14.282
R11326 a_27431_6965.n3 a_27431_6965.t4 14.282
R11327 a_27431_6965.t0 a_27431_6965.n3 14.282
R11328 a_27431_6965.n2 a_27431_6965.n0 2.546
R11329 a_27431_6965.n3 a_27431_6965.n2 2.367
R11330 a_27431_6965.n2 a_27431_6965.n1 0.001
R11331 a_30427_3858.n5 a_30427_3858.n4 465.933
R11332 a_30427_3858.t5 a_30427_3858.t4 415.315
R11333 a_30427_3858.n1 a_30427_3858.t15 394.151
R11334 a_30427_3858.n4 a_30427_3858.t14 294.653
R11335 a_30427_3858.n0 a_30427_3858.t7 269.523
R11336 a_30427_3858.t15 a_30427_3858.n0 269.523
R11337 a_30427_3858.n7 a_30427_3858.t5 220.285
R11338 a_30427_3858.n6 a_30427_3858.t12 214.335
R11339 a_30427_3858.t4 a_30427_3858.n6 214.335
R11340 a_30427_3858.n2 a_30427_3858.t6 198.043
R11341 a_30427_3858.n10 a_30427_3858.n9 192.754
R11342 a_30427_3858.n5 a_30427_3858.n3 163.88
R11343 a_30427_3858.n0 a_30427_3858.t10 160.666
R11344 a_30427_3858.n4 a_30427_3858.t11 111.663
R11345 a_30427_3858.n3 a_30427_3858.n1 97.816
R11346 a_30427_3858.n2 a_30427_3858.t13 93.989
R11347 a_30427_3858.n6 a_30427_3858.t8 80.333
R11348 a_30427_3858.n1 a_30427_3858.t9 80.333
R11349 a_30427_3858.n7 a_30427_3858.n5 61.538
R11350 a_30427_3858.n9 a_30427_3858.t2 28.568
R11351 a_30427_3858.n10 a_30427_3858.t1 28.565
R11352 a_30427_3858.t3 a_30427_3858.n10 28.565
R11353 a_30427_3858.n8 a_30427_3858.t0 18.824
R11354 a_30427_3858.n3 a_30427_3858.n2 6.615
R11355 a_30427_3858.n8 a_30427_3858.n7 4.769
R11356 a_30427_3858.n9 a_30427_3858.n8 1.105
R11357 a_n3606_8329.n1 a_n3606_8329.t7 318.119
R11358 a_n3606_8329.n1 a_n3606_8329.t4 269.919
R11359 a_n3606_8329.n0 a_n3606_8329.t5 267.853
R11360 a_n3606_8329.n0 a_n3606_8329.t6 267.853
R11361 a_n3606_8329.t7 a_n3606_8329.n0 160.666
R11362 a_n3606_8329.n2 a_n3606_8329.n1 107.263
R11363 a_n3606_8329.n3 a_n3606_8329.t2 29.444
R11364 a_n3606_8329.t3 a_n3606_8329.n4 28.565
R11365 a_n3606_8329.n4 a_n3606_8329.t1 28.565
R11366 a_n3606_8329.n2 a_n3606_8329.t0 18.145
R11367 a_n3606_8329.n3 a_n3606_8329.n2 2.878
R11368 a_n3606_8329.n4 a_n3606_8329.n3 0.764
R11369 a_29769_9285.n0 a_29769_9285.t9 214.335
R11370 a_29769_9285.t7 a_29769_9285.n0 214.335
R11371 a_29769_9285.n1 a_29769_9285.t7 143.851
R11372 a_29769_9285.n1 a_29769_9285.t8 135.658
R11373 a_29769_9285.n0 a_29769_9285.t10 80.333
R11374 a_29769_9285.n2 a_29769_9285.t4 28.565
R11375 a_29769_9285.n2 a_29769_9285.t6 28.565
R11376 a_29769_9285.n4 a_29769_9285.t5 28.565
R11377 a_29769_9285.n4 a_29769_9285.t1 28.565
R11378 a_29769_9285.t3 a_29769_9285.n7 28.565
R11379 a_29769_9285.n7 a_29769_9285.t2 28.565
R11380 a_29769_9285.n6 a_29769_9285.t0 9.714
R11381 a_29769_9285.n7 a_29769_9285.n6 1.003
R11382 a_29769_9285.n5 a_29769_9285.n3 0.833
R11383 a_29769_9285.n3 a_29769_9285.n2 0.653
R11384 a_29769_9285.n5 a_29769_9285.n4 0.653
R11385 a_29769_9285.n6 a_29769_9285.n5 0.341
R11386 a_29769_9285.n3 a_29769_9285.n1 0.032
R11387 a_25751_4129.n0 a_25751_4129.t4 14.282
R11388 a_25751_4129.t0 a_25751_4129.n0 14.282
R11389 a_25751_4129.n0 a_25751_4129.n9 0.999
R11390 a_25751_4129.n9 a_25751_4129.n6 0.575
R11391 a_25751_4129.n6 a_25751_4129.n8 0.2
R11392 a_25751_4129.n8 a_25751_4129.t2 16.058
R11393 a_25751_4129.n8 a_25751_4129.n7 0.999
R11394 a_25751_4129.n7 a_25751_4129.t1 14.282
R11395 a_25751_4129.n7 a_25751_4129.t3 14.282
R11396 a_25751_4129.n9 a_25751_4129.t5 16.058
R11397 a_25751_4129.n6 a_25751_4129.n4 0.227
R11398 a_25751_4129.n4 a_25751_4129.n5 1.511
R11399 a_25751_4129.n5 a_25751_4129.t6 14.282
R11400 a_25751_4129.n5 a_25751_4129.t7 14.282
R11401 a_25751_4129.n4 a_25751_4129.n1 0.669
R11402 a_25751_4129.n1 a_25751_4129.n2 0.001
R11403 a_25751_4129.n1 a_25751_4129.n3 267.767
R11404 a_25751_4129.n3 a_25751_4129.t11 14.282
R11405 a_25751_4129.n3 a_25751_4129.t9 14.282
R11406 a_25751_4129.n2 a_25751_4129.t8 14.282
R11407 a_25751_4129.n2 a_25751_4129.t10 14.282
R11408 a_23981_9703.n2 a_23981_9703.t7 214.335
R11409 a_23981_9703.t10 a_23981_9703.n2 214.335
R11410 a_23981_9703.n3 a_23981_9703.t10 143.851
R11411 a_23981_9703.n3 a_23981_9703.t8 135.658
R11412 a_23981_9703.n2 a_23981_9703.t9 80.333
R11413 a_23981_9703.n4 a_23981_9703.t5 28.565
R11414 a_23981_9703.n4 a_23981_9703.t4 28.565
R11415 a_23981_9703.n0 a_23981_9703.t3 28.565
R11416 a_23981_9703.n0 a_23981_9703.t1 28.565
R11417 a_23981_9703.n7 a_23981_9703.t6 28.565
R11418 a_23981_9703.t0 a_23981_9703.n7 28.565
R11419 a_23981_9703.n1 a_23981_9703.t2 9.714
R11420 a_23981_9703.n1 a_23981_9703.n0 1.003
R11421 a_23981_9703.n6 a_23981_9703.n5 0.833
R11422 a_23981_9703.n5 a_23981_9703.n4 0.653
R11423 a_23981_9703.n7 a_23981_9703.n6 0.653
R11424 a_23981_9703.n6 a_23981_9703.n1 0.341
R11425 a_23981_9703.n5 a_23981_9703.n3 0.032
R11426 a_24571_9266.t5 a_24571_9266.t4 574.43
R11427 a_24571_9266.n1 a_24571_9266.t7 285.109
R11428 a_24571_9266.n3 a_24571_9266.n2 197.217
R11429 a_24571_9266.n4 a_24571_9266.n0 192.754
R11430 a_24571_9266.n1 a_24571_9266.t6 160.666
R11431 a_24571_9266.n2 a_24571_9266.t5 160.666
R11432 a_24571_9266.n2 a_24571_9266.n1 114.829
R11433 a_24571_9266.t3 a_24571_9266.n4 28.568
R11434 a_24571_9266.n0 a_24571_9266.t2 28.565
R11435 a_24571_9266.n0 a_24571_9266.t1 28.565
R11436 a_24571_9266.n3 a_24571_9266.t0 18.838
R11437 a_24571_9266.n4 a_24571_9266.n3 1.129
R11438 a_n3608_1494.n1 a_n3608_1494.t7 318.119
R11439 a_n3608_1494.n1 a_n3608_1494.t4 269.919
R11440 a_n3608_1494.n0 a_n3608_1494.t5 267.256
R11441 a_n3608_1494.n0 a_n3608_1494.t6 267.256
R11442 a_n3608_1494.n4 a_n3608_1494.n3 193.227
R11443 a_n3608_1494.t7 a_n3608_1494.n0 160.666
R11444 a_n3608_1494.n2 a_n3608_1494.n1 106.999
R11445 a_n3608_1494.n3 a_n3608_1494.t2 28.568
R11446 a_n3608_1494.t3 a_n3608_1494.n4 28.565
R11447 a_n3608_1494.n4 a_n3608_1494.t1 28.565
R11448 a_n3608_1494.n2 a_n3608_1494.t0 18.149
R11449 a_n3608_1494.n3 a_n3608_1494.n2 3.726
R11450 a_26179_12829.t5 a_26179_12829.n2 404.877
R11451 a_26179_12829.n1 a_26179_12829.t8 210.902
R11452 a_26179_12829.n3 a_26179_12829.t5 136.943
R11453 a_26179_12829.n2 a_26179_12829.n1 107.801
R11454 a_26179_12829.n1 a_26179_12829.t7 80.333
R11455 a_26179_12829.n2 a_26179_12829.t6 80.333
R11456 a_26179_12829.n0 a_26179_12829.t4 17.4
R11457 a_26179_12829.n0 a_26179_12829.t2 17.4
R11458 a_26179_12829.n4 a_26179_12829.t3 15.032
R11459 a_26179_12829.t0 a_26179_12829.n5 14.282
R11460 a_26179_12829.n5 a_26179_12829.t1 14.282
R11461 a_26179_12829.n5 a_26179_12829.n4 1.65
R11462 a_26179_12829.n3 a_26179_12829.n0 0.672
R11463 a_26179_12829.n4 a_26179_12829.n3 0.665
R11464 a_9561_26713.n6 a_9561_26713.n5 501.28
R11465 a_9561_26713.t10 a_9561_26713.t7 437.233
R11466 a_9561_26713.t9 a_9561_26713.t11 415.315
R11467 a_9561_26713.t8 a_9561_26713.n3 313.873
R11468 a_9561_26713.n5 a_9561_26713.t19 294.986
R11469 a_9561_26713.n2 a_9561_26713.t13 272.288
R11470 a_9561_26713.n6 a_9561_26713.t15 236.01
R11471 a_9561_26713.n9 a_9561_26713.t10 216.627
R11472 a_9561_26713.n7 a_9561_26713.t9 216.111
R11473 a_9561_26713.n8 a_9561_26713.t4 214.686
R11474 a_9561_26713.t7 a_9561_26713.n8 214.686
R11475 a_9561_26713.n1 a_9561_26713.t18 214.335
R11476 a_9561_26713.t11 a_9561_26713.n1 214.335
R11477 a_9561_26713.n4 a_9561_26713.t8 190.152
R11478 a_9561_26713.n4 a_9561_26713.t17 190.152
R11479 a_9561_26713.n2 a_9561_26713.t14 160.666
R11480 a_9561_26713.n3 a_9561_26713.t16 160.666
R11481 a_9561_26713.n7 a_9561_26713.n6 148.428
R11482 a_9561_26713.n5 a_9561_26713.t5 110.859
R11483 a_9561_26713.n3 a_9561_26713.n2 96.129
R11484 a_9561_26713.n8 a_9561_26713.t6 80.333
R11485 a_9561_26713.n1 a_9561_26713.t12 80.333
R11486 a_9561_26713.t15 a_9561_26713.n4 80.333
R11487 a_9561_26713.n0 a_9561_26713.t1 28.57
R11488 a_9561_26713.t0 a_9561_26713.n11 28.565
R11489 a_9561_26713.n11 a_9561_26713.t2 28.565
R11490 a_9561_26713.n0 a_9561_26713.t3 17.638
R11491 a_9561_26713.n10 a_9561_26713.n9 5.375
R11492 a_9561_26713.n9 a_9561_26713.n7 2.923
R11493 a_9561_26713.n11 a_9561_26713.n10 0.69
R11494 a_9561_26713.n10 a_9561_26713.n0 0.6
R11495 a_5504_10602.n2 a_5504_10602.t6 318.922
R11496 a_5504_10602.n1 a_5504_10602.t7 273.935
R11497 a_5504_10602.n1 a_5504_10602.t4 273.935
R11498 a_5504_10602.n2 a_5504_10602.t5 269.116
R11499 a_5504_10602.n4 a_5504_10602.n0 193.227
R11500 a_5504_10602.t6 a_5504_10602.n1 179.142
R11501 a_5504_10602.n3 a_5504_10602.n2 106.999
R11502 a_5504_10602.t3 a_5504_10602.n4 28.568
R11503 a_5504_10602.n0 a_5504_10602.t1 28.565
R11504 a_5504_10602.n0 a_5504_10602.t2 28.565
R11505 a_5504_10602.n3 a_5504_10602.t0 18.149
R11506 a_5504_10602.n4 a_5504_10602.n3 3.726
R11507 a_16558_24431.n1 a_16558_24431.t5 318.922
R11508 a_16558_24431.n0 a_16558_24431.t4 274.739
R11509 a_16558_24431.n0 a_16558_24431.t6 274.739
R11510 a_16558_24431.n1 a_16558_24431.t7 269.116
R11511 a_16558_24431.t5 a_16558_24431.n0 179.946
R11512 a_16558_24431.n2 a_16558_24431.n1 105.178
R11513 a_16558_24431.n3 a_16558_24431.t1 29.444
R11514 a_16558_24431.n4 a_16558_24431.t2 28.565
R11515 a_16558_24431.t3 a_16558_24431.n4 28.565
R11516 a_16558_24431.n2 a_16558_24431.t0 18.145
R11517 a_16558_24431.n3 a_16558_24431.n2 2.878
R11518 a_16558_24431.n4 a_16558_24431.n3 0.764
R11519 a_6343_6961.t8 a_6343_6961.n2 404.877
R11520 a_6343_6961.n1 a_6343_6961.t7 210.902
R11521 a_6343_6961.n3 a_6343_6961.t8 136.943
R11522 a_6343_6961.n2 a_6343_6961.n1 107.801
R11523 a_6343_6961.n1 a_6343_6961.t6 80.333
R11524 a_6343_6961.n2 a_6343_6961.t5 80.333
R11525 a_6343_6961.n0 a_6343_6961.t4 17.4
R11526 a_6343_6961.n0 a_6343_6961.t2 17.4
R11527 a_6343_6961.n4 a_6343_6961.t3 15.032
R11528 a_6343_6961.n5 a_6343_6961.t1 14.282
R11529 a_6343_6961.t0 a_6343_6961.n5 14.282
R11530 a_6343_6961.n5 a_6343_6961.n4 1.65
R11531 a_6343_6961.n3 a_6343_6961.n0 0.672
R11532 a_6343_6961.n4 a_6343_6961.n3 0.665
R11533 a_6607_6378.t7 a_6607_6378.t4 800.071
R11534 a_6607_6378.n3 a_6607_6378.n2 672.951
R11535 a_6607_6378.n1 a_6607_6378.t5 285.109
R11536 a_6607_6378.n2 a_6607_6378.t7 193.602
R11537 a_6607_6378.n1 a_6607_6378.t6 160.666
R11538 a_6607_6378.n2 a_6607_6378.n1 91.507
R11539 a_6607_6378.t3 a_6607_6378.n4 28.57
R11540 a_6607_6378.n0 a_6607_6378.t1 28.565
R11541 a_6607_6378.n0 a_6607_6378.t2 28.565
R11542 a_6607_6378.n4 a_6607_6378.t0 17.638
R11543 a_6607_6378.n3 a_6607_6378.n0 0.69
R11544 a_6607_6378.n4 a_6607_6378.n3 0.6
R11545 a_n3604_11836.n1 a_n3604_11836.t7 318.119
R11546 a_n3604_11836.n1 a_n3604_11836.t4 269.919
R11547 a_n3604_11836.n0 a_n3604_11836.t5 267.256
R11548 a_n3604_11836.n0 a_n3604_11836.t6 267.256
R11549 a_n3604_11836.n4 a_n3604_11836.n3 193.227
R11550 a_n3604_11836.t7 a_n3604_11836.n0 160.666
R11551 a_n3604_11836.n2 a_n3604_11836.n1 106.999
R11552 a_n3604_11836.n3 a_n3604_11836.t1 28.568
R11553 a_n3604_11836.n4 a_n3604_11836.t2 28.565
R11554 a_n3604_11836.t3 a_n3604_11836.n4 28.565
R11555 a_n3604_11836.n2 a_n3604_11836.t0 18.149
R11556 a_n3604_11836.n3 a_n3604_11836.n2 3.726
R11557 a_n2379_11055.t0 a_n2379_11055.t1 379.845
R11558 a_15561_18528.n0 a_15561_18528.t7 214.335
R11559 a_15561_18528.t9 a_15561_18528.n0 214.335
R11560 a_15561_18528.n1 a_15561_18528.t9 143.851
R11561 a_15561_18528.n1 a_15561_18528.t10 135.658
R11562 a_15561_18528.n0 a_15561_18528.t8 80.333
R11563 a_15561_18528.n4 a_15561_18528.t1 28.565
R11564 a_15561_18528.n4 a_15561_18528.t2 28.565
R11565 a_15561_18528.n2 a_15561_18528.t6 28.565
R11566 a_15561_18528.n2 a_15561_18528.t4 28.565
R11567 a_15561_18528.t3 a_15561_18528.n7 28.565
R11568 a_15561_18528.n7 a_15561_18528.t5 28.565
R11569 a_15561_18528.n5 a_15561_18528.t0 9.714
R11570 a_15561_18528.n5 a_15561_18528.n4 1.003
R11571 a_15561_18528.n6 a_15561_18528.n3 0.833
R11572 a_15561_18528.n3 a_15561_18528.n2 0.653
R11573 a_15561_18528.n7 a_15561_18528.n6 0.653
R11574 a_15561_18528.n6 a_15561_18528.n5 0.341
R11575 a_15561_18528.n3 a_15561_18528.n1 0.032
R11576 a_10696_3833.n0 a_10696_3833.t10 214.335
R11577 a_10696_3833.t8 a_10696_3833.n0 214.335
R11578 a_10696_3833.n1 a_10696_3833.t8 143.851
R11579 a_10696_3833.n1 a_10696_3833.t9 135.658
R11580 a_10696_3833.n0 a_10696_3833.t7 80.333
R11581 a_10696_3833.n2 a_10696_3833.t4 28.565
R11582 a_10696_3833.n2 a_10696_3833.t6 28.565
R11583 a_10696_3833.n4 a_10696_3833.t5 28.565
R11584 a_10696_3833.n4 a_10696_3833.t1 28.565
R11585 a_10696_3833.t3 a_10696_3833.n7 28.565
R11586 a_10696_3833.n7 a_10696_3833.t2 28.565
R11587 a_10696_3833.n6 a_10696_3833.t0 9.714
R11588 a_10696_3833.n7 a_10696_3833.n6 1.003
R11589 a_10696_3833.n5 a_10696_3833.n3 0.833
R11590 a_10696_3833.n3 a_10696_3833.n2 0.653
R11591 a_10696_3833.n5 a_10696_3833.n4 0.653
R11592 a_10696_3833.n6 a_10696_3833.n5 0.341
R11593 a_10696_3833.n3 a_10696_3833.n1 0.032
R11594 a_29840_7365.n4 a_29840_7365.t8 214.335
R11595 a_29840_7365.t7 a_29840_7365.n4 214.335
R11596 a_29840_7365.n5 a_29840_7365.t7 143.851
R11597 a_29840_7365.n5 a_29840_7365.t9 135.658
R11598 a_29840_7365.n4 a_29840_7365.t10 80.333
R11599 a_29840_7365.n0 a_29840_7365.t6 28.565
R11600 a_29840_7365.n0 a_29840_7365.t5 28.565
R11601 a_29840_7365.n2 a_29840_7365.t1 28.565
R11602 a_29840_7365.n2 a_29840_7365.t4 28.565
R11603 a_29840_7365.n7 a_29840_7365.t0 28.565
R11604 a_29840_7365.t2 a_29840_7365.n7 28.565
R11605 a_29840_7365.n1 a_29840_7365.t3 9.714
R11606 a_29840_7365.n1 a_29840_7365.n0 1.003
R11607 a_29840_7365.n6 a_29840_7365.n3 0.833
R11608 a_29840_7365.n3 a_29840_7365.n2 0.653
R11609 a_29840_7365.n7 a_29840_7365.n6 0.653
R11610 a_29840_7365.n3 a_29840_7365.n1 0.341
R11611 a_29840_7365.n6 a_29840_7365.n5 0.032
R11612 a_13821_25150.n1 a_13821_25150.t5 318.922
R11613 a_13821_25150.n0 a_13821_25150.t4 273.935
R11614 a_13821_25150.n0 a_13821_25150.t6 273.935
R11615 a_13821_25150.n1 a_13821_25150.t7 269.116
R11616 a_13821_25150.n4 a_13821_25150.n3 193.227
R11617 a_13821_25150.t5 a_13821_25150.n0 179.142
R11618 a_13821_25150.n2 a_13821_25150.n1 106.999
R11619 a_13821_25150.n3 a_13821_25150.t2 28.568
R11620 a_13821_25150.t3 a_13821_25150.n4 28.565
R11621 a_13821_25150.n4 a_13821_25150.t1 28.565
R11622 a_13821_25150.n2 a_13821_25150.t0 18.149
R11623 a_13821_25150.n3 a_13821_25150.n2 3.726
R11624 a_33614_9753.t0 a_33614_9753.t1 17.4
R11625 B[6].n6 B[6].t4 5229.8
R11626 B[6].n12 B[6].n6 692.057
R11627 B[6].n11 B[6].n7 592.056
R11628 B[6].t6 B[6].t22 437.233
R11629 B[6].t10 B[6].t11 437.233
R11630 B[6].t4 B[6].t5 415.315
R11631 B[6].t16 B[6].t17 415.315
R11632 B[6].t21 B[6].n9 313.069
R11633 B[6].n7 B[6].t23 294.986
R11634 B[6].n8 B[6].t18 271.484
R11635 B[6].n4 B[6].t16 220.313
R11636 B[6].n5 B[6].t6 219.163
R11637 B[6].n4 B[6].t10 217.194
R11638 B[6].n1 B[6].t19 214.686
R11639 B[6].t22 B[6].n1 214.686
R11640 B[6].n3 B[6].t3 214.686
R11641 B[6].t11 B[6].n3 214.686
R11642 B[6].n0 B[6].t8 214.335
R11643 B[6].t5 B[6].n0 214.335
R11644 B[6].n2 B[6].t20 214.335
R11645 B[6].t17 B[6].n2 214.335
R11646 B[6].n11 B[6].t15 204.672
R11647 B[6].n10 B[6].t21 190.955
R11648 B[6].n10 B[6].t12 190.955
R11649 B[6].n9 B[6].t1 160.666
R11650 B[6].n8 B[6].t13 160.666
R11651 B[6].n7 B[6].t9 110.859
R11652 B[6].n9 B[6].n8 96.129
R11653 B[6].n0 B[6].t7 80.333
R11654 B[6].n1 B[6].t2 80.333
R11655 B[6].n2 B[6].t0 80.333
R11656 B[6].n3 B[6].t14 80.333
R11657 B[6].t15 B[6].n10 80.333
R11658 B[6].n12 B[6].n11 46.161
R11659 B[6] B[6].n12 33.336
R11660 B[6].n6 B[6].n5 23.931
R11661 B[6].n5 B[6].n4 11.749
R11662 a_38088_8192.t0 a_38088_8192.t1 17.4
R11663 a_36697_14478.n2 a_36697_14478.t6 448.381
R11664 a_36697_14478.n1 a_36697_14478.t7 287.241
R11665 a_36697_14478.n1 a_36697_14478.t4 287.241
R11666 a_36697_14478.n0 a_36697_14478.t5 247.733
R11667 a_36697_14478.n4 a_36697_14478.n3 182.117
R11668 a_36697_14478.t6 a_36697_14478.n1 160.666
R11669 a_36697_14478.n3 a_36697_14478.t1 28.568
R11670 a_36697_14478.n4 a_36697_14478.t2 28.565
R11671 a_36697_14478.t3 a_36697_14478.n4 28.565
R11672 a_36697_14478.n0 a_36697_14478.t0 18.127
R11673 a_36697_14478.n2 a_36697_14478.n0 4.036
R11674 a_36697_14478.n3 a_36697_14478.n2 0.937
R11675 a_5931_9909.n2 a_5931_9909.n0 267.767
R11676 a_5931_9909.n6 a_5931_9909.t6 16.058
R11677 a_5931_9909.n4 a_5931_9909.t3 16.058
R11678 a_5931_9909.n5 a_5931_9909.t8 14.282
R11679 a_5931_9909.n5 a_5931_9909.t7 14.282
R11680 a_5931_9909.n3 a_5931_9909.t5 14.282
R11681 a_5931_9909.n3 a_5931_9909.t4 14.282
R11682 a_5931_9909.n1 a_5931_9909.t11 14.282
R11683 a_5931_9909.n1 a_5931_9909.t0 14.282
R11684 a_5931_9909.n0 a_5931_9909.t9 14.282
R11685 a_5931_9909.n0 a_5931_9909.t10 14.282
R11686 a_5931_9909.n9 a_5931_9909.t1 14.282
R11687 a_5931_9909.t2 a_5931_9909.n9 14.282
R11688 a_5931_9909.n9 a_5931_9909.n8 1.511
R11689 a_5931_9909.n6 a_5931_9909.n5 0.999
R11690 a_5931_9909.n4 a_5931_9909.n3 0.999
R11691 a_5931_9909.n8 a_5931_9909.n2 0.669
R11692 a_5931_9909.n7 a_5931_9909.n6 0.575
R11693 a_5931_9909.n8 a_5931_9909.n7 0.227
R11694 a_5931_9909.n7 a_5931_9909.n4 0.2
R11695 a_5931_9909.n2 a_5931_9909.n1 0.001
R11696 a_29257_17925.t0 a_29257_17925.t1 17.4
R11697 a_7485_6965.t5 a_7485_6965.n3 404.877
R11698 a_7485_6965.n2 a_7485_6965.t8 210.902
R11699 a_7485_6965.n4 a_7485_6965.t5 136.943
R11700 a_7485_6965.n3 a_7485_6965.n2 107.801
R11701 a_7485_6965.n2 a_7485_6965.t7 80.333
R11702 a_7485_6965.n3 a_7485_6965.t6 80.333
R11703 a_7485_6965.n1 a_7485_6965.t0 17.4
R11704 a_7485_6965.n1 a_7485_6965.t2 17.4
R11705 a_7485_6965.t1 a_7485_6965.n5 15.032
R11706 a_7485_6965.n0 a_7485_6965.t4 14.282
R11707 a_7485_6965.n0 a_7485_6965.t3 14.282
R11708 a_7485_6965.n5 a_7485_6965.n0 1.65
R11709 a_7485_6965.n4 a_7485_6965.n1 0.672
R11710 a_7485_6965.n5 a_7485_6965.n4 0.665
R11711 a_7603_6965.n1 a_7603_6965.t0 14.282
R11712 a_7603_6965.n1 a_7603_6965.t4 14.282
R11713 a_7603_6965.n0 a_7603_6965.t3 14.282
R11714 a_7603_6965.n0 a_7603_6965.t5 14.282
R11715 a_7603_6965.t2 a_7603_6965.n3 14.282
R11716 a_7603_6965.n3 a_7603_6965.t1 14.282
R11717 a_7603_6965.n2 a_7603_6965.n0 2.546
R11718 a_7603_6965.n3 a_7603_6965.n2 2.367
R11719 a_7603_6965.n2 a_7603_6965.n1 0.001
R11720 a_29774_14889.n2 a_29774_14889.t7 214.335
R11721 a_29774_14889.t9 a_29774_14889.n2 214.335
R11722 a_29774_14889.n3 a_29774_14889.t9 143.851
R11723 a_29774_14889.n3 a_29774_14889.t8 135.658
R11724 a_29774_14889.n2 a_29774_14889.t10 80.333
R11725 a_29774_14889.n4 a_29774_14889.t0 28.565
R11726 a_29774_14889.n4 a_29774_14889.t1 28.565
R11727 a_29774_14889.n0 a_29774_14889.t5 28.565
R11728 a_29774_14889.n0 a_29774_14889.t6 28.565
R11729 a_29774_14889.t2 a_29774_14889.n7 28.565
R11730 a_29774_14889.n7 a_29774_14889.t4 28.565
R11731 a_29774_14889.n1 a_29774_14889.t3 9.714
R11732 a_29774_14889.n1 a_29774_14889.n0 1.003
R11733 a_29774_14889.n6 a_29774_14889.n5 0.833
R11734 a_29774_14889.n5 a_29774_14889.n4 0.653
R11735 a_29774_14889.n7 a_29774_14889.n6 0.653
R11736 a_29774_14889.n6 a_29774_14889.n1 0.341
R11737 a_29774_14889.n5 a_29774_14889.n3 0.032
R11738 a_30364_14452.n3 a_30364_14452.n2 2062.97
R11739 a_30364_14452.n2 a_30364_14452.t4 989.744
R11740 a_30364_14452.n2 a_30364_14452.t6 408.806
R11741 a_30364_14452.n1 a_30364_14452.t5 287.241
R11742 a_30364_14452.n1 a_30364_14452.t7 287.241
R11743 a_30364_14452.n4 a_30364_14452.n0 192.754
R11744 a_30364_14452.t4 a_30364_14452.n1 160.666
R11745 a_30364_14452.t3 a_30364_14452.n4 28.568
R11746 a_30364_14452.n0 a_30364_14452.t1 28.565
R11747 a_30364_14452.n0 a_30364_14452.t2 28.565
R11748 a_30364_14452.n3 a_30364_14452.t0 19.164
R11749 a_30364_14452.n4 a_30364_14452.n3 1.101
R11750 a_21381_3396.t0 a_21381_3396.t1 17.4
R11751 a_36751_16737.n0 a_36751_16737.t1 14.282
R11752 a_36751_16737.t0 a_36751_16737.n0 14.282
R11753 a_36751_16737.n0 a_36751_16737.n1 258.161
R11754 a_36751_16737.n1 a_36751_16737.t7 14.283
R11755 a_36751_16737.n1 a_36751_16737.n5 0.852
R11756 a_36751_16737.n5 a_36751_16737.n6 4.366
R11757 a_36751_16737.n6 a_36751_16737.n7 258.161
R11758 a_36751_16737.n7 a_36751_16737.t3 14.282
R11759 a_36751_16737.n7 a_36751_16737.t5 14.282
R11760 a_36751_16737.n6 a_36751_16737.t4 14.283
R11761 a_36751_16737.n5 a_36751_16737.n4 73.514
R11762 a_36751_16737.n4 a_36751_16737.t11 1551.5
R11763 a_36751_16737.t11 a_36751_16737.n3 656.576
R11764 a_36751_16737.n3 a_36751_16737.t2 8.7
R11765 a_36751_16737.n3 a_36751_16737.t6 8.7
R11766 a_36751_16737.n4 a_36751_16737.t10 224.129
R11767 a_36751_16737.t10 a_36751_16737.n2 207.225
R11768 a_36751_16737.n2 a_36751_16737.t9 207.225
R11769 a_36751_16737.n2 a_36751_16737.t8 80.333
R11770 a_38084_17682.t0 a_38084_17682.t1 17.4
R11771 a_11286_3396.t4 a_11286_3396.t6 574.43
R11772 a_11286_3396.n0 a_11286_3396.t7 285.109
R11773 a_11286_3396.n2 a_11286_3396.n1 197.217
R11774 a_11286_3396.n4 a_11286_3396.n3 192.754
R11775 a_11286_3396.n0 a_11286_3396.t5 160.666
R11776 a_11286_3396.n1 a_11286_3396.t4 160.666
R11777 a_11286_3396.n1 a_11286_3396.n0 114.829
R11778 a_11286_3396.n3 a_11286_3396.t1 28.568
R11779 a_11286_3396.t3 a_11286_3396.n4 28.565
R11780 a_11286_3396.n4 a_11286_3396.t2 28.565
R11781 a_11286_3396.n2 a_11286_3396.t0 18.838
R11782 a_11286_3396.n3 a_11286_3396.n2 1.129
R11783 a_13012_6959.n1 a_13012_6959.t0 14.282
R11784 a_13012_6959.n1 a_13012_6959.t3 14.282
R11785 a_13012_6959.n0 a_13012_6959.t4 14.282
R11786 a_13012_6959.n0 a_13012_6959.t5 14.282
R11787 a_13012_6959.t2 a_13012_6959.n3 14.282
R11788 a_13012_6959.n3 a_13012_6959.t1 14.282
R11789 a_13012_6959.n2 a_13012_6959.n0 2.546
R11790 a_13012_6959.n3 a_13012_6959.n2 2.367
R11791 a_13012_6959.n2 a_13012_6959.n1 0.001
R11792 a_36697_1856.n2 a_36697_1856.t4 448.381
R11793 a_36697_1856.n1 a_36697_1856.t6 287.241
R11794 a_36697_1856.n1 a_36697_1856.t7 287.241
R11795 a_36697_1856.n0 a_36697_1856.t5 247.733
R11796 a_36697_1856.n4 a_36697_1856.n3 182.117
R11797 a_36697_1856.t4 a_36697_1856.n1 160.666
R11798 a_36697_1856.n3 a_36697_1856.t2 28.568
R11799 a_36697_1856.t3 a_36697_1856.n4 28.565
R11800 a_36697_1856.n4 a_36697_1856.t1 28.565
R11801 a_36697_1856.n0 a_36697_1856.t0 18.127
R11802 a_36697_1856.n2 a_36697_1856.n0 4.036
R11803 a_36697_1856.n3 a_36697_1856.n2 0.937
R11804 a_30011_14252.t0 a_30011_14252.t1 17.4
R11805 a_24562_12520.t7 a_24562_12520.t4 800.071
R11806 a_24562_12520.n3 a_24562_12520.n2 659.097
R11807 a_24562_12520.n1 a_24562_12520.t6 285.109
R11808 a_24562_12520.n2 a_24562_12520.t7 193.602
R11809 a_24562_12520.n4 a_24562_12520.n0 192.754
R11810 a_24562_12520.n1 a_24562_12520.t5 160.666
R11811 a_24562_12520.n2 a_24562_12520.n1 91.507
R11812 a_24562_12520.t0 a_24562_12520.n4 28.568
R11813 a_24562_12520.n0 a_24562_12520.t3 28.565
R11814 a_24562_12520.n0 a_24562_12520.t1 28.565
R11815 a_24562_12520.n3 a_24562_12520.t2 19.061
R11816 a_24562_12520.n4 a_24562_12520.n3 1.005
R11817 a_19004_24158.n0 a_19004_24158.t10 214.335
R11818 a_19004_24158.t8 a_19004_24158.n0 214.335
R11819 a_19004_24158.n1 a_19004_24158.t8 143.851
R11820 a_19004_24158.n1 a_19004_24158.t7 135.658
R11821 a_19004_24158.n0 a_19004_24158.t9 80.333
R11822 a_19004_24158.n2 a_19004_24158.t5 28.565
R11823 a_19004_24158.n2 a_19004_24158.t6 28.565
R11824 a_19004_24158.n4 a_19004_24158.t4 28.565
R11825 a_19004_24158.n4 a_19004_24158.t2 28.565
R11826 a_19004_24158.t3 a_19004_24158.n7 28.565
R11827 a_19004_24158.n7 a_19004_24158.t1 28.565
R11828 a_19004_24158.n6 a_19004_24158.t0 9.714
R11829 a_19004_24158.n7 a_19004_24158.n6 1.003
R11830 a_19004_24158.n5 a_19004_24158.n3 0.833
R11831 a_19004_24158.n3 a_19004_24158.n2 0.653
R11832 a_19004_24158.n5 a_19004_24158.n4 0.653
R11833 a_19004_24158.n6 a_19004_24158.n5 0.341
R11834 a_19004_24158.n3 a_19004_24158.n1 0.032
R11835 a_19594_23721.t5 a_19594_23721.t4 574.43
R11836 a_19594_23721.n0 a_19594_23721.t7 285.109
R11837 a_19594_23721.n2 a_19594_23721.n1 197.217
R11838 a_19594_23721.n4 a_19594_23721.n3 192.754
R11839 a_19594_23721.n0 a_19594_23721.t6 160.666
R11840 a_19594_23721.n1 a_19594_23721.t5 160.666
R11841 a_19594_23721.n1 a_19594_23721.n0 114.829
R11842 a_19594_23721.n3 a_19594_23721.t1 28.568
R11843 a_19594_23721.n4 a_19594_23721.t2 28.565
R11844 a_19594_23721.t3 a_19594_23721.n4 28.565
R11845 a_19594_23721.n2 a_19594_23721.t0 18.838
R11846 a_19594_23721.n3 a_19594_23721.n2 1.129
R11847 a_28603_20140.n0 a_28603_20140.t7 214.335
R11848 a_28603_20140.t9 a_28603_20140.n0 214.335
R11849 a_28603_20140.n1 a_28603_20140.t9 143.851
R11850 a_28603_20140.n1 a_28603_20140.t10 135.658
R11851 a_28603_20140.n0 a_28603_20140.t8 80.333
R11852 a_28603_20140.n2 a_28603_20140.t4 28.565
R11853 a_28603_20140.n2 a_28603_20140.t5 28.565
R11854 a_28603_20140.n4 a_28603_20140.t6 28.565
R11855 a_28603_20140.n4 a_28603_20140.t1 28.565
R11856 a_28603_20140.t2 a_28603_20140.n7 28.565
R11857 a_28603_20140.n7 a_28603_20140.t0 28.565
R11858 a_28603_20140.n3 a_28603_20140.t3 9.714
R11859 a_28603_20140.n3 a_28603_20140.n2 1.003
R11860 a_28603_20140.n6 a_28603_20140.n5 0.833
R11861 a_28603_20140.n5 a_28603_20140.n4 0.653
R11862 a_28603_20140.n7 a_28603_20140.n6 0.653
R11863 a_28603_20140.n5 a_28603_20140.n3 0.341
R11864 a_28603_20140.n6 a_28603_20140.n1 0.032
R11865 a_n3606_13905.n1 a_n3606_13905.t6 318.119
R11866 a_n3606_13905.n1 a_n3606_13905.t5 269.919
R11867 a_n3606_13905.n0 a_n3606_13905.t7 267.256
R11868 a_n3606_13905.n0 a_n3606_13905.t4 267.256
R11869 a_n3606_13905.n4 a_n3606_13905.n3 193.227
R11870 a_n3606_13905.t6 a_n3606_13905.n0 160.666
R11871 a_n3606_13905.n2 a_n3606_13905.n1 106.999
R11872 a_n3606_13905.n3 a_n3606_13905.t2 28.568
R11873 a_n3606_13905.t3 a_n3606_13905.n4 28.565
R11874 a_n3606_13905.n4 a_n3606_13905.t1 28.565
R11875 a_n3606_13905.n2 a_n3606_13905.t0 18.149
R11876 a_n3606_13905.n3 a_n3606_13905.n2 3.726
R11877 a_20849_18121.t0 a_20849_18121.t1 17.4
R11878 a_33614_6258.t0 a_33614_6258.t1 17.4
R11879 a_20133_21659.t4 a_20133_21659.t5 800.071
R11880 a_20133_21659.n3 a_20133_21659.n2 659.095
R11881 a_20133_21659.n1 a_20133_21659.t6 285.109
R11882 a_20133_21659.n2 a_20133_21659.t4 193.602
R11883 a_20133_21659.n4 a_20133_21659.n0 192.754
R11884 a_20133_21659.n1 a_20133_21659.t7 160.666
R11885 a_20133_21659.n2 a_20133_21659.n1 91.507
R11886 a_20133_21659.t3 a_20133_21659.n4 28.568
R11887 a_20133_21659.n0 a_20133_21659.t1 28.565
R11888 a_20133_21659.n0 a_20133_21659.t2 28.565
R11889 a_20133_21659.n3 a_20133_21659.t0 19.063
R11890 a_20133_21659.n4 a_20133_21659.n3 1.005
R11891 a_22090_20137.n0 a_22090_20137.t10 214.335
R11892 a_22090_20137.t8 a_22090_20137.n0 214.335
R11893 a_22090_20137.n1 a_22090_20137.t8 143.851
R11894 a_22090_20137.n1 a_22090_20137.t9 135.658
R11895 a_22090_20137.n0 a_22090_20137.t7 80.333
R11896 a_22090_20137.n2 a_22090_20137.t5 28.565
R11897 a_22090_20137.n2 a_22090_20137.t6 28.565
R11898 a_22090_20137.n4 a_22090_20137.t1 28.565
R11899 a_22090_20137.n4 a_22090_20137.t4 28.565
R11900 a_22090_20137.t3 a_22090_20137.n7 28.565
R11901 a_22090_20137.n7 a_22090_20137.t2 28.565
R11902 a_22090_20137.n6 a_22090_20137.t0 9.714
R11903 a_22090_20137.n7 a_22090_20137.n6 1.003
R11904 a_22090_20137.n5 a_22090_20137.n3 0.833
R11905 a_22090_20137.n3 a_22090_20137.n2 0.653
R11906 a_22090_20137.n5 a_22090_20137.n4 0.653
R11907 a_22090_20137.n6 a_22090_20137.n5 0.341
R11908 a_22090_20137.n3 a_22090_20137.n1 0.032
R11909 a_4153_9615.n4 a_4153_9615.t8 214.335
R11910 a_4153_9615.t10 a_4153_9615.n4 214.335
R11911 a_4153_9615.n5 a_4153_9615.t10 143.851
R11912 a_4153_9615.n5 a_4153_9615.t9 135.658
R11913 a_4153_9615.n4 a_4153_9615.t7 80.333
R11914 a_4153_9615.n0 a_4153_9615.t3 28.565
R11915 a_4153_9615.n0 a_4153_9615.t4 28.565
R11916 a_4153_9615.n2 a_4153_9615.t6 28.565
R11917 a_4153_9615.n2 a_4153_9615.t5 28.565
R11918 a_4153_9615.n7 a_4153_9615.t1 28.565
R11919 a_4153_9615.t0 a_4153_9615.n7 28.565
R11920 a_4153_9615.n1 a_4153_9615.t2 9.714
R11921 a_4153_9615.n1 a_4153_9615.n0 1.003
R11922 a_4153_9615.n6 a_4153_9615.n3 0.833
R11923 a_4153_9615.n3 a_4153_9615.n2 0.653
R11924 a_4153_9615.n7 a_4153_9615.n6 0.653
R11925 a_4153_9615.n3 a_4153_9615.n1 0.341
R11926 a_4153_9615.n6 a_4153_9615.n5 0.032
R11927 a_4743_9178.t5 a_4743_9178.t4 574.43
R11928 a_4743_9178.n0 a_4743_9178.t7 285.109
R11929 a_4743_9178.n2 a_4743_9178.n1 197.217
R11930 a_4743_9178.n4 a_4743_9178.n3 192.754
R11931 a_4743_9178.n0 a_4743_9178.t6 160.666
R11932 a_4743_9178.n1 a_4743_9178.t5 160.666
R11933 a_4743_9178.n1 a_4743_9178.n0 114.829
R11934 a_4743_9178.n3 a_4743_9178.t2 28.568
R11935 a_4743_9178.t3 a_4743_9178.n4 28.565
R11936 a_4743_9178.n4 a_4743_9178.t1 28.565
R11937 a_4743_9178.n2 a_4743_9178.t0 18.838
R11938 a_4743_9178.n3 a_4743_9178.n2 1.129
R11939 a_19541_4102.n1 a_19541_4102.t7 318.922
R11940 a_19541_4102.n0 a_19541_4102.t4 274.739
R11941 a_19541_4102.n0 a_19541_4102.t5 274.739
R11942 a_19541_4102.n1 a_19541_4102.t6 269.116
R11943 a_19541_4102.t7 a_19541_4102.n0 179.946
R11944 a_19541_4102.n2 a_19541_4102.n1 107.263
R11945 a_19541_4102.t3 a_19541_4102.n4 29.444
R11946 a_19541_4102.n3 a_19541_4102.t1 28.565
R11947 a_19541_4102.n3 a_19541_4102.t2 28.565
R11948 a_19541_4102.n2 a_19541_4102.t0 18.145
R11949 a_19541_4102.n4 a_19541_4102.n2 2.878
R11950 a_19541_4102.n4 a_19541_4102.n3 0.764
R11951 a_19129_4128.n0 a_19129_4128.t7 14.282
R11952 a_19129_4128.t3 a_19129_4128.n0 14.282
R11953 a_19129_4128.n0 a_19129_4128.n9 0.999
R11954 a_19129_4128.n9 a_19129_4128.n6 0.575
R11955 a_19129_4128.n6 a_19129_4128.n8 0.2
R11956 a_19129_4128.n8 a_19129_4128.t5 16.058
R11957 a_19129_4128.n8 a_19129_4128.n7 0.999
R11958 a_19129_4128.n7 a_19129_4128.t6 14.282
R11959 a_19129_4128.n7 a_19129_4128.t4 14.282
R11960 a_19129_4128.n9 a_19129_4128.t8 16.058
R11961 a_19129_4128.n6 a_19129_4128.n4 0.227
R11962 a_19129_4128.n4 a_19129_4128.n5 1.511
R11963 a_19129_4128.n5 a_19129_4128.t1 14.282
R11964 a_19129_4128.n5 a_19129_4128.t2 14.282
R11965 a_19129_4128.n4 a_19129_4128.n1 0.669
R11966 a_19129_4128.n1 a_19129_4128.n2 0.001
R11967 a_19129_4128.n1 a_19129_4128.n3 267.767
R11968 a_19129_4128.n3 a_19129_4128.t9 14.282
R11969 a_19129_4128.n3 a_19129_4128.t10 14.282
R11970 a_19129_4128.n2 a_19129_4128.t0 14.282
R11971 a_19129_4128.n2 a_19129_4128.t11 14.282
R11972 a_29252_19529.t0 a_29252_19529.t1 17.4
R11973 a_29650_24430.n1 a_29650_24430.t6 318.922
R11974 a_29650_24430.n0 a_29650_24430.t5 274.739
R11975 a_29650_24430.n0 a_29650_24430.t7 274.739
R11976 a_29650_24430.n1 a_29650_24430.t4 269.116
R11977 a_29650_24430.t6 a_29650_24430.n0 179.946
R11978 a_29650_24430.n2 a_29650_24430.n1 105.178
R11979 a_29650_24430.n3 a_29650_24430.t2 29.444
R11980 a_29650_24430.t3 a_29650_24430.n4 28.565
R11981 a_29650_24430.n4 a_29650_24430.t1 28.565
R11982 a_29650_24430.n2 a_29650_24430.t0 18.145
R11983 a_29650_24430.n3 a_29650_24430.n2 2.878
R11984 a_29650_24430.n4 a_29650_24430.n3 0.764
R11985 a_9012_21786.n0 a_9012_21786.t9 214.335
R11986 a_9012_21786.t8 a_9012_21786.n0 214.335
R11987 a_9012_21786.n1 a_9012_21786.t8 143.851
R11988 a_9012_21786.n1 a_9012_21786.t7 135.658
R11989 a_9012_21786.n0 a_9012_21786.t10 80.333
R11990 a_9012_21786.n4 a_9012_21786.t5 28.565
R11991 a_9012_21786.n4 a_9012_21786.t6 28.565
R11992 a_9012_21786.n2 a_9012_21786.t2 28.565
R11993 a_9012_21786.n2 a_9012_21786.t3 28.565
R11994 a_9012_21786.t0 a_9012_21786.n7 28.565
R11995 a_9012_21786.n7 a_9012_21786.t1 28.565
R11996 a_9012_21786.n5 a_9012_21786.t4 9.714
R11997 a_9012_21786.n5 a_9012_21786.n4 1.003
R11998 a_9012_21786.n6 a_9012_21786.n3 0.833
R11999 a_9012_21786.n3 a_9012_21786.n2 0.653
R12000 a_9012_21786.n7 a_9012_21786.n6 0.653
R12001 a_9012_21786.n6 a_9012_21786.n5 0.341
R12002 a_9012_21786.n3 a_9012_21786.n1 0.032
R12003 a_7041_21658.t7 a_7041_21658.t5 800.071
R12004 a_7041_21658.n2 a_7041_21658.n1 659.095
R12005 a_7041_21658.n0 a_7041_21658.t4 285.109
R12006 a_7041_21658.n1 a_7041_21658.t7 193.602
R12007 a_7041_21658.n4 a_7041_21658.n3 192.754
R12008 a_7041_21658.n0 a_7041_21658.t6 160.666
R12009 a_7041_21658.n1 a_7041_21658.n0 91.507
R12010 a_7041_21658.n3 a_7041_21658.t2 28.568
R12011 a_7041_21658.t3 a_7041_21658.n4 28.565
R12012 a_7041_21658.n4 a_7041_21658.t1 28.565
R12013 a_7041_21658.n2 a_7041_21658.t0 19.063
R12014 a_7041_21658.n3 a_7041_21658.n2 1.005
R12015 a_10938_4800.t0 a_10938_4800.t1 17.4
R12016 a_n3113_2781.t0 a_n3113_2781.n0 14.282
R12017 a_n3113_2781.n0 a_n3113_2781.t7 14.282
R12018 a_n3113_2781.n0 a_n3113_2781.n16 90.436
R12019 a_n3113_2781.n16 a_n3113_2781.n2 74.302
R12020 a_n3113_2781.n2 a_n3113_2781.n4 50.575
R12021 a_n3113_2781.n4 a_n3113_2781.n5 110.084
R12022 a_n3113_2781.n16 a_n3113_2781.n6 691.471
R12023 a_n3113_2781.n6 a_n3113_2781.n8 16.411
R12024 a_n3113_2781.n8 a_n3113_2781.t9 198.921
R12025 a_n3113_2781.t9 a_n3113_2781.t22 415.315
R12026 a_n3113_2781.t22 a_n3113_2781.n15 214.335
R12027 a_n3113_2781.n15 a_n3113_2781.t21 80.333
R12028 a_n3113_2781.n15 a_n3113_2781.t19 214.335
R12029 a_n3113_2781.n8 a_n3113_2781.n14 861.987
R12030 a_n3113_2781.n14 a_n3113_2781.n9 560.726
R12031 a_n3113_2781.n14 a_n3113_2781.n13 65.07
R12032 a_n3113_2781.n13 a_n3113_2781.n12 6.615
R12033 a_n3113_2781.n12 a_n3113_2781.t14 93.989
R12034 a_n3113_2781.n12 a_n3113_2781.t12 198.043
R12035 a_n3113_2781.n13 a_n3113_2781.n11 97.816
R12036 a_n3113_2781.n11 a_n3113_2781.t11 80.333
R12037 a_n3113_2781.n11 a_n3113_2781.t20 394.151
R12038 a_n3113_2781.t20 a_n3113_2781.n10 269.523
R12039 a_n3113_2781.n10 a_n3113_2781.t18 160.666
R12040 a_n3113_2781.n10 a_n3113_2781.t17 269.523
R12041 a_n3113_2781.n9 a_n3113_2781.t10 294.653
R12042 a_n3113_2781.n9 a_n3113_2781.t8 111.663
R12043 a_n3113_2781.n6 a_n3113_2781.t23 217.716
R12044 a_n3113_2781.t23 a_n3113_2781.t15 415.315
R12045 a_n3113_2781.t15 a_n3113_2781.n7 214.335
R12046 a_n3113_2781.n7 a_n3113_2781.t13 80.333
R12047 a_n3113_2781.n7 a_n3113_2781.t16 214.335
R12048 a_n3113_2781.n5 a_n3113_2781.t4 14.282
R12049 a_n3113_2781.n5 a_n3113_2781.t6 14.282
R12050 a_n3113_2781.n4 a_n3113_2781.n3 157.665
R12051 a_n3113_2781.n3 a_n3113_2781.t1 8.7
R12052 a_n3113_2781.n3 a_n3113_2781.t3 8.7
R12053 a_n3113_2781.n2 a_n3113_2781.n1 90.416
R12054 a_n3113_2781.n1 a_n3113_2781.t2 14.282
R12055 a_n3113_2781.n1 a_n3113_2781.t5 14.282
R12056 a_14373_18822.n1 a_14373_18822.t7 318.922
R12057 a_14373_18822.n0 a_14373_18822.t6 273.935
R12058 a_14373_18822.n0 a_14373_18822.t5 273.935
R12059 a_14373_18822.n1 a_14373_18822.t4 269.116
R12060 a_14373_18822.n4 a_14373_18822.n3 193.227
R12061 a_14373_18822.t7 a_14373_18822.n0 179.142
R12062 a_14373_18822.n2 a_14373_18822.n1 106.999
R12063 a_14373_18822.n3 a_14373_18822.t2 28.568
R12064 a_14373_18822.n4 a_14373_18822.t1 28.565
R12065 a_14373_18822.t3 a_14373_18822.n4 28.565
R12066 a_14373_18822.n2 a_14373_18822.t0 18.149
R12067 a_14373_18822.n3 a_14373_18822.n2 3.726
R12068 Y[2].n1 Y[2].n0 185.55
R12069 Y[2].n1 Y[2].t1 28.568
R12070 Y[2].n0 Y[2].t2 28.565
R12071 Y[2].n0 Y[2].t3 28.565
R12072 Y[2].n2 Y[2].t0 20.393
R12073 Y[2].n2 Y[2].n1 1.834
R12074 Y[2].n3 Y[2].n2 1.049
R12075 Y[2] Y[2].n3 0.052
R12076 Y[2].n3 Y[2] 0.046
R12077 a_25324_4822.n1 a_25324_4822.t6 318.922
R12078 a_25324_4822.n0 a_25324_4822.t4 273.935
R12079 a_25324_4822.n0 a_25324_4822.t7 273.935
R12080 a_25324_4822.n1 a_25324_4822.t5 269.116
R12081 a_25324_4822.n4 a_25324_4822.n3 193.227
R12082 a_25324_4822.t6 a_25324_4822.n0 179.142
R12083 a_25324_4822.n2 a_25324_4822.n1 106.999
R12084 a_25324_4822.n3 a_25324_4822.t2 28.568
R12085 a_25324_4822.t3 a_25324_4822.n4 28.565
R12086 a_25324_4822.n4 a_25324_4822.t1 28.565
R12087 a_25324_4822.n2 a_25324_4822.t0 18.149
R12088 a_25324_4822.n3 a_25324_4822.n2 3.726
R12089 a_20900_23720.t0 a_20900_23720.t1 380.209
R12090 a_28024_26705.t4 a_28024_26705.t7 800.071
R12091 a_28024_26705.n3 a_28024_26705.n2 672.951
R12092 a_28024_26705.n1 a_28024_26705.t6 285.109
R12093 a_28024_26705.n2 a_28024_26705.t4 193.602
R12094 a_28024_26705.n1 a_28024_26705.t5 160.666
R12095 a_28024_26705.n2 a_28024_26705.n1 91.507
R12096 a_28024_26705.t3 a_28024_26705.n4 28.57
R12097 a_28024_26705.n0 a_28024_26705.t1 28.565
R12098 a_28024_26705.n0 a_28024_26705.t2 28.565
R12099 a_28024_26705.n4 a_28024_26705.t0 17.638
R12100 a_28024_26705.n3 a_28024_26705.n0 0.69
R12101 a_28024_26705.n4 a_28024_26705.n3 0.6
R12102 a_12053_10690.n2 a_12053_10690.t7 318.922
R12103 a_12053_10690.n1 a_12053_10690.t4 273.935
R12104 a_12053_10690.n1 a_12053_10690.t6 273.935
R12105 a_12053_10690.n2 a_12053_10690.t5 269.116
R12106 a_12053_10690.n4 a_12053_10690.n0 193.227
R12107 a_12053_10690.t7 a_12053_10690.n1 179.142
R12108 a_12053_10690.n3 a_12053_10690.n2 106.999
R12109 a_12053_10690.t3 a_12053_10690.n4 28.568
R12110 a_12053_10690.n0 a_12053_10690.t1 28.565
R12111 a_12053_10690.n0 a_12053_10690.t2 28.565
R12112 a_12053_10690.n3 a_12053_10690.t0 18.149
R12113 a_12053_10690.n4 a_12053_10690.n3 3.726
R12114 a_22680_24452.t3 a_22680_24452.n7 16.058
R12115 a_22680_24452.n7 a_22680_24452.n5 0.575
R12116 a_22680_24452.n5 a_22680_24452.n9 0.2
R12117 a_22680_24452.n9 a_22680_24452.t9 16.058
R12118 a_22680_24452.n9 a_22680_24452.n8 0.999
R12119 a_22680_24452.n8 a_22680_24452.t11 14.282
R12120 a_22680_24452.n8 a_22680_24452.t10 14.282
R12121 a_22680_24452.n7 a_22680_24452.n6 0.999
R12122 a_22680_24452.n6 a_22680_24452.t4 14.282
R12123 a_22680_24452.n6 a_22680_24452.t5 14.282
R12124 a_22680_24452.n5 a_22680_24452.n3 0.227
R12125 a_22680_24452.n3 a_22680_24452.n4 1.511
R12126 a_22680_24452.n4 a_22680_24452.t6 14.282
R12127 a_22680_24452.n4 a_22680_24452.t7 14.282
R12128 a_22680_24452.n3 a_22680_24452.n0 0.669
R12129 a_22680_24452.n0 a_22680_24452.n1 0.001
R12130 a_22680_24452.n0 a_22680_24452.n2 267.767
R12131 a_22680_24452.n2 a_22680_24452.t1 14.282
R12132 a_22680_24452.n2 a_22680_24452.t0 14.282
R12133 a_22680_24452.n1 a_22680_24452.t8 14.282
R12134 a_22680_24452.n1 a_22680_24452.t2 14.282
R12135 a_26443_12246.t4 a_26443_12246.t6 800.071
R12136 a_26443_12246.n3 a_26443_12246.n2 672.951
R12137 a_26443_12246.n1 a_26443_12246.t7 285.109
R12138 a_26443_12246.n2 a_26443_12246.t4 193.602
R12139 a_26443_12246.n1 a_26443_12246.t5 160.666
R12140 a_26443_12246.n2 a_26443_12246.n1 91.507
R12141 a_26443_12246.t3 a_26443_12246.n4 28.57
R12142 a_26443_12246.n0 a_26443_12246.t1 28.565
R12143 a_26443_12246.n0 a_26443_12246.t2 28.565
R12144 a_26443_12246.n4 a_26443_12246.t0 17.638
R12145 a_26443_12246.n3 a_26443_12246.n0 0.69
R12146 a_26443_12246.n4 a_26443_12246.n3 0.6
R12147 a_14790_9971.n1 a_14790_9971.t6 318.922
R12148 a_14790_9971.n0 a_14790_9971.t5 274.739
R12149 a_14790_9971.n0 a_14790_9971.t7 274.739
R12150 a_14790_9971.n1 a_14790_9971.t4 269.116
R12151 a_14790_9971.t6 a_14790_9971.n0 179.946
R12152 a_14790_9971.n2 a_14790_9971.n1 105.178
R12153 a_14790_9971.n3 a_14790_9971.t1 29.444
R12154 a_14790_9971.n4 a_14790_9971.t2 28.565
R12155 a_14790_9971.t3 a_14790_9971.n4 28.565
R12156 a_14790_9971.n2 a_14790_9971.t0 18.145
R12157 a_14790_9971.n3 a_14790_9971.n2 2.878
R12158 a_14790_9971.n4 a_14790_9971.n3 0.764
R12159 a_27222_4822.n1 a_27222_4822.t6 318.922
R12160 a_27222_4822.n0 a_27222_4822.t7 273.935
R12161 a_27222_4822.n0 a_27222_4822.t4 273.935
R12162 a_27222_4822.n1 a_27222_4822.t5 269.116
R12163 a_27222_4822.n4 a_27222_4822.n3 193.227
R12164 a_27222_4822.t6 a_27222_4822.n0 179.142
R12165 a_27222_4822.n2 a_27222_4822.n1 106.999
R12166 a_27222_4822.n3 a_27222_4822.t3 28.568
R12167 a_27222_4822.t0 a_27222_4822.n4 28.565
R12168 a_27222_4822.n4 a_27222_4822.t1 28.565
R12169 a_27222_4822.n2 a_27222_4822.t2 18.149
R12170 a_27222_4822.n3 a_27222_4822.n2 3.726
R12171 a_27767_4129.n2 a_27767_4129.t10 989.744
R12172 a_27767_4129.n2 a_27767_4129.t9 408.806
R12173 a_27767_4129.n1 a_27767_4129.t11 287.241
R12174 a_27767_4129.n1 a_27767_4129.t8 287.241
R12175 a_27767_4129.n3 a_27767_4129.n2 224.559
R12176 a_27767_4129.t10 a_27767_4129.n1 160.666
R12177 a_27767_4129.n6 a_27767_4129.n4 157.665
R12178 a_27767_4129.n6 a_27767_4129.n5 122.999
R12179 a_27767_4129.n3 a_27767_4129.n0 90.436
R12180 a_27767_4129.n8 a_27767_4129.n7 90.416
R12181 a_27767_4129.n7 a_27767_4129.n3 74.302
R12182 a_27767_4129.n7 a_27767_4129.n6 50.575
R12183 a_27767_4129.n0 a_27767_4129.t1 14.282
R12184 a_27767_4129.n0 a_27767_4129.t0 14.282
R12185 a_27767_4129.n5 a_27767_4129.t6 14.282
R12186 a_27767_4129.n5 a_27767_4129.t5 14.282
R12187 a_27767_4129.t2 a_27767_4129.n8 14.282
R12188 a_27767_4129.n8 a_27767_4129.t7 14.282
R12189 a_27767_4129.n4 a_27767_4129.t3 8.7
R12190 a_27767_4129.n4 a_27767_4129.t4 8.7
R12191 a_19009_25762.n2 a_19009_25762.t10 214.335
R12192 a_19009_25762.t8 a_19009_25762.n2 214.335
R12193 a_19009_25762.n3 a_19009_25762.t8 143.851
R12194 a_19009_25762.n3 a_19009_25762.t7 135.658
R12195 a_19009_25762.n2 a_19009_25762.t9 80.333
R12196 a_19009_25762.n4 a_19009_25762.t0 28.565
R12197 a_19009_25762.n4 a_19009_25762.t1 28.565
R12198 a_19009_25762.n0 a_19009_25762.t6 28.565
R12199 a_19009_25762.n0 a_19009_25762.t4 28.565
R12200 a_19009_25762.t2 a_19009_25762.n7 28.565
R12201 a_19009_25762.n7 a_19009_25762.t5 28.565
R12202 a_19009_25762.n1 a_19009_25762.t3 9.714
R12203 a_19009_25762.n1 a_19009_25762.n0 1.003
R12204 a_19009_25762.n6 a_19009_25762.n5 0.833
R12205 a_19009_25762.n5 a_19009_25762.n4 0.653
R12206 a_19009_25762.n7 a_19009_25762.n6 0.653
R12207 a_19009_25762.n6 a_19009_25762.n1 0.341
R12208 a_19009_25762.n5 a_19009_25762.n3 0.032
R12209 a_19599_25325.t5 a_19599_25325.t4 574.43
R12210 a_19599_25325.n0 a_19599_25325.t7 285.109
R12211 a_19599_25325.n2 a_19599_25325.n1 211.136
R12212 a_19599_25325.n4 a_19599_25325.n3 192.754
R12213 a_19599_25325.n0 a_19599_25325.t6 160.666
R12214 a_19599_25325.n1 a_19599_25325.t5 160.666
R12215 a_19599_25325.n1 a_19599_25325.n0 114.829
R12216 a_19599_25325.n3 a_19599_25325.t1 28.568
R12217 a_19599_25325.n4 a_19599_25325.t2 28.565
R12218 a_19599_25325.t3 a_19599_25325.n4 28.565
R12219 a_19599_25325.n2 a_19599_25325.t0 19.084
R12220 a_19599_25325.n3 a_19599_25325.n2 1.051
R12221 a_15057_14598.n4 a_15057_14598.n3 535.449
R12222 a_15057_14598.t5 a_15057_14598.t19 437.233
R12223 a_15057_14598.t10 a_15057_14598.t6 437.233
R12224 a_15057_14598.t11 a_15057_14598.n1 313.873
R12225 a_15057_14598.n3 a_15057_14598.t7 294.986
R12226 a_15057_14598.n0 a_15057_14598.t8 272.288
R12227 a_15057_14598.n4 a_15057_14598.t16 245.184
R12228 a_15057_14598.n6 a_15057_14598.t10 218.628
R12229 a_15057_14598.n8 a_15057_14598.t5 217.024
R12230 a_15057_14598.n7 a_15057_14598.t12 214.686
R12231 a_15057_14598.t19 a_15057_14598.n7 214.686
R12232 a_15057_14598.n5 a_15057_14598.t4 214.686
R12233 a_15057_14598.t6 a_15057_14598.n5 214.686
R12234 a_15057_14598.n11 a_15057_14598.n10 192.754
R12235 a_15057_14598.n2 a_15057_14598.t11 190.152
R12236 a_15057_14598.n2 a_15057_14598.t18 190.152
R12237 a_15057_14598.n0 a_15057_14598.t9 160.666
R12238 a_15057_14598.n1 a_15057_14598.t14 160.666
R12239 a_15057_14598.n3 a_15057_14598.t15 110.859
R12240 a_15057_14598.n1 a_15057_14598.n0 96.129
R12241 a_15057_14598.n7 a_15057_14598.t17 80.333
R12242 a_15057_14598.t16 a_15057_14598.n2 80.333
R12243 a_15057_14598.n5 a_15057_14598.t13 80.333
R12244 a_15057_14598.n10 a_15057_14598.t1 28.568
R12245 a_15057_14598.n11 a_15057_14598.t2 28.565
R12246 a_15057_14598.t3 a_15057_14598.n11 28.565
R12247 a_15057_14598.n9 a_15057_14598.t0 20.07
R12248 a_15057_14598.n6 a_15057_14598.n4 14.9
R12249 a_15057_14598.n9 a_15057_14598.n8 3.139
R12250 a_15057_14598.n8 a_15057_14598.n6 2.599
R12251 a_15057_14598.n10 a_15057_14598.n9 1.101
R12252 a_18916_21033.t5 a_18916_21033.n3 404.877
R12253 a_18916_21033.n2 a_18916_21033.t8 210.902
R12254 a_18916_21033.n4 a_18916_21033.t5 136.949
R12255 a_18916_21033.n3 a_18916_21033.n2 107.801
R12256 a_18916_21033.n2 a_18916_21033.t6 80.333
R12257 a_18916_21033.n3 a_18916_21033.t7 80.333
R12258 a_18916_21033.n1 a_18916_21033.t1 17.4
R12259 a_18916_21033.n1 a_18916_21033.t4 17.4
R12260 a_18916_21033.t0 a_18916_21033.n5 15.032
R12261 a_18916_21033.n0 a_18916_21033.t3 14.282
R12262 a_18916_21033.n0 a_18916_21033.t2 14.282
R12263 a_18916_21033.n5 a_18916_21033.n0 1.65
R12264 a_18916_21033.n4 a_18916_21033.n1 0.657
R12265 a_18916_21033.n5 a_18916_21033.n4 0.614
R12266 A[7].n4 A[7].n3 535.449
R12267 A[7].t4 A[7].t3 437.233
R12268 A[7].t5 A[7].t10 437.233
R12269 A[7].t15 A[7].n1 313.873
R12270 A[7].n3 A[7].t12 294.986
R12271 A[7].n0 A[7].t9 272.288
R12272 A[7].n4 A[7].t14 245.184
R12273 A[7].n6 A[7].t5 218.627
R12274 A[7].n8 A[7].t4 217.023
R12275 A[7].n7 A[7].t13 214.686
R12276 A[7].t3 A[7].n7 214.686
R12277 A[7].n5 A[7].t1 214.686
R12278 A[7].t10 A[7].n5 214.686
R12279 A[7].n2 A[7].t6 190.152
R12280 A[7].n2 A[7].t15 190.152
R12281 A[7].n0 A[7].t8 160.666
R12282 A[7].n1 A[7].t7 160.666
R12283 A[7].n3 A[7].t2 110.859
R12284 A[7].n1 A[7].n0 96.129
R12285 A[7].n7 A[7].t11 80.333
R12286 A[7].t14 A[7].n2 80.333
R12287 A[7].n5 A[7].t0 80.333
R12288 A[7] A[7].n8 32.3
R12289 A[7].n6 A[7].n4 14.9
R12290 A[7].n8 A[7].n6 2.599
R12291 a_9003_18532.n0 a_9003_18532.t7 214.335
R12292 a_9003_18532.t10 a_9003_18532.n0 214.335
R12293 a_9003_18532.n1 a_9003_18532.t10 143.851
R12294 a_9003_18532.n1 a_9003_18532.t9 135.658
R12295 a_9003_18532.n0 a_9003_18532.t8 80.333
R12296 a_9003_18532.n2 a_9003_18532.t5 28.565
R12297 a_9003_18532.n2 a_9003_18532.t6 28.565
R12298 a_9003_18532.n4 a_9003_18532.t1 28.565
R12299 a_9003_18532.n4 a_9003_18532.t4 28.565
R12300 a_9003_18532.n7 a_9003_18532.t2 28.565
R12301 a_9003_18532.t3 a_9003_18532.n7 28.565
R12302 a_9003_18532.n6 a_9003_18532.t0 9.714
R12303 a_9003_18532.n7 a_9003_18532.n6 1.003
R12304 a_9003_18532.n5 a_9003_18532.n3 0.833
R12305 a_9003_18532.n3 a_9003_18532.n2 0.653
R12306 a_9003_18532.n5 a_9003_18532.n4 0.653
R12307 a_9003_18532.n6 a_9003_18532.n5 0.341
R12308 a_9003_18532.n3 a_9003_18532.n1 0.032
R12309 a_25877_9997.n0 a_25877_9997.n12 122.999
R12310 a_25877_9997.t1 a_25877_9997.n0 14.282
R12311 a_25877_9997.n0 a_25877_9997.t3 14.282
R12312 a_25877_9997.n12 a_25877_9997.n10 50.575
R12313 a_25877_9997.n10 a_25877_9997.n8 74.302
R12314 a_25877_9997.n12 a_25877_9997.n11 157.665
R12315 a_25877_9997.n11 a_25877_9997.t0 8.7
R12316 a_25877_9997.n11 a_25877_9997.t5 8.7
R12317 a_25877_9997.n10 a_25877_9997.n9 90.416
R12318 a_25877_9997.n9 a_25877_9997.t2 14.282
R12319 a_25877_9997.n9 a_25877_9997.t6 14.282
R12320 a_25877_9997.n8 a_25877_9997.n7 90.436
R12321 a_25877_9997.n7 a_25877_9997.t4 14.282
R12322 a_25877_9997.n7 a_25877_9997.t7 14.282
R12323 a_25877_9997.n8 a_25877_9997.n1 342.688
R12324 a_25877_9997.n1 a_25877_9997.n6 126.566
R12325 a_25877_9997.n6 a_25877_9997.t12 294.653
R12326 a_25877_9997.n6 a_25877_9997.t13 111.663
R12327 a_25877_9997.n1 a_25877_9997.n5 552.333
R12328 a_25877_9997.n5 a_25877_9997.n4 6.615
R12329 a_25877_9997.n4 a_25877_9997.t8 93.989
R12330 a_25877_9997.n5 a_25877_9997.n3 97.816
R12331 a_25877_9997.n3 a_25877_9997.t9 80.333
R12332 a_25877_9997.n3 a_25877_9997.t10 394.151
R12333 a_25877_9997.t10 a_25877_9997.n2 269.523
R12334 a_25877_9997.n2 a_25877_9997.t11 160.666
R12335 a_25877_9997.n2 a_25877_9997.t15 269.523
R12336 a_25877_9997.n4 a_25877_9997.t14 198.043
R12337 a_27230_10690.n1 a_27230_10690.t4 318.922
R12338 a_27230_10690.n0 a_27230_10690.t5 273.935
R12339 a_27230_10690.n0 a_27230_10690.t7 273.935
R12340 a_27230_10690.n1 a_27230_10690.t6 269.116
R12341 a_27230_10690.n4 a_27230_10690.n3 193.227
R12342 a_27230_10690.t4 a_27230_10690.n0 179.142
R12343 a_27230_10690.n2 a_27230_10690.n1 106.999
R12344 a_27230_10690.n3 a_27230_10690.t1 28.568
R12345 a_27230_10690.n4 a_27230_10690.t2 28.565
R12346 a_27230_10690.t3 a_27230_10690.n4 28.565
R12347 a_27230_10690.n2 a_27230_10690.t0 18.149
R12348 a_27230_10690.n3 a_27230_10690.n2 3.726
R12349 a_4098_11193.n15 a_4098_11193.n14 3522.62
R12350 a_4098_11193.n6 a_4098_11193.n5 501.28
R12351 a_4098_11193.t7 a_4098_11193.t16 437.233
R12352 a_4098_11193.t6 a_4098_11193.t19 415.315
R12353 a_4098_11193.t14 a_4098_11193.n3 313.873
R12354 a_4098_11193.n5 a_4098_11193.t9 294.986
R12355 a_4098_11193.n2 a_4098_11193.t17 272.288
R12356 a_4098_11193.n6 a_4098_11193.t18 236.01
R12357 a_4098_11193.n9 a_4098_11193.t7 216.627
R12358 a_4098_11193.n7 a_4098_11193.t6 216.111
R12359 a_4098_11193.n8 a_4098_11193.t11 214.686
R12360 a_4098_11193.t16 a_4098_11193.n8 214.686
R12361 a_4098_11193.n1 a_4098_11193.t10 214.335
R12362 a_4098_11193.t19 a_4098_11193.n1 214.335
R12363 a_4098_11193.n17 a_4098_11193.n16 192.754
R12364 a_4098_11193.n4 a_4098_11193.t14 190.152
R12365 a_4098_11193.n4 a_4098_11193.t8 190.152
R12366 a_4098_11193.n2 a_4098_11193.t4 160.666
R12367 a_4098_11193.n3 a_4098_11193.t5 160.666
R12368 a_4098_11193.n7 a_4098_11193.n6 148.428
R12369 a_4098_11193.n5 a_4098_11193.t12 110.859
R12370 a_4098_11193.n3 a_4098_11193.n2 96.129
R12371 a_4098_11193.n8 a_4098_11193.t15 80.333
R12372 a_4098_11193.n1 a_4098_11193.t13 80.333
R12373 a_4098_11193.t18 a_4098_11193.n4 80.333
R12374 a_4098_11193.n16 a_4098_11193.t1 28.568
R12375 a_4098_11193.n17 a_4098_11193.t2 28.565
R12376 a_4098_11193.t3 a_4098_11193.n17 28.565
R12377 a_4098_11193.n15 a_4098_11193.t0 18.522
R12378 a_4098_11193.n14 a_4098_11193.n13 5.25
R12379 a_4098_11193.n13 a_4098_11193.n12 3.293
R12380 a_4098_11193.n9 a_4098_11193.n7 2.923
R12381 a_4098_11193.n16 a_4098_11193.n15 1.168
R12382 a_4098_11193.n10 a_4098_11193.n9 0.708
R12383 a_4098_11193.n13 a_4098_11193.n11 0.681
R12384 a_4098_11193.n11 a_4098_11193.n0 0.003
R12385 a_4098_11193.n11 a_4098_11193.n10 0.001
R12386 a_14704_14398.t0 a_14704_14398.t1 17.4
R12387 a_21711_14619.n4 a_21711_14619.n3 535.449
R12388 a_21711_14619.t15 a_21711_14619.t13 437.233
R12389 a_21711_14619.t16 a_21711_14619.t14 437.233
R12390 a_21711_14619.t4 a_21711_14619.n1 313.873
R12391 a_21711_14619.n3 a_21711_14619.t18 294.986
R12392 a_21711_14619.n0 a_21711_14619.t7 272.288
R12393 a_21711_14619.n4 a_21711_14619.t11 245.184
R12394 a_21711_14619.n6 a_21711_14619.t16 218.628
R12395 a_21711_14619.n8 a_21711_14619.t15 217.024
R12396 a_21711_14619.n7 a_21711_14619.t10 214.686
R12397 a_21711_14619.t13 a_21711_14619.n7 214.686
R12398 a_21711_14619.n5 a_21711_14619.t5 214.686
R12399 a_21711_14619.t14 a_21711_14619.n5 214.686
R12400 a_21711_14619.n11 a_21711_14619.n10 192.754
R12401 a_21711_14619.n2 a_21711_14619.t4 190.152
R12402 a_21711_14619.n2 a_21711_14619.t12 190.152
R12403 a_21711_14619.n0 a_21711_14619.t8 160.666
R12404 a_21711_14619.n1 a_21711_14619.t9 160.666
R12405 a_21711_14619.n3 a_21711_14619.t17 110.859
R12406 a_21711_14619.n1 a_21711_14619.n0 96.129
R12407 a_21711_14619.n7 a_21711_14619.t6 80.333
R12408 a_21711_14619.t11 a_21711_14619.n2 80.333
R12409 a_21711_14619.n5 a_21711_14619.t19 80.333
R12410 a_21711_14619.n10 a_21711_14619.t3 28.568
R12411 a_21711_14619.n11 a_21711_14619.t1 28.565
R12412 a_21711_14619.t0 a_21711_14619.n11 28.565
R12413 a_21711_14619.n9 a_21711_14619.t2 18.823
R12414 a_21711_14619.n6 a_21711_14619.n4 14.9
R12415 a_21711_14619.n9 a_21711_14619.n8 3.074
R12416 a_21711_14619.n8 a_21711_14619.n6 2.599
R12417 a_21711_14619.n10 a_21711_14619.n9 1.105
R12418 a_26171_9971.n1 a_26171_9971.t7 318.922
R12419 a_26171_9971.n0 a_26171_9971.t5 274.739
R12420 a_26171_9971.n0 a_26171_9971.t4 274.739
R12421 a_26171_9971.n1 a_26171_9971.t6 269.116
R12422 a_26171_9971.t7 a_26171_9971.n0 179.946
R12423 a_26171_9971.n2 a_26171_9971.n1 107.263
R12424 a_26171_9971.n3 a_26171_9971.t1 29.444
R12425 a_26171_9971.n4 a_26171_9971.t2 28.565
R12426 a_26171_9971.t3 a_26171_9971.n4 28.565
R12427 a_26171_9971.n2 a_26171_9971.t0 18.145
R12428 a_26171_9971.n3 a_26171_9971.n2 2.878
R12429 a_26171_9971.n4 a_26171_9971.n3 0.764
R12430 a_25228_18856.n0 a_25228_18856.t7 14.282
R12431 a_25228_18856.t0 a_25228_18856.n0 14.282
R12432 a_25228_18856.n0 a_25228_18856.n8 90.416
R12433 a_25228_18856.n8 a_25228_18856.n5 74.302
R12434 a_25228_18856.n8 a_25228_18856.n7 50.575
R12435 a_25228_18856.n7 a_25228_18856.n6 157.665
R12436 a_25228_18856.n6 a_25228_18856.t1 8.7
R12437 a_25228_18856.n6 a_25228_18856.t3 8.7
R12438 a_25228_18856.n5 a_25228_18856.n4 90.436
R12439 a_25228_18856.n4 a_25228_18856.t6 14.282
R12440 a_25228_18856.n4 a_25228_18856.t5 14.282
R12441 a_25228_18856.n7 a_25228_18856.n3 122.746
R12442 a_25228_18856.n3 a_25228_18856.t4 14.282
R12443 a_25228_18856.n3 a_25228_18856.t2 14.282
R12444 a_25228_18856.n5 a_25228_18856.n1 260.998
R12445 a_25228_18856.t11 a_25228_18856.n2 160.666
R12446 a_25228_18856.n1 a_25228_18856.t11 867.393
R12447 a_25228_18856.n2 a_25228_18856.t9 287.241
R12448 a_25228_18856.n2 a_25228_18856.t8 287.241
R12449 a_25228_18856.n1 a_25228_18856.t10 545.094
R12450 a_10045_24434.n1 a_10045_24434.t5 318.922
R12451 a_10045_24434.n0 a_10045_24434.t4 274.739
R12452 a_10045_24434.n0 a_10045_24434.t6 274.739
R12453 a_10045_24434.n1 a_10045_24434.t7 269.116
R12454 a_10045_24434.t5 a_10045_24434.n0 179.946
R12455 a_10045_24434.n2 a_10045_24434.n1 105.178
R12456 a_10045_24434.n3 a_10045_24434.t1 29.444
R12457 a_10045_24434.n4 a_10045_24434.t2 28.565
R12458 a_10045_24434.t3 a_10045_24434.n4 28.565
R12459 a_10045_24434.n2 a_10045_24434.t0 18.145
R12460 a_10045_24434.n3 a_10045_24434.n2 2.878
R12461 a_10045_24434.n4 a_10045_24434.n3 0.764
R12462 a_n3806_2724.t0 a_n3806_2724.n9 16.058
R12463 a_n3806_2724.n9 a_n3806_2724.n5 0.2
R12464 a_n3806_2724.n5 a_n3806_2724.n7 0.575
R12465 a_n3806_2724.n9 a_n3806_2724.n8 0.999
R12466 a_n3806_2724.n8 a_n3806_2724.t11 14.282
R12467 a_n3806_2724.n8 a_n3806_2724.t4 14.282
R12468 a_n3806_2724.n7 a_n3806_2724.n6 0.999
R12469 a_n3806_2724.n6 a_n3806_2724.t7 14.282
R12470 a_n3806_2724.n6 a_n3806_2724.t6 14.282
R12471 a_n3806_2724.n7 a_n3806_2724.t5 16.058
R12472 a_n3806_2724.n5 a_n3806_2724.n3 0.227
R12473 a_n3806_2724.n3 a_n3806_2724.n4 1.511
R12474 a_n3806_2724.n4 a_n3806_2724.t3 14.282
R12475 a_n3806_2724.n4 a_n3806_2724.t2 14.282
R12476 a_n3806_2724.n3 a_n3806_2724.n0 0.669
R12477 a_n3806_2724.n0 a_n3806_2724.n1 0.001
R12478 a_n3806_2724.n0 a_n3806_2724.n2 267.767
R12479 a_n3806_2724.n2 a_n3806_2724.t10 14.282
R12480 a_n3806_2724.n2 a_n3806_2724.t9 14.282
R12481 a_n3806_2724.n1 a_n3806_2724.t8 14.282
R12482 a_n3806_2724.n1 a_n3806_2724.t1 14.282
R12483 a_25553_27416.n0 a_25553_27416.t8 214.335
R12484 a_25553_27416.t10 a_25553_27416.n0 214.335
R12485 a_25553_27416.n1 a_25553_27416.t10 143.851
R12486 a_25553_27416.n1 a_25553_27416.t9 135.658
R12487 a_25553_27416.n0 a_25553_27416.t7 80.333
R12488 a_25553_27416.n2 a_25553_27416.t6 28.565
R12489 a_25553_27416.n2 a_25553_27416.t4 28.565
R12490 a_25553_27416.n4 a_25553_27416.t5 28.565
R12491 a_25553_27416.n4 a_25553_27416.t2 28.565
R12492 a_25553_27416.t3 a_25553_27416.n7 28.565
R12493 a_25553_27416.n7 a_25553_27416.t1 28.565
R12494 a_25553_27416.n6 a_25553_27416.t0 9.714
R12495 a_25553_27416.n7 a_25553_27416.n6 1.003
R12496 a_25553_27416.n5 a_25553_27416.n3 0.833
R12497 a_25553_27416.n3 a_25553_27416.n2 0.653
R12498 a_25553_27416.n5 a_25553_27416.n4 0.653
R12499 a_25553_27416.n6 a_25553_27416.n5 0.341
R12500 a_25553_27416.n3 a_25553_27416.n1 0.032
R12501 a_13953_21654.t7 a_13953_21654.t4 574.43
R12502 a_13953_21654.n1 a_13953_21654.t6 285.109
R12503 a_13953_21654.n3 a_13953_21654.n2 197.215
R12504 a_13953_21654.n4 a_13953_21654.n0 192.754
R12505 a_13953_21654.n1 a_13953_21654.t5 160.666
R12506 a_13953_21654.n2 a_13953_21654.t7 160.666
R12507 a_13953_21654.n2 a_13953_21654.n1 114.829
R12508 a_13953_21654.t3 a_13953_21654.n4 28.568
R12509 a_13953_21654.n0 a_13953_21654.t1 28.565
R12510 a_13953_21654.n0 a_13953_21654.t2 28.565
R12511 a_13953_21654.n3 a_13953_21654.t0 18.838
R12512 a_13953_21654.n4 a_13953_21654.n3 1.129
R12513 a_13524_21024.t8 a_13524_21024.n3 404.877
R12514 a_13524_21024.n2 a_13524_21024.t5 210.902
R12515 a_13524_21024.n4 a_13524_21024.t8 136.949
R12516 a_13524_21024.n3 a_13524_21024.n2 107.801
R12517 a_13524_21024.n2 a_13524_21024.t6 80.333
R12518 a_13524_21024.n3 a_13524_21024.t7 80.333
R12519 a_13524_21024.n1 a_13524_21024.t2 17.4
R12520 a_13524_21024.n1 a_13524_21024.t4 17.4
R12521 a_13524_21024.t0 a_13524_21024.n5 15.032
R12522 a_13524_21024.n0 a_13524_21024.t3 14.282
R12523 a_13524_21024.n0 a_13524_21024.t1 14.282
R12524 a_13524_21024.n5 a_13524_21024.n0 1.65
R12525 a_13524_21024.n4 a_13524_21024.n1 0.657
R12526 a_13524_21024.n5 a_13524_21024.n4 0.614
R12527 a_17598_10602.t0 a_17598_10602.t1 17.4
R12528 a_36751_4115.n2 a_36751_4115.t8 1551.5
R12529 a_36751_4115.t8 a_36751_4115.n0 656.576
R12530 a_36751_4115.n4 a_36751_4115.n3 258.161
R12531 a_36751_4115.n7 a_36751_4115.n6 258.161
R12532 a_36751_4115.n2 a_36751_4115.t9 224.129
R12533 a_36751_4115.n1 a_36751_4115.t11 207.225
R12534 a_36751_4115.t9 a_36751_4115.n1 207.225
R12535 a_36751_4115.n1 a_36751_4115.t10 80.333
R12536 a_36751_4115.n5 a_36751_4115.n2 73.514
R12537 a_36751_4115.n4 a_36751_4115.t5 14.283
R12538 a_36751_4115.t2 a_36751_4115.n7 14.283
R12539 a_36751_4115.n3 a_36751_4115.t3 14.282
R12540 a_36751_4115.n3 a_36751_4115.t4 14.282
R12541 a_36751_4115.n6 a_36751_4115.t1 14.282
R12542 a_36751_4115.n6 a_36751_4115.t0 14.282
R12543 a_36751_4115.n0 a_36751_4115.t7 8.7
R12544 a_36751_4115.n0 a_36751_4115.t6 8.7
R12545 a_36751_4115.n5 a_36751_4115.n4 4.366
R12546 a_36751_4115.n7 a_36751_4115.n5 0.852
R12547 Y[6].n1 Y[6].n0 185.55
R12548 Y[6].n1 Y[6].t3 28.568
R12549 Y[6].n0 Y[6].t1 28.565
R12550 Y[6].n0 Y[6].t2 28.565
R12551 Y[6].n2 Y[6].t0 20.393
R12552 Y[6].n2 Y[6].n1 1.836
R12553 Y[6].n3 Y[6].n2 1.049
R12554 Y[6] Y[6].n3 0.052
R12555 Y[6].n3 Y[6] 0.046
R12556 a_31466_10393.n2 a_31466_10393.t4 318.922
R12557 a_31466_10393.n1 a_31466_10393.t5 273.935
R12558 a_31466_10393.n1 a_31466_10393.t7 273.935
R12559 a_31466_10393.n2 a_31466_10393.t6 269.116
R12560 a_31466_10393.n4 a_31466_10393.n0 193.227
R12561 a_31466_10393.t4 a_31466_10393.n1 179.142
R12562 a_31466_10393.n3 a_31466_10393.n2 106.999
R12563 a_31466_10393.t3 a_31466_10393.n4 28.568
R12564 a_31466_10393.n0 a_31466_10393.t1 28.565
R12565 a_31466_10393.n0 a_31466_10393.t2 28.565
R12566 a_31466_10393.n3 a_31466_10393.t0 18.149
R12567 a_31466_10393.n4 a_31466_10393.n3 3.726
R12568 a_31893_9700.n8 a_31893_9700.n0 267.767
R12569 a_31893_9700.n4 a_31893_9700.t4 16.058
R12570 a_31893_9700.n2 a_31893_9700.t7 16.058
R12571 a_31893_9700.n3 a_31893_9700.t3 14.282
R12572 a_31893_9700.n3 a_31893_9700.t5 14.282
R12573 a_31893_9700.n1 a_31893_9700.t6 14.282
R12574 a_31893_9700.n1 a_31893_9700.t8 14.282
R12575 a_31893_9700.n6 a_31893_9700.t10 14.282
R12576 a_31893_9700.n6 a_31893_9700.t11 14.282
R12577 a_31893_9700.n0 a_31893_9700.t0 14.282
R12578 a_31893_9700.n0 a_31893_9700.t1 14.282
R12579 a_31893_9700.t2 a_31893_9700.n9 14.282
R12580 a_31893_9700.n9 a_31893_9700.t9 14.282
R12581 a_31893_9700.n7 a_31893_9700.n6 1.511
R12582 a_31893_9700.n4 a_31893_9700.n3 0.999
R12583 a_31893_9700.n2 a_31893_9700.n1 0.999
R12584 a_31893_9700.n8 a_31893_9700.n7 0.669
R12585 a_31893_9700.n5 a_31893_9700.n4 0.575
R12586 a_31893_9700.n7 a_31893_9700.n5 0.227
R12587 a_31893_9700.n5 a_31893_9700.n2 0.2
R12588 a_31893_9700.n9 a_31893_9700.n8 0.001
R12589 a_26913_25149.n1 a_26913_25149.t6 318.922
R12590 a_26913_25149.n0 a_26913_25149.t5 273.935
R12591 a_26913_25149.n0 a_26913_25149.t7 273.935
R12592 a_26913_25149.n1 a_26913_25149.t4 269.116
R12593 a_26913_25149.n4 a_26913_25149.n3 193.227
R12594 a_26913_25149.t6 a_26913_25149.n0 179.142
R12595 a_26913_25149.n2 a_26913_25149.n1 106.999
R12596 a_26913_25149.n3 a_26913_25149.t2 28.568
R12597 a_26913_25149.t3 a_26913_25149.n4 28.565
R12598 a_26913_25149.n4 a_26913_25149.t1 28.565
R12599 a_26913_25149.n2 a_26913_25149.t0 18.149
R12600 a_26913_25149.n3 a_26913_25149.n2 3.726
R12601 a_n3806_8930.n2 a_n3806_8930.n1 267.767
R12602 a_n3806_8930.n6 a_n3806_8930.t9 16.058
R12603 a_n3806_8930.n8 a_n3806_8930.t1 16.058
R12604 a_n3806_8930.n0 a_n3806_8930.t4 14.282
R12605 a_n3806_8930.n0 a_n3806_8930.t6 14.282
R12606 a_n3806_8930.n1 a_n3806_8930.t7 14.282
R12607 a_n3806_8930.n1 a_n3806_8930.t8 14.282
R12608 a_n3806_8930.n3 a_n3806_8930.t5 14.282
R12609 a_n3806_8930.n3 a_n3806_8930.t3 14.282
R12610 a_n3806_8930.n5 a_n3806_8930.t10 14.282
R12611 a_n3806_8930.n5 a_n3806_8930.t11 14.282
R12612 a_n3806_8930.t2 a_n3806_8930.n9 14.282
R12613 a_n3806_8930.n9 a_n3806_8930.t0 14.282
R12614 a_n3806_8930.n4 a_n3806_8930.n3 1.511
R12615 a_n3806_8930.n6 a_n3806_8930.n5 0.999
R12616 a_n3806_8930.n9 a_n3806_8930.n8 0.999
R12617 a_n3806_8930.n4 a_n3806_8930.n2 0.669
R12618 a_n3806_8930.n7 a_n3806_8930.n6 0.575
R12619 a_n3806_8930.n7 a_n3806_8930.n4 0.227
R12620 a_n3806_8930.n8 a_n3806_8930.n7 0.2
R12621 a_n3806_8930.n2 a_n3806_8930.n0 0.001
R12622 a_22798_24452.n5 a_22798_24452.n4 1467.36
R12623 a_22798_24452.n4 a_22798_24452.t11 867.393
R12624 a_22798_24452.n4 a_22798_24452.t10 545.094
R12625 a_22798_24452.n3 a_22798_24452.t8 287.241
R12626 a_22798_24452.n3 a_22798_24452.t9 287.241
R12627 a_22798_24452.t11 a_22798_24452.n3 160.666
R12628 a_22798_24452.n7 a_22798_24452.n0 157.665
R12629 a_22798_24452.n8 a_22798_24452.n7 122.999
R12630 a_22798_24452.n5 a_22798_24452.n2 90.436
R12631 a_22798_24452.n6 a_22798_24452.n1 90.416
R12632 a_22798_24452.n6 a_22798_24452.n5 74.302
R12633 a_22798_24452.n7 a_22798_24452.n6 50.575
R12634 a_22798_24452.n2 a_22798_24452.t5 14.282
R12635 a_22798_24452.n2 a_22798_24452.t6 14.282
R12636 a_22798_24452.n1 a_22798_24452.t7 14.282
R12637 a_22798_24452.n1 a_22798_24452.t1 14.282
R12638 a_22798_24452.n8 a_22798_24452.t2 14.282
R12639 a_22798_24452.t3 a_22798_24452.n8 14.282
R12640 a_22798_24452.n0 a_22798_24452.t4 8.7
R12641 a_22798_24452.n0 a_22798_24452.t0 8.7
R12642 a_32303_13765.n1 a_32303_13765.t5 318.922
R12643 a_32303_13765.n0 a_32303_13765.t4 274.739
R12644 a_32303_13765.n0 a_32303_13765.t6 274.739
R12645 a_32303_13765.n1 a_32303_13765.t7 269.116
R12646 a_32303_13765.t5 a_32303_13765.n0 179.946
R12647 a_32303_13765.n2 a_32303_13765.n1 107.263
R12648 a_32303_13765.n3 a_32303_13765.t1 29.444
R12649 a_32303_13765.n4 a_32303_13765.t2 28.565
R12650 a_32303_13765.t3 a_32303_13765.n4 28.565
R12651 a_32303_13765.n2 a_32303_13765.t0 18.145
R12652 a_32303_13765.n3 a_32303_13765.n2 2.878
R12653 a_32303_13765.n4 a_32303_13765.n3 0.764
R12654 a_23964_7089.n4 a_23964_7089.t10 214.335
R12655 a_23964_7089.t9 a_23964_7089.n4 214.335
R12656 a_23964_7089.n5 a_23964_7089.t9 143.851
R12657 a_23964_7089.n5 a_23964_7089.t7 135.658
R12658 a_23964_7089.n4 a_23964_7089.t8 80.333
R12659 a_23964_7089.n0 a_23964_7089.t4 28.565
R12660 a_23964_7089.n0 a_23964_7089.t5 28.565
R12661 a_23964_7089.n2 a_23964_7089.t0 28.565
R12662 a_23964_7089.n2 a_23964_7089.t6 28.565
R12663 a_23964_7089.t2 a_23964_7089.n7 28.565
R12664 a_23964_7089.n7 a_23964_7089.t1 28.565
R12665 a_23964_7089.n1 a_23964_7089.t3 9.714
R12666 a_23964_7089.n1 a_23964_7089.n0 1.003
R12667 a_23964_7089.n6 a_23964_7089.n3 0.833
R12668 a_23964_7089.n3 a_23964_7089.n2 0.653
R12669 a_23964_7089.n7 a_23964_7089.n6 0.653
R12670 a_23964_7089.n3 a_23964_7089.n1 0.341
R12671 a_23964_7089.n6 a_23964_7089.n5 0.032
R12672 a_24554_6652.t6 a_24554_6652.t4 800.071
R12673 a_24554_6652.n2 a_24554_6652.n1 659.097
R12674 a_24554_6652.n0 a_24554_6652.t5 285.109
R12675 a_24554_6652.n1 a_24554_6652.t6 193.602
R12676 a_24554_6652.n4 a_24554_6652.n3 192.754
R12677 a_24554_6652.n0 a_24554_6652.t7 160.666
R12678 a_24554_6652.n1 a_24554_6652.n0 91.507
R12679 a_24554_6652.n3 a_24554_6652.t1 28.568
R12680 a_24554_6652.t3 a_24554_6652.n4 28.565
R12681 a_24554_6652.n4 a_24554_6652.t2 28.565
R12682 a_24554_6652.n2 a_24554_6652.t0 19.061
R12683 a_24554_6652.n3 a_24554_6652.n2 1.005
R12684 a_18995_27412.n4 a_18995_27412.t10 214.335
R12685 a_18995_27412.t8 a_18995_27412.n4 214.335
R12686 a_18995_27412.n5 a_18995_27412.t8 143.851
R12687 a_18995_27412.n5 a_18995_27412.t7 135.658
R12688 a_18995_27412.n4 a_18995_27412.t9 80.333
R12689 a_18995_27412.n0 a_18995_27412.t6 28.565
R12690 a_18995_27412.n0 a_18995_27412.t4 28.565
R12691 a_18995_27412.n2 a_18995_27412.t0 28.565
R12692 a_18995_27412.n2 a_18995_27412.t5 28.565
R12693 a_18995_27412.n7 a_18995_27412.t1 28.565
R12694 a_18995_27412.t2 a_18995_27412.n7 28.565
R12695 a_18995_27412.n1 a_18995_27412.t3 9.714
R12696 a_18995_27412.n1 a_18995_27412.n0 1.003
R12697 a_18995_27412.n6 a_18995_27412.n3 0.833
R12698 a_18995_27412.n3 a_18995_27412.n2 0.653
R12699 a_18995_27412.n7 a_18995_27412.n6 0.653
R12700 a_18995_27412.n3 a_18995_27412.n1 0.341
R12701 a_18995_27412.n6 a_18995_27412.n5 0.032
R12702 a_19585_26975.t4 a_19585_26975.t7 800.071
R12703 a_19585_26975.n2 a_19585_26975.n1 659.097
R12704 a_19585_26975.n0 a_19585_26975.t6 285.109
R12705 a_19585_26975.n1 a_19585_26975.t4 193.602
R12706 a_19585_26975.n4 a_19585_26975.n3 192.754
R12707 a_19585_26975.n0 a_19585_26975.t5 160.666
R12708 a_19585_26975.n1 a_19585_26975.n0 91.507
R12709 a_19585_26975.n3 a_19585_26975.t1 28.568
R12710 a_19585_26975.n4 a_19585_26975.t2 28.565
R12711 a_19585_26975.t3 a_19585_26975.n4 28.565
R12712 a_19585_26975.n2 a_19585_26975.t0 19.061
R12713 a_19585_26975.n3 a_19585_26975.n2 1.005
R12714 a_26171_6961.t8 a_26171_6961.n2 404.877
R12715 a_26171_6961.n1 a_26171_6961.t5 210.902
R12716 a_26171_6961.n3 a_26171_6961.t8 136.943
R12717 a_26171_6961.n2 a_26171_6961.n1 107.801
R12718 a_26171_6961.n1 a_26171_6961.t6 80.333
R12719 a_26171_6961.n2 a_26171_6961.t7 80.333
R12720 a_26171_6961.n0 a_26171_6961.t4 17.4
R12721 a_26171_6961.n0 a_26171_6961.t2 17.4
R12722 a_26171_6961.n4 a_26171_6961.t3 15.032
R12723 a_26171_6961.n5 a_26171_6961.t1 14.282
R12724 a_26171_6961.t0 a_26171_6961.n5 14.282
R12725 a_26171_6961.n5 a_26171_6961.n4 1.65
R12726 a_26171_6961.n3 a_26171_6961.n0 0.672
R12727 a_26171_6961.n4 a_26171_6961.n3 0.665
R12728 a_26435_6378.t5 a_26435_6378.t6 800.071
R12729 a_26435_6378.n3 a_26435_6378.n2 672.951
R12730 a_26435_6378.n1 a_26435_6378.t7 285.109
R12731 a_26435_6378.n2 a_26435_6378.t5 193.602
R12732 a_26435_6378.n1 a_26435_6378.t4 160.666
R12733 a_26435_6378.n2 a_26435_6378.n1 91.507
R12734 a_26435_6378.n0 a_26435_6378.t1 28.57
R12735 a_26435_6378.t3 a_26435_6378.n4 28.565
R12736 a_26435_6378.n4 a_26435_6378.t2 28.565
R12737 a_26435_6378.n0 a_26435_6378.t0 17.638
R12738 a_26435_6378.n4 a_26435_6378.n3 0.69
R12739 a_26435_6378.n3 a_26435_6378.n0 0.6
R12740 a_18057_19546.n1 a_18057_19546.t5 318.922
R12741 a_18057_19546.n0 a_18057_19546.t4 274.739
R12742 a_18057_19546.n0 a_18057_19546.t6 274.739
R12743 a_18057_19546.n1 a_18057_19546.t7 269.116
R12744 a_18057_19546.t5 a_18057_19546.n0 179.946
R12745 a_18057_19546.n2 a_18057_19546.n1 105.178
R12746 a_18057_19546.t3 a_18057_19546.n4 29.444
R12747 a_18057_19546.n3 a_18057_19546.t1 28.565
R12748 a_18057_19546.n3 a_18057_19546.t2 28.565
R12749 a_18057_19546.n2 a_18057_19546.t0 18.145
R12750 a_18057_19546.n4 a_18057_19546.n2 2.878
R12751 a_18057_19546.n4 a_18057_19546.n3 0.764
R12752 a_18715_18853.n0 a_18715_18853.t2 14.282
R12753 a_18715_18853.t0 a_18715_18853.n0 14.282
R12754 a_18715_18853.n0 a_18715_18853.n8 122.747
R12755 a_18715_18853.n4 a_18715_18853.n6 74.302
R12756 a_18715_18853.n8 a_18715_18853.n4 50.575
R12757 a_18715_18853.n8 a_18715_18853.n7 157.665
R12758 a_18715_18853.n7 a_18715_18853.t3 8.7
R12759 a_18715_18853.n7 a_18715_18853.t1 8.7
R12760 a_18715_18853.n6 a_18715_18853.n5 90.436
R12761 a_18715_18853.n5 a_18715_18853.t6 14.282
R12762 a_18715_18853.n5 a_18715_18853.t5 14.282
R12763 a_18715_18853.n4 a_18715_18853.n3 90.416
R12764 a_18715_18853.n3 a_18715_18853.t4 14.282
R12765 a_18715_18853.n3 a_18715_18853.t7 14.282
R12766 a_18715_18853.n6 a_18715_18853.n1 275.913
R12767 a_18715_18853.t11 a_18715_18853.n2 160.666
R12768 a_18715_18853.n1 a_18715_18853.t11 867.393
R12769 a_18715_18853.n2 a_18715_18853.t9 287.241
R12770 a_18715_18853.n2 a_18715_18853.t8 287.241
R12771 a_18715_18853.n1 a_18715_18853.t10 545.094
R12772 a_n2379_15192.t0 a_n2379_15192.t1 379.845
R12773 a_21386_9197.t0 a_21386_9197.t1 17.4
R12774 a_19246_25125.t0 a_19246_25125.t1 17.4
R12775 a_25522_18830.n1 a_25522_18830.t5 318.922
R12776 a_25522_18830.n0 a_25522_18830.t4 273.935
R12777 a_25522_18830.n0 a_25522_18830.t6 273.935
R12778 a_25522_18830.n1 a_25522_18830.t7 269.116
R12779 a_25522_18830.n4 a_25522_18830.n3 193.227
R12780 a_25522_18830.t5 a_25522_18830.n0 179.142
R12781 a_25522_18830.n2 a_25522_18830.n1 106.999
R12782 a_25522_18830.n3 a_25522_18830.t2 28.568
R12783 a_25522_18830.t3 a_25522_18830.n4 28.565
R12784 a_25522_18830.n4 a_25522_18830.t1 28.565
R12785 a_25522_18830.n2 a_25522_18830.t0 18.149
R12786 a_25522_18830.n3 a_25522_18830.n2 3.726
R12787 a_19955_19546.n1 a_19955_19546.t5 318.922
R12788 a_19955_19546.n0 a_19955_19546.t4 274.739
R12789 a_19955_19546.n0 a_19955_19546.t6 274.739
R12790 a_19955_19546.n1 a_19955_19546.t7 269.116
R12791 a_19955_19546.t5 a_19955_19546.n0 179.946
R12792 a_19955_19546.n2 a_19955_19546.n1 107.263
R12793 a_19955_19546.n3 a_19955_19546.t2 29.444
R12794 a_19955_19546.t3 a_19955_19546.n4 28.565
R12795 a_19955_19546.n4 a_19955_19546.t1 28.565
R12796 a_19955_19546.n2 a_19955_19546.t0 18.145
R12797 a_19955_19546.n3 a_19955_19546.n2 2.878
R12798 a_19955_19546.n4 a_19955_19546.n3 0.764
R12799 a_8233_4103.n1 a_8233_4103.t7 318.922
R12800 a_8233_4103.n0 a_8233_4103.t4 274.739
R12801 a_8233_4103.n0 a_8233_4103.t5 274.739
R12802 a_8233_4103.n1 a_8233_4103.t6 269.116
R12803 a_8233_4103.t7 a_8233_4103.n0 179.946
R12804 a_8233_4103.n2 a_8233_4103.n1 105.178
R12805 a_8233_4103.n3 a_8233_4103.t2 29.444
R12806 a_8233_4103.n4 a_8233_4103.t1 28.565
R12807 a_8233_4103.t3 a_8233_4103.n4 28.565
R12808 a_8233_4103.n2 a_8233_4103.t0 18.145
R12809 a_8233_4103.n3 a_8233_4103.n2 2.878
R12810 a_8233_4103.n4 a_8233_4103.n3 0.764
R12811 a_31466_6898.n2 a_31466_6898.t6 318.922
R12812 a_31466_6898.n1 a_31466_6898.t7 273.935
R12813 a_31466_6898.n1 a_31466_6898.t4 273.935
R12814 a_31466_6898.n2 a_31466_6898.t5 269.116
R12815 a_31466_6898.n4 a_31466_6898.n0 193.227
R12816 a_31466_6898.t6 a_31466_6898.n1 179.142
R12817 a_31466_6898.n3 a_31466_6898.n2 106.999
R12818 a_31466_6898.t3 a_31466_6898.n4 28.568
R12819 a_31466_6898.n0 a_31466_6898.t2 28.565
R12820 a_31466_6898.n0 a_31466_6898.t1 28.565
R12821 a_31466_6898.n3 a_31466_6898.t0 18.149
R12822 a_31466_6898.n4 a_31466_6898.n3 3.726
R12823 a_32011_6205.n7 a_32011_6205.n1 1255.94
R12824 a_32011_6205.n1 a_32011_6205.t10 989.744
R12825 a_32011_6205.n1 a_32011_6205.t9 408.806
R12826 a_32011_6205.n0 a_32011_6205.t11 287.241
R12827 a_32011_6205.n0 a_32011_6205.t8 287.241
R12828 a_32011_6205.t10 a_32011_6205.n0 160.666
R12829 a_32011_6205.n5 a_32011_6205.n3 157.665
R12830 a_32011_6205.n5 a_32011_6205.n4 122.999
R12831 a_32011_6205.n8 a_32011_6205.n7 90.436
R12832 a_32011_6205.n6 a_32011_6205.n2 90.416
R12833 a_32011_6205.n7 a_32011_6205.n6 74.302
R12834 a_32011_6205.n6 a_32011_6205.n5 50.575
R12835 a_32011_6205.n2 a_32011_6205.t1 14.282
R12836 a_32011_6205.n2 a_32011_6205.t6 14.282
R12837 a_32011_6205.n4 a_32011_6205.t5 14.282
R12838 a_32011_6205.n4 a_32011_6205.t4 14.282
R12839 a_32011_6205.n8 a_32011_6205.t0 14.282
R12840 a_32011_6205.t2 a_32011_6205.n8 14.282
R12841 a_32011_6205.n3 a_32011_6205.t7 8.7
R12842 a_32011_6205.n3 a_32011_6205.t3 8.7
R12843 a_26706_21688.n1 a_26706_21688.t5 14.282
R12844 a_26706_21688.n1 a_26706_21688.t0 14.282
R12845 a_26706_21688.n0 a_26706_21688.t3 14.282
R12846 a_26706_21688.n0 a_26706_21688.t4 14.282
R12847 a_26706_21688.n3 a_26706_21688.t1 14.282
R12848 a_26706_21688.t2 a_26706_21688.n3 14.282
R12849 a_26706_21688.n2 a_26706_21688.n0 2.546
R12850 a_26706_21688.n3 a_26706_21688.n2 2.367
R12851 a_26706_21688.n2 a_26706_21688.n1 0.001
R12852 a_n2383_949.t0 a_n2383_949.t1 17.4
R12853 a_38084_4824.t0 a_38084_4824.t1 17.4
R12854 a_30434_1013.n6 a_30434_1013.n5 465.933
R12855 a_30434_1013.t12 a_30434_1013.t9 415.315
R12856 a_30434_1013.n2 a_30434_1013.t11 394.151
R12857 a_30434_1013.n5 a_30434_1013.t8 294.653
R12858 a_30434_1013.n1 a_30434_1013.t15 269.523
R12859 a_30434_1013.t11 a_30434_1013.n1 269.523
R12860 a_30434_1013.n8 a_30434_1013.t12 220.285
R12861 a_30434_1013.n7 a_30434_1013.t6 214.335
R12862 a_30434_1013.t9 a_30434_1013.n7 214.335
R12863 a_30434_1013.n3 a_30434_1013.t14 198.043
R12864 a_30434_1013.n10 a_30434_1013.n0 192.754
R12865 a_30434_1013.n6 a_30434_1013.n4 163.88
R12866 a_30434_1013.n1 a_30434_1013.t7 160.666
R12867 a_30434_1013.n5 a_30434_1013.t5 111.663
R12868 a_30434_1013.n4 a_30434_1013.n2 97.816
R12869 a_30434_1013.n3 a_30434_1013.t10 93.989
R12870 a_30434_1013.n7 a_30434_1013.t13 80.333
R12871 a_30434_1013.n2 a_30434_1013.t4 80.333
R12872 a_30434_1013.n8 a_30434_1013.n6 61.538
R12873 a_30434_1013.t0 a_30434_1013.n10 28.568
R12874 a_30434_1013.n0 a_30434_1013.t3 28.565
R12875 a_30434_1013.n0 a_30434_1013.t2 28.565
R12876 a_30434_1013.n9 a_30434_1013.t1 18.824
R12877 a_30434_1013.n4 a_30434_1013.n3 6.615
R12878 a_30434_1013.n9 a_30434_1013.n8 2.736
R12879 a_30434_1013.n10 a_30434_1013.n9 1.105
R12880 a_24201_6452.t0 a_24201_6452.t1 17.4
R12881 a_4390_8978.t0 a_4390_8978.t1 17.4
R12882 a_36751_13593.n2 a_36751_13593.t10 1551.5
R12883 a_36751_13593.t10 a_36751_13593.n0 656.576
R12884 a_36751_13593.n4 a_36751_13593.n3 258.161
R12885 a_36751_13593.n7 a_36751_13593.n6 258.161
R12886 a_36751_13593.n2 a_36751_13593.t11 224.129
R12887 a_36751_13593.n1 a_36751_13593.t9 207.225
R12888 a_36751_13593.t11 a_36751_13593.n1 207.225
R12889 a_36751_13593.n1 a_36751_13593.t8 80.333
R12890 a_36751_13593.n5 a_36751_13593.n2 73.514
R12891 a_36751_13593.n4 a_36751_13593.t4 14.283
R12892 a_36751_13593.n6 a_36751_13593.t1 14.283
R12893 a_36751_13593.n3 a_36751_13593.t5 14.282
R12894 a_36751_13593.n3 a_36751_13593.t6 14.282
R12895 a_36751_13593.t2 a_36751_13593.n7 14.282
R12896 a_36751_13593.n7 a_36751_13593.t0 14.282
R12897 a_36751_13593.n0 a_36751_13593.t7 8.7
R12898 a_36751_13593.n0 a_36751_13593.t3 8.7
R12899 a_36751_13593.n5 a_36751_13593.n4 4.366
R12900 a_36751_13593.n6 a_36751_13593.n5 0.852
R12901 a_4726_6652.t6 a_4726_6652.t5 800.071
R12902 a_4726_6652.n2 a_4726_6652.n1 659.097
R12903 a_4726_6652.n0 a_4726_6652.t7 285.109
R12904 a_4726_6652.n1 a_4726_6652.t6 193.602
R12905 a_4726_6652.n4 a_4726_6652.n3 192.754
R12906 a_4726_6652.n0 a_4726_6652.t4 160.666
R12907 a_4726_6652.n1 a_4726_6652.n0 91.507
R12908 a_4726_6652.n3 a_4726_6652.t2 28.568
R12909 a_4726_6652.t3 a_4726_6652.n4 28.565
R12910 a_4726_6652.n4 a_4726_6652.t1 28.565
R12911 a_4726_6652.n2 a_4726_6652.t0 19.061
R12912 a_4726_6652.n3 a_4726_6652.n2 1.005
R12913 a_20193_21685.n0 a_20193_21685.t0 14.282
R12914 a_20193_21685.n0 a_20193_21685.t1 14.282
R12915 a_20193_21685.n1 a_20193_21685.t3 14.282
R12916 a_20193_21685.n1 a_20193_21685.t4 14.282
R12917 a_20193_21685.t2 a_20193_21685.n3 14.282
R12918 a_20193_21685.n3 a_20193_21685.t5 14.282
R12919 a_20193_21685.n2 a_20193_21685.n0 2.546
R12920 a_20193_21685.n2 a_20193_21685.n1 2.367
R12921 a_20193_21685.n3 a_20193_21685.n2 0.001
R12922 a_11292_9266.t6 a_11292_9266.t7 574.43
R12923 a_11292_9266.n0 a_11292_9266.t5 285.109
R12924 a_11292_9266.n2 a_11292_9266.n1 197.217
R12925 a_11292_9266.n4 a_11292_9266.n3 192.754
R12926 a_11292_9266.n0 a_11292_9266.t4 160.666
R12927 a_11292_9266.n1 a_11292_9266.t6 160.666
R12928 a_11292_9266.n1 a_11292_9266.n0 114.829
R12929 a_11292_9266.n3 a_11292_9266.t2 28.568
R12930 a_11292_9266.n4 a_11292_9266.t1 28.565
R12931 a_11292_9266.t3 a_11292_9266.n4 28.565
R12932 a_11292_9266.n2 a_11292_9266.t0 18.838
R12933 a_11292_9266.n3 a_11292_9266.n2 1.129
R12934 a_24563_3398.t5 a_24563_3398.t6 574.43
R12935 a_24563_3398.n0 a_24563_3398.t7 285.109
R12936 a_24563_3398.n2 a_24563_3398.n1 197.217
R12937 a_24563_3398.n4 a_24563_3398.n3 192.754
R12938 a_24563_3398.n0 a_24563_3398.t4 160.666
R12939 a_24563_3398.n1 a_24563_3398.t5 160.666
R12940 a_24563_3398.n1 a_24563_3398.n0 114.829
R12941 a_24563_3398.n3 a_24563_3398.t2 28.568
R12942 a_24563_3398.n4 a_24563_3398.t1 28.565
R12943 a_24563_3398.t3 a_24563_3398.n4 28.565
R12944 a_24563_3398.n2 a_24563_3398.t0 18.838
R12945 a_24563_3398.n3 a_24563_3398.n2 1.129
R12946 a_26289_6961.n0 a_26289_6961.t4 14.282
R12947 a_26289_6961.n0 a_26289_6961.t0 14.282
R12948 a_26289_6961.n1 a_26289_6961.t5 14.282
R12949 a_26289_6961.n1 a_26289_6961.t3 14.282
R12950 a_26289_6961.t2 a_26289_6961.n3 14.282
R12951 a_26289_6961.n3 a_26289_6961.t1 14.282
R12952 a_26289_6961.n3 a_26289_6961.n2 2.546
R12953 a_26289_6961.n2 a_26289_6961.n1 2.367
R12954 a_26289_6961.n2 a_26289_6961.n0 0.001
R12955 a_4395_10582.t0 a_4395_10582.t1 17.4
R12956 a_8241_9883.n1 a_8241_9883.t7 318.922
R12957 a_8241_9883.n0 a_8241_9883.t4 274.739
R12958 a_8241_9883.n0 a_8241_9883.t5 274.739
R12959 a_8241_9883.n1 a_8241_9883.t6 269.116
R12960 a_8241_9883.t7 a_8241_9883.n0 179.946
R12961 a_8241_9883.n2 a_8241_9883.n1 105.178
R12962 a_8241_9883.t3 a_8241_9883.n4 29.444
R12963 a_8241_9883.n3 a_8241_9883.t1 28.565
R12964 a_8241_9883.n3 a_8241_9883.t2 28.565
R12965 a_8241_9883.n2 a_8241_9883.t0 18.145
R12966 a_8241_9883.n4 a_8241_9883.n2 2.878
R12967 a_8241_9883.n4 a_8241_9883.n3 0.764
R12968 a_19345_21663.t7 a_19345_21663.t4 574.43
R12969 a_19345_21663.n0 a_19345_21663.t5 285.109
R12970 a_19345_21663.n2 a_19345_21663.n1 211.134
R12971 a_19345_21663.n4 a_19345_21663.n3 192.754
R12972 a_19345_21663.n0 a_19345_21663.t6 160.666
R12973 a_19345_21663.n1 a_19345_21663.t7 160.666
R12974 a_19345_21663.n1 a_19345_21663.n0 114.829
R12975 a_19345_21663.n3 a_19345_21663.t1 28.568
R12976 a_19345_21663.n4 a_19345_21663.t2 28.565
R12977 a_19345_21663.t3 a_19345_21663.n4 28.565
R12978 a_19345_21663.n2 a_19345_21663.t0 19.087
R12979 a_19345_21663.n3 a_19345_21663.n2 1.051
R12980 a_25332_10690.n1 a_25332_10690.t5 318.922
R12981 a_25332_10690.n0 a_25332_10690.t7 273.935
R12982 a_25332_10690.n0 a_25332_10690.t6 273.935
R12983 a_25332_10690.n1 a_25332_10690.t4 269.116
R12984 a_25332_10690.n4 a_25332_10690.n3 193.227
R12985 a_25332_10690.t5 a_25332_10690.n0 179.142
R12986 a_25332_10690.n2 a_25332_10690.n1 106.999
R12987 a_25332_10690.n3 a_25332_10690.t1 28.568
R12988 a_25332_10690.n4 a_25332_10690.t2 28.565
R12989 a_25332_10690.t3 a_25332_10690.n4 28.565
R12990 a_25332_10690.n2 a_25332_10690.t0 18.149
R12991 a_25332_10690.n3 a_25332_10690.n2 3.726
R12992 a_8183_9177.t0 a_8183_9177.t1 17.4
R12993 a_27439_12833.n0 a_27439_12833.t0 14.282
R12994 a_27439_12833.n0 a_27439_12833.t1 14.282
R12995 a_27439_12833.n1 a_27439_12833.t3 14.282
R12996 a_27439_12833.n1 a_27439_12833.t4 14.282
R12997 a_27439_12833.n3 a_27439_12833.t5 14.282
R12998 a_27439_12833.t2 a_27439_12833.n3 14.282
R12999 a_27439_12833.n2 a_27439_12833.n0 2.546
R13000 a_27439_12833.n2 a_27439_12833.n1 2.367
R13001 a_27439_12833.n3 a_27439_12833.n2 0.001
R13002 a_38088_11336.t0 a_38088_11336.t1 17.4
R13003 a_20814_12765.n0 a_20814_12765.t5 14.282
R13004 a_20814_12765.n0 a_20814_12765.t2 14.282
R13005 a_20814_12765.n1 a_20814_12765.t3 14.282
R13006 a_20814_12765.n1 a_20814_12765.t4 14.282
R13007 a_20814_12765.t0 a_20814_12765.n3 14.282
R13008 a_20814_12765.n3 a_20814_12765.t1 14.282
R13009 a_20814_12765.n3 a_20814_12765.n2 2.546
R13010 a_20814_12765.n2 a_20814_12765.n1 2.367
R13011 a_20814_12765.n2 a_20814_12765.n0 0.001
R13012 a_38088_20814.t0 a_38088_20814.t1 17.4
R13013 a_10707_11307.n4 a_10707_11307.t9 214.335
R13014 a_10707_11307.t7 a_10707_11307.n4 214.335
R13015 a_10707_11307.n5 a_10707_11307.t7 143.851
R13016 a_10707_11307.n5 a_10707_11307.t10 135.658
R13017 a_10707_11307.n4 a_10707_11307.t8 80.333
R13018 a_10707_11307.n0 a_10707_11307.t5 28.565
R13019 a_10707_11307.n0 a_10707_11307.t6 28.565
R13020 a_10707_11307.n2 a_10707_11307.t0 28.565
R13021 a_10707_11307.n2 a_10707_11307.t4 28.565
R13022 a_10707_11307.n7 a_10707_11307.t1 28.565
R13023 a_10707_11307.t2 a_10707_11307.n7 28.565
R13024 a_10707_11307.n1 a_10707_11307.t3 9.714
R13025 a_10707_11307.n1 a_10707_11307.n0 1.003
R13026 a_10707_11307.n6 a_10707_11307.n3 0.833
R13027 a_10707_11307.n3 a_10707_11307.n2 0.653
R13028 a_10707_11307.n7 a_10707_11307.n6 0.653
R13029 a_10707_11307.n3 a_10707_11307.n1 0.341
R13030 a_10707_11307.n6 a_10707_11307.n5 0.032
R13031 a_10944_10670.t0 a_10944_10670.t1 17.4
R13032 a_13421_19541.n1 a_13421_19541.t6 318.922
R13033 a_13421_19541.n0 a_13421_19541.t5 274.739
R13034 a_13421_19541.n0 a_13421_19541.t7 274.739
R13035 a_13421_19541.n1 a_13421_19541.t4 269.116
R13036 a_13421_19541.t6 a_13421_19541.n0 179.946
R13037 a_13421_19541.n2 a_13421_19541.n1 107.263
R13038 a_13421_19541.t3 a_13421_19541.n4 29.444
R13039 a_13421_19541.n3 a_13421_19541.t1 28.565
R13040 a_13421_19541.n3 a_13421_19541.t2 28.565
R13041 a_13421_19541.n2 a_13421_19541.t0 18.145
R13042 a_13421_19541.n4 a_13421_19541.n2 2.878
R13043 a_13421_19541.n4 a_13421_19541.n3 0.764
R13044 a_14079_18116.t0 a_14079_18116.t1 380.209
R13045 a_12461_27417.n0 a_12461_27417.t10 214.335
R13046 a_12461_27417.t8 a_12461_27417.n0 214.335
R13047 a_12461_27417.n1 a_12461_27417.t8 143.851
R13048 a_12461_27417.n1 a_12461_27417.t7 135.658
R13049 a_12461_27417.n0 a_12461_27417.t9 80.333
R13050 a_12461_27417.n2 a_12461_27417.t4 28.565
R13051 a_12461_27417.n2 a_12461_27417.t5 28.565
R13052 a_12461_27417.n4 a_12461_27417.t6 28.565
R13053 a_12461_27417.n4 a_12461_27417.t2 28.565
R13054 a_12461_27417.t3 a_12461_27417.n7 28.565
R13055 a_12461_27417.n7 a_12461_27417.t1 28.565
R13056 a_12461_27417.n6 a_12461_27417.t0 9.714
R13057 a_12461_27417.n7 a_12461_27417.n6 1.003
R13058 a_12461_27417.n5 a_12461_27417.n3 0.833
R13059 a_12461_27417.n3 a_12461_27417.n2 0.653
R13060 a_12461_27417.n5 a_12461_27417.n4 0.653
R13061 a_12461_27417.n6 a_12461_27417.n5 0.341
R13062 a_12461_27417.n3 a_12461_27417.n1 0.032
R13063 a_29844_1450.n4 a_29844_1450.t8 214.335
R13064 a_29844_1450.t9 a_29844_1450.n4 214.335
R13065 a_29844_1450.n5 a_29844_1450.t9 143.851
R13066 a_29844_1450.n5 a_29844_1450.t10 135.658
R13067 a_29844_1450.n4 a_29844_1450.t7 80.333
R13068 a_29844_1450.n0 a_29844_1450.t4 28.565
R13069 a_29844_1450.n0 a_29844_1450.t6 28.565
R13070 a_29844_1450.n2 a_29844_1450.t0 28.565
R13071 a_29844_1450.n2 a_29844_1450.t5 28.565
R13072 a_29844_1450.t2 a_29844_1450.n7 28.565
R13073 a_29844_1450.n7 a_29844_1450.t1 28.565
R13074 a_29844_1450.n1 a_29844_1450.t3 9.714
R13075 a_29844_1450.n1 a_29844_1450.n0 1.003
R13076 a_29844_1450.n6 a_29844_1450.n3 0.833
R13077 a_29844_1450.n3 a_29844_1450.n2 0.653
R13078 a_29844_1450.n7 a_29844_1450.n6 0.653
R13079 a_29844_1450.n3 a_29844_1450.n1 0.341
R13080 a_29844_1450.n6 a_29844_1450.n5 0.032
R13081 a_17937_12452.t7 a_17937_12452.t5 800.071
R13082 a_17937_12452.n2 a_17937_12452.n1 659.097
R13083 a_17937_12452.n0 a_17937_12452.t6 285.109
R13084 a_17937_12452.n1 a_17937_12452.t7 193.602
R13085 a_17937_12452.n4 a_17937_12452.n3 192.754
R13086 a_17937_12452.n0 a_17937_12452.t4 160.666
R13087 a_17937_12452.n1 a_17937_12452.n0 91.507
R13088 a_17937_12452.n3 a_17937_12452.t1 28.568
R13089 a_17937_12452.t0 a_17937_12452.n4 28.565
R13090 a_17937_12452.n4 a_17937_12452.t2 28.565
R13091 a_17937_12452.n2 a_17937_12452.t3 19.061
R13092 a_17937_12452.n3 a_17937_12452.n2 1.005
R13093 a_19672_12761.n0 a_19672_12761.t3 14.282
R13094 a_19672_12761.n0 a_19672_12761.t0 14.282
R13095 a_19672_12761.n1 a_19672_12761.t4 14.282
R13096 a_19672_12761.n1 a_19672_12761.t5 14.282
R13097 a_19672_12761.n3 a_19672_12761.t1 14.282
R13098 a_19672_12761.t2 a_19672_12761.n3 14.282
R13099 a_19672_12761.n3 a_19672_12761.n2 2.546
R13100 a_19672_12761.n2 a_19672_12761.n1 2.367
R13101 a_19672_12761.n2 a_19672_12761.n0 0.001
R13102 Y[4].n1 Y[4].n0 185.55
R13103 Y[4].n1 Y[4].t3 28.568
R13104 Y[4].n0 Y[4].t1 28.565
R13105 Y[4].n0 Y[4].t2 28.565
R13106 Y[4].n2 Y[4].t0 20.393
R13107 Y[4].n2 Y[4].n1 1.835
R13108 Y[4].n3 Y[4].n2 1.048
R13109 Y[4] Y[4].n3 0.052
R13110 Y[4].n3 Y[4] 0.046
R13111 a_17593_8998.t0 a_17593_8998.t1 17.4
R13112 a_6461_6961.n0 a_6461_6961.t4 14.282
R13113 a_6461_6961.n0 a_6461_6961.t0 14.282
R13114 a_6461_6961.n1 a_6461_6961.t3 14.282
R13115 a_6461_6961.n1 a_6461_6961.t5 14.282
R13116 a_6461_6961.t2 a_6461_6961.n3 14.282
R13117 a_6461_6961.n3 a_6461_6961.t1 14.282
R13118 a_6461_6961.n3 a_6461_6961.n2 2.546
R13119 a_6461_6961.n2 a_6461_6961.n1 2.367
R13120 a_6461_6961.n2 a_6461_6961.n0 0.001
R13121 a_13018_12829.n1 a_13018_12829.t5 14.282
R13122 a_13018_12829.n1 a_13018_12829.t2 14.282
R13123 a_13018_12829.n0 a_13018_12829.t3 14.282
R13124 a_13018_12829.n0 a_13018_12829.t1 14.282
R13125 a_13018_12829.n3 a_13018_12829.t4 14.282
R13126 a_13018_12829.t0 a_13018_12829.n3 14.282
R13127 a_13018_12829.n2 a_13018_12829.n0 2.546
R13128 a_13018_12829.n3 a_13018_12829.n2 2.367
R13129 a_13018_12829.n2 a_13018_12829.n1 0.001
R13130 a_20691_6964.t8 a_20691_6964.n2 404.877
R13131 a_20691_6964.n1 a_20691_6964.t6 210.902
R13132 a_20691_6964.n3 a_20691_6964.t8 136.943
R13133 a_20691_6964.n2 a_20691_6964.n1 107.801
R13134 a_20691_6964.n1 a_20691_6964.t7 80.333
R13135 a_20691_6964.n2 a_20691_6964.t5 80.333
R13136 a_20691_6964.n0 a_20691_6964.t4 17.4
R13137 a_20691_6964.n0 a_20691_6964.t2 17.4
R13138 a_20691_6964.n4 a_20691_6964.t1 15.032
R13139 a_20691_6964.t0 a_20691_6964.n5 14.282
R13140 a_20691_6964.n5 a_20691_6964.t3 14.282
R13141 a_20691_6964.n5 a_20691_6964.n4 1.65
R13142 a_20691_6964.n3 a_20691_6964.n0 0.672
R13143 a_20691_6964.n4 a_20691_6964.n3 0.665
R13144 a_10933_3196.t0 a_10933_3196.t1 17.4
R13145 a_25869_4129.n8 a_25869_4129.n6 552.333
R13146 a_25869_4129.n4 a_25869_4129.t9 394.151
R13147 a_25869_4129.n9 a_25869_4129.n8 342.688
R13148 a_25869_4129.n7 a_25869_4129.t15 294.653
R13149 a_25869_4129.n3 a_25869_4129.t11 269.523
R13150 a_25869_4129.t9 a_25869_4129.n3 269.523
R13151 a_25869_4129.n5 a_25869_4129.t13 198.043
R13152 a_25869_4129.n3 a_25869_4129.t14 160.666
R13153 a_25869_4129.n11 a_25869_4129.n0 157.665
R13154 a_25869_4129.n8 a_25869_4129.n7 126.566
R13155 a_25869_4129.n12 a_25869_4129.n11 122.999
R13156 a_25869_4129.n7 a_25869_4129.t8 111.663
R13157 a_25869_4129.n6 a_25869_4129.n4 97.816
R13158 a_25869_4129.n5 a_25869_4129.t10 93.989
R13159 a_25869_4129.n9 a_25869_4129.n2 90.436
R13160 a_25869_4129.n10 a_25869_4129.n1 90.416
R13161 a_25869_4129.n4 a_25869_4129.t12 80.333
R13162 a_25869_4129.n10 a_25869_4129.n9 74.302
R13163 a_25869_4129.n11 a_25869_4129.n10 50.575
R13164 a_25869_4129.n2 a_25869_4129.t4 14.282
R13165 a_25869_4129.n2 a_25869_4129.t6 14.282
R13166 a_25869_4129.n1 a_25869_4129.t5 14.282
R13167 a_25869_4129.n1 a_25869_4129.t1 14.282
R13168 a_25869_4129.n12 a_25869_4129.t2 14.282
R13169 a_25869_4129.t3 a_25869_4129.n12 14.282
R13170 a_25869_4129.n0 a_25869_4129.t7 8.7
R13171 a_25869_4129.n0 a_25869_4129.t0 8.7
R13172 a_25869_4129.n6 a_25869_4129.n5 6.615
R13173 a_27657_9997.n2 a_27657_9997.n0 267.767
R13174 a_27657_9997.n8 a_27657_9997.t1 16.058
R13175 a_27657_9997.n6 a_27657_9997.t9 16.058
R13176 a_27657_9997.n1 a_27657_9997.t8 14.282
R13177 a_27657_9997.n1 a_27657_9997.t3 14.282
R13178 a_27657_9997.n0 a_27657_9997.t6 14.282
R13179 a_27657_9997.n0 a_27657_9997.t7 14.282
R13180 a_27657_9997.n3 a_27657_9997.t4 14.282
R13181 a_27657_9997.n3 a_27657_9997.t5 14.282
R13182 a_27657_9997.n5 a_27657_9997.t11 14.282
R13183 a_27657_9997.n5 a_27657_9997.t10 14.282
R13184 a_27657_9997.n9 a_27657_9997.t0 14.282
R13185 a_27657_9997.t2 a_27657_9997.n9 14.282
R13186 a_27657_9997.n4 a_27657_9997.n3 1.511
R13187 a_27657_9997.n6 a_27657_9997.n5 0.999
R13188 a_27657_9997.n9 a_27657_9997.n8 0.999
R13189 a_27657_9997.n4 a_27657_9997.n2 0.669
R13190 a_27657_9997.n8 a_27657_9997.n7 0.575
R13191 a_27657_9997.n7 a_27657_9997.n4 0.227
R13192 a_27657_9997.n7 a_27657_9997.n6 0.2
R13193 a_27657_9997.n2 a_27657_9997.n1 0.001
R13194 a_21358_14419.t0 a_21358_14419.t1 17.4
R13195 a_14315_18116.t0 a_14315_18116.t1 17.4
R13196 a_23972_12957.n0 a_23972_12957.t8 214.335
R13197 a_23972_12957.t10 a_23972_12957.n0 214.335
R13198 a_23972_12957.n1 a_23972_12957.t10 143.851
R13199 a_23972_12957.n1 a_23972_12957.t9 135.658
R13200 a_23972_12957.n0 a_23972_12957.t7 80.333
R13201 a_23972_12957.n2 a_23972_12957.t4 28.565
R13202 a_23972_12957.n2 a_23972_12957.t5 28.565
R13203 a_23972_12957.n4 a_23972_12957.t6 28.565
R13204 a_23972_12957.n4 a_23972_12957.t1 28.565
R13205 a_23972_12957.t3 a_23972_12957.n7 28.565
R13206 a_23972_12957.n7 a_23972_12957.t2 28.565
R13207 a_23972_12957.n6 a_23972_12957.t0 9.714
R13208 a_23972_12957.n7 a_23972_12957.n6 1.003
R13209 a_23972_12957.n5 a_23972_12957.n3 0.833
R13210 a_23972_12957.n3 a_23972_12957.n2 0.653
R13211 a_23972_12957.n5 a_23972_12957.n4 0.653
R13212 a_23972_12957.n6 a_23972_12957.n5 0.341
R13213 a_23972_12957.n3 a_23972_12957.n1 0.032
R13214 a_n3606_2123.n1 a_n3606_2123.t5 318.119
R13215 a_n3606_2123.n1 a_n3606_2123.t6 269.919
R13216 a_n3606_2123.n0 a_n3606_2123.t7 267.853
R13217 a_n3606_2123.n0 a_n3606_2123.t4 267.853
R13218 a_n3606_2123.t5 a_n3606_2123.n0 160.666
R13219 a_n3606_2123.n2 a_n3606_2123.n1 107.263
R13220 a_n3606_2123.t3 a_n3606_2123.n4 29.444
R13221 a_n3606_2123.n3 a_n3606_2123.t1 28.565
R13222 a_n3606_2123.n3 a_n3606_2123.t2 28.565
R13223 a_n3606_2123.n2 a_n3606_2123.t0 18.145
R13224 a_n3606_2123.n4 a_n3606_2123.n2 2.878
R13225 a_n3606_2123.n4 a_n3606_2123.n3 0.764
R13226 a_1464_6636.t0 a_1464_6636.t1 17.4
R13227 a_17347_12889.n4 a_17347_12889.t10 214.335
R13228 a_17347_12889.t8 a_17347_12889.n4 214.335
R13229 a_17347_12889.n5 a_17347_12889.t8 143.851
R13230 a_17347_12889.n5 a_17347_12889.t7 135.658
R13231 a_17347_12889.n4 a_17347_12889.t9 80.333
R13232 a_17347_12889.n0 a_17347_12889.t5 28.565
R13233 a_17347_12889.n0 a_17347_12889.t6 28.565
R13234 a_17347_12889.n2 a_17347_12889.t0 28.565
R13235 a_17347_12889.n2 a_17347_12889.t4 28.565
R13236 a_17347_12889.n7 a_17347_12889.t1 28.565
R13237 a_17347_12889.t2 a_17347_12889.n7 28.565
R13238 a_17347_12889.n1 a_17347_12889.t3 9.714
R13239 a_17347_12889.n1 a_17347_12889.n0 1.003
R13240 a_17347_12889.n6 a_17347_12889.n3 0.833
R13241 a_17347_12889.n3 a_17347_12889.n2 0.653
R13242 a_17347_12889.n7 a_17347_12889.n6 0.653
R13243 a_17347_12889.n3 a_17347_12889.n1 0.341
R13244 a_17347_12889.n6 a_17347_12889.n5 0.032
R13245 a_14366_24457.n8 a_14366_24457.n6 552.333
R13246 a_14366_24457.n4 a_14366_24457.t15 394.151
R13247 a_14366_24457.n9 a_14366_24457.n8 342.688
R13248 a_14366_24457.n7 a_14366_24457.t12 294.653
R13249 a_14366_24457.n3 a_14366_24457.t9 269.523
R13250 a_14366_24457.t15 a_14366_24457.n3 269.523
R13251 a_14366_24457.n5 a_14366_24457.t10 198.043
R13252 a_14366_24457.n3 a_14366_24457.t8 160.666
R13253 a_14366_24457.n11 a_14366_24457.n0 157.665
R13254 a_14366_24457.n8 a_14366_24457.n7 126.566
R13255 a_14366_24457.n12 a_14366_24457.n11 122.999
R13256 a_14366_24457.n7 a_14366_24457.t14 111.663
R13257 a_14366_24457.n6 a_14366_24457.n4 97.816
R13258 a_14366_24457.n5 a_14366_24457.t11 93.989
R13259 a_14366_24457.n9 a_14366_24457.n2 90.436
R13260 a_14366_24457.n10 a_14366_24457.n1 90.416
R13261 a_14366_24457.n4 a_14366_24457.t13 80.333
R13262 a_14366_24457.n10 a_14366_24457.n9 74.302
R13263 a_14366_24457.n11 a_14366_24457.n10 50.575
R13264 a_14366_24457.n2 a_14366_24457.t4 14.282
R13265 a_14366_24457.n2 a_14366_24457.t5 14.282
R13266 a_14366_24457.n1 a_14366_24457.t6 14.282
R13267 a_14366_24457.n1 a_14366_24457.t1 14.282
R13268 a_14366_24457.n12 a_14366_24457.t2 14.282
R13269 a_14366_24457.t3 a_14366_24457.n12 14.282
R13270 a_14366_24457.n0 a_14366_24457.t7 8.7
R13271 a_14366_24457.n0 a_14366_24457.t0 8.7
R13272 a_14366_24457.n6 a_14366_24457.n5 6.615
R13273 a_17584_12252.t0 a_17584_12252.t1 17.4
R13274 a_20782_24452.t3 a_20782_24452.n0 14.282
R13275 a_20782_24452.n0 a_20782_24452.t4 14.282
R13276 a_20782_24452.n0 a_20782_24452.n9 0.999
R13277 a_20782_24452.n6 a_20782_24452.n8 0.575
R13278 a_20782_24452.n9 a_20782_24452.n6 0.2
R13279 a_20782_24452.n9 a_20782_24452.t5 16.058
R13280 a_20782_24452.n8 a_20782_24452.n7 0.999
R13281 a_20782_24452.n7 a_20782_24452.t9 14.282
R13282 a_20782_24452.n7 a_20782_24452.t10 14.282
R13283 a_20782_24452.n8 a_20782_24452.t11 16.058
R13284 a_20782_24452.n6 a_20782_24452.n4 0.227
R13285 a_20782_24452.n4 a_20782_24452.n5 1.511
R13286 a_20782_24452.n5 a_20782_24452.t2 14.282
R13287 a_20782_24452.n5 a_20782_24452.t1 14.282
R13288 a_20782_24452.n4 a_20782_24452.n1 0.669
R13289 a_20782_24452.n1 a_20782_24452.n2 0.001
R13290 a_20782_24452.n1 a_20782_24452.n3 267.767
R13291 a_20782_24452.n3 a_20782_24452.t7 14.282
R13292 a_20782_24452.n3 a_20782_24452.t6 14.282
R13293 a_20782_24452.n2 a_20782_24452.t0 14.282
R13294 a_20782_24452.n2 a_20782_24452.t8 14.282
R13295 a_n2383_4850.t0 a_n2383_4850.t1 379.845
R13296 a_28011_9265.t0 a_28011_9265.t1 17.4
R13297 B[2].n4 B[2].n0 592.056
R13298 B[2].t1 B[2].n2 313.069
R13299 B[2].n0 B[2].t4 294.986
R13300 B[2].n1 B[2].t0 271.484
R13301 B[2].n4 B[2].t6 204.672
R13302 B[2].n3 B[2].t1 190.955
R13303 B[2].n3 B[2].t3 190.955
R13304 B[2].n2 B[2].t2 160.666
R13305 B[2].n1 B[2].t5 160.666
R13306 B[2].n0 B[2].t7 110.859
R13307 B[2].n2 B[2].n1 96.129
R13308 B[2].t6 B[2].n3 80.333
R13309 B[2] B[2].n4 60.44
R13310 a_16205_19521.t0 a_16205_19521.t1 17.4
R13311 a_29356_23724.t0 a_29356_23724.t1 380.209
R13312 a_12457_21658.t7 a_12457_21658.t4 800.071
R13313 a_12457_21658.n3 a_12457_21658.n2 672.95
R13314 a_12457_21658.n1 a_12457_21658.t5 285.109
R13315 a_12457_21658.n2 a_12457_21658.t7 193.602
R13316 a_12457_21658.n1 a_12457_21658.t6 160.666
R13317 a_12457_21658.n2 a_12457_21658.n1 91.507
R13318 a_12457_21658.n0 a_12457_21658.t1 28.57
R13319 a_12457_21658.n4 a_12457_21658.t2 28.565
R13320 a_12457_21658.t3 a_12457_21658.n4 28.565
R13321 a_12457_21658.n0 a_12457_21658.t0 17.638
R13322 a_12457_21658.n4 a_12457_21658.n3 0.693
R13323 a_12457_21658.n3 a_12457_21658.n0 0.597
R13324 a_6199_25133.t0 a_6199_25133.t1 17.4
R13325 a_25877_9265.t0 a_25877_9265.t1 380.209
R13326 a_9633_24460.n8 a_9633_24460.n0 267.767
R13327 a_9633_24460.n4 a_9633_24460.t6 16.058
R13328 a_9633_24460.n2 a_9633_24460.t9 16.058
R13329 a_9633_24460.n3 a_9633_24460.t7 14.282
R13330 a_9633_24460.n3 a_9633_24460.t8 14.282
R13331 a_9633_24460.n1 a_9633_24460.t10 14.282
R13332 a_9633_24460.n1 a_9633_24460.t11 14.282
R13333 a_9633_24460.n6 a_9633_24460.t4 14.282
R13334 a_9633_24460.n6 a_9633_24460.t5 14.282
R13335 a_9633_24460.n0 a_9633_24460.t0 14.282
R13336 a_9633_24460.n0 a_9633_24460.t1 14.282
R13337 a_9633_24460.t2 a_9633_24460.n9 14.282
R13338 a_9633_24460.n9 a_9633_24460.t3 14.282
R13339 a_9633_24460.n7 a_9633_24460.n6 1.511
R13340 a_9633_24460.n4 a_9633_24460.n3 0.999
R13341 a_9633_24460.n2 a_9633_24460.n1 0.999
R13342 a_9633_24460.n8 a_9633_24460.n7 0.669
R13343 a_9633_24460.n5 a_9633_24460.n4 0.575
R13344 a_9633_24460.n7 a_9633_24460.n5 0.227
R13345 a_9633_24460.n5 a_9633_24460.n2 0.2
R13346 a_9633_24460.n9 a_9633_24460.n8 0.001
R13347 a_14366_23725.t0 a_14366_23725.t1 380.209
R13348 a_38084_14302.t0 a_38084_14302.t1 17.4
R13349 a_32247_1125.t0 a_32247_1125.t1 17.4
R13350 a_19483_3396.t0 a_19483_3396.t1 17.4
R13351 a_26113_9265.t0 a_26113_9265.t1 17.4
R13352 a_11297_10870.t4 a_11297_10870.t5 574.43
R13353 a_11297_10870.n0 a_11297_10870.t7 285.109
R13354 a_11297_10870.n2 a_11297_10870.n1 211.136
R13355 a_11297_10870.n4 a_11297_10870.n3 192.754
R13356 a_11297_10870.n0 a_11297_10870.t6 160.666
R13357 a_11297_10870.n1 a_11297_10870.t4 160.666
R13358 a_11297_10870.n1 a_11297_10870.n0 114.829
R13359 a_11297_10870.n3 a_11297_10870.t1 28.568
R13360 a_11297_10870.n4 a_11297_10870.t2 28.565
R13361 a_11297_10870.t3 a_11297_10870.n4 28.565
R13362 a_11297_10870.n2 a_11297_10870.t0 19.084
R13363 a_11297_10870.n3 a_11297_10870.n2 1.051
R13364 a_14042_12833.t5 a_14042_12833.n2 404.877
R13365 a_14042_12833.n1 a_14042_12833.t8 210.902
R13366 a_14042_12833.n3 a_14042_12833.t5 136.943
R13367 a_14042_12833.n2 a_14042_12833.n1 107.801
R13368 a_14042_12833.n1 a_14042_12833.t7 80.333
R13369 a_14042_12833.n2 a_14042_12833.t6 80.333
R13370 a_14042_12833.n0 a_14042_12833.t0 17.4
R13371 a_14042_12833.n0 a_14042_12833.t2 17.4
R13372 a_14042_12833.n4 a_14042_12833.t3 15.032
R13373 a_14042_12833.t1 a_14042_12833.n5 14.282
R13374 a_14042_12833.n5 a_14042_12833.t4 14.282
R13375 a_14042_12833.n5 a_14042_12833.n4 1.65
R13376 a_14042_12833.n3 a_14042_12833.n0 0.672
R13377 a_14042_12833.n4 a_14042_12833.n3 0.665
R13378 a_14160_12833.n0 a_14160_12833.t4 14.282
R13379 a_14160_12833.n0 a_14160_12833.t5 14.282
R13380 a_14160_12833.n1 a_14160_12833.t0 14.282
R13381 a_14160_12833.n1 a_14160_12833.t1 14.282
R13382 a_14160_12833.t2 a_14160_12833.n3 14.282
R13383 a_14160_12833.n3 a_14160_12833.t3 14.282
R13384 a_14160_12833.n2 a_14160_12833.n0 2.546
R13385 a_14160_12833.n2 a_14160_12833.n1 2.367
R13386 a_14160_12833.n3 a_14160_12833.n2 0.001
R13387 a_11283_12520.t5 a_11283_12520.t4 800.071
R13388 a_11283_12520.n2 a_11283_12520.n1 659.097
R13389 a_11283_12520.n0 a_11283_12520.t7 285.109
R13390 a_11283_12520.n1 a_11283_12520.t5 193.602
R13391 a_11283_12520.n4 a_11283_12520.n3 192.754
R13392 a_11283_12520.n0 a_11283_12520.t6 160.666
R13393 a_11283_12520.n1 a_11283_12520.n0 91.507
R13394 a_11283_12520.n3 a_11283_12520.t1 28.568
R13395 a_11283_12520.n4 a_11283_12520.t2 28.565
R13396 a_11283_12520.t3 a_11283_12520.n4 28.565
R13397 a_11283_12520.n2 a_11283_12520.t0 19.061
R13398 a_11283_12520.n3 a_11283_12520.n2 1.005
R13399 a_6538_26983.t6 a_6538_26983.t4 800.071
R13400 a_6538_26983.n2 a_6538_26983.n1 659.097
R13401 a_6538_26983.n0 a_6538_26983.t5 285.109
R13402 a_6538_26983.n1 a_6538_26983.t6 193.602
R13403 a_6538_26983.n4 a_6538_26983.n3 192.754
R13404 a_6538_26983.n0 a_6538_26983.t7 160.666
R13405 a_6538_26983.n1 a_6538_26983.n0 91.507
R13406 a_6538_26983.n3 a_6538_26983.t1 28.568
R13407 a_6538_26983.n4 a_6538_26983.t2 28.565
R13408 a_6538_26983.t3 a_6538_26983.n4 28.565
R13409 a_6538_26983.n2 a_6538_26983.t0 19.061
R13410 a_6538_26983.n3 a_6538_26983.n2 1.005
R13411 a_6185_26783.t0 a_6185_26783.t1 17.4
R13412 a_5859_18120.t0 a_5859_18120.t1 17.4
R13413 a_27767_3397.t0 a_27767_3397.t1 380.209
R13414 a_7757_18120.t0 a_7757_18120.t1 17.4
R13415 a_4382_3198.t0 a_4382_3198.t1 17.4
R13416 a_18702_4821.n1 a_18702_4821.t7 318.922
R13417 a_18702_4821.n0 a_18702_4821.t4 273.935
R13418 a_18702_4821.n0 a_18702_4821.t5 273.935
R13419 a_18702_4821.n1 a_18702_4821.t6 269.116
R13420 a_18702_4821.n4 a_18702_4821.n3 193.227
R13421 a_18702_4821.t7 a_18702_4821.n0 179.142
R13422 a_18702_4821.n2 a_18702_4821.n1 106.999
R13423 a_18702_4821.n3 a_18702_4821.t2 28.568
R13424 a_18702_4821.n4 a_18702_4821.t1 28.565
R13425 a_18702_4821.t3 a_18702_4821.n4 28.565
R13426 a_18702_4821.n2 a_18702_4821.t0 18.149
R13427 a_18702_4821.n3 a_18702_4821.n2 3.726
R13428 a_17946_5001.t4 a_17946_5001.t6 574.43
R13429 a_17946_5001.n0 a_17946_5001.t5 285.109
R13430 a_17946_5001.n2 a_17946_5001.n1 211.136
R13431 a_17946_5001.n4 a_17946_5001.n3 192.754
R13432 a_17946_5001.n0 a_17946_5001.t7 160.666
R13433 a_17946_5001.n1 a_17946_5001.t4 160.666
R13434 a_17946_5001.n1 a_17946_5001.n0 114.829
R13435 a_17946_5001.n3 a_17946_5001.t1 28.568
R13436 a_17946_5001.t3 a_17946_5001.n4 28.565
R13437 a_17946_5001.n4 a_17946_5001.t2 28.565
R13438 a_17946_5001.n2 a_17946_5001.t0 19.084
R13439 a_17946_5001.n3 a_17946_5001.n2 1.051
R13440 a_9297_27296.t6 a_9297_27296.n3 404.877
R13441 a_9297_27296.n2 a_9297_27296.t8 210.902
R13442 a_9297_27296.n4 a_9297_27296.t6 136.943
R13443 a_9297_27296.n3 a_9297_27296.n2 107.801
R13444 a_9297_27296.n2 a_9297_27296.t7 80.333
R13445 a_9297_27296.n3 a_9297_27296.t5 80.333
R13446 a_9297_27296.n1 a_9297_27296.t0 17.4
R13447 a_9297_27296.n1 a_9297_27296.t1 17.4
R13448 a_9297_27296.t4 a_9297_27296.n5 15.032
R13449 a_9297_27296.n0 a_9297_27296.t2 14.282
R13450 a_9297_27296.n0 a_9297_27296.t3 14.282
R13451 a_9297_27296.n5 a_9297_27296.n0 1.65
R13452 a_9297_27296.n4 a_9297_27296.n1 0.672
R13453 a_9297_27296.n5 a_9297_27296.n4 0.665
R13454 Y[1].n1 Y[1].n0 185.55
R13455 Y[1].n1 Y[1].t1 28.568
R13456 Y[1].n0 Y[1].t2 28.565
R13457 Y[1].n0 Y[1].t3 28.565
R13458 Y[1].n2 Y[1].t0 20.393
R13459 Y[1].n2 Y[1].n1 1.835
R13460 Y[1].n3 Y[1].n2 1.048
R13461 Y[1] Y[1].n3 0.052
R13462 Y[1].n3 Y[1] 0.046
R13463 a_21121_15056.n0 a_21121_15056.t9 214.335
R13464 a_21121_15056.t7 a_21121_15056.n0 214.335
R13465 a_21121_15056.n1 a_21121_15056.t7 143.851
R13466 a_21121_15056.n1 a_21121_15056.t10 135.658
R13467 a_21121_15056.n0 a_21121_15056.t8 80.333
R13468 a_21121_15056.n2 a_21121_15056.t4 28.565
R13469 a_21121_15056.n2 a_21121_15056.t5 28.565
R13470 a_21121_15056.n4 a_21121_15056.t6 28.565
R13471 a_21121_15056.n4 a_21121_15056.t1 28.565
R13472 a_21121_15056.n7 a_21121_15056.t2 28.565
R13473 a_21121_15056.t3 a_21121_15056.n7 28.565
R13474 a_21121_15056.n6 a_21121_15056.t0 9.714
R13475 a_21121_15056.n7 a_21121_15056.n6 1.003
R13476 a_21121_15056.n5 a_21121_15056.n3 0.833
R13477 a_21121_15056.n3 a_21121_15056.n2 0.653
R13478 a_21121_15056.n5 a_21121_15056.n4 0.653
R13479 a_21121_15056.n6 a_21121_15056.n5 0.341
R13480 a_21121_15056.n3 a_21121_15056.n1 0.032
R13481 a_27458_23724.t0 a_27458_23724.t1 380.209
R13482 a_7918_15036.n2 a_7918_15036.t7 214.335
R13483 a_7918_15036.t9 a_7918_15036.n2 214.335
R13484 a_7918_15036.n3 a_7918_15036.t9 143.851
R13485 a_7918_15036.n3 a_7918_15036.t8 135.658
R13486 a_7918_15036.n2 a_7918_15036.t10 80.333
R13487 a_7918_15036.n4 a_7918_15036.t0 28.565
R13488 a_7918_15036.n4 a_7918_15036.t1 28.565
R13489 a_7918_15036.n0 a_7918_15036.t4 28.565
R13490 a_7918_15036.n0 a_7918_15036.t5 28.565
R13491 a_7918_15036.t2 a_7918_15036.n7 28.565
R13492 a_7918_15036.n7 a_7918_15036.t6 28.565
R13493 a_7918_15036.n1 a_7918_15036.t3 9.714
R13494 a_7918_15036.n1 a_7918_15036.n0 1.003
R13495 a_7918_15036.n6 a_7918_15036.n5 0.833
R13496 a_7918_15036.n5 a_7918_15036.n4 0.653
R13497 a_7918_15036.n7 a_7918_15036.n6 0.653
R13498 a_7918_15036.n6 a_7918_15036.n1 0.341
R13499 a_7918_15036.n5 a_7918_15036.n3 0.032
R13500 a_6049_9177.t0 a_6049_9177.t1 380.209
R13501 a_19051_21689.n0 a_19051_21689.t0 14.282
R13502 a_19051_21689.n0 a_19051_21689.t1 14.282
R13503 a_19051_21689.n1 a_19051_21689.t4 14.282
R13504 a_19051_21689.n1 a_19051_21689.t5 14.282
R13505 a_19051_21689.t2 a_19051_21689.n3 14.282
R13506 a_19051_21689.n3 a_19051_21689.t3 14.282
R13507 a_19051_21689.n2 a_19051_21689.n0 2.546
R13508 a_19051_21689.n2 a_19051_21689.n1 2.367
R13509 a_19051_21689.n3 a_19051_21689.n2 0.001
R13510 a_21320_27284.n0 a_21320_27284.t5 14.282
R13511 a_21320_27284.n0 a_21320_27284.t0 14.282
R13512 a_21320_27284.n1 a_21320_27284.t3 14.282
R13513 a_21320_27284.n1 a_21320_27284.t4 14.282
R13514 a_21320_27284.n3 a_21320_27284.t1 14.282
R13515 a_21320_27284.t2 a_21320_27284.n3 14.282
R13516 a_21320_27284.n3 a_21320_27284.n2 2.546
R13517 a_21320_27284.n2 a_21320_27284.n1 2.367
R13518 a_21320_27284.n2 a_21320_27284.n0 0.001
R13519 a_7815_18826.n1 a_7815_18826.t7 318.922
R13520 a_7815_18826.n0 a_7815_18826.t6 273.935
R13521 a_7815_18826.n0 a_7815_18826.t5 273.935
R13522 a_7815_18826.n1 a_7815_18826.t4 269.116
R13523 a_7815_18826.n4 a_7815_18826.n3 193.227
R13524 a_7815_18826.t7 a_7815_18826.n0 179.142
R13525 a_7815_18826.n2 a_7815_18826.n1 106.999
R13526 a_7815_18826.n3 a_7815_18826.t1 28.568
R13527 a_7815_18826.n4 a_7815_18826.t2 28.565
R13528 a_7815_18826.t3 a_7815_18826.n4 28.565
R13529 a_7815_18826.n2 a_7815_18826.t0 18.149
R13530 a_7815_18826.n3 a_7815_18826.n2 3.726
R13531 a_7521_18120.t0 a_7521_18120.t1 380.209
R13532 a_32009_13059.t0 a_32009_13059.t1 380.209
R13533 a_8175_3397.t0 a_8175_3397.t1 17.4
R13534 a_n2381_7154.t0 a_n2381_7154.t1 17.4
R13535 a_21393_1762.t0 a_21393_1762.t1 17.4
R13536 a_20696_12765.t5 a_20696_12765.n2 404.877
R13537 a_20696_12765.n1 a_20696_12765.t7 210.902
R13538 a_20696_12765.n3 a_20696_12765.t5 136.943
R13539 a_20696_12765.n2 a_20696_12765.n1 107.801
R13540 a_20696_12765.n1 a_20696_12765.t6 80.333
R13541 a_20696_12765.n2 a_20696_12765.t8 80.333
R13542 a_20696_12765.n0 a_20696_12765.t3 17.4
R13543 a_20696_12765.n0 a_20696_12765.t4 17.4
R13544 a_20696_12765.n4 a_20696_12765.t1 15.032
R13545 a_20696_12765.n5 a_20696_12765.t2 14.282
R13546 a_20696_12765.t0 a_20696_12765.n5 14.282
R13547 a_20696_12765.n5 a_20696_12765.n4 1.65
R13548 a_20696_12765.n3 a_20696_12765.n0 0.672
R13549 a_20696_12765.n4 a_20696_12765.n3 0.665
R13550 a_27694_23724.t0 a_27694_23724.t1 17.4
R13551 a_6547_23729.t5 a_6547_23729.t4 574.43
R13552 a_6547_23729.n0 a_6547_23729.t7 285.109
R13553 a_6547_23729.n2 a_6547_23729.n1 197.217
R13554 a_6547_23729.n4 a_6547_23729.n3 192.754
R13555 a_6547_23729.n0 a_6547_23729.t6 160.666
R13556 a_6547_23729.n1 a_6547_23729.t5 160.666
R13557 a_6547_23729.n1 a_6547_23729.n0 114.829
R13558 a_6547_23729.n3 a_6547_23729.t1 28.568
R13559 a_6547_23729.n4 a_6547_23729.t2 28.565
R13560 a_6547_23729.t3 a_6547_23729.n4 28.565
R13561 a_6547_23729.n2 a_6547_23729.t0 18.838
R13562 a_6547_23729.n3 a_6547_23729.n2 1.129
R13563 a_8155_27292.t7 a_8155_27292.n2 404.877
R13564 a_8155_27292.n1 a_8155_27292.t8 210.902
R13565 a_8155_27292.n3 a_8155_27292.t7 136.943
R13566 a_8155_27292.n2 a_8155_27292.n1 107.801
R13567 a_8155_27292.n1 a_8155_27292.t6 80.333
R13568 a_8155_27292.n2 a_8155_27292.t5 80.333
R13569 a_8155_27292.n0 a_8155_27292.t0 17.4
R13570 a_8155_27292.n0 a_8155_27292.t2 17.4
R13571 a_8155_27292.n4 a_8155_27292.t4 15.032
R13572 a_8155_27292.t1 a_8155_27292.n5 14.282
R13573 a_8155_27292.n5 a_8155_27292.t3 14.282
R13574 a_8155_27292.n5 a_8155_27292.n4 1.65
R13575 a_8155_27292.n3 a_8155_27292.n0 0.672
R13576 a_8155_27292.n4 a_8155_27292.n3 0.665
R13577 a_18951_18121.t0 a_18951_18121.t1 17.4
R13578 a_13659_21680.n0 a_13659_21680.t1 14.282
R13579 a_13659_21680.n0 a_13659_21680.t3 14.282
R13580 a_13659_21680.n1 a_13659_21680.t4 14.282
R13581 a_13659_21680.n1 a_13659_21680.t5 14.282
R13582 a_13659_21680.n3 a_13659_21680.t0 14.282
R13583 a_13659_21680.t2 a_13659_21680.n3 14.282
R13584 a_13659_21680.n3 a_13659_21680.n2 2.546
R13585 a_13659_21680.n2 a_13659_21680.n1 2.367
R13586 a_13659_21680.n2 a_13659_21680.n0 0.001
R13587 a_25429_21036.t8 a_25429_21036.n2 404.877
R13588 a_25429_21036.n1 a_25429_21036.t5 210.902
R13589 a_25429_21036.n3 a_25429_21036.t8 136.949
R13590 a_25429_21036.n2 a_25429_21036.n1 107.801
R13591 a_25429_21036.n1 a_25429_21036.t6 80.333
R13592 a_25429_21036.n2 a_25429_21036.t7 80.333
R13593 a_25429_21036.n0 a_25429_21036.t1 17.4
R13594 a_25429_21036.n0 a_25429_21036.t0 17.4
R13595 a_25429_21036.n4 a_25429_21036.t3 15.032
R13596 a_25429_21036.t2 a_25429_21036.n5 14.282
R13597 a_25429_21036.n5 a_25429_21036.t4 14.282
R13598 a_25429_21036.n5 a_25429_21036.n4 1.65
R13599 a_25429_21036.n3 a_25429_21036.n0 0.657
R13600 a_25429_21036.n4 a_25429_21036.n3 0.614
R13601 a_32245_13059.t0 a_32245_13059.t1 17.4
R13602 a_22753_21176.t0 a_22753_21176.t1 17.4
R13603 a_32247_8968.t0 a_32247_8968.t1 17.4
R13604 a_14732_9265.t0 a_14732_9265.t1 17.4
R13605 a_1480_3876.t0 a_1480_3876.t1 17.4
R13606 a_8273_27292.n1 a_8273_27292.t1 14.282
R13607 a_8273_27292.n1 a_8273_27292.t3 14.282
R13608 a_8273_27292.n0 a_8273_27292.t4 14.282
R13609 a_8273_27292.n0 a_8273_27292.t5 14.282
R13610 a_8273_27292.t2 a_8273_27292.n3 14.282
R13611 a_8273_27292.n3 a_8273_27292.t0 14.282
R13612 a_8273_27292.n2 a_8273_27292.n0 2.546
R13613 a_8273_27292.n3 a_8273_27292.n2 2.367
R13614 a_8273_27292.n2 a_8273_27292.n1 0.001
R13615 a_19009_18827.n1 a_19009_18827.t6 318.922
R13616 a_19009_18827.n0 a_19009_18827.t5 273.935
R13617 a_19009_18827.n0 a_19009_18827.t7 273.935
R13618 a_19009_18827.n1 a_19009_18827.t4 269.116
R13619 a_19009_18827.n4 a_19009_18827.n3 193.227
R13620 a_19009_18827.t6 a_19009_18827.n0 179.142
R13621 a_19009_18827.n2 a_19009_18827.n1 106.999
R13622 a_19009_18827.n3 a_19009_18827.t1 28.568
R13623 a_19009_18827.n4 a_19009_18827.t2 28.565
R13624 a_19009_18827.t3 a_19009_18827.n4 28.565
R13625 a_19009_18827.n2 a_19009_18827.t0 18.149
R13626 a_19009_18827.n3 a_19009_18827.n2 3.726
R13627 a_18715_18121.t0 a_18715_18121.t1 380.209
R13628 a_19247_3396.t0 a_19247_3396.t1 380.209
R13629 a_27585_12250.n2 a_27585_12250.t6 989.744
R13630 a_27585_12250.n3 a_27585_12250.n2 494.286
R13631 a_27585_12250.n2 a_27585_12250.t5 408.806
R13632 a_27585_12250.n1 a_27585_12250.t7 287.241
R13633 a_27585_12250.n1 a_27585_12250.t4 287.241
R13634 a_27585_12250.t6 a_27585_12250.n1 160.666
R13635 a_27585_12250.n0 a_27585_12250.t2 28.57
R13636 a_27585_12250.t3 a_27585_12250.n4 28.565
R13637 a_27585_12250.n4 a_27585_12250.t1 28.565
R13638 a_27585_12250.n0 a_27585_12250.t0 17.638
R13639 a_27585_12250.n4 a_27585_12250.n3 0.69
R13640 a_27585_12250.n3 a_27585_12250.n0 0.6
R13641 a_32011_1125.t0 a_32011_1125.t1 380.209
R13642 a_20605_10622.n2 a_20605_10622.t7 318.922
R13643 a_20605_10622.n1 a_20605_10622.t6 273.935
R13644 a_20605_10622.n1 a_20605_10622.t4 273.935
R13645 a_20605_10622.n2 a_20605_10622.t5 269.116
R13646 a_20605_10622.n4 a_20605_10622.n0 193.227
R13647 a_20605_10622.t7 a_20605_10622.n1 179.142
R13648 a_20605_10622.n3 a_20605_10622.n2 106.999
R13649 a_20605_10622.t3 a_20605_10622.n4 28.568
R13650 a_20605_10622.n0 a_20605_10622.t1 28.565
R13651 a_20605_10622.n0 a_20605_10622.t2 28.565
R13652 a_20605_10622.n3 a_20605_10622.t0 18.149
R13653 a_20605_10622.n4 a_20605_10622.n3 3.726
R13654 a_38084_14538.t0 a_38084_14538.t1 17.4
R13655 Cout.n1 Cout.t3 28.57
R13656 Cout.n0 Cout.t1 28.565
R13657 Cout.n0 Cout.t2 28.565
R13658 Cout.n1 Cout.t0 17.638
R13659 Cout Cout.n2 7.405
R13660 Cout.n2 Cout.n0 0.693
R13661 Cout.n2 Cout.n1 0.597
R13662 a_9652_17921.t0 a_9652_17921.t1 17.4
R13663 a_14744_1774.t0 a_14744_1774.t1 17.4
R13664 a_30081_813.t0 a_30081_813.t1 17.4
R13665 a_12707_23526.t0 a_12707_23526.t1 17.4
R13666 Y[3].n1 Y[3].n0 185.55
R13667 Y[3].n1 Y[3].t1 28.568
R13668 Y[3].n0 Y[3].t2 28.565
R13669 Y[3].n0 Y[3].t3 28.565
R13670 Y[3].n2 Y[3].t0 20.393
R13671 Y[3].n2 Y[3].n1 1.832
R13672 Y[3].n3 Y[3].n2 1.05
R13673 Y[3] Y[3].n3 0.052
R13674 Y[3].n3 Y[3] 0.046
R13675 a_10939_9066.t0 a_10939_9066.t1 17.4
R13676 a_38084_1916.t0 a_38084_1916.t1 17.4
R13677 a_26105_3397.t0 a_26105_3397.t1 17.4
R13678 a_19488_9197.t0 a_19488_9197.t1 17.4
R13679 a_32247_5473.t0 a_32247_5473.t1 17.4
R13680 a_25228_18124.t0 a_25228_18124.t1 380.209
R13681 a_n2381_3017.t0 a_n2381_3017.t1 17.4
R13682 a_6277_3397.t0 a_6277_3397.t1 17.4
R13683 a_27362_18124.t0 a_27362_18124.t1 17.4
R13684 a_20907_18827.n1 a_20907_18827.t5 318.922
R13685 a_20907_18827.n0 a_20907_18827.t7 273.935
R13686 a_20907_18827.n0 a_20907_18827.t6 273.935
R13687 a_20907_18827.n1 a_20907_18827.t4 269.116
R13688 a_20907_18827.n4 a_20907_18827.n3 193.227
R13689 a_20907_18827.t5 a_20907_18827.n0 179.142
R13690 a_20907_18827.n2 a_20907_18827.n1 106.999
R13691 a_20907_18827.n3 a_20907_18827.t1 28.568
R13692 a_20907_18827.n4 a_20907_18827.t2 28.565
R13693 a_20907_18827.t3 a_20907_18827.n4 28.565
R13694 a_20907_18827.n2 a_20907_18827.t0 18.149
R13695 a_20907_18827.n3 a_20907_18827.n2 3.726
R13696 a_20613_18121.t0 a_20613_18121.t1 380.209
R13697 a_12598_9265.t0 a_12598_9265.t1 380.209
R13698 a_32011_8968.t0 a_32011_8968.t1 380.209
R13699 a_8190_1769.t0 a_8190_1769.t1 17.4
R13700 a_30077_6728.t0 a_30077_6728.t1 17.4
R13701 a_21194_24426.n1 a_21194_24426.t6 318.922
R13702 a_21194_24426.n0 a_21194_24426.t5 274.739
R13703 a_21194_24426.n0 a_21194_24426.t7 274.739
R13704 a_21194_24426.n1 a_21194_24426.t4 269.116
R13705 a_21194_24426.t6 a_21194_24426.n0 179.946
R13706 a_21194_24426.n2 a_21194_24426.n1 107.263
R13707 a_21194_24426.n3 a_21194_24426.t1 29.444
R13708 a_21194_24426.n4 a_21194_24426.t2 28.565
R13709 a_21194_24426.t3 a_21194_24426.n4 28.565
R13710 a_21194_24426.n2 a_21194_24426.t0 18.145
R13711 a_21194_24426.n3 a_21194_24426.n2 2.878
R13712 a_21194_24426.n4 a_21194_24426.n3 0.764
R13713 a_9661_21175.t0 a_9661_21175.t1 17.4
R13714 a_12712_25130.t0 a_12712_25130.t1 17.4
R13715 a_1483_9914.t0 a_1483_9914.t1 17.4
R13716 a_n2381_13124.t0 a_n2381_13124.t1 379.845
R13717 a_8155_14399.t0 a_8155_14399.t1 17.4
R13718 a_4373_6452.t0 a_4373_6452.t1 17.4
R13719 a_38084_1680.t0 a_38084_1680.t1 17.4
R13720 a_30006_11681.t0 a_30006_11681.t1 17.4
R13721 a_17951_10802.t4 a_17951_10802.t7 574.43
R13722 a_17951_10802.n0 a_17951_10802.t6 285.109
R13723 a_17951_10802.n2 a_17951_10802.n1 211.136
R13724 a_17951_10802.n4 a_17951_10802.n3 192.754
R13725 a_17951_10802.n0 a_17951_10802.t5 160.666
R13726 a_17951_10802.n1 a_17951_10802.t4 160.666
R13727 a_17951_10802.n1 a_17951_10802.n0 114.829
R13728 a_17951_10802.n3 a_17951_10802.t1 28.568
R13729 a_17951_10802.n4 a_17951_10802.t2 28.565
R13730 a_17951_10802.t3 a_17951_10802.n4 28.565
R13731 a_17951_10802.n2 a_17951_10802.t0 19.084
R13732 a_17951_10802.n3 a_17951_10802.n2 1.051
R13733 a_25804_25129.t0 a_25804_25129.t1 17.4
R13734 a_9751_23728.t0 a_9751_23728.t1 380.209
R13735 a_n2381_9223.t0 a_n2381_9223.t1 17.4
R13736 a_24215_4802.t0 a_24215_4802.t1 17.4
R13737 a_21150_9197.t0 a_21150_9197.t1 380.209
R13738 a_38088_7956.t0 a_38088_7956.t1 17.4
R13739 a_25790_26779.t0 a_25790_26779.t1 17.4
R13740 a_9987_23728.t0 a_9987_23728.t1 17.4
R13741 a_38088_23958.t0 a_38088_23958.t1 17.4
R13742 a_26297_12829.n1 a_26297_12829.t0 14.282
R13743 a_26297_12829.n1 a_26297_12829.t3 14.282
R13744 a_26297_12829.n0 a_26297_12829.t4 14.282
R13745 a_26297_12829.n0 a_26297_12829.t5 14.282
R13746 a_26297_12829.n3 a_26297_12829.t1 14.282
R13747 a_26297_12829.t2 a_26297_12829.n3 14.282
R13748 a_26297_12829.n2 a_26297_12829.n0 2.546
R13749 a_26297_12829.n3 a_26297_12829.n2 2.367
R13750 a_26297_12829.n2 a_26297_12829.n1 0.001
R13751 a_4387_4802.t0 a_4387_4802.t1 17.4
R13752 a_25858_21666.t4 a_25858_21666.t5 574.43
R13753 a_25858_21666.n1 a_25858_21666.t6 285.109
R13754 a_25858_21666.n3 a_25858_21666.n2 211.134
R13755 a_25858_21666.n4 a_25858_21666.n0 192.754
R13756 a_25858_21666.n1 a_25858_21666.t7 160.666
R13757 a_25858_21666.n2 a_25858_21666.t4 160.666
R13758 a_25858_21666.n2 a_25858_21666.n1 114.829
R13759 a_25858_21666.t3 a_25858_21666.n4 28.568
R13760 a_25858_21666.n0 a_25858_21666.t1 28.565
R13761 a_25858_21666.n0 a_25858_21666.t2 28.565
R13762 a_25858_21666.n3 a_25858_21666.t0 19.087
R13763 a_25858_21666.n4 a_25858_21666.n3 1.051
R13764 a_25564_21692.n1 a_25564_21692.t4 14.282
R13765 a_25564_21692.n1 a_25564_21692.t0 14.282
R13766 a_25564_21692.n0 a_25564_21692.t5 14.282
R13767 a_25564_21692.n0 a_25564_21692.t3 14.282
R13768 a_25564_21692.n3 a_25564_21692.t1 14.282
R13769 a_25564_21692.t2 a_25564_21692.n3 14.282
R13770 a_25564_21692.n2 a_25564_21692.n0 2.546
R13771 a_25564_21692.n3 a_25564_21692.n2 2.367
R13772 a_25564_21692.n2 a_25564_21692.n1 0.001
R13773 a_17588_3197.t0 a_17588_3197.t1 17.4
R13774 a_7939_3397.t0 a_7939_3397.t1 380.209
R13775 a_24218_9066.t0 a_24218_9066.t1 17.4
R13776 a_n2381_2781.t0 a_n2381_2781.t1 379.845
R13777 a_6615_12158.t7 a_6615_12158.t4 800.071
R13778 a_6615_12158.n3 a_6615_12158.n2 672.951
R13779 a_6615_12158.n1 a_6615_12158.t6 285.109
R13780 a_6615_12158.n2 a_6615_12158.t7 193.602
R13781 a_6615_12158.n1 a_6615_12158.t5 160.666
R13782 a_6615_12158.n2 a_6615_12158.n1 91.507
R13783 a_6615_12158.t1 a_6615_12158.n4 28.57
R13784 a_6615_12158.n0 a_6615_12158.t3 28.565
R13785 a_6615_12158.n0 a_6615_12158.t2 28.565
R13786 a_6615_12158.n4 a_6615_12158.t0 17.638
R13787 a_6615_12158.n3 a_6615_12158.n0 0.69
R13788 a_6615_12158.n4 a_6615_12158.n3 0.6
R13789 a_6351_12741.t5 a_6351_12741.n3 404.877
R13790 a_6351_12741.n2 a_6351_12741.t6 210.902
R13791 a_6351_12741.n4 a_6351_12741.t5 136.943
R13792 a_6351_12741.n3 a_6351_12741.n2 107.801
R13793 a_6351_12741.n2 a_6351_12741.t8 80.333
R13794 a_6351_12741.n3 a_6351_12741.t7 80.333
R13795 a_6351_12741.n1 a_6351_12741.t4 17.4
R13796 a_6351_12741.n1 a_6351_12741.t1 17.4
R13797 a_6351_12741.t0 a_6351_12741.n5 15.032
R13798 a_6351_12741.n0 a_6351_12741.t2 14.282
R13799 a_6351_12741.n0 a_6351_12741.t3 14.282
R13800 a_6351_12741.n5 a_6351_12741.n0 1.65
R13801 a_6351_12741.n4 a_6351_12741.n1 0.672
R13802 a_6351_12741.n5 a_6351_12741.n4 0.665
R13803 a_12181_18116.t0 a_12181_18116.t1 380.209
R13804 a_38084_17446.t0 a_38084_17446.t1 17.4
R13805 a_16264_23725.t0 a_16264_23725.t1 380.209
R13806 a_12417_18116.t0 a_12417_18116.t1 17.4
R13807 a_22744_17922.t0 a_22744_17922.t1 17.4
R13808 a_14726_3395.t0 a_14726_3395.t1 17.4
R13809 a_6469_12741.n0 a_6469_12741.t5 14.282
R13810 a_6469_12741.n0 a_6469_12741.t0 14.282
R13811 a_6469_12741.n1 a_6469_12741.t3 14.282
R13812 a_6469_12741.n1 a_6469_12741.t4 14.282
R13813 a_6469_12741.n3 a_6469_12741.t1 14.282
R13814 a_6469_12741.t2 a_6469_12741.n3 14.282
R13815 a_6469_12741.n3 a_6469_12741.n2 2.546
R13816 a_6469_12741.n2 a_6469_12741.n1 2.367
R13817 a_6469_12741.n2 a_6469_12741.n0 0.001
R13818 a_7853_23728.t0 a_7853_23728.t1 380.209
R13819 a_16500_23725.t0 a_16500_23725.t1 17.4
R13820 a_7947_9177.t0 a_7947_9177.t1 380.209
R13821 a_n2379_11291.t0 a_n2379_11291.t1 17.4
R13822 a_6285_9177.t0 a_6285_9177.t1 17.4
R13823 a_30006_8648.t0 a_30006_8648.t1 17.4
R13824 a_1491_12499.t0 a_1491_12499.t1 17.4
R13825 a_16210_17917.t0 a_16210_17917.t1 17.4
R13826 a_38088_11100.t0 a_38088_11100.t1 17.4
R13827 a_33612_13844.t0 a_33612_13844.t1 17.4
R13828 a_12698_26780.t0 a_12698_26780.t1 17.4
R13829 a_25799_23525.t0 a_25799_23525.t1 17.4
R13830 a_23034_23720.t0 a_23034_23720.t1 17.4
R13831 a_24223_10670.t0 a_24223_10670.t1 17.4
R13832 a_25464_18124.t0 a_25464_18124.t1 17.4
R13833 a_14668_27289.t5 a_14668_27289.n3 404.877
R13834 a_14668_27289.n2 a_14668_27289.t8 210.902
R13835 a_14668_27289.n4 a_14668_27289.t5 136.943
R13836 a_14668_27289.n3 a_14668_27289.n2 107.801
R13837 a_14668_27289.n2 a_14668_27289.t7 80.333
R13838 a_14668_27289.n3 a_14668_27289.t6 80.333
R13839 a_14668_27289.n1 a_14668_27289.t0 17.4
R13840 a_14668_27289.n1 a_14668_27289.t4 17.4
R13841 a_14668_27289.t3 a_14668_27289.n5 15.032
R13842 a_14668_27289.n0 a_14668_27289.t1 14.282
R13843 a_14668_27289.n0 a_14668_27289.t2 14.282
R13844 a_14668_27289.n5 a_14668_27289.n0 1.65
R13845 a_14668_27289.n4 a_14668_27289.n1 0.672
R13846 a_14668_27289.n5 a_14668_27289.n4 0.665
R13847 a_8089_23728.t0 a_8089_23728.t1 17.4
R13848 a_12592_3395.t0 a_12592_3395.t1 380.209
R13849 a_38084_5060.t0 a_38084_5060.t1 17.4
R13850 a_27775_9265.t0 a_27775_9265.t1 380.209
R13851 a_24209_12320.t0 a_24209_12320.t1 17.4
R13852 a_19232_26775.t0 a_19232_26775.t1 17.4
R13853 a_29266_21179.t0 a_29266_21179.t1 17.4
R13854 a_n2381_6918.t0 a_n2381_6918.t1 379.845
R13855 a_22739_19526.t0 a_22739_19526.t1 17.4
R13856 a_6194_23529.t0 a_6194_23529.t1 17.4
R13857 a_28003_3397.t0 a_28003_3397.t1 17.4
R13858 a_29592_23724.t0 a_29592_23724.t1 17.4
R13859 a_14602_23725.t0 a_14602_23725.t1 17.4
C0 w_4929_19483# Cout 0.03fF
C1 w_12316_24101# opcode[0] 0.00fF
C2 w_6872_21039# A[1] 0.01fF
C3 w_5803_24104# VDD 0.34fF
C4 w_9261_27234# A[1] 0.00fF
C5 w_28523_21754# VDD 0.38fF
C6 w_14632_27227# w_15774_27231# 0.03fF
C7 A[2] opcode[0] 0.10fF
C8 VDD A[7] 1.94fF
C9 w_7271_25091# A[1] 0.07fF
C10 w_28866_27230# VDD 0.66fF
C11 VDD B[3] 3.54fF
C12 opcode[1] Y[1] 0.06fF
C13 A[7] A[5] 0.12fF
C14 A[6] B[1] 0.04fF
C15 A[5] B[3] 5.39fF
C16 A[4] B[6] 1.27fF
C17 opcode[1] Y[5] 0.06fF
C18 A[3] B[7] 0.01fF
C19 B[0] B[7] 0.00fF
C20 B[3] B[2] 5.48fF
C21 w_18850_24096# VDD 0.34fF
C22 w_12288_21039# A[7] 0.00fF
C23 w_18855_25700# w_18850_24096# 0.02fF
C24 w_25413_25704# w_25408_24100# 0.02fF
C25 w_14632_27227# A[1] 0.01fF
C26 w_6872_21039# A[2] 0.01fF
C27 w_5803_24104# A[0] 0.19fF
C28 w_21996_20101# VDD 0.37fF
C29 w_21996_20101# A[5] 0.08fF
C30 w_5730_21043# Cout 0.19fF
C31 w_19964_21040# A[3] 0.10fF
C32 w_22308_27226# VDD 0.66fF
C33 w_28523_21754# A[4] 0.07fF
C34 w_18822_21044# A[6] 0.00fF
C35 A[3] opcode[0] 0.21fF
C36 VDD Cout 2.57fF
C37 w_7271_25091# A[2] 0.00fF
C38 w_5730_21043# w_4929_19483# 0.01fF
C39 w_25335_21047# w_24534_19487# 0.01fF
C40 A[7] A[4] 0.14fF
C41 opcode[0] B[0] 0.32fF
C42 A[3] B[4] 1.84fF
C43 opcode[1] Y[2] 0.06fF
C44 VDD B[1] 1.16fF
C45 w_25335_21047# VDD 0.66fF
C46 B[0] B[4] 0.00fF
C47 opcode[0] B[7] 13.09fF
C48 A[5] B[1] 0.00fF
C49 A[4] B[3] 1.41fF
C50 opcode[1] Y[6] 0.06fF
C51 w_25335_21047# A[5] 0.00fF
C52 B[1] B[2] 2.00fF
C53 B[4] B[7] 0.09fF
C54 w_11487_19479# A[6] 0.59fF
C55 w_8918_21750# A[7] 0.07fF
C56 w_25413_25704# A[3] 0.08fF
C57 w_12307_27355# A[1] 0.06fF
C58 w_13430_21035# A[2] 0.00fF
C59 w_8904_20100# w_8909_18496# 0.02fF
C60 w_4929_19483# VDD 1.02fF
C61 w_5808_25708# opcode[0] 0.07fF
C62 w_6872_21039# A[3] 0.11fF
C63 w_5803_24104# A[1] 0.03fF
C64 w_25399_27354# VDD 0.39fF
C65 w_5794_27358# Cout 0.00fF
C66 w_28866_27230# w_26876_25087# 0.02fF
C67 w_20318_25083# A[2] 0.60fF
C68 w_18822_21044# VDD 0.63fF
C69 VDD A[6] 5.47fF
C70 A[0] Cout 0.22fF
C71 A[1] A[7] 0.00fF
C72 A[3] opcode[1] 0.11fF
C73 w_15476_21746# A[2] 0.00fF
C74 opcode[0] B[4] 1.24fF
C75 VDD Y[3] 0.73fF
C76 A[3] B[5] 53.99fF
C77 A[6] A[5] 43.72fF
C78 B[0] B[5] 0.00fF
C79 A[4] B[1] 0.00fF
C80 opcode[1] B[7] 0.00fF
C81 A[6] B[2] 0.07fF
C82 w_11487_19479# VDD 1.02fF
C83 w_27724_27226# w_28866_27230# 0.03fF
C84 B[5] B[7] 0.14fF
C85 w_13430_21035# A[3] 0.10fF
C86 w_12321_25705# VDD 0.37fF
C87 w_6872_21039# opcode[0] 0.01fF
C88 w_5803_24104# A[2] 0.01fF
C89 w_28523_21754# w_28509_20104# 0.01fF
C90 w_22010_21751# w_21996_20101# 0.01fF
C91 w_12288_21039# w_11487_19479# 0.01fF
C92 w_5730_21043# VDD 0.68fF
C93 w_9261_27234# opcode[0] 0.00fF
C94 w_15467_18492# A[6] 0.14fF
C95 w_20318_25083# A[3] 0.05fF
C96 w_8119_27230# VDD 0.53fF
C97 w_11487_19479# w_15467_18492# 0.00fF
C98 w_24534_19487# VDD 1.02fF
C99 w_24534_19487# A[5] 0.06fF
C100 A[2] A[7] 0.00fF
C101 A[1] Cout 0.08fF
C102 opcode[0] opcode[1] 4.50fF
C103 VDD A[5] 5.37fF
C104 w_7271_25091# opcode[0] 0.39fF
C105 opcode[1] B[4] 0.01fF
C106 A[6] A[4] 4.13fF
C107 VDD B[2] 0.96fF
C108 A[3] B[6] 25.77fF
C109 opcode[0] B[5] 0.74fF
C110 w_15476_21746# A[3] 0.08fF
C111 w_18855_25700# VDD 0.37fF
C112 B[4] B[5] 8.13fF
C113 opcode[1] Y[7] 0.02fF
C114 A[5] B[2] 0.01fF
C115 B[0] B[6] 0.00fF
C116 B[6] B[7] 6.39fF
C117 w_18850_24096# A[2] 0.20fF
C118 w_15476_21746# w_15462_20096# 0.01fF
C119 w_12288_21039# VDD 0.64fF
C120 w_8904_20100# A[7] 0.08fF
C121 w_5803_24104# A[3] 0.00fF
C122 w_5794_27358# VDD 0.39fF
C123 w_5730_21043# A[0] 0.03fF
C124 w_18021_19484# w_22001_18497# 0.00fF
C125 w_15467_18492# VDD 0.33fF
C126 w_9261_27234# w_7271_25091# 0.01fF
C127 w_21166_27222# w_22308_27226# 0.03fF
C128 w_8119_27230# A[0] 0.01fF
C129 w_13784_25088# VDD 0.92fF
C130 VDD A[0] 2.40fF
C131 w_24534_19487# A[4] 0.59fF
C132 A[3] A[7] 0.11fF
C133 VDD A[4] 6.19fF
C134 A[2] Cout 0.10fF
C135 A[1] A[6] 0.00fF
C136 w_5808_25708# w_5803_24104# 0.02fF
C137 opcode[1] B[5] 0.01fF
C138 opcode[0] B[6] 0.71fF
C139 A[3] B[3] 58.44fF
C140 VDD Y[4] 0.74fF
C141 A[5] A[4] 55.20fF
C142 A[4] B[2] 0.00fF
C143 B[0] B[3] 0.00fF
C144 B[4] B[6] 27.70fF
C145 w_8918_21750# VDD 0.36fF
C146 B[3] B[7] 0.16fF
C147 w_18850_24096# A[3] 0.00fF
C148 w_25408_24100# w_25335_21047# 0.00fF
C149 w_12321_25705# A[1] 0.08fF
C150 w_15774_27231# VDD 0.66fF
C151 w_24534_19487# w_28514_18500# 0.00fF
C152 w_28514_18500# VDD 0.33fF
C153 w_5803_24104# opcode[0] 0.20fF
C154 w_5794_27358# A[0] 0.06fF
C155 w_5730_21043# A[1] 0.01fF
C156 w_26876_25087# VDD 0.94fF
C157 w_12321_25705# w_12316_24101# 0.02fF
C158 w_22308_27226# A[3] 0.00fF
C159 w_18822_21044# A[2] 0.02fF
C160 w_22010_21751# VDD 0.36fF
C161 VDD A[1] 2.10fF
C162 w_22010_21751# A[5] 0.07fF
C163 A[1] A[5] 0.00fF
C164 A[2] A[6] 0.01fF
C165 A[0] A[4] 0.00fF
C166 opcode[1] Y[0] 0.06fF
C167 VDD Y[1] 0.73fF
C168 A[3] Cout 0.13fF
C169 opcode[0] A[7] 0.08fF
C170 A[7] B[4] 0.00fF
C171 opcode[1] B[6] 0.01fF
C172 VDD Y[5] 0.73fF
C173 opcode[0] B[3] 1.48fF
C174 w_25335_21047# w_26477_21043# 0.03fF
C175 w_25335_21047# A[3] 0.02fF
C176 w_5803_24104# w_6872_21039# 0.00fF
C177 w_27724_27226# VDD 0.53fF
C178 B[0] B[1] 0.28fF
C179 B[5] B[6] 8.44fF
C180 B[4] B[3] 8.68fF
C181 B[1] B[7] 0.00fF
C182 w_15774_27231# w_13784_25088# 0.01fF
C183 w_12288_21039# A[1] 0.02fF
C184 w_12316_24101# VDD 0.34fF
C185 w_5808_25708# Cout 0.00fF
C186 w_28514_18500# A[4] 0.14fF
C187 w_6872_21039# A[7] 0.01fF
C188 w_7271_25091# w_5803_24104# 0.00fF
C189 w_25399_27354# A[3] 0.06fF
C190 w_5730_21043# A[2] 0.01fF
C191 w_28509_20104# VDD 0.37fF
C192 w_8909_18496# A[7] 0.14fF
C193 w_12316_24101# w_12288_21039# 0.00fF
C194 w_18822_21044# A[3] 0.12fF
C195 w_13784_25088# A[1] 0.60fF
C196 w_21166_27222# VDD 0.53fF
C197 VDD A[2] 2.25fF
C198 A[0] A[1] 0.88fF
C199 opcode[1] A[7] 11.88fF
C200 A[3] A[6] 1.22fF
C201 opcode[0] Cout 0.25fF
C202 A[1] A[4] 0.01fF
C203 VDD Y[2] 0.74fF
C204 A[2] A[5] 0.01fF
C205 opcode[1] B[3] 0.01fF
C206 VDD Y[6] 0.73fF
C207 A[6] B[0] 0.00fF
C208 opcode[0] B[1] 0.48fF
C209 w_18855_25700# A[2] 0.08fF
C210 B[4] B[1] 0.00fF
C211 A[6] B[7] 0.28fF
C212 B[5] B[3] 0.30fF
C213 w_8918_21750# A[1] 0.01fF
C214 w_25408_24100# VDD 0.34fF
C215 w_15462_20096# A[6] 0.08fF
C216 w_13784_25088# w_12316_24101# 0.00fF
C217 w_12288_21039# A[2] 0.01fF
C218 w_8904_20100# VDD 0.37fF
C219 w_6872_21039# Cout 0.01fF
C220 w_5730_21043# A[3] 0.12fF
C221 w_18822_21044# w_19964_21040# 0.03fF
C222 w_18841_27350# VDD 0.40fF
C223 w_28509_20104# A[4] 0.08fF
C224 w_25399_27354# w_25413_25704# 0.01fF
C225 w_18841_27350# w_18855_25700# 0.01fF
C226 w_13784_25088# A[2] 0.06fF
C227 w_18822_21044# w_18021_19484# 0.01fF
C228 w_26477_21043# VDD 0.52fF
C229 A[0] A[2] 0.01fF
C230 VDD A[3] 11.72fF
C231 A[2] A[4] 0.01fF
C232 opcode[0] A[6] 0.95fF
C233 VDD B[0] 1.38fF
C234 A[3] A[5] 0.33fF
C235 w_18021_19484# A[6] 0.06fF
C236 A[3] B[2] 0.00fF
C237 A[6] B[4] 3.34fF
C238 VDD B[7] 0.93fF
C239 w_20318_25083# w_18850_24096# 0.00fF
C240 B[0] B[2] 0.00fF
C241 B[6] B[3] 0.22fF
C242 A[5] B[7] 0.08fF
C243 B[5] B[1] 0.00fF
C244 w_8918_21750# A[2] 0.01fF
C245 w_21996_20101# w_22001_18497# 0.02fF
C246 w_4929_19483# w_8909_18496# 0.00fF
C247 B[2] B[7] 0.00fF
C248 w_28509_20104# w_28514_18500# 0.02fF
C249 w_15462_20096# VDD 0.37fF
C250 w_15774_27231# A[2] 0.00fF
C251 w_12288_21039# A[3] 0.12fF
C252 w_12316_24101# A[1] 0.20fF
C253 w_5808_25708# VDD 0.37fF
C254 w_22308_27226# w_20318_25083# 0.01fF
C255 w_5730_21043# opcode[0] 0.02fF
C256 w_8918_21750# w_8904_20100# 0.01fF
C257 w_19964_21040# VDD 0.50fF
C258 w_19964_21040# A[5] 0.01fF
C259 w_26876_25087# w_25408_24100# 0.00fF
C260 A[0] A[3] 0.01fF
C261 VDD opcode[0] 7.03fF
C262 A[1] A[2] 18.01fF
C263 w_15462_20096# w_15467_18492# 0.02fF
C264 w_18021_19484# VDD 1.02fF
C265 w_26477_21043# A[4] 0.01fF
C266 A[3] A[4] 9.91fF
C267 VDD B[4] 6.06fF
C268 opcode[1] A[6] 1.37fF
C269 opcode[0] A[5] 0.45fF
C270 w_5794_27358# w_5808_25708# 0.01fF
C271 w_18021_19484# A[5] 0.59fF
C272 opcode[0] B[2] 0.50fF
C273 VDD Y[7] 0.67fF
C274 A[6] B[5] 18.85fF
C275 opcode[1] Y[3] 0.06fF
C276 A[5] B[4] 2.49fF
C277 A[4] B[7] 0.03fF
C278 B[4] B[2] 0.00fF
C279 B[6] B[1] 0.00fF
C280 w_5730_21043# w_6872_21039# 0.03fF
C281 w_8918_21750# A[3] 0.09fF
C282 w_25413_25704# VDD 0.37fF
C283 w_13430_21035# A[6] 0.01fF
C284 w_12316_24101# A[2] 0.01fF
C285 w_5808_25708# A[0] 0.07fF
C286 w_6872_21039# VDD 0.54fF
C287 w_8119_27230# w_9261_27234# 0.03fF
C288 w_5803_24104# Cout 0.00fF
C289 w_5794_27358# opcode[0] 0.00fF
C290 w_26876_25087# A[3] 0.60fF
C291 w_9261_27234# VDD 0.66fF
C292 w_8909_18496# VDD 0.33fF
C293 w_21166_27222# A[2] 0.01fF
C294 w_22010_21751# A[3] 0.08fF
C295 VDD opcode[1] 16.29fF
C296 A[0] opcode[0] 0.85fF
C297 A[1] A[3] 0.08fF
C298 w_7271_25091# VDD 0.93fF
C299 opcode[0] A[4] 0.30fF
C300 opcode[1] A[5] 0.77fF
C301 VDD B[5] 9.32fF
C302 A[6] B[6] 12.43fF
C303 A[4] B[4] 25.38fF
C304 A[5] B[5] 27.51fF
C305 w_15476_21746# A[6] 0.07fF
C306 w_27724_27226# A[3] 0.01fF
C307 B[5] B[2] 0.00fF
C308 B[3] B[1] 0.00fF
C309 w_8918_21750# opcode[0] 0.00fF
C310 w_13430_21035# VDD 0.50fF
C311 w_4929_19483# A[7] 0.59fF
C312 w_12316_24101# A[3] 0.00fF
C313 w_14632_27227# VDD 0.53fF
C314 w_22001_18497# VDD 0.33fF
C315 w_12307_27355# w_12321_25705# 0.01fF
C316 w_22001_18497# A[5] 0.14fF
C317 w_18841_27350# A[2] 0.06fF
C318 w_12288_21039# w_13430_21035# 0.03fF
C319 w_20318_25083# VDD 0.92fF
C320 A[2] A[3] 23.65fF
C321 w_7271_25091# A[0] 0.60fF
C322 A[1] opcode[0] 5.93fF
C323 VDD Y[0] 0.73fF
C324 A[7] A[6] 16.20fF
C325 VDD B[6] 7.09fF
C326 w_15476_21746# VDD 0.36fF
C327 opcode[1] A[4] 0.57fF
C328 A[6] B[3] 4.20fF
C329 A[4] B[5] 1.71fF
C330 A[5] B[6] 1.32fF
C331 opcode[1] Y[4] 0.06fF
C332 B[6] B[2] 0.00fF
C333 w_11487_19479# A[7] 0.05fF
C334 w_25408_24100# w_26477_21043# 0.00fF
C335 w_25408_24100# A[3] 0.20fF
C336 w_5803_24104# w_5730_21043# 0.00fF
C337 w_18850_24096# w_18822_21044# 0.00fF
C338 w_12307_27355# VDD 0.39fF
.ends

