magic
tech sky130B
timestamp 1735993133
<< nwell >>
rect 0 0 242 274
<< nmos >>
rect 106 -162 136 -62
<< pmos >>
rect 47 31 77 131
rect 106 31 136 131
rect 165 31 195 131
<< ndiff >>
rect 77 -68 106 -62
rect 77 -156 83 -68
rect 100 -156 106 -68
rect 77 -162 106 -156
rect 136 -68 165 -62
rect 136 -156 142 -68
rect 159 -156 165 -68
rect 136 -162 165 -156
<< pdiff >>
rect 18 125 47 131
rect 18 37 24 125
rect 41 37 47 125
rect 18 31 47 37
rect 77 125 106 131
rect 77 37 83 125
rect 100 37 106 125
rect 77 31 106 37
rect 136 125 165 131
rect 136 37 142 125
rect 159 37 165 125
rect 136 31 165 37
rect 195 125 224 131
rect 195 37 201 125
rect 218 37 224 125
rect 195 31 224 37
<< ndiffc >>
rect 83 -156 100 -68
rect 142 -156 159 -68
<< pdiffc >>
rect 24 37 41 125
rect 83 37 100 125
rect 142 37 159 125
rect 201 37 218 125
<< psubdiff >>
rect 22 -214 152 -191
rect 22 -249 53 -214
rect 125 -249 152 -214
rect 22 -266 152 -249
<< nsubdiff >>
rect 47 226 195 233
rect 47 195 86 226
rect 156 195 195 226
rect 47 167 195 195
<< psubdiffcont >>
rect 53 -249 125 -214
<< nsubdiffcont >>
rect 86 195 156 226
<< poly >>
rect 47 131 77 144
rect 106 131 136 144
rect 165 131 195 144
rect 47 21 77 31
rect 106 21 136 31
rect 165 21 195 31
rect 47 3 195 21
rect 106 -18 136 3
rect 106 -35 112 -18
rect 129 -35 136 -18
rect 106 -62 136 -35
rect 106 -175 136 -162
<< polycont >>
rect 112 -35 129 -18
<< locali >>
rect 69 226 176 228
rect 69 195 86 226
rect 156 195 176 226
rect 69 186 176 195
rect 83 151 218 168
rect 24 125 41 133
rect 24 29 41 37
rect 83 125 100 151
rect 83 29 100 37
rect 142 125 159 133
rect 142 29 159 37
rect 201 125 218 151
rect 201 29 218 37
rect 104 -35 112 -18
rect 129 -35 137 -18
rect 83 -68 100 -60
rect 83 -164 100 -156
rect 142 -68 159 -60
rect 142 -164 159 -156
rect 43 -214 135 -204
rect 43 -249 53 -214
rect 125 -249 135 -214
rect 43 -252 135 -249
<< viali >>
rect 96 198 144 216
rect 24 37 41 125
rect 83 37 100 125
rect 142 37 159 125
rect 201 37 218 125
rect 112 -35 129 -18
rect 83 -156 100 -68
rect 142 -156 159 -68
rect 71 -245 110 -218
<< metal1 >>
rect 98 219 103 226
rect 83 216 103 219
rect 141 219 146 226
rect 141 216 162 219
rect 83 198 96 216
rect 144 198 162 216
rect 83 189 103 198
rect 141 189 162 198
rect 83 169 162 189
rect 21 146 162 169
rect 21 125 44 146
rect 21 37 24 125
rect 41 37 44 125
rect 21 31 44 37
rect 80 125 103 131
rect 80 37 83 125
rect 100 37 103 125
rect 80 31 103 37
rect 139 125 162 146
rect 139 37 142 125
rect 159 37 162 125
rect 139 31 162 37
rect 198 125 221 131
rect 198 37 201 125
rect 218 37 221 125
rect 198 34 221 37
rect 20 -15 39 -12
rect 198 -13 222 34
rect 20 -18 135 -15
rect 20 -35 112 -18
rect 129 -35 135 -18
rect 196 -32 224 -13
rect 20 -38 135 -35
rect 20 -40 39 -38
rect 198 -62 222 -32
rect 80 -68 103 -62
rect 80 -156 83 -68
rect 100 -156 103 -68
rect 80 -215 103 -156
rect 139 -68 222 -62
rect 139 -156 142 -68
rect 159 -77 222 -68
rect 159 -156 162 -77
rect 139 -162 162 -156
rect 60 -248 65 -215
rect 116 -248 121 -215
<< via1 >>
rect 103 216 141 226
rect 103 198 141 216
rect 103 189 141 198
rect 65 -218 116 -215
rect 65 -245 71 -218
rect 71 -245 110 -218
rect 110 -245 116 -218
rect 65 -248 116 -245
<< metal2 >>
rect 99 231 146 236
rect 99 184 146 189
rect 65 -213 116 -210
rect 65 -215 117 -213
rect 116 -248 117 -215
rect 65 -252 117 -248
rect 65 -253 116 -252
<< via2 >>
rect 99 226 146 231
rect 99 189 103 226
rect 103 189 141 226
rect 141 189 146 226
rect 73 -247 106 -218
<< metal3 >>
rect 21 238 218 241
rect 21 184 95 238
rect 150 184 218 238
rect 21 166 218 184
rect 50 -208 130 -207
rect 50 -213 65 -208
rect 49 -254 65 -213
rect 50 -258 65 -254
rect 116 -258 130 -208
rect 50 -261 130 -258
<< via3 >>
rect 95 231 150 238
rect 95 189 99 231
rect 99 189 146 231
rect 146 189 150 231
rect 95 184 150 189
rect 65 -218 116 -208
rect 65 -247 73 -218
rect 73 -247 106 -218
rect 106 -247 116 -218
rect 65 -258 116 -247
<< metal4 >>
rect 2 238 225 257
rect 2 184 95 238
rect 150 184 225 238
rect 2 181 225 184
rect 12 -208 160 -187
rect 12 -258 65 -208
rect 116 -258 160 -208
rect 12 -269 160 -258
<< labels >>
flabel metal1 20 -40 39 -12 1 FreeSerif 160 0 0 0 IN
port 1 n
flabel metal1 196 -32 224 -13 1 FreeSerif 160 0 0 0 OUT
port 2 n
flabel metal4 66 184 183 238 1 FreeSerif 240 0 0 0 VDD
port 3 n
flabel metal4 45 -258 130 -203 1 FreeSerif 240 0 0 0 VSS
port 4 n
<< end >>
