magic
tech sky130B
magscale 1 2
timestamp 1736777825
<< nwell >>
rect -471 524 1306 814
rect 2673 524 4450 814
rect 5805 528 7582 818
rect 8949 528 10726 818
rect -471 324 1307 524
rect 2673 324 4451 524
rect 5805 328 7583 528
rect 8949 328 10727 528
rect 12151 524 13928 814
rect 15295 524 17072 814
rect 18427 528 20204 818
rect 21571 528 23348 818
rect -912 0 1780 324
rect 2232 0 4924 324
rect 5364 4 8056 328
rect 8508 4 11200 328
rect 12151 324 13929 524
rect 15295 324 17073 524
rect 18427 328 20205 528
rect 21571 328 23349 528
rect 11710 0 14402 324
rect 14854 0 17546 324
rect 17986 4 20678 328
rect 21130 4 23822 328
<< nmos >>
rect 16 -1071 76 -871
rect 208 -1271 268 -871
rect 326 -1271 386 -871
rect 444 -1271 504 -871
rect 562 -1271 622 -871
rect 758 -1071 818 -871
rect 3160 -1071 3220 -871
rect 3352 -1271 3412 -871
rect 3470 -1271 3530 -871
rect 3588 -1271 3648 -871
rect 3706 -1271 3766 -871
rect 3902 -1071 3962 -871
rect 6292 -1067 6352 -867
rect 6484 -1267 6544 -867
rect 6602 -1267 6662 -867
rect 6720 -1267 6780 -867
rect 6838 -1267 6898 -867
rect 7034 -1067 7094 -867
rect 9436 -1067 9496 -867
rect 9628 -1267 9688 -867
rect 9746 -1267 9806 -867
rect 9864 -1267 9924 -867
rect 9982 -1267 10042 -867
rect 10178 -1067 10238 -867
rect 12638 -1071 12698 -871
rect 12830 -1271 12890 -871
rect 12948 -1271 13008 -871
rect 13066 -1271 13126 -871
rect 13184 -1271 13244 -871
rect 13380 -1071 13440 -871
rect 15782 -1071 15842 -871
rect 15974 -1271 16034 -871
rect 16092 -1271 16152 -871
rect 16210 -1271 16270 -871
rect 16328 -1271 16388 -871
rect 16524 -1071 16584 -871
rect 18914 -1067 18974 -867
rect 19106 -1267 19166 -867
rect 19224 -1267 19284 -867
rect 19342 -1267 19402 -867
rect 19460 -1267 19520 -867
rect 19656 -1067 19716 -867
rect 22058 -1067 22118 -867
rect 22250 -1267 22310 -867
rect 22368 -1267 22428 -867
rect 22486 -1267 22546 -867
rect 22604 -1267 22664 -867
rect 22800 -1067 22860 -867
<< pmos >>
rect -818 62 -758 262
rect -700 62 -640 262
rect -582 62 -522 262
rect -377 62 -317 462
rect -259 62 -199 462
rect -141 62 -81 462
rect 90 62 150 462
rect 208 62 268 462
rect 326 62 386 462
rect 444 62 504 462
rect 562 62 622 462
rect 680 62 740 462
rect 917 62 977 462
rect 1035 62 1095 462
rect 1153 62 1213 462
rect 1390 62 1450 262
rect 1508 62 1568 262
rect 1626 62 1686 262
rect 2326 62 2386 262
rect 2444 62 2504 262
rect 2562 62 2622 262
rect 2767 62 2827 462
rect 2885 62 2945 462
rect 3003 62 3063 462
rect 3234 62 3294 462
rect 3352 62 3412 462
rect 3470 62 3530 462
rect 3588 62 3648 462
rect 3706 62 3766 462
rect 3824 62 3884 462
rect 4061 62 4121 462
rect 4179 62 4239 462
rect 4297 62 4357 462
rect 4534 62 4594 262
rect 4652 62 4712 262
rect 4770 62 4830 262
rect 5458 66 5518 266
rect 5576 66 5636 266
rect 5694 66 5754 266
rect 5899 66 5959 466
rect 6017 66 6077 466
rect 6135 66 6195 466
rect 6366 66 6426 466
rect 6484 66 6544 466
rect 6602 66 6662 466
rect 6720 66 6780 466
rect 6838 66 6898 466
rect 6956 66 7016 466
rect 7193 66 7253 466
rect 7311 66 7371 466
rect 7429 66 7489 466
rect 7666 66 7726 266
rect 7784 66 7844 266
rect 7902 66 7962 266
rect 8602 66 8662 266
rect 8720 66 8780 266
rect 8838 66 8898 266
rect 9043 66 9103 466
rect 9161 66 9221 466
rect 9279 66 9339 466
rect 9510 66 9570 466
rect 9628 66 9688 466
rect 9746 66 9806 466
rect 9864 66 9924 466
rect 9982 66 10042 466
rect 10100 66 10160 466
rect 10337 66 10397 466
rect 10455 66 10515 466
rect 10573 66 10633 466
rect 10810 66 10870 266
rect 10928 66 10988 266
rect 11046 66 11106 266
rect 11804 62 11864 262
rect 11922 62 11982 262
rect 12040 62 12100 262
rect 12245 62 12305 462
rect 12363 62 12423 462
rect 12481 62 12541 462
rect 12712 62 12772 462
rect 12830 62 12890 462
rect 12948 62 13008 462
rect 13066 62 13126 462
rect 13184 62 13244 462
rect 13302 62 13362 462
rect 13539 62 13599 462
rect 13657 62 13717 462
rect 13775 62 13835 462
rect 14012 62 14072 262
rect 14130 62 14190 262
rect 14248 62 14308 262
rect 14948 62 15008 262
rect 15066 62 15126 262
rect 15184 62 15244 262
rect 15389 62 15449 462
rect 15507 62 15567 462
rect 15625 62 15685 462
rect 15856 62 15916 462
rect 15974 62 16034 462
rect 16092 62 16152 462
rect 16210 62 16270 462
rect 16328 62 16388 462
rect 16446 62 16506 462
rect 16683 62 16743 462
rect 16801 62 16861 462
rect 16919 62 16979 462
rect 17156 62 17216 262
rect 17274 62 17334 262
rect 17392 62 17452 262
rect 18080 66 18140 266
rect 18198 66 18258 266
rect 18316 66 18376 266
rect 18521 66 18581 466
rect 18639 66 18699 466
rect 18757 66 18817 466
rect 18988 66 19048 466
rect 19106 66 19166 466
rect 19224 66 19284 466
rect 19342 66 19402 466
rect 19460 66 19520 466
rect 19578 66 19638 466
rect 19815 66 19875 466
rect 19933 66 19993 466
rect 20051 66 20111 466
rect 20288 66 20348 266
rect 20406 66 20466 266
rect 20524 66 20584 266
rect 21224 66 21284 266
rect 21342 66 21402 266
rect 21460 66 21520 266
rect 21665 66 21725 466
rect 21783 66 21843 466
rect 21901 66 21961 466
rect 22132 66 22192 466
rect 22250 66 22310 466
rect 22368 66 22428 466
rect 22486 66 22546 466
rect 22604 66 22664 466
rect 22722 66 22782 466
rect 22959 66 23019 466
rect 23077 66 23137 466
rect 23195 66 23255 466
rect 23432 66 23492 266
rect 23550 66 23610 266
rect 23668 66 23728 266
<< ndiff >>
rect -42 -883 16 -871
rect -42 -1059 -30 -883
rect 4 -1059 16 -883
rect -42 -1071 16 -1059
rect 76 -883 208 -871
rect 76 -1059 88 -883
rect 122 -1059 162 -883
rect 76 -1071 162 -1059
rect 150 -1259 162 -1071
rect 196 -1259 208 -883
rect 150 -1271 208 -1259
rect 268 -883 326 -871
rect 268 -1259 280 -883
rect 314 -1259 326 -883
rect 268 -1271 326 -1259
rect 386 -883 444 -871
rect 386 -1259 398 -883
rect 432 -1259 444 -883
rect 386 -1271 444 -1259
rect 504 -883 562 -871
rect 504 -1259 516 -883
rect 550 -1259 562 -883
rect 504 -1271 562 -1259
rect 622 -883 758 -871
rect 622 -1259 634 -883
rect 668 -1059 712 -883
rect 746 -1059 758 -883
rect 668 -1071 758 -1059
rect 818 -883 876 -871
rect 818 -1059 830 -883
rect 864 -1059 876 -883
rect 818 -1071 876 -1059
rect 3102 -883 3160 -871
rect 3102 -1059 3114 -883
rect 3148 -1059 3160 -883
rect 3102 -1071 3160 -1059
rect 3220 -883 3352 -871
rect 3220 -1059 3232 -883
rect 3266 -1059 3306 -883
rect 3220 -1071 3306 -1059
rect 668 -1259 680 -1071
rect 622 -1271 680 -1259
rect 3294 -1259 3306 -1071
rect 3340 -1259 3352 -883
rect 3294 -1271 3352 -1259
rect 3412 -883 3470 -871
rect 3412 -1259 3424 -883
rect 3458 -1259 3470 -883
rect 3412 -1271 3470 -1259
rect 3530 -883 3588 -871
rect 3530 -1259 3542 -883
rect 3576 -1259 3588 -883
rect 3530 -1271 3588 -1259
rect 3648 -883 3706 -871
rect 3648 -1259 3660 -883
rect 3694 -1259 3706 -883
rect 3648 -1271 3706 -1259
rect 3766 -883 3902 -871
rect 3766 -1259 3778 -883
rect 3812 -1059 3856 -883
rect 3890 -1059 3902 -883
rect 3812 -1071 3902 -1059
rect 3962 -883 4020 -871
rect 3962 -1059 3974 -883
rect 4008 -1059 4020 -883
rect 3962 -1071 4020 -1059
rect 6234 -879 6292 -867
rect 6234 -1055 6246 -879
rect 6280 -1055 6292 -879
rect 6234 -1067 6292 -1055
rect 6352 -879 6484 -867
rect 6352 -1055 6364 -879
rect 6398 -1055 6438 -879
rect 6352 -1067 6438 -1055
rect 3812 -1259 3824 -1071
rect 3766 -1271 3824 -1259
rect 6426 -1255 6438 -1067
rect 6472 -1255 6484 -879
rect 6426 -1267 6484 -1255
rect 6544 -879 6602 -867
rect 6544 -1255 6556 -879
rect 6590 -1255 6602 -879
rect 6544 -1267 6602 -1255
rect 6662 -879 6720 -867
rect 6662 -1255 6674 -879
rect 6708 -1255 6720 -879
rect 6662 -1267 6720 -1255
rect 6780 -879 6838 -867
rect 6780 -1255 6792 -879
rect 6826 -1255 6838 -879
rect 6780 -1267 6838 -1255
rect 6898 -879 7034 -867
rect 6898 -1255 6910 -879
rect 6944 -1055 6988 -879
rect 7022 -1055 7034 -879
rect 6944 -1067 7034 -1055
rect 7094 -879 7152 -867
rect 7094 -1055 7106 -879
rect 7140 -1055 7152 -879
rect 7094 -1067 7152 -1055
rect 9378 -879 9436 -867
rect 9378 -1055 9390 -879
rect 9424 -1055 9436 -879
rect 9378 -1067 9436 -1055
rect 9496 -879 9628 -867
rect 9496 -1055 9508 -879
rect 9542 -1055 9582 -879
rect 9496 -1067 9582 -1055
rect 6944 -1255 6956 -1067
rect 6898 -1267 6956 -1255
rect 9570 -1255 9582 -1067
rect 9616 -1255 9628 -879
rect 9570 -1267 9628 -1255
rect 9688 -879 9746 -867
rect 9688 -1255 9700 -879
rect 9734 -1255 9746 -879
rect 9688 -1267 9746 -1255
rect 9806 -879 9864 -867
rect 9806 -1255 9818 -879
rect 9852 -1255 9864 -879
rect 9806 -1267 9864 -1255
rect 9924 -879 9982 -867
rect 9924 -1255 9936 -879
rect 9970 -1255 9982 -879
rect 9924 -1267 9982 -1255
rect 10042 -879 10178 -867
rect 10042 -1255 10054 -879
rect 10088 -1055 10132 -879
rect 10166 -1055 10178 -879
rect 10088 -1067 10178 -1055
rect 10238 -879 10296 -867
rect 10238 -1055 10250 -879
rect 10284 -1055 10296 -879
rect 10238 -1067 10296 -1055
rect 12580 -883 12638 -871
rect 12580 -1059 12592 -883
rect 12626 -1059 12638 -883
rect 10088 -1255 10100 -1067
rect 10042 -1267 10100 -1255
rect 12580 -1071 12638 -1059
rect 12698 -883 12830 -871
rect 12698 -1059 12710 -883
rect 12744 -1059 12784 -883
rect 12698 -1071 12784 -1059
rect 12772 -1259 12784 -1071
rect 12818 -1259 12830 -883
rect 12772 -1271 12830 -1259
rect 12890 -883 12948 -871
rect 12890 -1259 12902 -883
rect 12936 -1259 12948 -883
rect 12890 -1271 12948 -1259
rect 13008 -883 13066 -871
rect 13008 -1259 13020 -883
rect 13054 -1259 13066 -883
rect 13008 -1271 13066 -1259
rect 13126 -883 13184 -871
rect 13126 -1259 13138 -883
rect 13172 -1259 13184 -883
rect 13126 -1271 13184 -1259
rect 13244 -883 13380 -871
rect 13244 -1259 13256 -883
rect 13290 -1059 13334 -883
rect 13368 -1059 13380 -883
rect 13290 -1071 13380 -1059
rect 13440 -883 13498 -871
rect 13440 -1059 13452 -883
rect 13486 -1059 13498 -883
rect 13440 -1071 13498 -1059
rect 15724 -883 15782 -871
rect 15724 -1059 15736 -883
rect 15770 -1059 15782 -883
rect 15724 -1071 15782 -1059
rect 15842 -883 15974 -871
rect 15842 -1059 15854 -883
rect 15888 -1059 15928 -883
rect 15842 -1071 15928 -1059
rect 13290 -1259 13302 -1071
rect 13244 -1271 13302 -1259
rect 15916 -1259 15928 -1071
rect 15962 -1259 15974 -883
rect 15916 -1271 15974 -1259
rect 16034 -883 16092 -871
rect 16034 -1259 16046 -883
rect 16080 -1259 16092 -883
rect 16034 -1271 16092 -1259
rect 16152 -883 16210 -871
rect 16152 -1259 16164 -883
rect 16198 -1259 16210 -883
rect 16152 -1271 16210 -1259
rect 16270 -883 16328 -871
rect 16270 -1259 16282 -883
rect 16316 -1259 16328 -883
rect 16270 -1271 16328 -1259
rect 16388 -883 16524 -871
rect 16388 -1259 16400 -883
rect 16434 -1059 16478 -883
rect 16512 -1059 16524 -883
rect 16434 -1071 16524 -1059
rect 16584 -883 16642 -871
rect 16584 -1059 16596 -883
rect 16630 -1059 16642 -883
rect 16584 -1071 16642 -1059
rect 18856 -879 18914 -867
rect 18856 -1055 18868 -879
rect 18902 -1055 18914 -879
rect 18856 -1067 18914 -1055
rect 18974 -879 19106 -867
rect 18974 -1055 18986 -879
rect 19020 -1055 19060 -879
rect 18974 -1067 19060 -1055
rect 16434 -1259 16446 -1071
rect 16388 -1271 16446 -1259
rect 19048 -1255 19060 -1067
rect 19094 -1255 19106 -879
rect 19048 -1267 19106 -1255
rect 19166 -879 19224 -867
rect 19166 -1255 19178 -879
rect 19212 -1255 19224 -879
rect 19166 -1267 19224 -1255
rect 19284 -879 19342 -867
rect 19284 -1255 19296 -879
rect 19330 -1255 19342 -879
rect 19284 -1267 19342 -1255
rect 19402 -879 19460 -867
rect 19402 -1255 19414 -879
rect 19448 -1255 19460 -879
rect 19402 -1267 19460 -1255
rect 19520 -879 19656 -867
rect 19520 -1255 19532 -879
rect 19566 -1055 19610 -879
rect 19644 -1055 19656 -879
rect 19566 -1067 19656 -1055
rect 19716 -879 19774 -867
rect 19716 -1055 19728 -879
rect 19762 -1055 19774 -879
rect 19716 -1067 19774 -1055
rect 22000 -879 22058 -867
rect 22000 -1055 22012 -879
rect 22046 -1055 22058 -879
rect 22000 -1067 22058 -1055
rect 22118 -879 22250 -867
rect 22118 -1055 22130 -879
rect 22164 -1055 22204 -879
rect 22118 -1067 22204 -1055
rect 19566 -1255 19578 -1067
rect 19520 -1267 19578 -1255
rect 22192 -1255 22204 -1067
rect 22238 -1255 22250 -879
rect 22192 -1267 22250 -1255
rect 22310 -879 22368 -867
rect 22310 -1255 22322 -879
rect 22356 -1255 22368 -879
rect 22310 -1267 22368 -1255
rect 22428 -879 22486 -867
rect 22428 -1255 22440 -879
rect 22474 -1255 22486 -879
rect 22428 -1267 22486 -1255
rect 22546 -879 22604 -867
rect 22546 -1255 22558 -879
rect 22592 -1255 22604 -879
rect 22546 -1267 22604 -1255
rect 22664 -879 22800 -867
rect 22664 -1255 22676 -879
rect 22710 -1055 22754 -879
rect 22788 -1055 22800 -879
rect 22710 -1067 22800 -1055
rect 22860 -879 22918 -867
rect 22860 -1055 22872 -879
rect 22906 -1055 22918 -879
rect 22860 -1067 22918 -1055
rect 22710 -1255 22722 -1067
rect 22664 -1267 22722 -1255
<< pdiff >>
rect -435 450 -377 462
rect -435 262 -423 450
rect -876 250 -818 262
rect -876 74 -864 250
rect -830 74 -818 250
rect -876 62 -818 74
rect -758 250 -700 262
rect -758 74 -746 250
rect -712 74 -700 250
rect -758 62 -700 74
rect -640 250 -582 262
rect -640 74 -628 250
rect -594 74 -582 250
rect -640 62 -582 74
rect -522 250 -423 262
rect -522 74 -510 250
rect -476 74 -423 250
rect -389 74 -377 450
rect -522 62 -377 74
rect -317 450 -259 462
rect -317 74 -305 450
rect -271 74 -259 450
rect -317 62 -259 74
rect -199 450 -141 462
rect -199 74 -187 450
rect -153 74 -141 450
rect -199 62 -141 74
rect -81 450 -23 462
rect -81 74 -69 450
rect -35 74 -23 450
rect -81 62 -23 74
rect 32 450 90 462
rect 32 74 44 450
rect 78 74 90 450
rect 32 62 90 74
rect 150 450 208 462
rect 150 74 162 450
rect 196 74 208 450
rect 150 62 208 74
rect 268 450 326 462
rect 268 74 280 450
rect 314 74 326 450
rect 268 62 326 74
rect 386 450 444 462
rect 386 74 398 450
rect 432 74 444 450
rect 386 62 444 74
rect 504 450 562 462
rect 504 74 516 450
rect 550 74 562 450
rect 504 62 562 74
rect 622 450 680 462
rect 622 74 634 450
rect 668 74 680 450
rect 622 62 680 74
rect 740 450 798 462
rect 740 74 752 450
rect 786 74 798 450
rect 740 62 798 74
rect 859 450 917 462
rect 859 74 871 450
rect 905 74 917 450
rect 859 62 917 74
rect 977 450 1035 462
rect 977 74 989 450
rect 1023 74 1035 450
rect 977 62 1035 74
rect 1095 450 1153 462
rect 1095 74 1107 450
rect 1141 74 1153 450
rect 1095 62 1153 74
rect 1213 450 1271 462
rect 1213 74 1225 450
rect 1259 74 1271 450
rect 2709 450 2767 462
rect 2709 262 2721 450
rect 1213 62 1271 74
rect 1332 250 1390 262
rect 1332 74 1344 250
rect 1378 74 1390 250
rect 1332 62 1390 74
rect 1450 250 1508 262
rect 1450 74 1462 250
rect 1496 74 1508 250
rect 1450 62 1508 74
rect 1568 250 1626 262
rect 1568 74 1580 250
rect 1614 74 1626 250
rect 1568 62 1626 74
rect 1686 250 1744 262
rect 1686 74 1698 250
rect 1732 74 1744 250
rect 1686 62 1744 74
rect 2268 250 2326 262
rect 2268 74 2280 250
rect 2314 74 2326 250
rect 2268 62 2326 74
rect 2386 250 2444 262
rect 2386 74 2398 250
rect 2432 74 2444 250
rect 2386 62 2444 74
rect 2504 250 2562 262
rect 2504 74 2516 250
rect 2550 74 2562 250
rect 2504 62 2562 74
rect 2622 250 2721 262
rect 2622 74 2634 250
rect 2668 74 2721 250
rect 2755 74 2767 450
rect 2622 62 2767 74
rect 2827 450 2885 462
rect 2827 74 2839 450
rect 2873 74 2885 450
rect 2827 62 2885 74
rect 2945 450 3003 462
rect 2945 74 2957 450
rect 2991 74 3003 450
rect 2945 62 3003 74
rect 3063 450 3121 462
rect 3063 74 3075 450
rect 3109 74 3121 450
rect 3063 62 3121 74
rect 3176 450 3234 462
rect 3176 74 3188 450
rect 3222 74 3234 450
rect 3176 62 3234 74
rect 3294 450 3352 462
rect 3294 74 3306 450
rect 3340 74 3352 450
rect 3294 62 3352 74
rect 3412 450 3470 462
rect 3412 74 3424 450
rect 3458 74 3470 450
rect 3412 62 3470 74
rect 3530 450 3588 462
rect 3530 74 3542 450
rect 3576 74 3588 450
rect 3530 62 3588 74
rect 3648 450 3706 462
rect 3648 74 3660 450
rect 3694 74 3706 450
rect 3648 62 3706 74
rect 3766 450 3824 462
rect 3766 74 3778 450
rect 3812 74 3824 450
rect 3766 62 3824 74
rect 3884 450 3942 462
rect 3884 74 3896 450
rect 3930 74 3942 450
rect 3884 62 3942 74
rect 4003 450 4061 462
rect 4003 74 4015 450
rect 4049 74 4061 450
rect 4003 62 4061 74
rect 4121 450 4179 462
rect 4121 74 4133 450
rect 4167 74 4179 450
rect 4121 62 4179 74
rect 4239 450 4297 462
rect 4239 74 4251 450
rect 4285 74 4297 450
rect 4239 62 4297 74
rect 4357 450 4415 462
rect 4357 74 4369 450
rect 4403 74 4415 450
rect 5841 454 5899 466
rect 5841 266 5853 454
rect 4357 62 4415 74
rect 4476 250 4534 262
rect 4476 74 4488 250
rect 4522 74 4534 250
rect 4476 62 4534 74
rect 4594 250 4652 262
rect 4594 74 4606 250
rect 4640 74 4652 250
rect 4594 62 4652 74
rect 4712 250 4770 262
rect 4712 74 4724 250
rect 4758 74 4770 250
rect 4712 62 4770 74
rect 4830 250 4888 262
rect 4830 74 4842 250
rect 4876 74 4888 250
rect 4830 62 4888 74
rect 5400 254 5458 266
rect 5400 78 5412 254
rect 5446 78 5458 254
rect 5400 66 5458 78
rect 5518 254 5576 266
rect 5518 78 5530 254
rect 5564 78 5576 254
rect 5518 66 5576 78
rect 5636 254 5694 266
rect 5636 78 5648 254
rect 5682 78 5694 254
rect 5636 66 5694 78
rect 5754 254 5853 266
rect 5754 78 5766 254
rect 5800 78 5853 254
rect 5887 78 5899 454
rect 5754 66 5899 78
rect 5959 454 6017 466
rect 5959 78 5971 454
rect 6005 78 6017 454
rect 5959 66 6017 78
rect 6077 454 6135 466
rect 6077 78 6089 454
rect 6123 78 6135 454
rect 6077 66 6135 78
rect 6195 454 6253 466
rect 6195 78 6207 454
rect 6241 78 6253 454
rect 6195 66 6253 78
rect 6308 454 6366 466
rect 6308 78 6320 454
rect 6354 78 6366 454
rect 6308 66 6366 78
rect 6426 454 6484 466
rect 6426 78 6438 454
rect 6472 78 6484 454
rect 6426 66 6484 78
rect 6544 454 6602 466
rect 6544 78 6556 454
rect 6590 78 6602 454
rect 6544 66 6602 78
rect 6662 454 6720 466
rect 6662 78 6674 454
rect 6708 78 6720 454
rect 6662 66 6720 78
rect 6780 454 6838 466
rect 6780 78 6792 454
rect 6826 78 6838 454
rect 6780 66 6838 78
rect 6898 454 6956 466
rect 6898 78 6910 454
rect 6944 78 6956 454
rect 6898 66 6956 78
rect 7016 454 7074 466
rect 7016 78 7028 454
rect 7062 78 7074 454
rect 7016 66 7074 78
rect 7135 454 7193 466
rect 7135 78 7147 454
rect 7181 78 7193 454
rect 7135 66 7193 78
rect 7253 454 7311 466
rect 7253 78 7265 454
rect 7299 78 7311 454
rect 7253 66 7311 78
rect 7371 454 7429 466
rect 7371 78 7383 454
rect 7417 78 7429 454
rect 7371 66 7429 78
rect 7489 454 7547 466
rect 7489 78 7501 454
rect 7535 78 7547 454
rect 8985 454 9043 466
rect 8985 266 8997 454
rect 7489 66 7547 78
rect 7608 254 7666 266
rect 7608 78 7620 254
rect 7654 78 7666 254
rect 7608 66 7666 78
rect 7726 254 7784 266
rect 7726 78 7738 254
rect 7772 78 7784 254
rect 7726 66 7784 78
rect 7844 254 7902 266
rect 7844 78 7856 254
rect 7890 78 7902 254
rect 7844 66 7902 78
rect 7962 254 8020 266
rect 7962 78 7974 254
rect 8008 78 8020 254
rect 7962 66 8020 78
rect 8544 254 8602 266
rect 8544 78 8556 254
rect 8590 78 8602 254
rect 8544 66 8602 78
rect 8662 254 8720 266
rect 8662 78 8674 254
rect 8708 78 8720 254
rect 8662 66 8720 78
rect 8780 254 8838 266
rect 8780 78 8792 254
rect 8826 78 8838 254
rect 8780 66 8838 78
rect 8898 254 8997 266
rect 8898 78 8910 254
rect 8944 78 8997 254
rect 9031 78 9043 454
rect 8898 66 9043 78
rect 9103 454 9161 466
rect 9103 78 9115 454
rect 9149 78 9161 454
rect 9103 66 9161 78
rect 9221 454 9279 466
rect 9221 78 9233 454
rect 9267 78 9279 454
rect 9221 66 9279 78
rect 9339 454 9397 466
rect 9339 78 9351 454
rect 9385 78 9397 454
rect 9339 66 9397 78
rect 9452 454 9510 466
rect 9452 78 9464 454
rect 9498 78 9510 454
rect 9452 66 9510 78
rect 9570 454 9628 466
rect 9570 78 9582 454
rect 9616 78 9628 454
rect 9570 66 9628 78
rect 9688 454 9746 466
rect 9688 78 9700 454
rect 9734 78 9746 454
rect 9688 66 9746 78
rect 9806 454 9864 466
rect 9806 78 9818 454
rect 9852 78 9864 454
rect 9806 66 9864 78
rect 9924 454 9982 466
rect 9924 78 9936 454
rect 9970 78 9982 454
rect 9924 66 9982 78
rect 10042 454 10100 466
rect 10042 78 10054 454
rect 10088 78 10100 454
rect 10042 66 10100 78
rect 10160 454 10218 466
rect 10160 78 10172 454
rect 10206 78 10218 454
rect 10160 66 10218 78
rect 10279 454 10337 466
rect 10279 78 10291 454
rect 10325 78 10337 454
rect 10279 66 10337 78
rect 10397 454 10455 466
rect 10397 78 10409 454
rect 10443 78 10455 454
rect 10397 66 10455 78
rect 10515 454 10573 466
rect 10515 78 10527 454
rect 10561 78 10573 454
rect 10515 66 10573 78
rect 10633 454 10691 466
rect 10633 78 10645 454
rect 10679 78 10691 454
rect 12187 450 12245 462
rect 10633 66 10691 78
rect 10752 254 10810 266
rect 10752 78 10764 254
rect 10798 78 10810 254
rect 10752 66 10810 78
rect 10870 254 10928 266
rect 10870 78 10882 254
rect 10916 78 10928 254
rect 10870 66 10928 78
rect 10988 254 11046 266
rect 10988 78 11000 254
rect 11034 78 11046 254
rect 10988 66 11046 78
rect 11106 254 11164 266
rect 12187 262 12199 450
rect 11106 78 11118 254
rect 11152 78 11164 254
rect 11106 66 11164 78
rect 11746 250 11804 262
rect 11746 74 11758 250
rect 11792 74 11804 250
rect 11746 62 11804 74
rect 11864 250 11922 262
rect 11864 74 11876 250
rect 11910 74 11922 250
rect 11864 62 11922 74
rect 11982 250 12040 262
rect 11982 74 11994 250
rect 12028 74 12040 250
rect 11982 62 12040 74
rect 12100 250 12199 262
rect 12100 74 12112 250
rect 12146 74 12199 250
rect 12233 74 12245 450
rect 12100 62 12245 74
rect 12305 450 12363 462
rect 12305 74 12317 450
rect 12351 74 12363 450
rect 12305 62 12363 74
rect 12423 450 12481 462
rect 12423 74 12435 450
rect 12469 74 12481 450
rect 12423 62 12481 74
rect 12541 450 12599 462
rect 12541 74 12553 450
rect 12587 74 12599 450
rect 12541 62 12599 74
rect 12654 450 12712 462
rect 12654 74 12666 450
rect 12700 74 12712 450
rect 12654 62 12712 74
rect 12772 450 12830 462
rect 12772 74 12784 450
rect 12818 74 12830 450
rect 12772 62 12830 74
rect 12890 450 12948 462
rect 12890 74 12902 450
rect 12936 74 12948 450
rect 12890 62 12948 74
rect 13008 450 13066 462
rect 13008 74 13020 450
rect 13054 74 13066 450
rect 13008 62 13066 74
rect 13126 450 13184 462
rect 13126 74 13138 450
rect 13172 74 13184 450
rect 13126 62 13184 74
rect 13244 450 13302 462
rect 13244 74 13256 450
rect 13290 74 13302 450
rect 13244 62 13302 74
rect 13362 450 13420 462
rect 13362 74 13374 450
rect 13408 74 13420 450
rect 13362 62 13420 74
rect 13481 450 13539 462
rect 13481 74 13493 450
rect 13527 74 13539 450
rect 13481 62 13539 74
rect 13599 450 13657 462
rect 13599 74 13611 450
rect 13645 74 13657 450
rect 13599 62 13657 74
rect 13717 450 13775 462
rect 13717 74 13729 450
rect 13763 74 13775 450
rect 13717 62 13775 74
rect 13835 450 13893 462
rect 13835 74 13847 450
rect 13881 74 13893 450
rect 15331 450 15389 462
rect 15331 262 15343 450
rect 13835 62 13893 74
rect 13954 250 14012 262
rect 13954 74 13966 250
rect 14000 74 14012 250
rect 13954 62 14012 74
rect 14072 250 14130 262
rect 14072 74 14084 250
rect 14118 74 14130 250
rect 14072 62 14130 74
rect 14190 250 14248 262
rect 14190 74 14202 250
rect 14236 74 14248 250
rect 14190 62 14248 74
rect 14308 250 14366 262
rect 14308 74 14320 250
rect 14354 74 14366 250
rect 14308 62 14366 74
rect 14890 250 14948 262
rect 14890 74 14902 250
rect 14936 74 14948 250
rect 14890 62 14948 74
rect 15008 250 15066 262
rect 15008 74 15020 250
rect 15054 74 15066 250
rect 15008 62 15066 74
rect 15126 250 15184 262
rect 15126 74 15138 250
rect 15172 74 15184 250
rect 15126 62 15184 74
rect 15244 250 15343 262
rect 15244 74 15256 250
rect 15290 74 15343 250
rect 15377 74 15389 450
rect 15244 62 15389 74
rect 15449 450 15507 462
rect 15449 74 15461 450
rect 15495 74 15507 450
rect 15449 62 15507 74
rect 15567 450 15625 462
rect 15567 74 15579 450
rect 15613 74 15625 450
rect 15567 62 15625 74
rect 15685 450 15743 462
rect 15685 74 15697 450
rect 15731 74 15743 450
rect 15685 62 15743 74
rect 15798 450 15856 462
rect 15798 74 15810 450
rect 15844 74 15856 450
rect 15798 62 15856 74
rect 15916 450 15974 462
rect 15916 74 15928 450
rect 15962 74 15974 450
rect 15916 62 15974 74
rect 16034 450 16092 462
rect 16034 74 16046 450
rect 16080 74 16092 450
rect 16034 62 16092 74
rect 16152 450 16210 462
rect 16152 74 16164 450
rect 16198 74 16210 450
rect 16152 62 16210 74
rect 16270 450 16328 462
rect 16270 74 16282 450
rect 16316 74 16328 450
rect 16270 62 16328 74
rect 16388 450 16446 462
rect 16388 74 16400 450
rect 16434 74 16446 450
rect 16388 62 16446 74
rect 16506 450 16564 462
rect 16506 74 16518 450
rect 16552 74 16564 450
rect 16506 62 16564 74
rect 16625 450 16683 462
rect 16625 74 16637 450
rect 16671 74 16683 450
rect 16625 62 16683 74
rect 16743 450 16801 462
rect 16743 74 16755 450
rect 16789 74 16801 450
rect 16743 62 16801 74
rect 16861 450 16919 462
rect 16861 74 16873 450
rect 16907 74 16919 450
rect 16861 62 16919 74
rect 16979 450 17037 462
rect 16979 74 16991 450
rect 17025 74 17037 450
rect 18463 454 18521 466
rect 18463 266 18475 454
rect 16979 62 17037 74
rect 17098 250 17156 262
rect 17098 74 17110 250
rect 17144 74 17156 250
rect 17098 62 17156 74
rect 17216 250 17274 262
rect 17216 74 17228 250
rect 17262 74 17274 250
rect 17216 62 17274 74
rect 17334 250 17392 262
rect 17334 74 17346 250
rect 17380 74 17392 250
rect 17334 62 17392 74
rect 17452 250 17510 262
rect 17452 74 17464 250
rect 17498 74 17510 250
rect 17452 62 17510 74
rect 18022 254 18080 266
rect 18022 78 18034 254
rect 18068 78 18080 254
rect 18022 66 18080 78
rect 18140 254 18198 266
rect 18140 78 18152 254
rect 18186 78 18198 254
rect 18140 66 18198 78
rect 18258 254 18316 266
rect 18258 78 18270 254
rect 18304 78 18316 254
rect 18258 66 18316 78
rect 18376 254 18475 266
rect 18376 78 18388 254
rect 18422 78 18475 254
rect 18509 78 18521 454
rect 18376 66 18521 78
rect 18581 454 18639 466
rect 18581 78 18593 454
rect 18627 78 18639 454
rect 18581 66 18639 78
rect 18699 454 18757 466
rect 18699 78 18711 454
rect 18745 78 18757 454
rect 18699 66 18757 78
rect 18817 454 18875 466
rect 18817 78 18829 454
rect 18863 78 18875 454
rect 18817 66 18875 78
rect 18930 454 18988 466
rect 18930 78 18942 454
rect 18976 78 18988 454
rect 18930 66 18988 78
rect 19048 454 19106 466
rect 19048 78 19060 454
rect 19094 78 19106 454
rect 19048 66 19106 78
rect 19166 454 19224 466
rect 19166 78 19178 454
rect 19212 78 19224 454
rect 19166 66 19224 78
rect 19284 454 19342 466
rect 19284 78 19296 454
rect 19330 78 19342 454
rect 19284 66 19342 78
rect 19402 454 19460 466
rect 19402 78 19414 454
rect 19448 78 19460 454
rect 19402 66 19460 78
rect 19520 454 19578 466
rect 19520 78 19532 454
rect 19566 78 19578 454
rect 19520 66 19578 78
rect 19638 454 19696 466
rect 19638 78 19650 454
rect 19684 78 19696 454
rect 19638 66 19696 78
rect 19757 454 19815 466
rect 19757 78 19769 454
rect 19803 78 19815 454
rect 19757 66 19815 78
rect 19875 454 19933 466
rect 19875 78 19887 454
rect 19921 78 19933 454
rect 19875 66 19933 78
rect 19993 454 20051 466
rect 19993 78 20005 454
rect 20039 78 20051 454
rect 19993 66 20051 78
rect 20111 454 20169 466
rect 20111 78 20123 454
rect 20157 78 20169 454
rect 21607 454 21665 466
rect 21607 266 21619 454
rect 20111 66 20169 78
rect 20230 254 20288 266
rect 20230 78 20242 254
rect 20276 78 20288 254
rect 20230 66 20288 78
rect 20348 254 20406 266
rect 20348 78 20360 254
rect 20394 78 20406 254
rect 20348 66 20406 78
rect 20466 254 20524 266
rect 20466 78 20478 254
rect 20512 78 20524 254
rect 20466 66 20524 78
rect 20584 254 20642 266
rect 20584 78 20596 254
rect 20630 78 20642 254
rect 20584 66 20642 78
rect 21166 254 21224 266
rect 21166 78 21178 254
rect 21212 78 21224 254
rect 21166 66 21224 78
rect 21284 254 21342 266
rect 21284 78 21296 254
rect 21330 78 21342 254
rect 21284 66 21342 78
rect 21402 254 21460 266
rect 21402 78 21414 254
rect 21448 78 21460 254
rect 21402 66 21460 78
rect 21520 254 21619 266
rect 21520 78 21532 254
rect 21566 78 21619 254
rect 21653 78 21665 454
rect 21520 66 21665 78
rect 21725 454 21783 466
rect 21725 78 21737 454
rect 21771 78 21783 454
rect 21725 66 21783 78
rect 21843 454 21901 466
rect 21843 78 21855 454
rect 21889 78 21901 454
rect 21843 66 21901 78
rect 21961 454 22019 466
rect 21961 78 21973 454
rect 22007 78 22019 454
rect 21961 66 22019 78
rect 22074 454 22132 466
rect 22074 78 22086 454
rect 22120 78 22132 454
rect 22074 66 22132 78
rect 22192 454 22250 466
rect 22192 78 22204 454
rect 22238 78 22250 454
rect 22192 66 22250 78
rect 22310 454 22368 466
rect 22310 78 22322 454
rect 22356 78 22368 454
rect 22310 66 22368 78
rect 22428 454 22486 466
rect 22428 78 22440 454
rect 22474 78 22486 454
rect 22428 66 22486 78
rect 22546 454 22604 466
rect 22546 78 22558 454
rect 22592 78 22604 454
rect 22546 66 22604 78
rect 22664 454 22722 466
rect 22664 78 22676 454
rect 22710 78 22722 454
rect 22664 66 22722 78
rect 22782 454 22840 466
rect 22782 78 22794 454
rect 22828 78 22840 454
rect 22782 66 22840 78
rect 22901 454 22959 466
rect 22901 78 22913 454
rect 22947 78 22959 454
rect 22901 66 22959 78
rect 23019 454 23077 466
rect 23019 78 23031 454
rect 23065 78 23077 454
rect 23019 66 23077 78
rect 23137 454 23195 466
rect 23137 78 23149 454
rect 23183 78 23195 454
rect 23137 66 23195 78
rect 23255 454 23313 466
rect 23255 78 23267 454
rect 23301 78 23313 454
rect 23255 66 23313 78
rect 23374 254 23432 266
rect 23374 78 23386 254
rect 23420 78 23432 254
rect 23374 66 23432 78
rect 23492 254 23550 266
rect 23492 78 23504 254
rect 23538 78 23550 254
rect 23492 66 23550 78
rect 23610 254 23668 266
rect 23610 78 23622 254
rect 23656 78 23668 254
rect 23610 66 23668 78
rect 23728 254 23786 266
rect 23728 78 23740 254
rect 23774 78 23786 254
rect 23728 66 23786 78
<< ndiffc >>
rect -30 -1059 4 -883
rect 88 -1059 122 -883
rect 162 -1259 196 -883
rect 280 -1259 314 -883
rect 398 -1259 432 -883
rect 516 -1259 550 -883
rect 634 -1259 668 -883
rect 712 -1059 746 -883
rect 830 -1059 864 -883
rect 3114 -1059 3148 -883
rect 3232 -1059 3266 -883
rect 3306 -1259 3340 -883
rect 3424 -1259 3458 -883
rect 3542 -1259 3576 -883
rect 3660 -1259 3694 -883
rect 3778 -1259 3812 -883
rect 3856 -1059 3890 -883
rect 3974 -1059 4008 -883
rect 6246 -1055 6280 -879
rect 6364 -1055 6398 -879
rect 6438 -1255 6472 -879
rect 6556 -1255 6590 -879
rect 6674 -1255 6708 -879
rect 6792 -1255 6826 -879
rect 6910 -1255 6944 -879
rect 6988 -1055 7022 -879
rect 7106 -1055 7140 -879
rect 9390 -1055 9424 -879
rect 9508 -1055 9542 -879
rect 9582 -1255 9616 -879
rect 9700 -1255 9734 -879
rect 9818 -1255 9852 -879
rect 9936 -1255 9970 -879
rect 10054 -1255 10088 -879
rect 10132 -1055 10166 -879
rect 10250 -1055 10284 -879
rect 12592 -1059 12626 -883
rect 12710 -1059 12744 -883
rect 12784 -1259 12818 -883
rect 12902 -1259 12936 -883
rect 13020 -1259 13054 -883
rect 13138 -1259 13172 -883
rect 13256 -1259 13290 -883
rect 13334 -1059 13368 -883
rect 13452 -1059 13486 -883
rect 15736 -1059 15770 -883
rect 15854 -1059 15888 -883
rect 15928 -1259 15962 -883
rect 16046 -1259 16080 -883
rect 16164 -1259 16198 -883
rect 16282 -1259 16316 -883
rect 16400 -1259 16434 -883
rect 16478 -1059 16512 -883
rect 16596 -1059 16630 -883
rect 18868 -1055 18902 -879
rect 18986 -1055 19020 -879
rect 19060 -1255 19094 -879
rect 19178 -1255 19212 -879
rect 19296 -1255 19330 -879
rect 19414 -1255 19448 -879
rect 19532 -1255 19566 -879
rect 19610 -1055 19644 -879
rect 19728 -1055 19762 -879
rect 22012 -1055 22046 -879
rect 22130 -1055 22164 -879
rect 22204 -1255 22238 -879
rect 22322 -1255 22356 -879
rect 22440 -1255 22474 -879
rect 22558 -1255 22592 -879
rect 22676 -1255 22710 -879
rect 22754 -1055 22788 -879
rect 22872 -1055 22906 -879
<< pdiffc >>
rect -864 74 -830 250
rect -746 74 -712 250
rect -628 74 -594 250
rect -510 74 -476 250
rect -423 74 -389 450
rect -305 74 -271 450
rect -187 74 -153 450
rect -69 74 -35 450
rect 44 74 78 450
rect 162 74 196 450
rect 280 74 314 450
rect 398 74 432 450
rect 516 74 550 450
rect 634 74 668 450
rect 752 74 786 450
rect 871 74 905 450
rect 989 74 1023 450
rect 1107 74 1141 450
rect 1225 74 1259 450
rect 1344 74 1378 250
rect 1462 74 1496 250
rect 1580 74 1614 250
rect 1698 74 1732 250
rect 2280 74 2314 250
rect 2398 74 2432 250
rect 2516 74 2550 250
rect 2634 74 2668 250
rect 2721 74 2755 450
rect 2839 74 2873 450
rect 2957 74 2991 450
rect 3075 74 3109 450
rect 3188 74 3222 450
rect 3306 74 3340 450
rect 3424 74 3458 450
rect 3542 74 3576 450
rect 3660 74 3694 450
rect 3778 74 3812 450
rect 3896 74 3930 450
rect 4015 74 4049 450
rect 4133 74 4167 450
rect 4251 74 4285 450
rect 4369 74 4403 450
rect 4488 74 4522 250
rect 4606 74 4640 250
rect 4724 74 4758 250
rect 4842 74 4876 250
rect 5412 78 5446 254
rect 5530 78 5564 254
rect 5648 78 5682 254
rect 5766 78 5800 254
rect 5853 78 5887 454
rect 5971 78 6005 454
rect 6089 78 6123 454
rect 6207 78 6241 454
rect 6320 78 6354 454
rect 6438 78 6472 454
rect 6556 78 6590 454
rect 6674 78 6708 454
rect 6792 78 6826 454
rect 6910 78 6944 454
rect 7028 78 7062 454
rect 7147 78 7181 454
rect 7265 78 7299 454
rect 7383 78 7417 454
rect 7501 78 7535 454
rect 7620 78 7654 254
rect 7738 78 7772 254
rect 7856 78 7890 254
rect 7974 78 8008 254
rect 8556 78 8590 254
rect 8674 78 8708 254
rect 8792 78 8826 254
rect 8910 78 8944 254
rect 8997 78 9031 454
rect 9115 78 9149 454
rect 9233 78 9267 454
rect 9351 78 9385 454
rect 9464 78 9498 454
rect 9582 78 9616 454
rect 9700 78 9734 454
rect 9818 78 9852 454
rect 9936 78 9970 454
rect 10054 78 10088 454
rect 10172 78 10206 454
rect 10291 78 10325 454
rect 10409 78 10443 454
rect 10527 78 10561 454
rect 10645 78 10679 454
rect 10764 78 10798 254
rect 10882 78 10916 254
rect 11000 78 11034 254
rect 11118 78 11152 254
rect 11758 74 11792 250
rect 11876 74 11910 250
rect 11994 74 12028 250
rect 12112 74 12146 250
rect 12199 74 12233 450
rect 12317 74 12351 450
rect 12435 74 12469 450
rect 12553 74 12587 450
rect 12666 74 12700 450
rect 12784 74 12818 450
rect 12902 74 12936 450
rect 13020 74 13054 450
rect 13138 74 13172 450
rect 13256 74 13290 450
rect 13374 74 13408 450
rect 13493 74 13527 450
rect 13611 74 13645 450
rect 13729 74 13763 450
rect 13847 74 13881 450
rect 13966 74 14000 250
rect 14084 74 14118 250
rect 14202 74 14236 250
rect 14320 74 14354 250
rect 14902 74 14936 250
rect 15020 74 15054 250
rect 15138 74 15172 250
rect 15256 74 15290 250
rect 15343 74 15377 450
rect 15461 74 15495 450
rect 15579 74 15613 450
rect 15697 74 15731 450
rect 15810 74 15844 450
rect 15928 74 15962 450
rect 16046 74 16080 450
rect 16164 74 16198 450
rect 16282 74 16316 450
rect 16400 74 16434 450
rect 16518 74 16552 450
rect 16637 74 16671 450
rect 16755 74 16789 450
rect 16873 74 16907 450
rect 16991 74 17025 450
rect 17110 74 17144 250
rect 17228 74 17262 250
rect 17346 74 17380 250
rect 17464 74 17498 250
rect 18034 78 18068 254
rect 18152 78 18186 254
rect 18270 78 18304 254
rect 18388 78 18422 254
rect 18475 78 18509 454
rect 18593 78 18627 454
rect 18711 78 18745 454
rect 18829 78 18863 454
rect 18942 78 18976 454
rect 19060 78 19094 454
rect 19178 78 19212 454
rect 19296 78 19330 454
rect 19414 78 19448 454
rect 19532 78 19566 454
rect 19650 78 19684 454
rect 19769 78 19803 454
rect 19887 78 19921 454
rect 20005 78 20039 454
rect 20123 78 20157 454
rect 20242 78 20276 254
rect 20360 78 20394 254
rect 20478 78 20512 254
rect 20596 78 20630 254
rect 21178 78 21212 254
rect 21296 78 21330 254
rect 21414 78 21448 254
rect 21532 78 21566 254
rect 21619 78 21653 454
rect 21737 78 21771 454
rect 21855 78 21889 454
rect 21973 78 22007 454
rect 22086 78 22120 454
rect 22204 78 22238 454
rect 22322 78 22356 454
rect 22440 78 22474 454
rect 22558 78 22592 454
rect 22676 78 22710 454
rect 22794 78 22828 454
rect 22913 78 22947 454
rect 23031 78 23065 454
rect 23149 78 23183 454
rect 23267 78 23301 454
rect 23386 78 23420 254
rect 23504 78 23538 254
rect 23622 78 23656 254
rect 23740 78 23774 254
<< psubdiff >>
rect 338 -1526 524 -1502
rect 338 -1572 380 -1526
rect 484 -1572 524 -1526
rect 338 -1608 524 -1572
rect 3482 -1526 3668 -1502
rect 3482 -1572 3524 -1526
rect 3628 -1572 3668 -1526
rect 3482 -1608 3668 -1572
rect 6614 -1522 6800 -1498
rect 6614 -1568 6656 -1522
rect 6760 -1568 6800 -1522
rect 6614 -1604 6800 -1568
rect 9758 -1522 9944 -1498
rect 9758 -1568 9800 -1522
rect 9904 -1568 9944 -1522
rect 9758 -1604 9944 -1568
rect 12960 -1526 13146 -1502
rect 12960 -1572 13002 -1526
rect 13106 -1572 13146 -1526
rect 12960 -1608 13146 -1572
rect 16104 -1526 16290 -1502
rect 16104 -1572 16146 -1526
rect 16250 -1572 16290 -1526
rect 16104 -1608 16290 -1572
rect 19236 -1522 19422 -1498
rect 19236 -1568 19278 -1522
rect 19382 -1568 19422 -1522
rect 19236 -1604 19422 -1568
rect 22380 -1522 22566 -1498
rect 22380 -1568 22422 -1522
rect 22526 -1568 22566 -1522
rect 22380 -1604 22566 -1568
<< nsubdiff >>
rect 268 720 572 776
rect 268 644 322 720
rect 518 644 572 720
rect 268 630 572 644
rect 3412 720 3716 776
rect 3412 644 3466 720
rect 3662 644 3716 720
rect 3412 630 3716 644
rect 6544 724 6848 780
rect 6544 648 6598 724
rect 6794 648 6848 724
rect 6544 634 6848 648
rect 9688 724 9992 780
rect 9688 648 9742 724
rect 9938 648 9992 724
rect 9688 634 9992 648
rect 12890 720 13194 776
rect 12890 644 12944 720
rect 13140 644 13194 720
rect 12890 630 13194 644
rect 16034 720 16338 776
rect 16034 644 16088 720
rect 16284 644 16338 720
rect 16034 630 16338 644
rect 19166 724 19470 780
rect 19166 648 19220 724
rect 19416 648 19470 724
rect 19166 634 19470 648
rect 22310 724 22614 780
rect 22310 648 22364 724
rect 22560 648 22614 724
rect 22310 634 22614 648
<< psubdiffcont >>
rect 380 -1572 484 -1526
rect 3524 -1572 3628 -1526
rect 6656 -1568 6760 -1522
rect 9800 -1568 9904 -1522
rect 13002 -1572 13106 -1526
rect 16146 -1572 16250 -1526
rect 19278 -1568 19382 -1522
rect 22422 -1568 22526 -1522
<< nsubdiffcont >>
rect 322 644 518 720
rect 3466 644 3662 720
rect 6598 648 6794 724
rect 9742 648 9938 724
rect 12944 644 13140 720
rect 16088 644 16284 720
rect 19220 648 19416 724
rect 22364 648 22560 724
<< poly >>
rect -377 477 -81 516
rect -377 462 -317 477
rect -259 462 -199 477
rect -141 462 -81 477
rect 90 477 386 516
rect 90 462 150 477
rect 208 462 268 477
rect 326 462 386 477
rect 444 477 740 516
rect 444 462 504 477
rect 562 462 622 477
rect 680 462 740 477
rect 917 477 1213 516
rect 917 462 977 477
rect 1035 462 1095 477
rect 1153 462 1213 477
rect 2767 477 3063 516
rect 2767 462 2827 477
rect 2885 462 2945 477
rect 3003 462 3063 477
rect 3234 477 3530 516
rect 3234 462 3294 477
rect 3352 462 3412 477
rect 3470 462 3530 477
rect 3588 477 3884 516
rect 3588 462 3648 477
rect 3706 462 3766 477
rect 3824 462 3884 477
rect 4061 477 4357 516
rect 4061 462 4121 477
rect 4179 462 4239 477
rect 4297 462 4357 477
rect 5899 481 6195 520
rect 5899 466 5959 481
rect 6017 466 6077 481
rect 6135 466 6195 481
rect 6366 481 6662 520
rect 6366 466 6426 481
rect 6484 466 6544 481
rect 6602 466 6662 481
rect 6720 481 7016 520
rect 6720 466 6780 481
rect 6838 466 6898 481
rect 6956 466 7016 481
rect 7193 481 7489 520
rect 7193 466 7253 481
rect 7311 466 7371 481
rect 7429 466 7489 481
rect 9043 481 9339 520
rect 9043 466 9103 481
rect 9161 466 9221 481
rect 9279 466 9339 481
rect 9510 481 9806 520
rect 9510 466 9570 481
rect 9628 466 9688 481
rect 9746 466 9806 481
rect 9864 481 10160 520
rect 9864 466 9924 481
rect 9982 466 10042 481
rect 10100 466 10160 481
rect 10337 481 10633 520
rect 10337 466 10397 481
rect 10455 466 10515 481
rect 10573 466 10633 481
rect 12245 477 12541 516
rect -818 278 -522 317
rect -818 262 -758 278
rect -700 262 -640 278
rect -582 262 -522 278
rect 1390 278 1686 317
rect 1390 262 1450 278
rect 1508 262 1568 278
rect 1626 262 1686 278
rect 2326 278 2622 317
rect 2326 262 2386 278
rect 2444 262 2504 278
rect 2562 262 2622 278
rect 4534 278 4830 317
rect 4534 262 4594 278
rect 4652 262 4712 278
rect 4770 262 4830 278
rect 5458 282 5754 321
rect 5458 266 5518 282
rect 5576 266 5636 282
rect 5694 266 5754 282
rect 7666 282 7962 321
rect 7666 266 7726 282
rect 7784 266 7844 282
rect 7902 266 7962 282
rect 8602 282 8898 321
rect 8602 266 8662 282
rect 8720 266 8780 282
rect 8838 266 8898 282
rect 12245 462 12305 477
rect 12363 462 12423 477
rect 12481 462 12541 477
rect 12712 477 13008 516
rect 12712 462 12772 477
rect 12830 462 12890 477
rect 12948 462 13008 477
rect 13066 477 13362 516
rect 13066 462 13126 477
rect 13184 462 13244 477
rect 13302 462 13362 477
rect 13539 477 13835 516
rect 13539 462 13599 477
rect 13657 462 13717 477
rect 13775 462 13835 477
rect 15389 477 15685 516
rect 15389 462 15449 477
rect 15507 462 15567 477
rect 15625 462 15685 477
rect 15856 477 16152 516
rect 15856 462 15916 477
rect 15974 462 16034 477
rect 16092 462 16152 477
rect 16210 477 16506 516
rect 16210 462 16270 477
rect 16328 462 16388 477
rect 16446 462 16506 477
rect 16683 477 16979 516
rect 16683 462 16743 477
rect 16801 462 16861 477
rect 16919 462 16979 477
rect 18521 481 18817 520
rect 18521 466 18581 481
rect 18639 466 18699 481
rect 18757 466 18817 481
rect 18988 481 19284 520
rect 18988 466 19048 481
rect 19106 466 19166 481
rect 19224 466 19284 481
rect 19342 481 19638 520
rect 19342 466 19402 481
rect 19460 466 19520 481
rect 19578 466 19638 481
rect 19815 481 20111 520
rect 19815 466 19875 481
rect 19933 466 19993 481
rect 20051 466 20111 481
rect 21665 481 21961 520
rect 21665 466 21725 481
rect 21783 466 21843 481
rect 21901 466 21961 481
rect 22132 481 22428 520
rect 22132 466 22192 481
rect 22250 466 22310 481
rect 22368 466 22428 481
rect 22486 481 22782 520
rect 22486 466 22546 481
rect 22604 466 22664 481
rect 22722 466 22782 481
rect 22959 481 23255 520
rect 22959 466 23019 481
rect 23077 466 23137 481
rect 23195 466 23255 481
rect 10810 282 11106 321
rect 10810 266 10870 282
rect 10928 266 10988 282
rect 11046 266 11106 282
rect 11804 278 12100 317
rect 11804 262 11864 278
rect 11922 262 11982 278
rect 12040 262 12100 278
rect -818 -224 -758 62
rect -700 36 -640 62
rect -582 36 -522 62
rect -377 36 -317 62
rect -818 -241 -682 -224
rect -818 -296 -759 -241
rect -701 -296 -682 -241
rect -818 -311 -682 -296
rect -818 -623 -758 -311
rect -259 -356 -199 62
rect -141 36 -81 62
rect 90 36 150 62
rect 208 36 268 62
rect 326 36 386 62
rect 444 36 504 62
rect 209 -124 268 36
rect 209 -125 272 -124
rect 206 -141 272 -125
rect 206 -175 222 -141
rect 256 -175 272 -141
rect 206 -191 272 -175
rect 309 -240 404 -225
rect 309 -295 328 -240
rect 386 -263 404 -240
rect 562 -263 622 62
rect 680 36 740 62
rect 917 36 977 62
rect 386 -295 622 -263
rect 309 -312 622 -295
rect -259 -413 268 -356
rect 208 -512 268 -413
rect 197 -525 278 -512
rect 197 -580 210 -525
rect 268 -580 278 -525
rect 197 -591 278 -580
rect -818 -668 76 -623
rect 16 -871 76 -668
rect 208 -871 268 -591
rect 326 -871 386 -312
rect 1035 -354 1095 62
rect 1153 36 1213 62
rect 1390 36 1450 62
rect 1508 36 1568 62
rect 1516 -87 1582 -84
rect 1626 -87 1686 62
rect 1516 -100 1686 -87
rect 1516 -134 1532 -100
rect 1566 -134 1686 -100
rect 1516 -147 1686 -134
rect 1516 -150 1582 -147
rect 557 -371 1095 -354
rect 557 -405 576 -371
rect 610 -405 1095 -371
rect 557 -411 1095 -405
rect 557 -421 626 -411
rect 557 -423 622 -421
rect 441 -761 507 -745
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect 444 -871 504 -811
rect 562 -871 622 -423
rect 1626 -623 1686 -147
rect 758 -668 1686 -623
rect 2326 -224 2386 62
rect 2444 36 2504 62
rect 2562 36 2622 62
rect 2767 36 2827 62
rect 2326 -241 2462 -224
rect 2326 -296 2385 -241
rect 2443 -296 2462 -241
rect 2326 -311 2462 -296
rect 2326 -623 2386 -311
rect 2885 -356 2945 62
rect 3003 36 3063 62
rect 3234 36 3294 62
rect 3352 36 3412 62
rect 3470 36 3530 62
rect 3588 36 3648 62
rect 3353 -124 3412 36
rect 3353 -125 3416 -124
rect 3350 -141 3416 -125
rect 3350 -175 3366 -141
rect 3400 -175 3416 -141
rect 3350 -191 3416 -175
rect 3453 -240 3548 -225
rect 3453 -295 3472 -240
rect 3530 -263 3548 -240
rect 3706 -263 3766 62
rect 3824 36 3884 62
rect 4061 36 4121 62
rect 3530 -295 3766 -263
rect 3453 -312 3766 -295
rect 2885 -413 3412 -356
rect 3352 -512 3412 -413
rect 3341 -525 3422 -512
rect 3341 -580 3354 -525
rect 3412 -580 3422 -525
rect 3341 -591 3422 -580
rect 2326 -668 3220 -623
rect 758 -871 818 -668
rect 3160 -871 3220 -668
rect 3352 -871 3412 -591
rect 3470 -871 3530 -312
rect 4179 -354 4239 62
rect 4297 36 4357 62
rect 4534 36 4594 62
rect 4652 36 4712 62
rect 4660 -87 4726 -84
rect 4770 -87 4830 62
rect 4660 -100 4830 -87
rect 4660 -134 4676 -100
rect 4710 -134 4830 -100
rect 4660 -147 4830 -134
rect 4660 -150 4726 -147
rect 3701 -371 4239 -354
rect 3701 -405 3720 -371
rect 3754 -405 4239 -371
rect 3701 -411 4239 -405
rect 3701 -421 3770 -411
rect 3701 -423 3766 -421
rect 3585 -761 3651 -745
rect 3585 -795 3601 -761
rect 3635 -795 3651 -761
rect 3585 -811 3651 -795
rect 3588 -871 3648 -811
rect 3706 -871 3766 -423
rect 4770 -623 4830 -147
rect 3902 -668 4830 -623
rect 5458 -220 5518 66
rect 5576 40 5636 66
rect 5694 40 5754 66
rect 5899 40 5959 66
rect 5458 -237 5594 -220
rect 5458 -292 5517 -237
rect 5575 -292 5594 -237
rect 5458 -307 5594 -292
rect 5458 -619 5518 -307
rect 6017 -352 6077 66
rect 6135 40 6195 66
rect 6366 40 6426 66
rect 6484 40 6544 66
rect 6602 40 6662 66
rect 6720 40 6780 66
rect 6485 -120 6544 40
rect 6485 -121 6548 -120
rect 6482 -137 6548 -121
rect 6482 -171 6498 -137
rect 6532 -171 6548 -137
rect 6482 -187 6548 -171
rect 6585 -236 6680 -221
rect 6585 -291 6604 -236
rect 6662 -259 6680 -236
rect 6838 -259 6898 66
rect 6956 40 7016 66
rect 7193 40 7253 66
rect 6662 -291 6898 -259
rect 6585 -308 6898 -291
rect 6017 -409 6544 -352
rect 6484 -508 6544 -409
rect 6473 -521 6554 -508
rect 6473 -576 6486 -521
rect 6544 -576 6554 -521
rect 6473 -587 6554 -576
rect 5458 -664 6352 -619
rect 3902 -871 3962 -668
rect 6292 -867 6352 -664
rect 6484 -867 6544 -587
rect 6602 -867 6662 -308
rect 7311 -350 7371 66
rect 7429 40 7489 66
rect 7666 40 7726 66
rect 7784 40 7844 66
rect 7792 -83 7858 -80
rect 7902 -83 7962 66
rect 7792 -96 7962 -83
rect 7792 -130 7808 -96
rect 7842 -130 7962 -96
rect 7792 -143 7962 -130
rect 7792 -146 7858 -143
rect 6833 -367 7371 -350
rect 6833 -401 6852 -367
rect 6886 -401 7371 -367
rect 6833 -407 7371 -401
rect 6833 -417 6902 -407
rect 6833 -419 6898 -417
rect 6717 -757 6783 -741
rect 6717 -791 6733 -757
rect 6767 -791 6783 -757
rect 6717 -807 6783 -791
rect 6720 -867 6780 -807
rect 6838 -867 6898 -419
rect 7902 -619 7962 -143
rect 7034 -664 7962 -619
rect 8602 -220 8662 66
rect 8720 40 8780 66
rect 8838 40 8898 66
rect 9043 40 9103 66
rect 8602 -237 8738 -220
rect 8602 -292 8661 -237
rect 8719 -292 8738 -237
rect 8602 -307 8738 -292
rect 8602 -619 8662 -307
rect 9161 -352 9221 66
rect 9279 40 9339 66
rect 9510 40 9570 66
rect 9628 40 9688 66
rect 9746 40 9806 66
rect 9864 40 9924 66
rect 9629 -120 9688 40
rect 9629 -121 9692 -120
rect 9626 -137 9692 -121
rect 9626 -171 9642 -137
rect 9676 -171 9692 -137
rect 9626 -187 9692 -171
rect 9729 -236 9824 -221
rect 9729 -291 9748 -236
rect 9806 -259 9824 -236
rect 9982 -259 10042 66
rect 10100 40 10160 66
rect 10337 40 10397 66
rect 9806 -291 10042 -259
rect 9729 -308 10042 -291
rect 9161 -409 9688 -352
rect 9628 -508 9688 -409
rect 9617 -521 9698 -508
rect 9617 -576 9630 -521
rect 9688 -576 9698 -521
rect 9617 -587 9698 -576
rect 8602 -664 9496 -619
rect 7034 -867 7094 -664
rect 9436 -867 9496 -664
rect 9628 -867 9688 -587
rect 9746 -867 9806 -308
rect 10455 -350 10515 66
rect 10573 40 10633 66
rect 10810 40 10870 66
rect 10928 40 10988 66
rect 10936 -83 11002 -80
rect 11046 -83 11106 66
rect 14012 278 14308 317
rect 14012 262 14072 278
rect 14130 262 14190 278
rect 14248 262 14308 278
rect 14948 278 15244 317
rect 14948 262 15008 278
rect 15066 262 15126 278
rect 15184 262 15244 278
rect 17156 278 17452 317
rect 17156 262 17216 278
rect 17274 262 17334 278
rect 17392 262 17452 278
rect 18080 282 18376 321
rect 18080 266 18140 282
rect 18198 266 18258 282
rect 18316 266 18376 282
rect 20288 282 20584 321
rect 20288 266 20348 282
rect 20406 266 20466 282
rect 20524 266 20584 282
rect 21224 282 21520 321
rect 21224 266 21284 282
rect 21342 266 21402 282
rect 21460 266 21520 282
rect 23432 282 23728 321
rect 23432 266 23492 282
rect 23550 266 23610 282
rect 23668 266 23728 282
rect 10936 -96 11106 -83
rect 10936 -130 10952 -96
rect 10986 -130 11106 -96
rect 10936 -143 11106 -130
rect 10936 -146 11002 -143
rect 9977 -367 10515 -350
rect 9977 -401 9996 -367
rect 10030 -401 10515 -367
rect 9977 -407 10515 -401
rect 9977 -417 10046 -407
rect 9977 -419 10042 -417
rect 9861 -757 9927 -741
rect 9861 -791 9877 -757
rect 9911 -791 9927 -757
rect 9861 -807 9927 -791
rect 9864 -867 9924 -807
rect 9982 -867 10042 -419
rect 11046 -619 11106 -143
rect 10178 -664 11106 -619
rect 11804 -224 11864 62
rect 11922 36 11982 62
rect 12040 36 12100 62
rect 12245 36 12305 62
rect 11804 -241 11940 -224
rect 11804 -296 11863 -241
rect 11921 -296 11940 -241
rect 11804 -311 11940 -296
rect 11804 -623 11864 -311
rect 12363 -356 12423 62
rect 12481 36 12541 62
rect 12712 36 12772 62
rect 12830 36 12890 62
rect 12948 36 13008 62
rect 13066 36 13126 62
rect 12831 -124 12890 36
rect 12831 -125 12894 -124
rect 12828 -141 12894 -125
rect 12828 -175 12844 -141
rect 12878 -175 12894 -141
rect 12828 -191 12894 -175
rect 12931 -240 13026 -225
rect 12931 -295 12950 -240
rect 13008 -263 13026 -240
rect 13184 -263 13244 62
rect 13302 36 13362 62
rect 13539 36 13599 62
rect 13008 -295 13244 -263
rect 12931 -312 13244 -295
rect 12363 -413 12890 -356
rect 12830 -512 12890 -413
rect 12819 -525 12900 -512
rect 12819 -580 12832 -525
rect 12890 -580 12900 -525
rect 12819 -591 12900 -580
rect 10178 -867 10238 -664
rect 11804 -668 12698 -623
rect 16 -1097 76 -1071
rect 208 -1297 268 -1271
rect 326 -1297 386 -1271
rect 444 -1297 504 -1271
rect 562 -1297 622 -1271
rect 383 -1352 449 -1344
rect 758 -1352 818 -1071
rect 3160 -1097 3220 -1071
rect 3352 -1297 3412 -1271
rect 3470 -1297 3530 -1271
rect 3588 -1297 3648 -1271
rect 3706 -1297 3766 -1271
rect 383 -1360 818 -1352
rect 383 -1394 399 -1360
rect 433 -1394 818 -1360
rect 383 -1403 818 -1394
rect 3527 -1352 3593 -1344
rect 3902 -1352 3962 -1071
rect 6292 -1093 6352 -1067
rect 6484 -1293 6544 -1267
rect 6602 -1293 6662 -1267
rect 6720 -1293 6780 -1267
rect 6838 -1293 6898 -1267
rect 3527 -1360 3962 -1352
rect 3527 -1394 3543 -1360
rect 3577 -1394 3962 -1360
rect 3527 -1403 3962 -1394
rect 6659 -1348 6725 -1340
rect 7034 -1348 7094 -1067
rect 9436 -1093 9496 -1067
rect 12638 -871 12698 -668
rect 12830 -871 12890 -591
rect 12948 -871 13008 -312
rect 13657 -354 13717 62
rect 13775 36 13835 62
rect 14012 36 14072 62
rect 14130 36 14190 62
rect 14138 -87 14204 -84
rect 14248 -87 14308 62
rect 14138 -100 14308 -87
rect 14138 -134 14154 -100
rect 14188 -134 14308 -100
rect 14138 -147 14308 -134
rect 14138 -150 14204 -147
rect 13179 -371 13717 -354
rect 13179 -405 13198 -371
rect 13232 -405 13717 -371
rect 13179 -411 13717 -405
rect 13179 -421 13248 -411
rect 13179 -423 13244 -421
rect 13063 -761 13129 -745
rect 13063 -795 13079 -761
rect 13113 -795 13129 -761
rect 13063 -811 13129 -795
rect 13066 -871 13126 -811
rect 13184 -871 13244 -423
rect 14248 -623 14308 -147
rect 13380 -668 14308 -623
rect 14948 -224 15008 62
rect 15066 36 15126 62
rect 15184 36 15244 62
rect 15389 36 15449 62
rect 14948 -241 15084 -224
rect 14948 -296 15007 -241
rect 15065 -296 15084 -241
rect 14948 -311 15084 -296
rect 14948 -623 15008 -311
rect 15507 -356 15567 62
rect 15625 36 15685 62
rect 15856 36 15916 62
rect 15974 36 16034 62
rect 16092 36 16152 62
rect 16210 36 16270 62
rect 15975 -124 16034 36
rect 15975 -125 16038 -124
rect 15972 -141 16038 -125
rect 15972 -175 15988 -141
rect 16022 -175 16038 -141
rect 15972 -191 16038 -175
rect 16075 -240 16170 -225
rect 16075 -295 16094 -240
rect 16152 -263 16170 -240
rect 16328 -263 16388 62
rect 16446 36 16506 62
rect 16683 36 16743 62
rect 16152 -295 16388 -263
rect 16075 -312 16388 -295
rect 15507 -413 16034 -356
rect 15974 -512 16034 -413
rect 15963 -525 16044 -512
rect 15963 -580 15976 -525
rect 16034 -580 16044 -525
rect 15963 -591 16044 -580
rect 14948 -668 15842 -623
rect 13380 -871 13440 -668
rect 15782 -871 15842 -668
rect 15974 -871 16034 -591
rect 16092 -871 16152 -312
rect 16801 -354 16861 62
rect 16919 36 16979 62
rect 17156 36 17216 62
rect 17274 36 17334 62
rect 17282 -87 17348 -84
rect 17392 -87 17452 62
rect 17282 -100 17452 -87
rect 17282 -134 17298 -100
rect 17332 -134 17452 -100
rect 17282 -147 17452 -134
rect 17282 -150 17348 -147
rect 16323 -371 16861 -354
rect 16323 -405 16342 -371
rect 16376 -405 16861 -371
rect 16323 -411 16861 -405
rect 16323 -421 16392 -411
rect 16323 -423 16388 -421
rect 16207 -761 16273 -745
rect 16207 -795 16223 -761
rect 16257 -795 16273 -761
rect 16207 -811 16273 -795
rect 16210 -871 16270 -811
rect 16328 -871 16388 -423
rect 17392 -623 17452 -147
rect 16524 -668 17452 -623
rect 18080 -220 18140 66
rect 18198 40 18258 66
rect 18316 40 18376 66
rect 18521 40 18581 66
rect 18080 -237 18216 -220
rect 18080 -292 18139 -237
rect 18197 -292 18216 -237
rect 18080 -307 18216 -292
rect 18080 -619 18140 -307
rect 18639 -352 18699 66
rect 18757 40 18817 66
rect 18988 40 19048 66
rect 19106 40 19166 66
rect 19224 40 19284 66
rect 19342 40 19402 66
rect 19107 -120 19166 40
rect 19107 -121 19170 -120
rect 19104 -137 19170 -121
rect 19104 -171 19120 -137
rect 19154 -171 19170 -137
rect 19104 -187 19170 -171
rect 19207 -236 19302 -221
rect 19207 -291 19226 -236
rect 19284 -259 19302 -236
rect 19460 -259 19520 66
rect 19578 40 19638 66
rect 19815 40 19875 66
rect 19284 -291 19520 -259
rect 19207 -308 19520 -291
rect 18639 -409 19166 -352
rect 19106 -508 19166 -409
rect 19095 -521 19176 -508
rect 19095 -576 19108 -521
rect 19166 -576 19176 -521
rect 19095 -587 19176 -576
rect 18080 -664 18974 -619
rect 16524 -871 16584 -668
rect 18914 -867 18974 -664
rect 19106 -867 19166 -587
rect 19224 -867 19284 -308
rect 19933 -350 19993 66
rect 20051 40 20111 66
rect 20288 40 20348 66
rect 20406 40 20466 66
rect 20414 -83 20480 -80
rect 20524 -83 20584 66
rect 20414 -96 20584 -83
rect 20414 -130 20430 -96
rect 20464 -130 20584 -96
rect 20414 -143 20584 -130
rect 20414 -146 20480 -143
rect 19455 -367 19993 -350
rect 19455 -401 19474 -367
rect 19508 -401 19993 -367
rect 19455 -407 19993 -401
rect 19455 -417 19524 -407
rect 19455 -419 19520 -417
rect 19339 -757 19405 -741
rect 19339 -791 19355 -757
rect 19389 -791 19405 -757
rect 19339 -807 19405 -791
rect 19342 -867 19402 -807
rect 19460 -867 19520 -419
rect 20524 -619 20584 -143
rect 19656 -664 20584 -619
rect 21224 -220 21284 66
rect 21342 40 21402 66
rect 21460 40 21520 66
rect 21665 40 21725 66
rect 21224 -237 21360 -220
rect 21224 -292 21283 -237
rect 21341 -292 21360 -237
rect 21224 -307 21360 -292
rect 21224 -619 21284 -307
rect 21783 -352 21843 66
rect 21901 40 21961 66
rect 22132 40 22192 66
rect 22250 40 22310 66
rect 22368 40 22428 66
rect 22486 40 22546 66
rect 22251 -120 22310 40
rect 22251 -121 22314 -120
rect 22248 -137 22314 -121
rect 22248 -171 22264 -137
rect 22298 -171 22314 -137
rect 22248 -187 22314 -171
rect 22351 -236 22446 -221
rect 22351 -291 22370 -236
rect 22428 -259 22446 -236
rect 22604 -259 22664 66
rect 22722 40 22782 66
rect 22959 40 23019 66
rect 22428 -291 22664 -259
rect 22351 -308 22664 -291
rect 21783 -409 22310 -352
rect 22250 -508 22310 -409
rect 22239 -521 22320 -508
rect 22239 -576 22252 -521
rect 22310 -576 22320 -521
rect 22239 -587 22320 -576
rect 21224 -664 22118 -619
rect 19656 -867 19716 -664
rect 22058 -867 22118 -664
rect 22250 -867 22310 -587
rect 22368 -867 22428 -308
rect 23077 -350 23137 66
rect 23195 40 23255 66
rect 23432 40 23492 66
rect 23550 40 23610 66
rect 23558 -83 23624 -80
rect 23668 -83 23728 66
rect 23558 -96 23728 -83
rect 23558 -130 23574 -96
rect 23608 -130 23728 -96
rect 23558 -143 23728 -130
rect 23558 -146 23624 -143
rect 22599 -367 23137 -350
rect 22599 -401 22618 -367
rect 22652 -401 23137 -367
rect 22599 -407 23137 -401
rect 22599 -417 22668 -407
rect 22599 -419 22664 -417
rect 22483 -757 22549 -741
rect 22483 -791 22499 -757
rect 22533 -791 22549 -757
rect 22483 -807 22549 -791
rect 22486 -867 22546 -807
rect 22604 -867 22664 -419
rect 23668 -619 23728 -143
rect 22800 -664 23728 -619
rect 22800 -867 22860 -664
rect 9628 -1293 9688 -1267
rect 9746 -1293 9806 -1267
rect 9864 -1293 9924 -1267
rect 9982 -1293 10042 -1267
rect 6659 -1356 7094 -1348
rect 6659 -1390 6675 -1356
rect 6709 -1390 7094 -1356
rect 6659 -1399 7094 -1390
rect 9803 -1348 9869 -1340
rect 10178 -1348 10238 -1067
rect 12638 -1097 12698 -1071
rect 12830 -1297 12890 -1271
rect 12948 -1297 13008 -1271
rect 13066 -1297 13126 -1271
rect 13184 -1297 13244 -1271
rect 9803 -1356 10238 -1348
rect 9803 -1390 9819 -1356
rect 9853 -1390 10238 -1356
rect 9803 -1399 10238 -1390
rect 13005 -1352 13071 -1344
rect 13380 -1352 13440 -1071
rect 15782 -1097 15842 -1071
rect 15974 -1297 16034 -1271
rect 16092 -1297 16152 -1271
rect 16210 -1297 16270 -1271
rect 16328 -1297 16388 -1271
rect 13005 -1360 13440 -1352
rect 13005 -1394 13021 -1360
rect 13055 -1394 13440 -1360
rect 383 -1410 449 -1403
rect 3527 -1410 3593 -1403
rect 6659 -1406 6725 -1399
rect 9803 -1406 9869 -1399
rect 13005 -1403 13440 -1394
rect 16149 -1352 16215 -1344
rect 16524 -1352 16584 -1071
rect 18914 -1093 18974 -1067
rect 19106 -1293 19166 -1267
rect 19224 -1293 19284 -1267
rect 19342 -1293 19402 -1267
rect 19460 -1293 19520 -1267
rect 16149 -1360 16584 -1352
rect 16149 -1394 16165 -1360
rect 16199 -1394 16584 -1360
rect 16149 -1403 16584 -1394
rect 19281 -1348 19347 -1340
rect 19656 -1348 19716 -1067
rect 22058 -1093 22118 -1067
rect 22250 -1293 22310 -1267
rect 22368 -1293 22428 -1267
rect 22486 -1293 22546 -1267
rect 22604 -1293 22664 -1267
rect 19281 -1356 19716 -1348
rect 19281 -1390 19297 -1356
rect 19331 -1390 19716 -1356
rect 19281 -1399 19716 -1390
rect 22425 -1348 22491 -1340
rect 22800 -1348 22860 -1067
rect 22425 -1356 22860 -1348
rect 22425 -1390 22441 -1356
rect 22475 -1390 22860 -1356
rect 22425 -1399 22860 -1390
rect 13005 -1410 13071 -1403
rect 16149 -1410 16215 -1403
rect 19281 -1406 19347 -1399
rect 22425 -1406 22491 -1399
<< polycont >>
rect -759 -296 -701 -241
rect 222 -175 256 -141
rect 328 -295 386 -240
rect 210 -580 268 -525
rect 1532 -134 1566 -100
rect 576 -405 610 -371
rect 457 -795 491 -761
rect 2385 -296 2443 -241
rect 3366 -175 3400 -141
rect 3472 -295 3530 -240
rect 3354 -580 3412 -525
rect 4676 -134 4710 -100
rect 3720 -405 3754 -371
rect 3601 -795 3635 -761
rect 5517 -292 5575 -237
rect 6498 -171 6532 -137
rect 6604 -291 6662 -236
rect 6486 -576 6544 -521
rect 7808 -130 7842 -96
rect 6852 -401 6886 -367
rect 6733 -791 6767 -757
rect 8661 -292 8719 -237
rect 9642 -171 9676 -137
rect 9748 -291 9806 -236
rect 9630 -576 9688 -521
rect 10952 -130 10986 -96
rect 9996 -401 10030 -367
rect 9877 -791 9911 -757
rect 11863 -296 11921 -241
rect 12844 -175 12878 -141
rect 12950 -295 13008 -240
rect 12832 -580 12890 -525
rect 399 -1394 433 -1360
rect 3543 -1394 3577 -1360
rect 14154 -134 14188 -100
rect 13198 -405 13232 -371
rect 13079 -795 13113 -761
rect 15007 -296 15065 -241
rect 15988 -175 16022 -141
rect 16094 -295 16152 -240
rect 15976 -580 16034 -525
rect 17298 -134 17332 -100
rect 16342 -405 16376 -371
rect 16223 -795 16257 -761
rect 18139 -292 18197 -237
rect 19120 -171 19154 -137
rect 19226 -291 19284 -236
rect 19108 -576 19166 -521
rect 20430 -130 20464 -96
rect 19474 -401 19508 -367
rect 19355 -791 19389 -757
rect 21283 -292 21341 -237
rect 22264 -171 22298 -137
rect 22370 -291 22428 -236
rect 22252 -576 22310 -521
rect 23574 -130 23608 -96
rect 22618 -401 22652 -367
rect 22499 -791 22533 -757
rect 6675 -1390 6709 -1356
rect 9819 -1390 9853 -1356
rect 13021 -1394 13055 -1360
rect 16165 -1394 16199 -1360
rect 19297 -1390 19331 -1356
rect 22441 -1390 22475 -1356
<< locali >>
rect 306 720 534 738
rect 306 644 322 720
rect 518 644 534 720
rect 306 628 534 644
rect 3450 720 3678 738
rect 3450 644 3466 720
rect 3662 644 3678 720
rect 3450 628 3678 644
rect 6582 724 6810 742
rect 6582 648 6598 724
rect 6794 648 6810 724
rect 6582 632 6810 648
rect 9726 724 9954 742
rect 9726 648 9742 724
rect 9938 648 9954 724
rect 9726 632 9954 648
rect 12928 720 13156 738
rect 12928 644 12944 720
rect 13140 644 13156 720
rect 12928 628 13156 644
rect 16072 720 16300 738
rect 16072 644 16088 720
rect 16284 644 16300 720
rect 16072 628 16300 644
rect 19204 724 19432 742
rect 19204 648 19220 724
rect 19416 648 19432 724
rect 19204 632 19432 648
rect 22348 724 22576 742
rect 22348 648 22364 724
rect 22560 648 22576 724
rect 22348 632 22576 648
rect -423 503 -153 542
rect -423 450 -389 503
rect -864 301 -594 340
rect -864 250 -830 301
rect -864 58 -830 74
rect -746 250 -712 266
rect -746 23 -712 74
rect -628 250 -594 301
rect -628 58 -594 74
rect -510 250 -476 266
rect -510 23 -476 74
rect -423 58 -389 74
rect -305 450 -271 466
rect -746 -16 -476 23
rect -305 23 -271 74
rect -187 450 -153 503
rect 44 502 314 541
rect -187 58 -153 74
rect -69 450 -35 466
rect -69 23 -35 74
rect 44 450 78 502
rect 44 58 78 74
rect 162 450 196 466
rect 162 23 196 74
rect 280 450 314 502
rect 516 502 786 541
rect 280 58 314 74
rect 398 450 432 466
rect 398 23 432 74
rect 516 450 550 502
rect 516 58 550 74
rect 634 450 668 466
rect 634 23 668 74
rect 752 450 786 502
rect 989 502 1259 541
rect 752 58 786 74
rect 871 450 905 466
rect 871 23 905 74
rect 989 450 1023 502
rect 989 58 1023 74
rect 1107 450 1141 466
rect 1107 23 1141 74
rect 1225 450 1259 502
rect 2721 503 2991 542
rect 2721 450 2755 503
rect 1462 300 1732 337
rect 1225 58 1259 74
rect 1344 250 1378 266
rect -305 -16 1141 23
rect 1344 20 1378 74
rect 1462 250 1496 300
rect 1462 58 1496 74
rect 1580 250 1614 266
rect 1580 20 1614 74
rect 1698 250 1732 300
rect 1698 58 1732 74
rect 2280 301 2550 340
rect 2280 250 2314 301
rect 2280 58 2314 74
rect 2398 250 2432 266
rect 1344 -19 1614 20
rect 2398 23 2432 74
rect 2516 250 2550 301
rect 2516 58 2550 74
rect 2634 250 2668 266
rect 2634 23 2668 74
rect 2721 58 2755 74
rect 2839 450 2873 466
rect 2398 -16 2668 23
rect 2839 23 2873 74
rect 2957 450 2991 503
rect 3188 502 3458 541
rect 2957 58 2991 74
rect 3075 450 3109 466
rect 3075 23 3109 74
rect 3188 450 3222 502
rect 3188 58 3222 74
rect 3306 450 3340 466
rect 3306 23 3340 74
rect 3424 450 3458 502
rect 3660 502 3930 541
rect 3424 58 3458 74
rect 3542 450 3576 466
rect 3542 23 3576 74
rect 3660 450 3694 502
rect 3660 58 3694 74
rect 3778 450 3812 466
rect 3778 23 3812 74
rect 3896 450 3930 502
rect 4133 502 4403 541
rect 3896 58 3930 74
rect 4015 450 4049 466
rect 4015 23 4049 74
rect 4133 450 4167 502
rect 4133 58 4167 74
rect 4251 450 4285 466
rect 4251 23 4285 74
rect 4369 450 4403 502
rect 5853 507 6123 546
rect 5853 454 5887 507
rect 4606 300 4876 337
rect 4369 58 4403 74
rect 4488 250 4522 266
rect 2839 -16 4285 23
rect 4488 20 4522 74
rect 4606 250 4640 300
rect 4606 58 4640 74
rect 4724 250 4758 266
rect 4724 20 4758 74
rect 4842 250 4876 300
rect 4842 58 4876 74
rect 5412 305 5682 344
rect 5412 254 5446 305
rect 5412 62 5446 78
rect 5530 254 5564 270
rect 4488 -19 4758 20
rect 5530 27 5564 78
rect 5648 254 5682 305
rect 5648 62 5682 78
rect 5766 254 5800 270
rect 5766 27 5800 78
rect 5853 62 5887 78
rect 5971 454 6005 470
rect 5530 -12 5800 27
rect 5971 27 6005 78
rect 6089 454 6123 507
rect 6320 506 6590 545
rect 6089 62 6123 78
rect 6207 454 6241 470
rect 6207 27 6241 78
rect 6320 454 6354 506
rect 6320 62 6354 78
rect 6438 454 6472 470
rect 6438 27 6472 78
rect 6556 454 6590 506
rect 6792 506 7062 545
rect 6556 62 6590 78
rect 6674 454 6708 470
rect 6674 27 6708 78
rect 6792 454 6826 506
rect 6792 62 6826 78
rect 6910 454 6944 470
rect 6910 27 6944 78
rect 7028 454 7062 506
rect 7265 506 7535 545
rect 7028 62 7062 78
rect 7147 454 7181 470
rect 7147 27 7181 78
rect 7265 454 7299 506
rect 7265 62 7299 78
rect 7383 454 7417 470
rect 7383 27 7417 78
rect 7501 454 7535 506
rect 8997 507 9267 546
rect 8997 454 9031 507
rect 7738 304 8008 341
rect 7501 62 7535 78
rect 7620 254 7654 270
rect 5971 -12 7417 27
rect 7620 24 7654 78
rect 7738 254 7772 304
rect 7738 62 7772 78
rect 7856 254 7890 270
rect 7856 24 7890 78
rect 7974 254 8008 304
rect 7974 62 8008 78
rect 8556 305 8826 344
rect 8556 254 8590 305
rect 8556 62 8590 78
rect 8674 254 8708 270
rect 7620 -15 7890 24
rect 8674 27 8708 78
rect 8792 254 8826 305
rect 8792 62 8826 78
rect 8910 254 8944 270
rect 8910 27 8944 78
rect 8997 62 9031 78
rect 9115 454 9149 470
rect 8674 -12 8944 27
rect 9115 27 9149 78
rect 9233 454 9267 507
rect 9464 506 9734 545
rect 9233 62 9267 78
rect 9351 454 9385 470
rect 9351 27 9385 78
rect 9464 454 9498 506
rect 9464 62 9498 78
rect 9582 454 9616 470
rect 9582 27 9616 78
rect 9700 454 9734 506
rect 9936 506 10206 545
rect 9700 62 9734 78
rect 9818 454 9852 470
rect 9818 27 9852 78
rect 9936 454 9970 506
rect 9936 62 9970 78
rect 10054 454 10088 470
rect 10054 27 10088 78
rect 10172 454 10206 506
rect 10409 506 10679 545
rect 10172 62 10206 78
rect 10291 454 10325 470
rect 10291 27 10325 78
rect 10409 454 10443 506
rect 10409 62 10443 78
rect 10527 454 10561 470
rect 10527 27 10561 78
rect 10645 454 10679 506
rect 12199 503 12469 542
rect 12199 450 12233 503
rect 10882 304 11152 341
rect 10645 62 10679 78
rect 10764 254 10798 270
rect 9115 -12 10561 27
rect 10764 24 10798 78
rect 10882 254 10916 304
rect 10882 62 10916 78
rect 11000 254 11034 270
rect 11000 24 11034 78
rect 11118 254 11152 304
rect 11118 62 11152 78
rect 11758 301 12028 340
rect 11758 250 11792 301
rect 11758 58 11792 74
rect 11876 250 11910 266
rect 10764 -15 11034 24
rect 11876 23 11910 74
rect 11994 250 12028 301
rect 11994 58 12028 74
rect 12112 250 12146 266
rect 12112 23 12146 74
rect 12199 58 12233 74
rect 12317 450 12351 466
rect 11876 -16 12146 23
rect 12317 23 12351 74
rect 12435 450 12469 503
rect 12666 502 12936 541
rect 12435 58 12469 74
rect 12553 450 12587 466
rect 12553 23 12587 74
rect 12666 450 12700 502
rect 12666 58 12700 74
rect 12784 450 12818 466
rect 12784 23 12818 74
rect 12902 450 12936 502
rect 13138 502 13408 541
rect 12902 58 12936 74
rect 13020 450 13054 466
rect 13020 23 13054 74
rect 13138 450 13172 502
rect 13138 58 13172 74
rect 13256 450 13290 466
rect 13256 23 13290 74
rect 13374 450 13408 502
rect 13611 502 13881 541
rect 13374 58 13408 74
rect 13493 450 13527 466
rect 13493 23 13527 74
rect 13611 450 13645 502
rect 13611 58 13645 74
rect 13729 450 13763 466
rect 13729 23 13763 74
rect 13847 450 13881 502
rect 15343 503 15613 542
rect 15343 450 15377 503
rect 14084 300 14354 337
rect 13847 58 13881 74
rect 13966 250 14000 266
rect 12317 -16 13763 23
rect 13966 20 14000 74
rect 14084 250 14118 300
rect 14084 58 14118 74
rect 14202 250 14236 266
rect 14202 20 14236 74
rect 14320 250 14354 300
rect 14320 58 14354 74
rect 14902 301 15172 340
rect 14902 250 14936 301
rect 14902 58 14936 74
rect 15020 250 15054 266
rect 13966 -19 14236 20
rect 15020 23 15054 74
rect 15138 250 15172 301
rect 15138 58 15172 74
rect 15256 250 15290 266
rect 15256 23 15290 74
rect 15343 58 15377 74
rect 15461 450 15495 466
rect 15020 -16 15290 23
rect 15461 23 15495 74
rect 15579 450 15613 503
rect 15810 502 16080 541
rect 15579 58 15613 74
rect 15697 450 15731 466
rect 15697 23 15731 74
rect 15810 450 15844 502
rect 15810 58 15844 74
rect 15928 450 15962 466
rect 15928 23 15962 74
rect 16046 450 16080 502
rect 16282 502 16552 541
rect 16046 58 16080 74
rect 16164 450 16198 466
rect 16164 23 16198 74
rect 16282 450 16316 502
rect 16282 58 16316 74
rect 16400 450 16434 466
rect 16400 23 16434 74
rect 16518 450 16552 502
rect 16755 502 17025 541
rect 16518 58 16552 74
rect 16637 450 16671 466
rect 16637 23 16671 74
rect 16755 450 16789 502
rect 16755 58 16789 74
rect 16873 450 16907 466
rect 16873 23 16907 74
rect 16991 450 17025 502
rect 18475 507 18745 546
rect 18475 454 18509 507
rect 17228 300 17498 337
rect 16991 58 17025 74
rect 17110 250 17144 266
rect 15461 -16 16907 23
rect 17110 20 17144 74
rect 17228 250 17262 300
rect 17228 58 17262 74
rect 17346 250 17380 266
rect 17346 20 17380 74
rect 17464 250 17498 300
rect 17464 58 17498 74
rect 18034 305 18304 344
rect 18034 254 18068 305
rect 18034 62 18068 78
rect 18152 254 18186 270
rect 17110 -19 17380 20
rect 18152 27 18186 78
rect 18270 254 18304 305
rect 18270 62 18304 78
rect 18388 254 18422 270
rect 18388 27 18422 78
rect 18475 62 18509 78
rect 18593 454 18627 470
rect 18152 -12 18422 27
rect 18593 27 18627 78
rect 18711 454 18745 507
rect 18942 506 19212 545
rect 18711 62 18745 78
rect 18829 454 18863 470
rect 18829 27 18863 78
rect 18942 454 18976 506
rect 18942 62 18976 78
rect 19060 454 19094 470
rect 19060 27 19094 78
rect 19178 454 19212 506
rect 19414 506 19684 545
rect 19178 62 19212 78
rect 19296 454 19330 470
rect 19296 27 19330 78
rect 19414 454 19448 506
rect 19414 62 19448 78
rect 19532 454 19566 470
rect 19532 27 19566 78
rect 19650 454 19684 506
rect 19887 506 20157 545
rect 19650 62 19684 78
rect 19769 454 19803 470
rect 19769 27 19803 78
rect 19887 454 19921 506
rect 19887 62 19921 78
rect 20005 454 20039 470
rect 20005 27 20039 78
rect 20123 454 20157 506
rect 21619 507 21889 546
rect 21619 454 21653 507
rect 20360 304 20630 341
rect 20123 62 20157 78
rect 20242 254 20276 270
rect 18593 -12 20039 27
rect 20242 24 20276 78
rect 20360 254 20394 304
rect 20360 62 20394 78
rect 20478 254 20512 270
rect 20478 24 20512 78
rect 20596 254 20630 304
rect 20596 62 20630 78
rect 21178 305 21448 344
rect 21178 254 21212 305
rect 21178 62 21212 78
rect 21296 254 21330 270
rect 20242 -15 20512 24
rect 21296 27 21330 78
rect 21414 254 21448 305
rect 21414 62 21448 78
rect 21532 254 21566 270
rect 21532 27 21566 78
rect 21619 62 21653 78
rect 21737 454 21771 470
rect 21296 -12 21566 27
rect 21737 27 21771 78
rect 21855 454 21889 507
rect 22086 506 22356 545
rect 21855 62 21889 78
rect 21973 454 22007 470
rect 21973 27 22007 78
rect 22086 454 22120 506
rect 22086 62 22120 78
rect 22204 454 22238 470
rect 22204 27 22238 78
rect 22322 454 22356 506
rect 22558 506 22828 545
rect 22322 62 22356 78
rect 22440 454 22474 470
rect 22440 27 22474 78
rect 22558 454 22592 506
rect 22558 62 22592 78
rect 22676 454 22710 470
rect 22676 27 22710 78
rect 22794 454 22828 506
rect 23031 506 23301 545
rect 22794 62 22828 78
rect 22913 454 22947 470
rect 22913 27 22947 78
rect 23031 454 23065 506
rect 23031 62 23065 78
rect 23149 454 23183 470
rect 23149 27 23183 78
rect 23267 454 23301 506
rect 23504 304 23774 341
rect 23267 62 23301 78
rect 23386 254 23420 270
rect 21737 -12 23183 27
rect 23386 24 23420 78
rect 23504 254 23538 304
rect 23504 62 23538 78
rect 23622 254 23656 270
rect 23622 24 23656 78
rect 23740 254 23774 304
rect 23740 62 23774 78
rect 23386 -15 23656 24
rect 222 -141 256 -125
rect 1516 -134 1532 -100
rect 1566 -134 1582 -100
rect 222 -191 256 -175
rect 3366 -141 3400 -125
rect 4660 -134 4676 -100
rect 4710 -134 4726 -100
rect 3366 -191 3400 -175
rect 6498 -137 6532 -121
rect 7792 -130 7808 -96
rect 7842 -130 7858 -96
rect 6498 -187 6532 -171
rect 9642 -137 9676 -121
rect 10936 -130 10952 -96
rect 10986 -130 11002 -96
rect 9642 -187 9676 -171
rect 12844 -141 12878 -125
rect 14138 -134 14154 -100
rect 14188 -134 14204 -100
rect 12844 -191 12878 -175
rect 15988 -141 16022 -125
rect 17282 -134 17298 -100
rect 17332 -134 17348 -100
rect 15988 -191 16022 -175
rect 19120 -137 19154 -121
rect 20414 -130 20430 -96
rect 20464 -130 20480 -96
rect 19120 -187 19154 -171
rect 22264 -137 22298 -121
rect 23558 -130 23574 -96
rect 23608 -130 23624 -96
rect 22264 -187 22298 -171
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -775 -241 -683 -224
rect -775 -296 -759 -241
rect -699 -296 -683 -241
rect -775 -309 -683 -296
rect 310 -240 402 -227
rect 310 -295 326 -240
rect 386 -295 402 -240
rect 310 -312 402 -295
rect 2369 -241 2461 -224
rect 2369 -296 2385 -241
rect 2445 -296 2461 -241
rect 2369 -309 2461 -296
rect 3454 -240 3546 -227
rect 3454 -295 3470 -240
rect 3530 -295 3546 -240
rect 3454 -312 3546 -295
rect 5501 -237 5593 -220
rect 5501 -292 5517 -237
rect 5577 -292 5593 -237
rect 5501 -305 5593 -292
rect 6586 -236 6678 -223
rect 6586 -291 6602 -236
rect 6662 -291 6678 -236
rect 6586 -308 6678 -291
rect 8645 -237 8737 -220
rect 8645 -292 8661 -237
rect 8721 -292 8737 -237
rect 8645 -305 8737 -292
rect 9730 -236 9822 -223
rect 9730 -291 9746 -236
rect 9806 -291 9822 -236
rect 9730 -308 9822 -291
rect 11847 -241 11939 -224
rect 11847 -296 11863 -241
rect 11923 -296 11939 -241
rect 11847 -309 11939 -296
rect 12932 -240 13024 -227
rect 12932 -295 12948 -240
rect 13008 -295 13024 -240
rect 12932 -312 13024 -295
rect 14991 -241 15083 -224
rect 14991 -296 15007 -241
rect 15067 -296 15083 -241
rect 14991 -309 15083 -296
rect 16076 -240 16168 -227
rect 16076 -295 16092 -240
rect 16152 -295 16168 -240
rect 16076 -312 16168 -295
rect 18123 -237 18215 -220
rect 18123 -292 18139 -237
rect 18199 -292 18215 -237
rect 18123 -305 18215 -292
rect 19208 -236 19300 -223
rect 19208 -291 19224 -236
rect 19284 -291 19300 -236
rect 19208 -308 19300 -291
rect 21267 -237 21359 -220
rect 21267 -292 21283 -237
rect 21343 -292 21359 -237
rect 21267 -305 21359 -292
rect 22352 -236 22444 -223
rect 22352 -291 22368 -236
rect 22428 -291 22444 -236
rect 22352 -308 22444 -291
rect 576 -371 610 -355
rect 576 -421 610 -405
rect 2137 -356 2194 -352
rect 2137 -416 2141 -356
rect 2190 -416 2194 -356
rect 2137 -420 2194 -416
rect 3720 -371 3754 -355
rect 3720 -421 3754 -405
rect 6852 -367 6886 -351
rect 6852 -417 6886 -401
rect 8287 -352 8482 -348
rect 8287 -412 8417 -352
rect 8466 -412 8482 -352
rect 8287 -420 8482 -412
rect 9996 -367 10030 -351
rect 14538 -352 14792 -351
rect 17891 -352 17948 -348
rect 9996 -417 10030 -401
rect 13198 -371 13232 -355
rect 8287 -423 8345 -420
rect 13198 -421 13232 -405
rect 14538 -356 14816 -352
rect 14538 -416 14763 -356
rect 14812 -416 14816 -356
rect 14538 -420 14816 -416
rect 16342 -371 16376 -355
rect 8114 -480 8345 -423
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect 192 -525 284 -512
rect 192 -580 208 -525
rect 268 -580 284 -525
rect 192 -597 284 -580
rect 2137 -524 2194 -520
rect 2137 -584 2141 -524
rect 2190 -584 2194 -524
rect 2137 -588 2194 -584
rect 3336 -525 4743 -512
rect 3336 -580 3352 -525
rect 3412 -580 4743 -525
rect 3336 -597 4743 -580
rect 5269 -520 5326 -516
rect 5269 -580 5273 -520
rect 5322 -580 5326 -520
rect 5269 -584 5326 -580
rect 6468 -521 6560 -508
rect 6468 -576 6484 -521
rect 6544 -576 6560 -521
rect 6468 -593 6560 -576
rect 4663 -654 4743 -597
rect 8114 -654 8191 -480
rect 8413 -520 8470 -516
rect 8413 -580 8417 -520
rect 8466 -580 8470 -520
rect 8413 -584 8470 -580
rect 9612 -521 10484 -508
rect 9612 -576 9628 -521
rect 9688 -576 10484 -521
rect 9612 -593 10484 -576
rect 11615 -524 11672 -520
rect 11615 -584 11619 -524
rect 11668 -584 11672 -524
rect 11615 -588 11672 -584
rect 12814 -525 12906 -512
rect 12814 -580 12830 -525
rect 12890 -580 12906 -525
rect 4663 -707 8191 -654
rect 10407 -648 10484 -593
rect 12814 -597 12906 -580
rect 14538 -648 14606 -420
rect 16342 -421 16376 -405
rect 17891 -412 17895 -352
rect 17944 -412 17948 -352
rect 17891 -416 17948 -412
rect 19474 -367 19508 -351
rect 19474 -417 19508 -401
rect 20841 -352 21092 -348
rect 20841 -412 21039 -352
rect 21088 -412 21092 -352
rect 20841 -416 21092 -412
rect 22618 -367 22652 -351
rect 14759 -524 14816 -520
rect 14759 -584 14763 -524
rect 14812 -584 14816 -524
rect 14759 -588 14816 -584
rect 15958 -525 16895 -512
rect 15958 -580 15974 -525
rect 16034 -580 16895 -525
rect 15958 -597 16895 -580
rect 17891 -520 17948 -516
rect 17891 -580 17895 -520
rect 17944 -580 17948 -520
rect 17891 -584 17948 -580
rect 19090 -521 19182 -508
rect 19090 -576 19106 -521
rect 19166 -576 19182 -521
rect 19090 -593 19182 -576
rect 10407 -710 14606 -648
rect 16820 -642 16895 -597
rect 20841 -642 20898 -416
rect 22618 -417 22652 -401
rect 22234 -521 22326 -508
rect 22234 -576 22250 -521
rect 22310 -576 22326 -521
rect 22234 -593 22326 -576
rect 16820 -707 20898 -642
rect 457 -761 491 -745
rect 457 -811 491 -795
rect 3601 -761 3635 -745
rect 3601 -811 3635 -795
rect 6733 -757 6767 -741
rect 6733 -807 6767 -791
rect 9877 -757 9911 -741
rect 9877 -807 9911 -791
rect 13079 -761 13113 -745
rect 13079 -811 13113 -795
rect 16223 -761 16257 -745
rect 16223 -811 16257 -795
rect 19355 -757 19389 -741
rect 19355 -807 19389 -791
rect 22499 -757 22533 -741
rect 22499 -807 22533 -791
rect -30 -883 4 -867
rect -30 -1075 4 -1059
rect 88 -871 122 -867
rect 162 -871 196 -867
rect 88 -883 196 -871
rect 122 -1059 162 -883
rect 88 -1071 162 -1059
rect 88 -1075 122 -1071
rect 162 -1275 196 -1259
rect 280 -883 314 -867
rect 280 -1275 314 -1259
rect 398 -883 432 -867
rect 398 -1275 432 -1259
rect 516 -883 550 -867
rect 516 -1275 550 -1259
rect 634 -871 668 -867
rect 712 -871 746 -867
rect 634 -883 746 -871
rect 668 -1059 712 -883
rect 668 -1071 746 -1059
rect 712 -1075 746 -1071
rect 830 -883 864 -867
rect 830 -1075 864 -1059
rect 3114 -883 3148 -867
rect 3114 -1075 3148 -1059
rect 3232 -871 3266 -867
rect 3306 -871 3340 -867
rect 3232 -883 3340 -871
rect 3266 -1059 3306 -883
rect 3232 -1071 3306 -1059
rect 3232 -1075 3266 -1071
rect 634 -1275 668 -1259
rect 3306 -1275 3340 -1259
rect 3424 -883 3458 -867
rect 3424 -1275 3458 -1259
rect 3542 -883 3576 -867
rect 3542 -1275 3576 -1259
rect 3660 -883 3694 -867
rect 3660 -1275 3694 -1259
rect 3778 -871 3812 -867
rect 3856 -871 3890 -867
rect 3778 -883 3890 -871
rect 3812 -1059 3856 -883
rect 3812 -1071 3890 -1059
rect 3856 -1075 3890 -1071
rect 3974 -883 4008 -867
rect 3974 -1075 4008 -1059
rect 6246 -879 6280 -863
rect 6246 -1071 6280 -1055
rect 6364 -867 6398 -863
rect 6438 -867 6472 -863
rect 6364 -879 6472 -867
rect 6398 -1055 6438 -879
rect 6364 -1067 6438 -1055
rect 6364 -1071 6398 -1067
rect 3778 -1275 3812 -1259
rect 6438 -1271 6472 -1255
rect 6556 -879 6590 -863
rect 6556 -1271 6590 -1255
rect 6674 -879 6708 -863
rect 6674 -1271 6708 -1255
rect 6792 -879 6826 -863
rect 6792 -1271 6826 -1255
rect 6910 -867 6944 -863
rect 6988 -867 7022 -863
rect 6910 -879 7022 -867
rect 6944 -1055 6988 -879
rect 6944 -1067 7022 -1055
rect 6988 -1071 7022 -1067
rect 7106 -879 7140 -863
rect 7106 -1071 7140 -1055
rect 9390 -879 9424 -863
rect 9390 -1071 9424 -1055
rect 9508 -867 9542 -863
rect 9582 -867 9616 -863
rect 9508 -879 9616 -867
rect 9542 -1055 9582 -879
rect 9508 -1067 9582 -1055
rect 9508 -1071 9542 -1067
rect 6910 -1271 6944 -1255
rect 9582 -1271 9616 -1255
rect 9700 -879 9734 -863
rect 9700 -1271 9734 -1255
rect 9818 -879 9852 -863
rect 9818 -1271 9852 -1255
rect 9936 -879 9970 -863
rect 9936 -1271 9970 -1255
rect 10054 -867 10088 -863
rect 10132 -867 10166 -863
rect 10054 -879 10166 -867
rect 10088 -1055 10132 -879
rect 10088 -1067 10166 -1055
rect 10132 -1071 10166 -1067
rect 10250 -879 10284 -863
rect 10250 -1071 10284 -1055
rect 12592 -883 12626 -867
rect 12592 -1075 12626 -1059
rect 12710 -871 12744 -867
rect 12784 -871 12818 -867
rect 12710 -883 12818 -871
rect 12744 -1059 12784 -883
rect 12710 -1071 12784 -1059
rect 12710 -1075 12744 -1071
rect 10054 -1271 10088 -1255
rect 12784 -1275 12818 -1259
rect 12902 -883 12936 -867
rect 12902 -1275 12936 -1259
rect 13020 -883 13054 -867
rect 13020 -1275 13054 -1259
rect 13138 -883 13172 -867
rect 13138 -1275 13172 -1259
rect 13256 -871 13290 -867
rect 13334 -871 13368 -867
rect 13256 -883 13368 -871
rect 13290 -1059 13334 -883
rect 13290 -1071 13368 -1059
rect 13334 -1075 13368 -1071
rect 13452 -883 13486 -867
rect 13452 -1075 13486 -1059
rect 15736 -883 15770 -867
rect 15736 -1075 15770 -1059
rect 15854 -871 15888 -867
rect 15928 -871 15962 -867
rect 15854 -883 15962 -871
rect 15888 -1059 15928 -883
rect 15854 -1071 15928 -1059
rect 15854 -1075 15888 -1071
rect 13256 -1275 13290 -1259
rect 15928 -1275 15962 -1259
rect 16046 -883 16080 -867
rect 16046 -1275 16080 -1259
rect 16164 -883 16198 -867
rect 16164 -1275 16198 -1259
rect 16282 -883 16316 -867
rect 16282 -1275 16316 -1259
rect 16400 -871 16434 -867
rect 16478 -871 16512 -867
rect 16400 -883 16512 -871
rect 16434 -1059 16478 -883
rect 16434 -1071 16512 -1059
rect 16478 -1075 16512 -1071
rect 16596 -883 16630 -867
rect 16596 -1075 16630 -1059
rect 18868 -879 18902 -863
rect 18868 -1071 18902 -1055
rect 18986 -867 19020 -863
rect 19060 -867 19094 -863
rect 18986 -879 19094 -867
rect 19020 -1055 19060 -879
rect 18986 -1067 19060 -1055
rect 18986 -1071 19020 -1067
rect 16400 -1275 16434 -1259
rect 19060 -1271 19094 -1255
rect 19178 -879 19212 -863
rect 19178 -1271 19212 -1255
rect 19296 -879 19330 -863
rect 19296 -1271 19330 -1255
rect 19414 -879 19448 -863
rect 19414 -1271 19448 -1255
rect 19532 -867 19566 -863
rect 19610 -867 19644 -863
rect 19532 -879 19644 -867
rect 19566 -1055 19610 -879
rect 19566 -1067 19644 -1055
rect 19610 -1071 19644 -1067
rect 19728 -879 19762 -863
rect 19728 -1071 19762 -1055
rect 22012 -879 22046 -863
rect 22012 -1071 22046 -1055
rect 22130 -867 22164 -863
rect 22204 -867 22238 -863
rect 22130 -879 22238 -867
rect 22164 -1055 22204 -879
rect 22130 -1067 22204 -1055
rect 22130 -1071 22164 -1067
rect 19532 -1271 19566 -1255
rect 22204 -1271 22238 -1255
rect 22322 -879 22356 -863
rect 22322 -1271 22356 -1255
rect 22440 -879 22474 -863
rect 22440 -1271 22474 -1255
rect 22558 -879 22592 -863
rect 22558 -1271 22592 -1255
rect 22676 -867 22710 -863
rect 22754 -867 22788 -863
rect 22676 -879 22788 -867
rect 22710 -1055 22754 -879
rect 22710 -1067 22788 -1055
rect 22754 -1071 22788 -1067
rect 22872 -879 22906 -863
rect 22872 -1071 22906 -1055
rect 22676 -1271 22710 -1255
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 3527 -1394 3543 -1360
rect 3577 -1394 3593 -1360
rect 6659 -1390 6675 -1356
rect 6709 -1390 6725 -1356
rect 9803 -1390 9819 -1356
rect 9853 -1390 9869 -1356
rect 13005 -1394 13021 -1360
rect 13055 -1394 13071 -1360
rect 16149 -1394 16165 -1360
rect 16199 -1394 16215 -1360
rect 19281 -1390 19297 -1356
rect 19331 -1390 19347 -1356
rect 22425 -1390 22441 -1356
rect 22475 -1390 22491 -1356
rect 6640 -1508 6776 -1504
rect 364 -1512 500 -1508
rect 364 -1526 402 -1512
rect 460 -1526 500 -1512
rect 364 -1572 380 -1526
rect 484 -1572 500 -1526
rect 364 -1594 500 -1572
rect 3508 -1512 3644 -1508
rect 3508 -1526 3546 -1512
rect 3604 -1526 3644 -1512
rect 3508 -1572 3524 -1526
rect 3628 -1572 3644 -1526
rect 3508 -1594 3644 -1572
rect 6640 -1522 6678 -1508
rect 6736 -1522 6776 -1508
rect 6640 -1568 6656 -1522
rect 6760 -1568 6776 -1522
rect 6640 -1590 6776 -1568
rect 9784 -1508 9920 -1504
rect 19262 -1508 19398 -1504
rect 9784 -1522 9822 -1508
rect 9880 -1522 9920 -1508
rect 9784 -1568 9800 -1522
rect 9904 -1568 9920 -1522
rect 9784 -1590 9920 -1568
rect 12986 -1512 13122 -1508
rect 12986 -1526 13024 -1512
rect 13082 -1526 13122 -1512
rect 12986 -1572 13002 -1526
rect 13106 -1572 13122 -1526
rect 12986 -1594 13122 -1572
rect 16130 -1512 16266 -1508
rect 16130 -1526 16168 -1512
rect 16226 -1526 16266 -1512
rect 16130 -1572 16146 -1526
rect 16250 -1572 16266 -1526
rect 16130 -1594 16266 -1572
rect 19262 -1522 19300 -1508
rect 19358 -1522 19398 -1508
rect 19262 -1568 19278 -1522
rect 19382 -1568 19398 -1522
rect 19262 -1590 19398 -1568
rect 22406 -1508 22542 -1504
rect 22406 -1522 22444 -1508
rect 22502 -1522 22542 -1508
rect 22406 -1568 22422 -1522
rect 22526 -1568 22542 -1522
rect 22406 -1590 22542 -1568
<< viali >>
rect 388 646 460 700
rect 3532 646 3604 700
rect 6664 650 6736 704
rect 9808 650 9880 704
rect 13010 646 13082 700
rect 16154 646 16226 700
rect 19286 650 19358 704
rect 22430 650 22502 704
rect -864 74 -830 250
rect -746 74 -712 250
rect -628 74 -594 250
rect -510 74 -476 250
rect -423 74 -389 450
rect -305 74 -271 450
rect -187 74 -153 450
rect -69 74 -35 450
rect 44 74 78 450
rect 162 74 196 450
rect 280 74 314 450
rect 398 74 432 450
rect 516 74 550 450
rect 634 74 668 450
rect 752 74 786 450
rect 871 74 905 450
rect 989 74 1023 450
rect 1107 74 1141 450
rect 1225 74 1259 450
rect 1344 74 1378 250
rect 1462 74 1496 250
rect 1580 74 1614 250
rect 1698 74 1732 250
rect 2280 74 2314 250
rect 2398 74 2432 250
rect 2516 74 2550 250
rect 2634 74 2668 250
rect 2721 74 2755 450
rect 2839 74 2873 450
rect 2957 74 2991 450
rect 3075 74 3109 450
rect 3188 74 3222 450
rect 3306 74 3340 450
rect 3424 74 3458 450
rect 3542 74 3576 450
rect 3660 74 3694 450
rect 3778 74 3812 450
rect 3896 74 3930 450
rect 4015 74 4049 450
rect 4133 74 4167 450
rect 4251 74 4285 450
rect 4369 74 4403 450
rect 4488 74 4522 250
rect 4606 74 4640 250
rect 4724 74 4758 250
rect 4842 74 4876 250
rect 5412 78 5446 254
rect 5530 78 5564 254
rect 5648 78 5682 254
rect 5766 78 5800 254
rect 5853 78 5887 454
rect 5971 78 6005 454
rect 6089 78 6123 454
rect 6207 78 6241 454
rect 6320 78 6354 454
rect 6438 78 6472 454
rect 6556 78 6590 454
rect 6674 78 6708 454
rect 6792 78 6826 454
rect 6910 78 6944 454
rect 7028 78 7062 454
rect 7147 78 7181 454
rect 7265 78 7299 454
rect 7383 78 7417 454
rect 7501 78 7535 454
rect 7620 78 7654 254
rect 7738 78 7772 254
rect 7856 78 7890 254
rect 7974 78 8008 254
rect 8556 78 8590 254
rect 8674 78 8708 254
rect 8792 78 8826 254
rect 8910 78 8944 254
rect 8997 78 9031 454
rect 9115 78 9149 454
rect 9233 78 9267 454
rect 9351 78 9385 454
rect 9464 78 9498 454
rect 9582 78 9616 454
rect 9700 78 9734 454
rect 9818 78 9852 454
rect 9936 78 9970 454
rect 10054 78 10088 454
rect 10172 78 10206 454
rect 10291 78 10325 454
rect 10409 78 10443 454
rect 10527 78 10561 454
rect 10645 78 10679 454
rect 10764 78 10798 254
rect 10882 78 10916 254
rect 11000 78 11034 254
rect 11118 78 11152 254
rect 11758 74 11792 250
rect 11876 74 11910 250
rect 11994 74 12028 250
rect 12112 74 12146 250
rect 12199 74 12233 450
rect 12317 74 12351 450
rect 12435 74 12469 450
rect 12553 74 12587 450
rect 12666 74 12700 450
rect 12784 74 12818 450
rect 12902 74 12936 450
rect 13020 74 13054 450
rect 13138 74 13172 450
rect 13256 74 13290 450
rect 13374 74 13408 450
rect 13493 74 13527 450
rect 13611 74 13645 450
rect 13729 74 13763 450
rect 13847 74 13881 450
rect 13966 74 14000 250
rect 14084 74 14118 250
rect 14202 74 14236 250
rect 14320 74 14354 250
rect 14902 74 14936 250
rect 15020 74 15054 250
rect 15138 74 15172 250
rect 15256 74 15290 250
rect 15343 74 15377 450
rect 15461 74 15495 450
rect 15579 74 15613 450
rect 15697 74 15731 450
rect 15810 74 15844 450
rect 15928 74 15962 450
rect 16046 74 16080 450
rect 16164 74 16198 450
rect 16282 74 16316 450
rect 16400 74 16434 450
rect 16518 74 16552 450
rect 16637 74 16671 450
rect 16755 74 16789 450
rect 16873 74 16907 450
rect 16991 74 17025 450
rect 17110 74 17144 250
rect 17228 74 17262 250
rect 17346 74 17380 250
rect 17464 74 17498 250
rect 18034 78 18068 254
rect 18152 78 18186 254
rect 18270 78 18304 254
rect 18388 78 18422 254
rect 18475 78 18509 454
rect 18593 78 18627 454
rect 18711 78 18745 454
rect 18829 78 18863 454
rect 18942 78 18976 454
rect 19060 78 19094 454
rect 19178 78 19212 454
rect 19296 78 19330 454
rect 19414 78 19448 454
rect 19532 78 19566 454
rect 19650 78 19684 454
rect 19769 78 19803 454
rect 19887 78 19921 454
rect 20005 78 20039 454
rect 20123 78 20157 454
rect 20242 78 20276 254
rect 20360 78 20394 254
rect 20478 78 20512 254
rect 20596 78 20630 254
rect 21178 78 21212 254
rect 21296 78 21330 254
rect 21414 78 21448 254
rect 21532 78 21566 254
rect 21619 78 21653 454
rect 21737 78 21771 454
rect 21855 78 21889 454
rect 21973 78 22007 454
rect 22086 78 22120 454
rect 22204 78 22238 454
rect 22322 78 22356 454
rect 22440 78 22474 454
rect 22558 78 22592 454
rect 22676 78 22710 454
rect 22794 78 22828 454
rect 22913 78 22947 454
rect 23031 78 23065 454
rect 23149 78 23183 454
rect 23267 78 23301 454
rect 23386 78 23420 254
rect 23504 78 23538 254
rect 23622 78 23656 254
rect 23740 78 23774 254
rect 1532 -134 1566 -100
rect 222 -175 256 -141
rect 4676 -134 4710 -100
rect 3366 -175 3400 -141
rect 7808 -130 7842 -96
rect 6498 -171 6532 -137
rect 10952 -130 10986 -96
rect 9642 -171 9676 -137
rect 14154 -134 14188 -100
rect 12844 -175 12878 -141
rect 17298 -134 17332 -100
rect 15988 -175 16022 -141
rect 20430 -130 20464 -96
rect 19120 -171 19154 -137
rect 23574 -130 23608 -96
rect 22264 -171 22298 -137
rect -1003 -300 -954 -240
rect -759 -296 -701 -241
rect -701 -296 -699 -241
rect 326 -295 328 -240
rect 328 -295 386 -240
rect 2385 -296 2443 -241
rect 2443 -296 2445 -241
rect 3470 -295 3472 -240
rect 3472 -295 3530 -240
rect 5517 -292 5575 -237
rect 5575 -292 5577 -237
rect 6602 -291 6604 -236
rect 6604 -291 6662 -236
rect 8661 -292 8719 -237
rect 8719 -292 8721 -237
rect 9746 -291 9748 -236
rect 9748 -291 9806 -236
rect 11863 -296 11921 -241
rect 11921 -296 11923 -241
rect 12948 -295 12950 -240
rect 12950 -295 13008 -240
rect 15007 -296 15065 -241
rect 15065 -296 15067 -241
rect 16092 -295 16094 -240
rect 16094 -295 16152 -240
rect 18139 -292 18197 -237
rect 18197 -292 18199 -237
rect 19224 -291 19226 -236
rect 19226 -291 19284 -236
rect 21283 -292 21341 -237
rect 21341 -292 21343 -237
rect 22368 -291 22370 -236
rect 22370 -291 22428 -236
rect 576 -405 610 -371
rect 2141 -416 2190 -356
rect 3720 -405 3754 -371
rect 6852 -401 6886 -367
rect 8417 -412 8466 -352
rect 9996 -401 10030 -367
rect 13198 -405 13232 -371
rect 14763 -416 14812 -356
rect 16342 -405 16376 -371
rect -1003 -584 -954 -524
rect 208 -580 210 -525
rect 210 -580 268 -525
rect 2141 -584 2190 -524
rect 3352 -580 3354 -525
rect 3354 -580 3412 -525
rect 5273 -580 5322 -520
rect 6484 -576 6486 -521
rect 6486 -576 6544 -521
rect 8417 -580 8466 -520
rect 9628 -576 9630 -521
rect 9630 -576 9688 -521
rect 11619 -584 11668 -524
rect 12830 -580 12832 -525
rect 12832 -580 12890 -525
rect 17895 -412 17944 -352
rect 19474 -401 19508 -367
rect 21039 -412 21088 -352
rect 22618 -401 22652 -367
rect 14763 -584 14812 -524
rect 15974 -580 15976 -525
rect 15976 -580 16034 -525
rect 17895 -580 17944 -520
rect 19106 -576 19108 -521
rect 19108 -576 19166 -521
rect 22250 -576 22252 -521
rect 22252 -576 22310 -521
rect 457 -795 491 -761
rect 3601 -795 3635 -761
rect 6733 -791 6767 -757
rect 9877 -791 9911 -757
rect 13079 -795 13113 -761
rect 16223 -795 16257 -761
rect 19355 -791 19389 -757
rect 22499 -791 22533 -757
rect -30 -1059 4 -883
rect 88 -1059 122 -883
rect 162 -1259 196 -883
rect 280 -1259 314 -883
rect 398 -1259 432 -883
rect 516 -1259 550 -883
rect 634 -1259 668 -883
rect 712 -1059 746 -883
rect 830 -1059 864 -883
rect 3114 -1059 3148 -883
rect 3232 -1059 3266 -883
rect 3306 -1259 3340 -883
rect 3424 -1259 3458 -883
rect 3542 -1259 3576 -883
rect 3660 -1259 3694 -883
rect 3778 -1259 3812 -883
rect 3856 -1059 3890 -883
rect 3974 -1059 4008 -883
rect 6246 -1055 6280 -879
rect 6364 -1055 6398 -879
rect 6438 -1255 6472 -879
rect 6556 -1255 6590 -879
rect 6674 -1255 6708 -879
rect 6792 -1255 6826 -879
rect 6910 -1255 6944 -879
rect 6988 -1055 7022 -879
rect 7106 -1055 7140 -879
rect 9390 -1055 9424 -879
rect 9508 -1055 9542 -879
rect 9582 -1255 9616 -879
rect 9700 -1255 9734 -879
rect 9818 -1255 9852 -879
rect 9936 -1255 9970 -879
rect 10054 -1255 10088 -879
rect 10132 -1055 10166 -879
rect 10250 -1055 10284 -879
rect 12592 -1059 12626 -883
rect 12710 -1059 12744 -883
rect 12784 -1259 12818 -883
rect 12902 -1259 12936 -883
rect 13020 -1259 13054 -883
rect 13138 -1259 13172 -883
rect 13256 -1259 13290 -883
rect 13334 -1059 13368 -883
rect 13452 -1059 13486 -883
rect 15736 -1059 15770 -883
rect 15854 -1059 15888 -883
rect 15928 -1259 15962 -883
rect 16046 -1259 16080 -883
rect 16164 -1259 16198 -883
rect 16282 -1259 16316 -883
rect 16400 -1259 16434 -883
rect 16478 -1059 16512 -883
rect 16596 -1059 16630 -883
rect 18868 -1055 18902 -879
rect 18986 -1055 19020 -879
rect 19060 -1255 19094 -879
rect 19178 -1255 19212 -879
rect 19296 -1255 19330 -879
rect 19414 -1255 19448 -879
rect 19532 -1255 19566 -879
rect 19610 -1055 19644 -879
rect 19728 -1055 19762 -879
rect 22012 -1055 22046 -879
rect 22130 -1055 22164 -879
rect 22204 -1255 22238 -879
rect 22322 -1255 22356 -879
rect 22440 -1255 22474 -879
rect 22558 -1255 22592 -879
rect 22676 -1255 22710 -879
rect 22754 -1055 22788 -879
rect 22872 -1055 22906 -879
rect 399 -1394 433 -1360
rect 3543 -1394 3577 -1360
rect 6675 -1390 6709 -1356
rect 9819 -1390 9853 -1356
rect 13021 -1394 13055 -1360
rect 16165 -1394 16199 -1360
rect 19297 -1390 19331 -1356
rect 22441 -1390 22475 -1356
rect 402 -1526 460 -1512
rect 402 -1558 460 -1526
rect 3546 -1526 3604 -1512
rect 3546 -1558 3604 -1526
rect 6678 -1522 6736 -1508
rect 6678 -1554 6736 -1522
rect 9822 -1522 9880 -1508
rect 9822 -1554 9880 -1522
rect 13024 -1526 13082 -1512
rect 13024 -1558 13082 -1526
rect 16168 -1526 16226 -1512
rect 16168 -1558 16226 -1526
rect 19300 -1522 19358 -1508
rect 19300 -1554 19358 -1522
rect 22444 -1522 22502 -1508
rect 22444 -1554 22502 -1522
<< metal1 >>
rect 374 646 384 706
rect 464 646 474 706
rect 374 606 474 646
rect 3518 646 3528 706
rect 3608 646 3618 706
rect 3518 606 3618 646
rect 6650 650 6660 710
rect 6740 650 6750 710
rect 6650 610 6750 650
rect 9794 650 9804 710
rect 9884 650 9894 710
rect 9794 610 9894 650
rect 12996 646 13006 706
rect 13086 646 13096 706
rect -423 549 1380 606
rect -423 462 -389 549
rect 752 462 786 549
rect -429 450 -383 462
rect -429 262 -423 450
rect -870 250 -824 262
rect -870 74 -864 250
rect -830 74 -824 250
rect -870 62 -824 74
rect -752 250 -706 262
rect -752 74 -746 250
rect -712 74 -706 250
rect -752 62 -706 74
rect -634 250 -588 262
rect -634 74 -628 250
rect -594 74 -588 250
rect -634 62 -588 74
rect -516 250 -423 262
rect -516 74 -510 250
rect -476 74 -423 250
rect -389 74 -383 450
rect -516 62 -383 74
rect -311 450 -265 462
rect -311 74 -305 450
rect -271 74 -265 450
rect -311 62 -265 74
rect -193 450 -147 462
rect -193 74 -187 450
rect -153 74 -147 450
rect -193 62 -147 74
rect -75 450 -29 462
rect -75 74 -69 450
rect -35 74 -29 450
rect -75 62 -29 74
rect 38 450 84 462
rect 38 74 44 450
rect 78 74 84 450
rect 38 62 84 74
rect 156 450 202 462
rect 156 74 162 450
rect 196 74 202 450
rect 156 62 202 74
rect 274 450 320 462
rect 274 74 280 450
rect 314 74 320 450
rect 274 62 320 74
rect 392 450 438 462
rect 392 74 398 450
rect 432 74 438 450
rect 392 62 438 74
rect 510 450 556 462
rect 510 74 516 450
rect 550 74 556 450
rect 510 62 556 74
rect 628 450 674 462
rect 628 74 634 450
rect 668 74 674 450
rect 628 62 674 74
rect 746 450 792 462
rect 746 74 752 450
rect 786 74 792 450
rect 746 62 792 74
rect 865 450 911 462
rect 865 74 871 450
rect 905 74 911 450
rect 865 62 911 74
rect 983 450 1029 462
rect 983 74 989 450
rect 1023 74 1029 450
rect 983 62 1029 74
rect 1101 450 1147 462
rect 1101 74 1107 450
rect 1141 74 1147 450
rect 1101 62 1147 74
rect 1219 450 1265 462
rect 1219 74 1225 450
rect 1259 74 1265 450
rect 1343 262 1380 549
rect 2721 549 4524 606
rect 2721 462 2755 549
rect 3896 462 3930 549
rect 2715 450 2761 462
rect 2715 262 2721 450
rect 1219 62 1265 74
rect 1338 250 1384 262
rect 1338 74 1344 250
rect 1378 74 1384 250
rect 1338 62 1384 74
rect 1456 250 1502 262
rect 1456 74 1462 250
rect 1496 74 1502 250
rect 1456 62 1502 74
rect 1574 250 1620 262
rect 1574 74 1580 250
rect 1614 74 1620 250
rect 1574 62 1620 74
rect 1692 250 1738 262
rect 1692 74 1698 250
rect 1732 74 1738 250
rect 1692 62 1738 74
rect 2274 250 2320 262
rect 2274 74 2280 250
rect 2314 74 2320 250
rect 2274 62 2320 74
rect 2392 250 2438 262
rect 2392 74 2398 250
rect 2432 74 2438 250
rect 2392 62 2438 74
rect 2510 250 2556 262
rect 2510 74 2516 250
rect 2550 74 2556 250
rect 2510 62 2556 74
rect 2628 250 2721 262
rect 2628 74 2634 250
rect 2668 74 2721 250
rect 2755 74 2761 450
rect 2628 62 2761 74
rect 2833 450 2879 462
rect 2833 74 2839 450
rect 2873 74 2879 450
rect 2833 62 2879 74
rect 2951 450 2997 462
rect 2951 74 2957 450
rect 2991 74 2997 450
rect 2951 62 2997 74
rect 3069 450 3115 462
rect 3069 74 3075 450
rect 3109 74 3115 450
rect 3069 62 3115 74
rect 3182 450 3228 462
rect 3182 74 3188 450
rect 3222 74 3228 450
rect 3182 62 3228 74
rect 3300 450 3346 462
rect 3300 74 3306 450
rect 3340 74 3346 450
rect 3300 62 3346 74
rect 3418 450 3464 462
rect 3418 74 3424 450
rect 3458 74 3464 450
rect 3418 62 3464 74
rect 3536 450 3582 462
rect 3536 74 3542 450
rect 3576 74 3582 450
rect 3536 62 3582 74
rect 3654 450 3700 462
rect 3654 74 3660 450
rect 3694 74 3700 450
rect 3654 62 3700 74
rect 3772 450 3818 462
rect 3772 74 3778 450
rect 3812 74 3818 450
rect 3772 62 3818 74
rect 3890 450 3936 462
rect 3890 74 3896 450
rect 3930 74 3936 450
rect 3890 62 3936 74
rect 4009 450 4055 462
rect 4009 74 4015 450
rect 4049 74 4055 450
rect 4009 62 4055 74
rect 4127 450 4173 462
rect 4127 74 4133 450
rect 4167 74 4173 450
rect 4127 62 4173 74
rect 4245 450 4291 462
rect 4245 74 4251 450
rect 4285 74 4291 450
rect 4245 62 4291 74
rect 4363 450 4409 462
rect 4363 74 4369 450
rect 4403 74 4409 450
rect 4487 262 4524 549
rect 5853 553 7656 610
rect 5853 466 5887 553
rect 7028 466 7062 553
rect 5847 454 5893 466
rect 5847 266 5853 454
rect 4363 62 4409 74
rect 4482 250 4528 262
rect 4482 74 4488 250
rect 4522 74 4528 250
rect 4482 62 4528 74
rect 4600 250 4646 262
rect 4600 74 4606 250
rect 4640 74 4646 250
rect 4600 62 4646 74
rect 4718 250 4764 262
rect 4718 74 4724 250
rect 4758 74 4764 250
rect 4718 62 4764 74
rect 4836 250 4882 262
rect 4836 74 4842 250
rect 4876 74 4882 250
rect 4836 62 4882 74
rect 5406 254 5452 266
rect 5406 78 5412 254
rect 5446 78 5452 254
rect 5406 66 5452 78
rect 5524 254 5570 266
rect 5524 78 5530 254
rect 5564 78 5570 254
rect 5524 66 5570 78
rect 5642 254 5688 266
rect 5642 78 5648 254
rect 5682 78 5688 254
rect 5642 66 5688 78
rect 5760 254 5853 266
rect 5760 78 5766 254
rect 5800 78 5853 254
rect 5887 78 5893 454
rect 5760 66 5893 78
rect 5965 454 6011 466
rect 5965 78 5971 454
rect 6005 78 6011 454
rect 5965 66 6011 78
rect 6083 454 6129 466
rect 6083 78 6089 454
rect 6123 78 6129 454
rect 6083 66 6129 78
rect 6201 454 6247 466
rect 6201 78 6207 454
rect 6241 78 6247 454
rect 6201 66 6247 78
rect 6314 454 6360 466
rect 6314 78 6320 454
rect 6354 78 6360 454
rect 6314 66 6360 78
rect 6432 454 6478 466
rect 6432 78 6438 454
rect 6472 78 6478 454
rect 6432 66 6478 78
rect 6550 454 6596 466
rect 6550 78 6556 454
rect 6590 78 6596 454
rect 6550 66 6596 78
rect 6668 454 6714 466
rect 6668 78 6674 454
rect 6708 78 6714 454
rect 6668 66 6714 78
rect 6786 454 6832 466
rect 6786 78 6792 454
rect 6826 78 6832 454
rect 6786 66 6832 78
rect 6904 454 6950 466
rect 6904 78 6910 454
rect 6944 78 6950 454
rect 6904 66 6950 78
rect 7022 454 7068 466
rect 7022 78 7028 454
rect 7062 78 7068 454
rect 7022 66 7068 78
rect 7141 454 7187 466
rect 7141 78 7147 454
rect 7181 78 7187 454
rect 7141 66 7187 78
rect 7259 454 7305 466
rect 7259 78 7265 454
rect 7299 78 7305 454
rect 7259 66 7305 78
rect 7377 454 7423 466
rect 7377 78 7383 454
rect 7417 78 7423 454
rect 7377 66 7423 78
rect 7495 454 7541 466
rect 7495 78 7501 454
rect 7535 78 7541 454
rect 7619 266 7656 553
rect 8997 553 10800 610
rect 12996 606 13096 646
rect 16140 646 16150 706
rect 16230 646 16240 706
rect 16140 606 16240 646
rect 19272 650 19282 710
rect 19362 650 19372 710
rect 19272 610 19372 650
rect 22416 650 22426 710
rect 22506 650 22516 710
rect 22416 610 22516 650
rect 8997 466 9031 553
rect 10172 466 10206 553
rect 8991 454 9037 466
rect 8991 266 8997 454
rect 7495 66 7541 78
rect 7614 254 7660 266
rect 7614 78 7620 254
rect 7654 78 7660 254
rect 7614 66 7660 78
rect 7732 254 7778 266
rect 7732 78 7738 254
rect 7772 78 7778 254
rect 7732 66 7778 78
rect 7850 254 7896 266
rect 7850 78 7856 254
rect 7890 78 7896 254
rect 7850 66 7896 78
rect 7968 254 8014 266
rect 7968 78 7974 254
rect 8008 78 8014 254
rect 7968 66 8014 78
rect 8550 254 8596 266
rect 8550 78 8556 254
rect 8590 78 8596 254
rect 8550 66 8596 78
rect 8668 254 8714 266
rect 8668 78 8674 254
rect 8708 78 8714 254
rect 8668 66 8714 78
rect 8786 254 8832 266
rect 8786 78 8792 254
rect 8826 78 8832 254
rect 8786 66 8832 78
rect 8904 254 8997 266
rect 8904 78 8910 254
rect 8944 78 8997 254
rect 9031 78 9037 454
rect 8904 66 9037 78
rect 9109 454 9155 466
rect 9109 78 9115 454
rect 9149 78 9155 454
rect 9109 66 9155 78
rect 9227 454 9273 466
rect 9227 78 9233 454
rect 9267 78 9273 454
rect 9227 66 9273 78
rect 9345 454 9391 466
rect 9345 78 9351 454
rect 9385 78 9391 454
rect 9345 66 9391 78
rect 9458 454 9504 466
rect 9458 78 9464 454
rect 9498 78 9504 454
rect 9458 66 9504 78
rect 9576 454 9622 466
rect 9576 78 9582 454
rect 9616 78 9622 454
rect 9576 66 9622 78
rect 9694 454 9740 466
rect 9694 78 9700 454
rect 9734 78 9740 454
rect 9694 66 9740 78
rect 9812 454 9858 466
rect 9812 78 9818 454
rect 9852 78 9858 454
rect 9812 66 9858 78
rect 9930 454 9976 466
rect 9930 78 9936 454
rect 9970 78 9976 454
rect 9930 66 9976 78
rect 10048 454 10094 466
rect 10048 78 10054 454
rect 10088 78 10094 454
rect 10048 66 10094 78
rect 10166 454 10212 466
rect 10166 78 10172 454
rect 10206 78 10212 454
rect 10166 66 10212 78
rect 10285 454 10331 466
rect 10285 78 10291 454
rect 10325 78 10331 454
rect 10285 66 10331 78
rect 10403 454 10449 466
rect 10403 78 10409 454
rect 10443 78 10449 454
rect 10403 66 10449 78
rect 10521 454 10567 466
rect 10521 78 10527 454
rect 10561 78 10567 454
rect 10521 66 10567 78
rect 10639 454 10685 466
rect 10639 78 10645 454
rect 10679 78 10685 454
rect 10763 266 10800 553
rect 12199 549 14002 606
rect 12199 462 12233 549
rect 13374 462 13408 549
rect 12193 450 12239 462
rect 10639 66 10685 78
rect 10758 254 10804 266
rect 10758 78 10764 254
rect 10798 78 10804 254
rect 10758 66 10804 78
rect 10876 254 10922 266
rect 10876 78 10882 254
rect 10916 78 10922 254
rect 10876 66 10922 78
rect 10994 254 11040 266
rect 10994 78 11000 254
rect 11034 78 11040 254
rect 10994 66 11040 78
rect 11112 254 11158 266
rect 12193 262 12199 450
rect 11112 78 11118 254
rect 11152 78 11158 254
rect 11112 66 11158 78
rect 11752 250 11798 262
rect 11752 74 11758 250
rect 11792 74 11798 250
rect -1269 -87 -942 -86
rect -1269 -149 -1006 -87
rect -952 -149 -942 -87
rect -865 -124 -830 62
rect 44 -22 78 62
rect 1225 -22 1259 62
rect 44 -64 1259 -22
rect 1225 -84 1259 -64
rect 1225 -100 1582 -84
rect -865 -141 272 -124
rect -865 -175 222 -141
rect 256 -175 272 -141
rect 1225 -134 1532 -100
rect 1566 -134 1582 -100
rect 1225 -150 1582 -134
rect -865 -191 272 -175
rect -1270 -236 -948 -228
rect -1270 -304 -1007 -236
rect -950 -304 -940 -236
rect -1270 -312 -948 -304
rect -1270 -512 -1105 -511
rect -1270 -520 -948 -512
rect -1270 -588 -1007 -520
rect -950 -588 -940 -520
rect -1270 -596 -948 -588
rect -1270 -597 -1105 -596
rect -865 -701 -830 -191
rect -775 -237 -683 -224
rect -775 -300 -763 -237
rect -692 -300 -683 -237
rect -775 -309 -683 -300
rect 310 -237 402 -227
rect 310 -299 322 -237
rect 392 -299 402 -237
rect 310 -312 402 -299
rect 1698 -292 1733 62
rect 2279 -124 2314 62
rect 3188 -22 3222 62
rect 4369 -22 4403 62
rect 3188 -64 4403 -22
rect 4369 -84 4403 -64
rect 4369 -100 4726 -84
rect 2012 -187 2022 -134
rect 2082 -187 2092 -134
rect 2279 -141 3416 -124
rect 2279 -175 3366 -141
rect 3400 -175 3416 -141
rect 4369 -134 4676 -100
rect 4710 -134 4726 -100
rect 4369 -150 4726 -134
rect 557 -354 622 -351
rect 557 -357 626 -354
rect 557 -417 563 -357
rect 622 -417 632 -357
rect 1698 -410 1879 -292
rect 2020 -344 2083 -187
rect 2279 -191 3416 -175
rect 2020 -352 2196 -344
rect 557 -421 626 -417
rect 557 -423 622 -421
rect 1698 -438 1880 -410
rect 2020 -420 2137 -352
rect 2194 -420 2204 -352
rect 2020 -428 2196 -420
rect 192 -520 284 -512
rect 192 -585 204 -520
rect 272 -585 284 -520
rect 192 -597 284 -585
rect 1698 -700 1733 -438
rect -865 -748 507 -701
rect 829 -747 1733 -700
rect -1270 -762 -943 -761
rect -1270 -824 -1007 -762
rect -953 -824 -943 -762
rect -31 -871 3 -748
rect 441 -761 507 -748
rect 441 -795 457 -761
rect 491 -795 507 -761
rect 441 -811 507 -795
rect 830 -871 864 -747
rect -36 -883 10 -871
rect -1270 -897 -943 -896
rect -1270 -959 -1007 -897
rect -953 -959 -943 -897
rect -1268 -1009 -941 -1008
rect -1268 -1071 -1005 -1009
rect -951 -1071 -941 -1009
rect -36 -1059 -30 -883
rect 4 -1059 10 -883
rect -36 -1071 10 -1059
rect 82 -883 202 -871
rect 82 -1059 88 -883
rect 122 -1059 162 -883
rect 82 -1071 162 -1059
rect -1268 -1134 -941 -1133
rect -1268 -1196 -1005 -1134
rect -951 -1196 -941 -1134
rect -1263 -1375 -936 -1374
rect -1263 -1437 -1000 -1375
rect -946 -1437 -936 -1375
rect 88 -1438 122 -1071
rect 156 -1259 162 -1071
rect 196 -1259 202 -883
rect 156 -1271 202 -1259
rect 274 -883 320 -871
rect 274 -1259 280 -883
rect 314 -1259 320 -883
rect 274 -1271 320 -1259
rect 392 -883 438 -871
rect 392 -1259 398 -883
rect 432 -1259 438 -883
rect 392 -1271 438 -1259
rect 510 -883 556 -871
rect 510 -1259 516 -883
rect 550 -1259 556 -883
rect 510 -1271 556 -1259
rect 628 -883 752 -871
rect 628 -1259 634 -883
rect 668 -1059 712 -883
rect 746 -1059 752 -883
rect 668 -1071 752 -1059
rect 824 -883 870 -871
rect 824 -1059 830 -883
rect 864 -1059 870 -883
rect 824 -1071 870 -1059
rect 668 -1259 674 -1071
rect 628 -1271 674 -1259
rect 398 -1344 432 -1271
rect 383 -1360 449 -1344
rect 383 -1394 399 -1360
rect 433 -1394 449 -1360
rect 383 -1410 449 -1394
rect 712 -1438 746 -1071
rect 88 -1490 746 -1438
rect 386 -1512 478 -1490
rect 386 -1564 398 -1512
rect 464 -1564 478 -1512
rect 386 -1568 478 -1564
rect -1266 -1597 -939 -1596
rect -1266 -1659 -1003 -1597
rect -949 -1659 -939 -1597
rect 1819 -1648 1880 -438
rect 2020 -520 2196 -512
rect 2020 -588 2137 -520
rect 2194 -588 2204 -520
rect 2020 -596 2196 -588
rect 2020 -758 2109 -596
rect 2279 -701 2314 -191
rect 2369 -237 2461 -224
rect 2369 -300 2381 -237
rect 2452 -300 2461 -237
rect 2369 -309 2461 -300
rect 3454 -237 3546 -227
rect 3454 -299 3466 -237
rect 3536 -299 3546 -237
rect 3454 -312 3546 -299
rect 4842 -292 4877 62
rect 5411 -120 5446 66
rect 6320 -18 6354 66
rect 7501 -18 7535 66
rect 6320 -60 7535 -18
rect 7501 -80 7535 -60
rect 7501 -96 7858 -80
rect 5411 -137 6548 -120
rect 5411 -171 6498 -137
rect 6532 -171 6548 -137
rect 7501 -130 7808 -96
rect 7842 -130 7858 -96
rect 7501 -146 7858 -130
rect 5411 -187 6548 -171
rect 3701 -354 3766 -351
rect 3701 -357 3770 -354
rect 3701 -417 3707 -357
rect 3766 -417 3776 -357
rect 3701 -421 3770 -417
rect 3701 -423 3766 -421
rect 4842 -438 5023 -292
rect 3336 -520 3428 -512
rect 3336 -585 3348 -520
rect 3416 -585 3428 -520
rect 3336 -597 3428 -585
rect 4842 -700 4877 -438
rect 2279 -748 3651 -701
rect 3973 -747 4877 -700
rect 2020 -818 2032 -758
rect 2102 -818 2112 -758
rect 2020 -825 2109 -818
rect 3113 -871 3147 -748
rect 3585 -761 3651 -748
rect 3585 -795 3601 -761
rect 3635 -795 3651 -761
rect 3585 -811 3651 -795
rect 3974 -871 4008 -747
rect 3108 -883 3154 -871
rect 3108 -1059 3114 -883
rect 3148 -1059 3154 -883
rect 3108 -1071 3154 -1059
rect 3226 -883 3346 -871
rect 3226 -1059 3232 -883
rect 3266 -1059 3306 -883
rect 3226 -1071 3306 -1059
rect 3232 -1438 3266 -1071
rect 3300 -1259 3306 -1071
rect 3340 -1259 3346 -883
rect 3300 -1271 3346 -1259
rect 3418 -883 3464 -871
rect 3418 -1259 3424 -883
rect 3458 -1259 3464 -883
rect 3418 -1271 3464 -1259
rect 3536 -883 3582 -871
rect 3536 -1259 3542 -883
rect 3576 -1259 3582 -883
rect 3536 -1271 3582 -1259
rect 3654 -883 3700 -871
rect 3654 -1259 3660 -883
rect 3694 -1259 3700 -883
rect 3654 -1271 3700 -1259
rect 3772 -883 3896 -871
rect 3772 -1259 3778 -883
rect 3812 -1059 3856 -883
rect 3890 -1059 3896 -883
rect 3812 -1071 3896 -1059
rect 3968 -883 4014 -871
rect 3968 -1059 3974 -883
rect 4008 -1059 4014 -883
rect 3968 -1071 4014 -1059
rect 3812 -1259 3818 -1071
rect 3772 -1271 3818 -1259
rect 3542 -1344 3576 -1271
rect 3527 -1360 3593 -1344
rect 3527 -1394 3543 -1360
rect 3577 -1394 3593 -1360
rect 3527 -1410 3593 -1394
rect 3856 -1438 3890 -1071
rect 4935 -1368 5023 -438
rect 5152 -516 5328 -508
rect 5152 -584 5269 -516
rect 5326 -584 5336 -516
rect 5152 -592 5328 -584
rect 5172 -899 5249 -592
rect 5411 -697 5446 -187
rect 5501 -233 5593 -220
rect 5501 -296 5513 -233
rect 5584 -296 5593 -233
rect 5501 -305 5593 -296
rect 6586 -233 6678 -223
rect 6586 -295 6598 -233
rect 6668 -295 6678 -233
rect 6586 -308 6678 -295
rect 7974 -288 8009 66
rect 8555 -120 8590 66
rect 9464 -18 9498 66
rect 10645 -18 10679 66
rect 9464 -60 10679 -18
rect 10645 -80 10679 -60
rect 10645 -96 11002 -80
rect 8555 -137 9692 -120
rect 8555 -171 9642 -137
rect 9676 -171 9692 -137
rect 10645 -130 10952 -96
rect 10986 -130 11002 -96
rect 10645 -146 11002 -130
rect 8555 -187 9692 -171
rect 6833 -350 6898 -347
rect 6833 -353 6902 -350
rect 6833 -413 6839 -353
rect 6898 -413 6908 -353
rect 6833 -417 6902 -413
rect 6833 -419 6898 -417
rect 7974 -434 8155 -288
rect 8401 -348 8472 -340
rect 8401 -416 8413 -348
rect 8470 -416 8480 -348
rect 8401 -424 8472 -416
rect 6468 -516 6560 -508
rect 6468 -581 6480 -516
rect 6548 -581 6560 -516
rect 6468 -593 6560 -581
rect 7974 -696 8009 -434
rect 5411 -744 6783 -697
rect 7105 -743 8009 -696
rect 6245 -867 6279 -744
rect 6717 -757 6783 -744
rect 6717 -791 6733 -757
rect 6767 -791 6783 -757
rect 6717 -807 6783 -791
rect 7106 -867 7140 -743
rect 6240 -879 6286 -867
rect 5172 -956 5182 -899
rect 5246 -956 5256 -899
rect 5172 -960 5249 -956
rect 6240 -1055 6246 -879
rect 6280 -1055 6286 -879
rect 6240 -1067 6286 -1055
rect 6358 -879 6478 -867
rect 6358 -1055 6364 -879
rect 6398 -1055 6438 -879
rect 6358 -1067 6438 -1055
rect 4904 -1434 4914 -1368
rect 4973 -1434 5023 -1368
rect 6364 -1434 6398 -1067
rect 6432 -1255 6438 -1067
rect 6472 -1255 6478 -879
rect 6432 -1267 6478 -1255
rect 6550 -879 6596 -867
rect 6550 -1255 6556 -879
rect 6590 -1255 6596 -879
rect 6550 -1267 6596 -1255
rect 6668 -879 6714 -867
rect 6668 -1255 6674 -879
rect 6708 -1255 6714 -879
rect 6668 -1267 6714 -1255
rect 6786 -879 6832 -867
rect 6786 -1255 6792 -879
rect 6826 -1255 6832 -879
rect 6786 -1267 6832 -1255
rect 6904 -879 7028 -867
rect 6904 -1255 6910 -879
rect 6944 -1055 6988 -879
rect 7022 -1055 7028 -879
rect 6944 -1067 7028 -1055
rect 7100 -879 7146 -867
rect 7100 -1055 7106 -879
rect 7140 -1055 7146 -879
rect 7100 -1067 7146 -1055
rect 6944 -1255 6950 -1067
rect 6904 -1267 6950 -1255
rect 6674 -1340 6708 -1267
rect 6659 -1356 6725 -1340
rect 6659 -1390 6675 -1356
rect 6709 -1390 6725 -1356
rect 6659 -1406 6725 -1390
rect 6988 -1434 7022 -1067
rect 8058 -1251 8155 -434
rect 8296 -516 8472 -508
rect 8296 -584 8413 -516
rect 8470 -584 8480 -516
rect 8296 -592 8472 -584
rect 8301 -1004 8389 -592
rect 8555 -697 8590 -187
rect 8645 -233 8737 -220
rect 8645 -296 8657 -233
rect 8728 -296 8737 -233
rect 8645 -305 8737 -296
rect 9730 -233 9822 -223
rect 9730 -295 9742 -233
rect 9812 -295 9822 -233
rect 9730 -308 9822 -295
rect 11118 -288 11153 66
rect 11752 62 11798 74
rect 11870 250 11916 262
rect 11870 74 11876 250
rect 11910 74 11916 250
rect 11870 62 11916 74
rect 11988 250 12034 262
rect 11988 74 11994 250
rect 12028 74 12034 250
rect 11988 62 12034 74
rect 12106 250 12199 262
rect 12106 74 12112 250
rect 12146 74 12199 250
rect 12233 74 12239 450
rect 12106 62 12239 74
rect 12311 450 12357 462
rect 12311 74 12317 450
rect 12351 74 12357 450
rect 12311 62 12357 74
rect 12429 450 12475 462
rect 12429 74 12435 450
rect 12469 74 12475 450
rect 12429 62 12475 74
rect 12547 450 12593 462
rect 12547 74 12553 450
rect 12587 74 12593 450
rect 12547 62 12593 74
rect 12660 450 12706 462
rect 12660 74 12666 450
rect 12700 74 12706 450
rect 12660 62 12706 74
rect 12778 450 12824 462
rect 12778 74 12784 450
rect 12818 74 12824 450
rect 12778 62 12824 74
rect 12896 450 12942 462
rect 12896 74 12902 450
rect 12936 74 12942 450
rect 12896 62 12942 74
rect 13014 450 13060 462
rect 13014 74 13020 450
rect 13054 74 13060 450
rect 13014 62 13060 74
rect 13132 450 13178 462
rect 13132 74 13138 450
rect 13172 74 13178 450
rect 13132 62 13178 74
rect 13250 450 13296 462
rect 13250 74 13256 450
rect 13290 74 13296 450
rect 13250 62 13296 74
rect 13368 450 13414 462
rect 13368 74 13374 450
rect 13408 74 13414 450
rect 13368 62 13414 74
rect 13487 450 13533 462
rect 13487 74 13493 450
rect 13527 74 13533 450
rect 13487 62 13533 74
rect 13605 450 13651 462
rect 13605 74 13611 450
rect 13645 74 13651 450
rect 13605 62 13651 74
rect 13723 450 13769 462
rect 13723 74 13729 450
rect 13763 74 13769 450
rect 13723 62 13769 74
rect 13841 450 13887 462
rect 13841 74 13847 450
rect 13881 74 13887 450
rect 13965 262 14002 549
rect 15343 549 17146 606
rect 15343 462 15377 549
rect 16518 462 16552 549
rect 15337 450 15383 462
rect 15337 262 15343 450
rect 13841 62 13887 74
rect 13960 250 14006 262
rect 13960 74 13966 250
rect 14000 74 14006 250
rect 13960 62 14006 74
rect 14078 250 14124 262
rect 14078 74 14084 250
rect 14118 74 14124 250
rect 14078 62 14124 74
rect 14196 250 14242 262
rect 14196 74 14202 250
rect 14236 74 14242 250
rect 14196 62 14242 74
rect 14314 250 14360 262
rect 14314 74 14320 250
rect 14354 74 14360 250
rect 14314 62 14360 74
rect 14896 250 14942 262
rect 14896 74 14902 250
rect 14936 74 14942 250
rect 14896 62 14942 74
rect 15014 250 15060 262
rect 15014 74 15020 250
rect 15054 74 15060 250
rect 15014 62 15060 74
rect 15132 250 15178 262
rect 15132 74 15138 250
rect 15172 74 15178 250
rect 15132 62 15178 74
rect 15250 250 15343 262
rect 15250 74 15256 250
rect 15290 74 15343 250
rect 15377 74 15383 450
rect 15250 62 15383 74
rect 15455 450 15501 462
rect 15455 74 15461 450
rect 15495 74 15501 450
rect 15455 62 15501 74
rect 15573 450 15619 462
rect 15573 74 15579 450
rect 15613 74 15619 450
rect 15573 62 15619 74
rect 15691 450 15737 462
rect 15691 74 15697 450
rect 15731 74 15737 450
rect 15691 62 15737 74
rect 15804 450 15850 462
rect 15804 74 15810 450
rect 15844 74 15850 450
rect 15804 62 15850 74
rect 15922 450 15968 462
rect 15922 74 15928 450
rect 15962 74 15968 450
rect 15922 62 15968 74
rect 16040 450 16086 462
rect 16040 74 16046 450
rect 16080 74 16086 450
rect 16040 62 16086 74
rect 16158 450 16204 462
rect 16158 74 16164 450
rect 16198 74 16204 450
rect 16158 62 16204 74
rect 16276 450 16322 462
rect 16276 74 16282 450
rect 16316 74 16322 450
rect 16276 62 16322 74
rect 16394 450 16440 462
rect 16394 74 16400 450
rect 16434 74 16440 450
rect 16394 62 16440 74
rect 16512 450 16558 462
rect 16512 74 16518 450
rect 16552 74 16558 450
rect 16512 62 16558 74
rect 16631 450 16677 462
rect 16631 74 16637 450
rect 16671 74 16677 450
rect 16631 62 16677 74
rect 16749 450 16795 462
rect 16749 74 16755 450
rect 16789 74 16795 450
rect 16749 62 16795 74
rect 16867 450 16913 462
rect 16867 74 16873 450
rect 16907 74 16913 450
rect 16867 62 16913 74
rect 16985 450 17031 462
rect 16985 74 16991 450
rect 17025 74 17031 450
rect 17109 262 17146 549
rect 18475 553 20278 610
rect 18475 466 18509 553
rect 19650 466 19684 553
rect 18469 454 18515 466
rect 18469 266 18475 454
rect 16985 62 17031 74
rect 17104 250 17150 262
rect 17104 74 17110 250
rect 17144 74 17150 250
rect 17104 62 17150 74
rect 17222 250 17268 262
rect 17222 74 17228 250
rect 17262 74 17268 250
rect 17222 62 17268 74
rect 17340 250 17386 262
rect 17340 74 17346 250
rect 17380 74 17386 250
rect 17340 62 17386 74
rect 17458 250 17504 262
rect 17458 74 17464 250
rect 17498 74 17504 250
rect 17458 62 17504 74
rect 18028 254 18074 266
rect 18028 78 18034 254
rect 18068 78 18074 254
rect 18028 66 18074 78
rect 18146 254 18192 266
rect 18146 78 18152 254
rect 18186 78 18192 254
rect 18146 66 18192 78
rect 18264 254 18310 266
rect 18264 78 18270 254
rect 18304 78 18310 254
rect 18264 66 18310 78
rect 18382 254 18475 266
rect 18382 78 18388 254
rect 18422 78 18475 254
rect 18509 78 18515 454
rect 18382 66 18515 78
rect 18587 454 18633 466
rect 18587 78 18593 454
rect 18627 78 18633 454
rect 18587 66 18633 78
rect 18705 454 18751 466
rect 18705 78 18711 454
rect 18745 78 18751 454
rect 18705 66 18751 78
rect 18823 454 18869 466
rect 18823 78 18829 454
rect 18863 78 18869 454
rect 18823 66 18869 78
rect 18936 454 18982 466
rect 18936 78 18942 454
rect 18976 78 18982 454
rect 18936 66 18982 78
rect 19054 454 19100 466
rect 19054 78 19060 454
rect 19094 78 19100 454
rect 19054 66 19100 78
rect 19172 454 19218 466
rect 19172 78 19178 454
rect 19212 78 19218 454
rect 19172 66 19218 78
rect 19290 454 19336 466
rect 19290 78 19296 454
rect 19330 78 19336 454
rect 19290 66 19336 78
rect 19408 454 19454 466
rect 19408 78 19414 454
rect 19448 78 19454 454
rect 19408 66 19454 78
rect 19526 454 19572 466
rect 19526 78 19532 454
rect 19566 78 19572 454
rect 19526 66 19572 78
rect 19644 454 19690 466
rect 19644 78 19650 454
rect 19684 78 19690 454
rect 19644 66 19690 78
rect 19763 454 19809 466
rect 19763 78 19769 454
rect 19803 78 19809 454
rect 19763 66 19809 78
rect 19881 454 19927 466
rect 19881 78 19887 454
rect 19921 78 19927 454
rect 19881 66 19927 78
rect 19999 454 20045 466
rect 19999 78 20005 454
rect 20039 78 20045 454
rect 19999 66 20045 78
rect 20117 454 20163 466
rect 20117 78 20123 454
rect 20157 78 20163 454
rect 20241 266 20278 553
rect 21619 553 23422 610
rect 21619 466 21653 553
rect 22794 466 22828 553
rect 21613 454 21659 466
rect 21613 266 21619 454
rect 20117 66 20163 78
rect 20236 254 20282 266
rect 20236 78 20242 254
rect 20276 78 20282 254
rect 20236 66 20282 78
rect 20354 254 20400 266
rect 20354 78 20360 254
rect 20394 78 20400 254
rect 20354 66 20400 78
rect 20472 254 20518 266
rect 20472 78 20478 254
rect 20512 78 20518 254
rect 20472 66 20518 78
rect 20590 254 20636 266
rect 20590 78 20596 254
rect 20630 78 20636 254
rect 20590 66 20636 78
rect 21172 254 21218 266
rect 21172 78 21178 254
rect 21212 78 21218 254
rect 21172 66 21218 78
rect 21290 254 21336 266
rect 21290 78 21296 254
rect 21330 78 21336 254
rect 21290 66 21336 78
rect 21408 254 21454 266
rect 21408 78 21414 254
rect 21448 78 21454 254
rect 21408 66 21454 78
rect 21526 254 21619 266
rect 21526 78 21532 254
rect 21566 78 21619 254
rect 21653 78 21659 454
rect 21526 66 21659 78
rect 21731 454 21777 466
rect 21731 78 21737 454
rect 21771 78 21777 454
rect 21731 66 21777 78
rect 21849 454 21895 466
rect 21849 78 21855 454
rect 21889 78 21895 454
rect 21849 66 21895 78
rect 21967 454 22013 466
rect 21967 78 21973 454
rect 22007 78 22013 454
rect 21967 66 22013 78
rect 22080 454 22126 466
rect 22080 78 22086 454
rect 22120 78 22126 454
rect 22080 66 22126 78
rect 22198 454 22244 466
rect 22198 78 22204 454
rect 22238 78 22244 454
rect 22198 66 22244 78
rect 22316 454 22362 466
rect 22316 78 22322 454
rect 22356 78 22362 454
rect 22316 66 22362 78
rect 22434 454 22480 466
rect 22434 78 22440 454
rect 22474 78 22480 454
rect 22434 66 22480 78
rect 22552 454 22598 466
rect 22552 78 22558 454
rect 22592 78 22598 454
rect 22552 66 22598 78
rect 22670 454 22716 466
rect 22670 78 22676 454
rect 22710 78 22716 454
rect 22670 66 22716 78
rect 22788 454 22834 466
rect 22788 78 22794 454
rect 22828 78 22834 454
rect 22788 66 22834 78
rect 22907 454 22953 466
rect 22907 78 22913 454
rect 22947 78 22953 454
rect 22907 66 22953 78
rect 23025 454 23071 466
rect 23025 78 23031 454
rect 23065 78 23071 454
rect 23025 66 23071 78
rect 23143 454 23189 466
rect 23143 78 23149 454
rect 23183 78 23189 454
rect 23143 66 23189 78
rect 23261 454 23307 466
rect 23261 78 23267 454
rect 23301 78 23307 454
rect 23385 266 23422 553
rect 23261 66 23307 78
rect 23380 254 23426 266
rect 23380 78 23386 254
rect 23420 78 23426 254
rect 23380 66 23426 78
rect 23498 254 23544 266
rect 23498 78 23504 254
rect 23538 78 23544 254
rect 23498 66 23544 78
rect 23616 254 23662 266
rect 23616 78 23622 254
rect 23656 78 23662 254
rect 23616 66 23662 78
rect 23734 254 23780 266
rect 23734 78 23740 254
rect 23774 78 23780 254
rect 23734 66 23780 78
rect 11757 -124 11792 62
rect 12666 -22 12700 62
rect 13847 -22 13881 62
rect 12666 -64 13881 -22
rect 13847 -84 13881 -64
rect 13847 -100 14204 -84
rect 11757 -141 12894 -124
rect 11757 -175 12844 -141
rect 12878 -175 12894 -141
rect 13847 -134 14154 -100
rect 14188 -134 14204 -100
rect 13847 -150 14204 -134
rect 11757 -191 12894 -175
rect 9977 -350 10042 -347
rect 9977 -353 10046 -350
rect 9977 -413 9983 -353
rect 10042 -413 10052 -353
rect 9977 -417 10046 -413
rect 9977 -419 10042 -417
rect 11118 -434 11299 -288
rect 9612 -516 9704 -508
rect 9612 -581 9624 -516
rect 9692 -581 9704 -516
rect 9612 -593 9704 -581
rect 11118 -696 11153 -434
rect 8555 -744 9927 -697
rect 10249 -743 11153 -696
rect 9389 -867 9423 -744
rect 9861 -757 9927 -744
rect 9861 -791 9877 -757
rect 9911 -791 9927 -757
rect 9861 -807 9927 -791
rect 10250 -867 10284 -743
rect 8301 -1062 8324 -1004
rect 8378 -1062 8389 -1004
rect 8301 -1072 8389 -1062
rect 9384 -879 9430 -867
rect 9384 -1055 9390 -879
rect 9424 -1055 9430 -879
rect 9384 -1067 9430 -1055
rect 9502 -879 9622 -867
rect 9502 -1055 9508 -879
rect 9542 -1055 9582 -879
rect 9502 -1067 9582 -1055
rect 8030 -1308 8040 -1251
rect 8099 -1308 8155 -1251
rect 8030 -1309 8155 -1308
rect 3232 -1490 3890 -1438
rect 6364 -1486 7022 -1434
rect 9508 -1434 9542 -1067
rect 9576 -1255 9582 -1067
rect 9616 -1255 9622 -879
rect 9576 -1267 9622 -1255
rect 9694 -879 9740 -867
rect 9694 -1255 9700 -879
rect 9734 -1255 9740 -879
rect 9694 -1267 9740 -1255
rect 9812 -879 9858 -867
rect 9812 -1255 9818 -879
rect 9852 -1255 9858 -879
rect 9812 -1267 9858 -1255
rect 9930 -879 9976 -867
rect 9930 -1255 9936 -879
rect 9970 -1255 9976 -879
rect 9930 -1267 9976 -1255
rect 10048 -879 10172 -867
rect 10048 -1255 10054 -879
rect 10088 -1055 10132 -879
rect 10166 -1055 10172 -879
rect 10088 -1067 10172 -1055
rect 10244 -879 10290 -867
rect 10244 -1055 10250 -879
rect 10284 -1055 10290 -879
rect 10244 -1067 10290 -1055
rect 10088 -1255 10094 -1067
rect 10048 -1267 10094 -1255
rect 9818 -1340 9852 -1267
rect 9803 -1356 9869 -1340
rect 9803 -1390 9819 -1356
rect 9853 -1390 9869 -1356
rect 9803 -1406 9869 -1390
rect 10132 -1434 10166 -1067
rect 11205 -1103 11298 -434
rect 11205 -1171 11215 -1103
rect 11277 -1171 11298 -1103
rect 11205 -1176 11298 -1171
rect 11498 -520 11674 -512
rect 11498 -588 11615 -520
rect 11672 -588 11682 -520
rect 11498 -596 11674 -588
rect 11498 -1228 11564 -596
rect 11757 -701 11792 -191
rect 11847 -237 11939 -224
rect 11847 -300 11859 -237
rect 11930 -300 11939 -237
rect 11847 -309 11939 -300
rect 12932 -237 13024 -227
rect 12932 -299 12944 -237
rect 13014 -299 13024 -237
rect 12932 -312 13024 -299
rect 14320 -292 14355 62
rect 14901 -124 14936 62
rect 15810 -22 15844 62
rect 16991 -22 17025 62
rect 15810 -64 17025 -22
rect 16991 -84 17025 -64
rect 16991 -100 17348 -84
rect 14901 -141 16038 -124
rect 14901 -175 15988 -141
rect 16022 -175 16038 -141
rect 16991 -134 17298 -100
rect 17332 -134 17348 -100
rect 16991 -150 17348 -134
rect 14901 -191 16038 -175
rect 13179 -354 13244 -351
rect 13179 -357 13248 -354
rect 13179 -417 13185 -357
rect 13244 -417 13254 -357
rect 13179 -421 13248 -417
rect 13179 -423 13244 -421
rect 14320 -438 14501 -292
rect 14747 -352 14818 -347
rect 14747 -420 14759 -352
rect 14816 -420 14826 -352
rect 14747 -426 14818 -420
rect 12814 -520 12906 -512
rect 12814 -585 12826 -520
rect 12894 -585 12906 -520
rect 12814 -597 12906 -585
rect 14320 -700 14355 -438
rect 11757 -748 13129 -701
rect 13451 -747 14355 -700
rect 12591 -871 12625 -748
rect 13063 -761 13129 -748
rect 13063 -795 13079 -761
rect 13113 -795 13129 -761
rect 13063 -811 13129 -795
rect 13452 -871 13486 -747
rect 12586 -883 12632 -871
rect 12586 -1059 12592 -883
rect 12626 -1059 12632 -883
rect 12586 -1071 12632 -1059
rect 12704 -883 12824 -871
rect 12704 -1059 12710 -883
rect 12744 -1059 12784 -883
rect 12704 -1071 12784 -1059
rect 11484 -1289 11494 -1228
rect 11563 -1289 11573 -1228
rect 11484 -1297 11573 -1289
rect 9508 -1486 10166 -1434
rect 12710 -1438 12744 -1071
rect 12778 -1259 12784 -1071
rect 12818 -1259 12824 -883
rect 12778 -1271 12824 -1259
rect 12896 -883 12942 -871
rect 12896 -1259 12902 -883
rect 12936 -1259 12942 -883
rect 12896 -1271 12942 -1259
rect 13014 -883 13060 -871
rect 13014 -1259 13020 -883
rect 13054 -1259 13060 -883
rect 13014 -1271 13060 -1259
rect 13132 -883 13178 -871
rect 13132 -1259 13138 -883
rect 13172 -1259 13178 -883
rect 13132 -1271 13178 -1259
rect 13250 -883 13374 -871
rect 13250 -1259 13256 -883
rect 13290 -1059 13334 -883
rect 13368 -1059 13374 -883
rect 13290 -1071 13374 -1059
rect 13446 -883 13492 -871
rect 13446 -1059 13452 -883
rect 13486 -1059 13492 -883
rect 14431 -952 14501 -438
rect 14642 -520 14818 -512
rect 14642 -588 14759 -520
rect 14816 -588 14826 -520
rect 14642 -596 14818 -588
rect 14430 -1021 14440 -952
rect 14496 -1021 14506 -952
rect 14431 -1027 14501 -1021
rect 13446 -1071 13492 -1059
rect 13290 -1259 13296 -1071
rect 13250 -1271 13296 -1259
rect 13020 -1344 13054 -1271
rect 13005 -1360 13071 -1344
rect 13005 -1394 13021 -1360
rect 13055 -1394 13071 -1360
rect 13005 -1410 13071 -1394
rect 13334 -1438 13368 -1071
rect 14642 -1363 14725 -596
rect 14901 -701 14936 -191
rect 14991 -237 15083 -224
rect 14991 -300 15003 -237
rect 15074 -300 15083 -237
rect 14991 -309 15083 -300
rect 16076 -237 16168 -227
rect 16076 -299 16088 -237
rect 16158 -299 16168 -237
rect 16076 -312 16168 -299
rect 17464 -292 17499 62
rect 18033 -120 18068 66
rect 18942 -18 18976 66
rect 20123 -18 20157 66
rect 18942 -60 20157 -18
rect 20123 -80 20157 -60
rect 20123 -96 20480 -80
rect 18033 -137 19170 -120
rect 18033 -171 19120 -137
rect 19154 -171 19170 -137
rect 20123 -130 20430 -96
rect 20464 -130 20480 -96
rect 20123 -146 20480 -130
rect 18033 -187 19170 -171
rect 16323 -354 16388 -351
rect 16323 -357 16392 -354
rect 16323 -417 16329 -357
rect 16388 -417 16398 -357
rect 16323 -421 16392 -417
rect 16323 -423 16388 -421
rect 17464 -438 17645 -292
rect 17880 -348 17950 -343
rect 17880 -416 17891 -348
rect 17948 -416 17958 -348
rect 17880 -422 17950 -416
rect 15958 -520 16050 -512
rect 15958 -585 15970 -520
rect 16038 -585 16050 -520
rect 15958 -597 16050 -585
rect 17464 -700 17499 -438
rect 14901 -748 16273 -701
rect 16595 -747 17499 -700
rect 15735 -871 15769 -748
rect 16207 -761 16273 -748
rect 16207 -795 16223 -761
rect 16257 -795 16273 -761
rect 16207 -811 16273 -795
rect 16596 -871 16630 -747
rect 17573 -799 17645 -438
rect 17774 -516 17950 -508
rect 17774 -584 17891 -516
rect 17948 -584 17958 -516
rect 17774 -592 17950 -584
rect 17566 -858 17576 -799
rect 17640 -858 17650 -799
rect 15730 -883 15776 -871
rect 15730 -1059 15736 -883
rect 15770 -1059 15776 -883
rect 15730 -1071 15776 -1059
rect 15848 -883 15968 -871
rect 15848 -1059 15854 -883
rect 15888 -1059 15928 -883
rect 15848 -1071 15928 -1059
rect 14635 -1430 14645 -1363
rect 14702 -1427 14725 -1363
rect 14702 -1430 14712 -1427
rect 3530 -1512 3622 -1490
rect 3530 -1564 3542 -1512
rect 3608 -1564 3622 -1512
rect 6662 -1508 6754 -1486
rect 6662 -1560 6674 -1508
rect 6740 -1560 6754 -1508
rect 6662 -1564 6754 -1560
rect 9806 -1508 9898 -1486
rect 12710 -1490 13368 -1438
rect 15854 -1438 15888 -1071
rect 15922 -1259 15928 -1071
rect 15962 -1259 15968 -883
rect 15922 -1271 15968 -1259
rect 16040 -883 16086 -871
rect 16040 -1259 16046 -883
rect 16080 -1259 16086 -883
rect 16040 -1271 16086 -1259
rect 16158 -883 16204 -871
rect 16158 -1259 16164 -883
rect 16198 -1259 16204 -883
rect 16158 -1271 16204 -1259
rect 16276 -883 16322 -871
rect 16276 -1259 16282 -883
rect 16316 -1259 16322 -883
rect 16276 -1271 16322 -1259
rect 16394 -883 16518 -871
rect 16394 -1259 16400 -883
rect 16434 -1059 16478 -883
rect 16512 -1059 16518 -883
rect 16434 -1071 16518 -1059
rect 16590 -883 16636 -871
rect 16590 -1059 16596 -883
rect 16630 -1059 16636 -883
rect 16590 -1071 16636 -1059
rect 16434 -1259 16440 -1071
rect 16394 -1271 16440 -1259
rect 16164 -1344 16198 -1271
rect 16149 -1360 16215 -1344
rect 16149 -1394 16165 -1360
rect 16199 -1394 16215 -1360
rect 16149 -1410 16215 -1394
rect 16478 -1438 16512 -1071
rect 15854 -1490 16512 -1438
rect 9806 -1560 9818 -1508
rect 9884 -1560 9898 -1508
rect 9806 -1564 9898 -1560
rect 13008 -1512 13100 -1490
rect 13008 -1564 13020 -1512
rect 13086 -1564 13100 -1512
rect 3530 -1568 3622 -1564
rect 13008 -1568 13100 -1564
rect 16152 -1512 16244 -1490
rect 16152 -1564 16164 -1512
rect 16230 -1564 16244 -1512
rect 16152 -1568 16244 -1564
rect 17774 -1579 17847 -592
rect 18033 -697 18068 -187
rect 18123 -233 18215 -220
rect 18123 -296 18135 -233
rect 18206 -296 18215 -233
rect 18123 -305 18215 -296
rect 19208 -233 19300 -223
rect 19208 -295 19220 -233
rect 19290 -295 19300 -233
rect 19208 -308 19300 -295
rect 20596 -288 20631 66
rect 21177 -120 21212 66
rect 22086 -18 22120 66
rect 23267 -18 23301 66
rect 22086 -60 23301 -18
rect 23267 -80 23301 -60
rect 23267 -96 23624 -80
rect 21177 -137 22314 -120
rect 21177 -171 22264 -137
rect 22298 -171 22314 -137
rect 23267 -130 23574 -96
rect 23608 -130 23624 -96
rect 23267 -146 23624 -130
rect 21177 -187 22314 -171
rect 19455 -350 19520 -347
rect 19455 -353 19524 -350
rect 19455 -413 19461 -353
rect 19520 -413 19530 -353
rect 20596 -383 20777 -288
rect 21024 -348 21094 -343
rect 19455 -417 19524 -413
rect 19455 -419 19520 -417
rect 20596 -434 20778 -383
rect 21024 -416 21035 -348
rect 21092 -416 21102 -348
rect 21024 -422 21094 -416
rect 19090 -516 19182 -508
rect 19090 -581 19102 -516
rect 19170 -581 19182 -516
rect 19090 -593 19182 -581
rect 20596 -696 20631 -434
rect 18033 -744 19405 -697
rect 19727 -743 20631 -696
rect 20683 -672 20778 -434
rect 20683 -729 20721 -672
rect 20774 -729 20784 -672
rect 21177 -697 21212 -187
rect 21267 -233 21359 -220
rect 21267 -296 21279 -233
rect 21350 -296 21359 -233
rect 21267 -305 21359 -296
rect 22352 -233 22444 -223
rect 22352 -295 22364 -233
rect 22434 -295 22444 -233
rect 22352 -308 22444 -295
rect 23740 -288 23775 66
rect 22599 -350 22664 -347
rect 22599 -353 22668 -350
rect 22599 -413 22605 -353
rect 22664 -413 22674 -353
rect 23740 -376 24354 -288
rect 22599 -417 22668 -413
rect 22599 -419 22664 -417
rect 22234 -516 22326 -508
rect 22234 -581 22246 -516
rect 22314 -581 22326 -516
rect 22234 -593 22326 -581
rect 23740 -696 23775 -376
rect 20683 -737 20778 -729
rect 18867 -867 18901 -744
rect 19339 -757 19405 -744
rect 19339 -791 19355 -757
rect 19389 -791 19405 -757
rect 19339 -807 19405 -791
rect 19728 -867 19762 -743
rect 21177 -744 22549 -697
rect 22871 -743 23775 -696
rect 24206 -664 24355 -652
rect 24206 -735 24219 -664
rect 24290 -735 24355 -664
rect 22011 -867 22045 -744
rect 22483 -757 22549 -744
rect 22483 -791 22499 -757
rect 22533 -791 22549 -757
rect 22483 -807 22549 -791
rect 22872 -867 22906 -743
rect 24206 -746 24355 -735
rect 24197 -800 24356 -789
rect 24197 -860 24207 -800
rect 24273 -860 24356 -800
rect 18862 -879 18908 -867
rect 18862 -1055 18868 -879
rect 18902 -1055 18908 -879
rect 18862 -1067 18908 -1055
rect 18980 -879 19100 -867
rect 18980 -1055 18986 -879
rect 19020 -1055 19060 -879
rect 18980 -1067 19060 -1055
rect 18986 -1434 19020 -1067
rect 19054 -1255 19060 -1067
rect 19094 -1255 19100 -879
rect 19054 -1267 19100 -1255
rect 19172 -879 19218 -867
rect 19172 -1255 19178 -879
rect 19212 -1255 19218 -879
rect 19172 -1267 19218 -1255
rect 19290 -879 19336 -867
rect 19290 -1255 19296 -879
rect 19330 -1255 19336 -879
rect 19290 -1267 19336 -1255
rect 19408 -879 19454 -867
rect 19408 -1255 19414 -879
rect 19448 -1255 19454 -879
rect 19408 -1267 19454 -1255
rect 19526 -879 19650 -867
rect 19526 -1255 19532 -879
rect 19566 -1055 19610 -879
rect 19644 -1055 19650 -879
rect 19566 -1067 19650 -1055
rect 19722 -879 19768 -867
rect 19722 -1055 19728 -879
rect 19762 -1055 19768 -879
rect 19722 -1067 19768 -1055
rect 22006 -879 22052 -867
rect 22006 -1055 22012 -879
rect 22046 -1055 22052 -879
rect 22006 -1067 22052 -1055
rect 22124 -879 22244 -867
rect 22124 -1055 22130 -879
rect 22164 -1055 22204 -879
rect 22124 -1067 22204 -1055
rect 19566 -1255 19572 -1067
rect 19526 -1267 19572 -1255
rect 19296 -1340 19330 -1267
rect 19281 -1356 19347 -1340
rect 19281 -1390 19297 -1356
rect 19331 -1390 19347 -1356
rect 19281 -1406 19347 -1390
rect 19610 -1434 19644 -1067
rect 18986 -1486 19644 -1434
rect 22130 -1434 22164 -1067
rect 22198 -1255 22204 -1067
rect 22238 -1255 22244 -879
rect 22198 -1267 22244 -1255
rect 22316 -879 22362 -867
rect 22316 -1255 22322 -879
rect 22356 -1255 22362 -879
rect 22316 -1267 22362 -1255
rect 22434 -879 22480 -867
rect 22434 -1255 22440 -879
rect 22474 -1255 22480 -879
rect 22434 -1267 22480 -1255
rect 22552 -879 22598 -867
rect 22552 -1255 22558 -879
rect 22592 -1255 22598 -879
rect 22552 -1267 22598 -1255
rect 22670 -879 22794 -867
rect 22670 -1255 22676 -879
rect 22710 -1055 22754 -879
rect 22788 -1055 22794 -879
rect 22710 -1067 22794 -1055
rect 22866 -879 22912 -867
rect 24197 -871 24356 -860
rect 22866 -1055 22872 -879
rect 22906 -1055 22912 -879
rect 24186 -958 24356 -947
rect 24186 -1027 24197 -958
rect 24261 -1027 24356 -958
rect 24186 -1038 24356 -1027
rect 22866 -1067 22912 -1055
rect 22710 -1255 22716 -1067
rect 22670 -1267 22716 -1255
rect 22440 -1340 22474 -1267
rect 22425 -1356 22491 -1340
rect 22425 -1390 22441 -1356
rect 22475 -1390 22491 -1356
rect 22425 -1406 22491 -1390
rect 22754 -1434 22788 -1067
rect 24186 -1104 24356 -1093
rect 24186 -1173 24197 -1104
rect 24261 -1173 24356 -1104
rect 24186 -1184 24356 -1173
rect 24186 -1244 24356 -1233
rect 24186 -1313 24197 -1244
rect 24261 -1313 24356 -1244
rect 24186 -1324 24356 -1313
rect 22130 -1486 22788 -1434
rect 24185 -1383 24355 -1372
rect 24185 -1452 24196 -1383
rect 24260 -1452 24355 -1383
rect 24185 -1463 24355 -1452
rect 19284 -1508 19376 -1486
rect 19284 -1560 19296 -1508
rect 19362 -1560 19376 -1508
rect 19284 -1564 19376 -1560
rect 22428 -1508 22520 -1486
rect 22428 -1560 22440 -1508
rect 22506 -1560 22520 -1508
rect 22428 -1564 22520 -1560
rect 1771 -1729 1781 -1648
rect 1854 -1729 1880 -1648
rect 17764 -1655 17774 -1579
rect 17844 -1655 17854 -1579
rect 24185 -1651 24355 -1640
rect 1819 -1730 1880 -1729
rect 24185 -1720 24196 -1651
rect 24260 -1720 24355 -1651
rect 24185 -1731 24355 -1720
<< via1 >>
rect 384 700 464 706
rect 384 646 388 700
rect 388 646 460 700
rect 460 646 464 700
rect 3528 700 3608 706
rect 3528 646 3532 700
rect 3532 646 3604 700
rect 3604 646 3608 700
rect 6660 704 6740 710
rect 6660 650 6664 704
rect 6664 650 6736 704
rect 6736 650 6740 704
rect 9804 704 9884 710
rect 9804 650 9808 704
rect 9808 650 9880 704
rect 9880 650 9884 704
rect 13006 700 13086 706
rect 13006 646 13010 700
rect 13010 646 13082 700
rect 13082 646 13086 700
rect 16150 700 16230 706
rect 16150 646 16154 700
rect 16154 646 16226 700
rect 16226 646 16230 700
rect 19282 704 19362 710
rect 19282 650 19286 704
rect 19286 650 19358 704
rect 19358 650 19362 704
rect 22426 704 22506 710
rect 22426 650 22430 704
rect 22430 650 22502 704
rect 22502 650 22506 704
rect -1006 -149 -952 -87
rect -1007 -240 -950 -236
rect -1007 -300 -1003 -240
rect -1003 -300 -954 -240
rect -954 -300 -950 -240
rect -1007 -304 -950 -300
rect -1007 -524 -950 -520
rect -1007 -584 -1003 -524
rect -1003 -584 -954 -524
rect -954 -584 -950 -524
rect -1007 -588 -950 -584
rect -763 -241 -692 -237
rect -763 -296 -759 -241
rect -759 -296 -699 -241
rect -699 -296 -692 -241
rect -763 -300 -692 -296
rect 322 -240 392 -237
rect 322 -295 326 -240
rect 326 -295 386 -240
rect 386 -295 392 -240
rect 322 -299 392 -295
rect 2022 -187 2082 -134
rect 563 -371 622 -357
rect 563 -405 576 -371
rect 576 -405 610 -371
rect 610 -405 622 -371
rect 563 -417 622 -405
rect 2137 -356 2194 -352
rect 2137 -416 2141 -356
rect 2141 -416 2190 -356
rect 2190 -416 2194 -356
rect 2137 -420 2194 -416
rect 204 -525 272 -520
rect 204 -580 208 -525
rect 208 -580 268 -525
rect 268 -580 272 -525
rect 204 -585 272 -580
rect -1007 -824 -953 -762
rect -1007 -959 -953 -897
rect -1005 -1071 -951 -1009
rect -1005 -1196 -951 -1134
rect -1000 -1437 -946 -1375
rect 398 -1558 402 -1512
rect 402 -1558 460 -1512
rect 460 -1558 464 -1512
rect 398 -1564 464 -1558
rect -1003 -1659 -949 -1597
rect 2137 -524 2194 -520
rect 2137 -584 2141 -524
rect 2141 -584 2190 -524
rect 2190 -584 2194 -524
rect 2137 -588 2194 -584
rect 2381 -241 2452 -237
rect 2381 -296 2385 -241
rect 2385 -296 2445 -241
rect 2445 -296 2452 -241
rect 2381 -300 2452 -296
rect 3466 -240 3536 -237
rect 3466 -295 3470 -240
rect 3470 -295 3530 -240
rect 3530 -295 3536 -240
rect 3466 -299 3536 -295
rect 3707 -371 3766 -357
rect 3707 -405 3720 -371
rect 3720 -405 3754 -371
rect 3754 -405 3766 -371
rect 3707 -417 3766 -405
rect 3348 -525 3416 -520
rect 3348 -580 3352 -525
rect 3352 -580 3412 -525
rect 3412 -580 3416 -525
rect 3348 -585 3416 -580
rect 2032 -818 2102 -758
rect 5269 -520 5326 -516
rect 5269 -580 5273 -520
rect 5273 -580 5322 -520
rect 5322 -580 5326 -520
rect 5269 -584 5326 -580
rect 5513 -237 5584 -233
rect 5513 -292 5517 -237
rect 5517 -292 5577 -237
rect 5577 -292 5584 -237
rect 5513 -296 5584 -292
rect 6598 -236 6668 -233
rect 6598 -291 6602 -236
rect 6602 -291 6662 -236
rect 6662 -291 6668 -236
rect 6598 -295 6668 -291
rect 6839 -367 6898 -353
rect 6839 -401 6852 -367
rect 6852 -401 6886 -367
rect 6886 -401 6898 -367
rect 6839 -413 6898 -401
rect 8413 -352 8470 -348
rect 8413 -412 8417 -352
rect 8417 -412 8466 -352
rect 8466 -412 8470 -352
rect 8413 -416 8470 -412
rect 6480 -521 6548 -516
rect 6480 -576 6484 -521
rect 6484 -576 6544 -521
rect 6544 -576 6548 -521
rect 6480 -581 6548 -576
rect 5182 -956 5246 -899
rect 4914 -1434 4973 -1368
rect 8413 -520 8470 -516
rect 8413 -580 8417 -520
rect 8417 -580 8466 -520
rect 8466 -580 8470 -520
rect 8413 -584 8470 -580
rect 8657 -237 8728 -233
rect 8657 -292 8661 -237
rect 8661 -292 8721 -237
rect 8721 -292 8728 -237
rect 8657 -296 8728 -292
rect 9742 -236 9812 -233
rect 9742 -291 9746 -236
rect 9746 -291 9806 -236
rect 9806 -291 9812 -236
rect 9742 -295 9812 -291
rect 9983 -367 10042 -353
rect 9983 -401 9996 -367
rect 9996 -401 10030 -367
rect 10030 -401 10042 -367
rect 9983 -413 10042 -401
rect 9624 -521 9692 -516
rect 9624 -576 9628 -521
rect 9628 -576 9688 -521
rect 9688 -576 9692 -521
rect 9624 -581 9692 -576
rect 8324 -1062 8378 -1004
rect 8040 -1308 8099 -1251
rect 11215 -1171 11277 -1103
rect 11615 -524 11672 -520
rect 11615 -584 11619 -524
rect 11619 -584 11668 -524
rect 11668 -584 11672 -524
rect 11615 -588 11672 -584
rect 11859 -241 11930 -237
rect 11859 -296 11863 -241
rect 11863 -296 11923 -241
rect 11923 -296 11930 -241
rect 11859 -300 11930 -296
rect 12944 -240 13014 -237
rect 12944 -295 12948 -240
rect 12948 -295 13008 -240
rect 13008 -295 13014 -240
rect 12944 -299 13014 -295
rect 13185 -371 13244 -357
rect 13185 -405 13198 -371
rect 13198 -405 13232 -371
rect 13232 -405 13244 -371
rect 13185 -417 13244 -405
rect 14759 -356 14816 -352
rect 14759 -416 14763 -356
rect 14763 -416 14812 -356
rect 14812 -416 14816 -356
rect 14759 -420 14816 -416
rect 12826 -525 12894 -520
rect 12826 -580 12830 -525
rect 12830 -580 12890 -525
rect 12890 -580 12894 -525
rect 12826 -585 12894 -580
rect 11494 -1289 11563 -1228
rect 14759 -524 14816 -520
rect 14759 -584 14763 -524
rect 14763 -584 14812 -524
rect 14812 -584 14816 -524
rect 14759 -588 14816 -584
rect 14440 -1021 14496 -952
rect 15003 -241 15074 -237
rect 15003 -296 15007 -241
rect 15007 -296 15067 -241
rect 15067 -296 15074 -241
rect 15003 -300 15074 -296
rect 16088 -240 16158 -237
rect 16088 -295 16092 -240
rect 16092 -295 16152 -240
rect 16152 -295 16158 -240
rect 16088 -299 16158 -295
rect 16329 -371 16388 -357
rect 16329 -405 16342 -371
rect 16342 -405 16376 -371
rect 16376 -405 16388 -371
rect 16329 -417 16388 -405
rect 17891 -352 17948 -348
rect 17891 -412 17895 -352
rect 17895 -412 17944 -352
rect 17944 -412 17948 -352
rect 17891 -416 17948 -412
rect 15970 -525 16038 -520
rect 15970 -580 15974 -525
rect 15974 -580 16034 -525
rect 16034 -580 16038 -525
rect 15970 -585 16038 -580
rect 17891 -520 17948 -516
rect 17891 -580 17895 -520
rect 17895 -580 17944 -520
rect 17944 -580 17948 -520
rect 17891 -584 17948 -580
rect 17576 -858 17640 -799
rect 14645 -1430 14702 -1363
rect 3542 -1558 3546 -1512
rect 3546 -1558 3604 -1512
rect 3604 -1558 3608 -1512
rect 3542 -1564 3608 -1558
rect 6674 -1554 6678 -1508
rect 6678 -1554 6736 -1508
rect 6736 -1554 6740 -1508
rect 6674 -1560 6740 -1554
rect 9818 -1554 9822 -1508
rect 9822 -1554 9880 -1508
rect 9880 -1554 9884 -1508
rect 9818 -1560 9884 -1554
rect 13020 -1558 13024 -1512
rect 13024 -1558 13082 -1512
rect 13082 -1558 13086 -1512
rect 13020 -1564 13086 -1558
rect 16164 -1558 16168 -1512
rect 16168 -1558 16226 -1512
rect 16226 -1558 16230 -1512
rect 16164 -1564 16230 -1558
rect 18135 -237 18206 -233
rect 18135 -292 18139 -237
rect 18139 -292 18199 -237
rect 18199 -292 18206 -237
rect 18135 -296 18206 -292
rect 19220 -236 19290 -233
rect 19220 -291 19224 -236
rect 19224 -291 19284 -236
rect 19284 -291 19290 -236
rect 19220 -295 19290 -291
rect 19461 -367 19520 -353
rect 19461 -401 19474 -367
rect 19474 -401 19508 -367
rect 19508 -401 19520 -367
rect 19461 -413 19520 -401
rect 21035 -352 21092 -348
rect 21035 -412 21039 -352
rect 21039 -412 21088 -352
rect 21088 -412 21092 -352
rect 21035 -416 21092 -412
rect 19102 -521 19170 -516
rect 19102 -576 19106 -521
rect 19106 -576 19166 -521
rect 19166 -576 19170 -521
rect 19102 -581 19170 -576
rect 20721 -729 20774 -672
rect 21279 -237 21350 -233
rect 21279 -292 21283 -237
rect 21283 -292 21343 -237
rect 21343 -292 21350 -237
rect 21279 -296 21350 -292
rect 22364 -236 22434 -233
rect 22364 -291 22368 -236
rect 22368 -291 22428 -236
rect 22428 -291 22434 -236
rect 22364 -295 22434 -291
rect 22605 -367 22664 -353
rect 22605 -401 22618 -367
rect 22618 -401 22652 -367
rect 22652 -401 22664 -367
rect 22605 -413 22664 -401
rect 22246 -521 22314 -516
rect 22246 -576 22250 -521
rect 22250 -576 22310 -521
rect 22310 -576 22314 -521
rect 22246 -581 22314 -576
rect 24219 -735 24290 -664
rect 24207 -860 24273 -800
rect 24197 -1027 24261 -958
rect 24197 -1173 24261 -1104
rect 24197 -1313 24261 -1244
rect 24196 -1452 24260 -1383
rect 19296 -1554 19300 -1508
rect 19300 -1554 19358 -1508
rect 19358 -1554 19362 -1508
rect 19296 -1560 19362 -1554
rect 22440 -1554 22444 -1508
rect 22444 -1554 22502 -1508
rect 22502 -1554 22506 -1508
rect 22440 -1560 22506 -1554
rect 1781 -1729 1854 -1648
rect 17774 -1655 17844 -1579
rect 24196 -1720 24260 -1651
<< metal2 >>
rect 372 734 472 744
rect 372 632 472 642
rect 3516 734 3616 744
rect 3516 632 3616 642
rect 6648 738 6748 748
rect 6648 636 6748 646
rect 9792 738 9892 748
rect 9792 636 9892 646
rect 12994 734 13094 744
rect 12994 632 13094 642
rect 16138 734 16238 744
rect 16138 632 16238 642
rect 19270 738 19370 748
rect 19270 636 19370 646
rect 22414 738 22514 748
rect 22414 636 22514 646
rect -1006 -85 -952 -77
rect -1017 -87 2082 -85
rect -1017 -149 -1006 -87
rect -952 -134 2082 -87
rect -952 -149 2022 -134
rect -1017 -150 -938 -149
rect -1006 -159 -952 -150
rect 2022 -197 2082 -187
rect 5502 -223 5595 -221
rect 8646 -223 8739 -221
rect 18124 -223 18217 -221
rect 21268 -223 21361 -221
rect -1007 -227 -950 -226
rect -774 -227 -681 -225
rect 2370 -227 2463 -225
rect 3413 -227 9821 -223
rect 11848 -227 11941 -225
rect 14992 -227 15085 -225
rect 16076 -227 22443 -223
rect -1015 -228 401 -227
rect 2196 -228 22443 -227
rect -1018 -233 22443 -228
rect -1018 -236 5513 -233
rect -1018 -304 -1007 -236
rect -950 -237 5513 -236
rect -950 -300 -763 -237
rect -692 -299 322 -237
rect 392 -299 2381 -237
rect -692 -300 2381 -299
rect 2452 -299 3466 -237
rect 3536 -296 5513 -237
rect 5584 -295 6598 -233
rect 6668 -295 8657 -233
rect 5584 -296 8657 -295
rect 8728 -295 9742 -233
rect 9812 -237 18135 -233
rect 9812 -295 11859 -237
rect 8728 -296 11859 -295
rect 3536 -299 11859 -296
rect 2452 -300 11859 -299
rect 11930 -299 12944 -237
rect 13014 -299 15003 -237
rect 11930 -300 15003 -299
rect 15074 -299 16088 -237
rect 16158 -296 18135 -237
rect 18206 -295 19220 -233
rect 19290 -295 21279 -233
rect 18206 -296 21279 -295
rect 21350 -295 22364 -233
rect 22434 -295 22443 -233
rect 21350 -296 22443 -295
rect 16158 -299 22443 -296
rect 15074 -300 22443 -299
rect -950 -304 22443 -300
rect -1018 -307 22443 -304
rect -1018 -308 5336 -307
rect -1018 -311 5226 -308
rect 11604 -311 17955 -307
rect -1018 -312 -940 -311
rect 358 -312 2204 -311
rect 12932 -312 14826 -311
rect -1007 -314 -950 -312
rect 8413 -340 8470 -338
rect 2137 -344 2194 -342
rect 8402 -343 8498 -340
rect 2126 -347 2222 -344
rect -1018 -357 622 -347
rect -1018 -361 563 -357
rect -1018 -417 -1008 -361
rect -952 -417 563 -361
rect -1018 -426 622 -417
rect -1008 -427 -952 -426
rect 563 -427 622 -426
rect 2126 -352 3766 -347
rect 2126 -420 2137 -352
rect 2194 -357 3766 -352
rect 2194 -417 3707 -357
rect 2194 -420 3766 -417
rect 2126 -426 3766 -420
rect 2126 -429 2222 -426
rect 3707 -427 3766 -426
rect 5080 -353 6898 -343
rect 5080 -413 6839 -353
rect 5080 -422 6898 -413
rect 2137 -430 2194 -429
rect 5080 -466 5137 -422
rect 6839 -423 6898 -422
rect 8402 -348 10042 -343
rect 8402 -416 8413 -348
rect 8470 -353 10042 -348
rect 8470 -413 9983 -353
rect 8470 -416 10042 -413
rect 8402 -422 10042 -416
rect 8402 -425 8498 -422
rect 9983 -423 10042 -422
rect 11337 -357 13244 -347
rect 11337 -417 13185 -357
rect 8413 -426 8470 -425
rect 11337 -426 13244 -417
rect 14748 -352 16388 -347
rect 14748 -420 14759 -352
rect 14816 -357 16388 -352
rect 14816 -417 16329 -357
rect 14816 -420 16388 -417
rect 14748 -426 16388 -420
rect -1007 -511 -950 -510
rect 2137 -511 2194 -510
rect 4922 -511 5137 -466
rect 5269 -507 5326 -506
rect 8413 -507 8470 -506
rect 5258 -508 5354 -507
rect 8402 -508 8498 -507
rect -1018 -512 -922 -511
rect 2126 -512 2222 -511
rect -1018 -520 1815 -512
rect -1018 -588 -1007 -520
rect -950 -585 204 -520
rect 272 -585 1815 -520
rect -950 -588 1815 -585
rect -1018 -596 1815 -588
rect 2126 -520 3427 -512
rect 2126 -588 2137 -520
rect 2194 -585 3348 -520
rect 3416 -585 3427 -520
rect 2194 -588 3427 -585
rect 2126 -596 3427 -588
rect -1007 -598 -950 -596
rect 1740 -637 1815 -596
rect 2137 -598 2194 -596
rect 4922 -637 4994 -511
rect 5258 -516 8036 -508
rect 5258 -584 5269 -516
rect 5326 -581 6480 -516
rect 6548 -581 8036 -516
rect 5326 -584 8036 -581
rect 5258 -592 8036 -584
rect 8402 -516 9703 -508
rect 8402 -584 8413 -516
rect 8470 -581 9624 -516
rect 9692 -581 9703 -516
rect 8470 -584 9703 -581
rect 8402 -592 9703 -584
rect 5269 -594 5326 -592
rect 1740 -702 4994 -637
rect 7957 -675 8036 -592
rect 8413 -594 8470 -592
rect 11337 -675 11427 -426
rect 13185 -427 13244 -426
rect 16329 -427 16388 -426
rect 17658 -348 19520 -343
rect 17658 -416 17891 -348
rect 17948 -353 19520 -348
rect 17948 -413 19461 -353
rect 17948 -416 19520 -413
rect 17658 -422 19520 -416
rect 21024 -348 22664 -343
rect 21024 -416 21035 -348
rect 21092 -353 22664 -348
rect 21092 -413 22605 -353
rect 21092 -416 22664 -413
rect 21024 -422 22664 -416
rect 11615 -511 11672 -510
rect 14759 -511 14816 -510
rect 11604 -512 11700 -511
rect 14748 -512 14844 -511
rect 11604 -520 12906 -512
rect 11604 -588 11615 -520
rect 11672 -585 12826 -520
rect 12894 -585 12906 -520
rect 11672 -588 12906 -585
rect 11604 -596 12906 -588
rect 14748 -520 16049 -512
rect 14748 -588 14759 -520
rect 14816 -585 15970 -520
rect 16038 -585 16049 -520
rect 14816 -588 16049 -585
rect 14748 -596 16049 -588
rect 11615 -598 11672 -596
rect 7957 -743 11427 -675
rect 12825 -653 12906 -596
rect 14759 -598 14816 -596
rect 17658 -653 17739 -422
rect 19461 -423 19520 -422
rect 22605 -423 22664 -422
rect 21024 -506 21103 -496
rect 17891 -507 17948 -506
rect 17880 -508 17976 -507
rect 17880 -516 19181 -508
rect 17880 -584 17891 -516
rect 17948 -581 19102 -516
rect 19170 -581 19181 -516
rect 17948 -584 19181 -581
rect 17880 -592 19181 -584
rect 17891 -594 17948 -592
rect 21103 -508 21120 -507
rect 21103 -516 22325 -508
rect 21103 -581 22246 -516
rect 22314 -581 22325 -516
rect 21103 -592 22325 -581
rect 21024 -605 21103 -595
rect 12825 -732 17739 -653
rect 20721 -654 24255 -653
rect 20721 -664 24290 -654
rect 20721 -672 24219 -664
rect 20774 -729 24219 -672
rect 20721 -735 24219 -729
rect 20721 -743 24290 -735
rect 24219 -745 24290 -743
rect -1007 -761 -953 -752
rect 2032 -758 2102 -748
rect -1018 -762 2032 -761
rect -1018 -824 -1007 -762
rect -953 -818 2032 -762
rect 2102 -818 2109 -761
rect -953 -824 2109 -818
rect -1018 -825 2109 -824
rect 17576 -799 17640 -789
rect -1007 -834 -953 -825
rect 2032 -828 2102 -825
rect 17576 -868 17640 -858
rect 24207 -800 24273 -790
rect 24207 -870 24273 -860
rect -1007 -896 -953 -887
rect 5182 -896 5246 -889
rect -1018 -897 5246 -896
rect -1018 -959 -1007 -897
rect -953 -899 5246 -897
rect -953 -956 5182 -899
rect -953 -959 5246 -956
rect -1018 -960 5246 -959
rect -1007 -969 -953 -960
rect 5182 -966 5246 -960
rect 14440 -952 14496 -942
rect -1005 -1008 -951 -999
rect 8324 -1004 8378 -994
rect -1016 -1009 8324 -1008
rect -1016 -1071 -1005 -1009
rect -951 -1062 8324 -1009
rect 14440 -1031 14496 -1021
rect 24197 -958 24261 -948
rect 24197 -1037 24261 -1027
rect -951 -1071 8378 -1062
rect -1016 -1072 8378 -1071
rect -1005 -1081 -951 -1072
rect 11215 -1103 11277 -1093
rect -1005 -1133 -951 -1124
rect -1016 -1134 -789 -1133
rect -1016 -1196 -1005 -1134
rect -951 -1196 11091 -1134
rect 11215 -1181 11277 -1171
rect 24197 -1104 24261 -1094
rect 24197 -1183 24261 -1173
rect -1016 -1197 11091 -1196
rect -1005 -1206 -951 -1197
rect 11023 -1232 11091 -1197
rect 11494 -1228 11563 -1218
rect 8040 -1251 8099 -1241
rect 4688 -1327 5135 -1263
rect 11023 -1289 11494 -1232
rect 11023 -1296 11563 -1289
rect 11494 -1299 11563 -1296
rect 24197 -1244 24261 -1234
rect 8040 -1318 8099 -1308
rect 24197 -1323 24261 -1313
rect -1000 -1367 -946 -1365
rect 4688 -1367 4752 -1327
rect -1017 -1375 4752 -1367
rect -1017 -1432 -1000 -1375
rect -1011 -1437 -1000 -1432
rect -946 -1432 4752 -1375
rect 4914 -1368 4973 -1358
rect -946 -1437 -935 -1432
rect -1011 -1438 -935 -1437
rect 5071 -1368 5135 -1327
rect 14645 -1363 14702 -1353
rect 5071 -1430 14645 -1368
rect 5071 -1432 14702 -1430
rect -1000 -1447 -946 -1438
rect 4914 -1444 4973 -1434
rect 14645 -1440 14702 -1432
rect 24196 -1383 24260 -1373
rect 24196 -1462 24260 -1452
rect 392 -1510 468 -1500
rect 392 -1578 468 -1568
rect 3536 -1510 3612 -1500
rect 3536 -1578 3612 -1568
rect 6668 -1506 6744 -1496
rect 6668 -1574 6744 -1564
rect 9812 -1506 9888 -1496
rect 9812 -1574 9888 -1564
rect 13014 -1510 13090 -1500
rect 13014 -1578 13090 -1568
rect 16158 -1510 16234 -1500
rect 16158 -1578 16234 -1568
rect 19290 -1506 19366 -1496
rect 17774 -1579 17844 -1569
rect 19290 -1574 19366 -1564
rect 22434 -1506 22510 -1496
rect 22434 -1574 22510 -1564
rect -1003 -1596 -949 -1589
rect -1014 -1597 -896 -1596
rect -1014 -1659 -1003 -1597
rect -949 -1607 -896 -1597
rect -949 -1659 1642 -1607
rect -1014 -1660 1642 -1659
rect -1003 -1669 -949 -1660
rect 1578 -1768 1642 -1660
rect 1781 -1648 1854 -1638
rect 1913 -1655 17774 -1606
rect 1913 -1660 17844 -1655
rect 1913 -1665 1976 -1660
rect 17774 -1665 17844 -1660
rect 24196 -1651 24260 -1641
rect 1781 -1739 1854 -1729
rect 1912 -1768 1976 -1665
rect 24196 -1730 24260 -1720
rect 1578 -1796 1976 -1768
<< via2 >>
rect 372 706 472 734
rect 372 646 384 706
rect 384 646 464 706
rect 464 646 472 706
rect 372 642 472 646
rect 3516 706 3616 734
rect 3516 646 3528 706
rect 3528 646 3608 706
rect 3608 646 3616 706
rect 3516 642 3616 646
rect 6648 710 6748 738
rect 6648 650 6660 710
rect 6660 650 6740 710
rect 6740 650 6748 710
rect 6648 646 6748 650
rect 9792 710 9892 738
rect 9792 650 9804 710
rect 9804 650 9884 710
rect 9884 650 9892 710
rect 9792 646 9892 650
rect 12994 706 13094 734
rect 12994 646 13006 706
rect 13006 646 13086 706
rect 13086 646 13094 706
rect 12994 642 13094 646
rect 16138 706 16238 734
rect 16138 646 16150 706
rect 16150 646 16230 706
rect 16230 646 16238 706
rect 16138 642 16238 646
rect 19270 710 19370 738
rect 19270 650 19282 710
rect 19282 650 19362 710
rect 19362 650 19370 710
rect 19270 646 19370 650
rect 22414 710 22514 738
rect 22414 650 22426 710
rect 22426 650 22506 710
rect 22506 650 22514 710
rect 22414 646 22514 650
rect -1008 -417 -952 -361
rect 21024 -595 21103 -506
rect 17576 -858 17640 -799
rect 24207 -860 24273 -800
rect 14440 -1021 14496 -952
rect 24197 -1027 24261 -958
rect 11215 -1171 11277 -1103
rect 24197 -1173 24261 -1104
rect 8040 -1308 8099 -1251
rect 24197 -1313 24261 -1244
rect 4914 -1434 4973 -1368
rect 24196 -1452 24260 -1383
rect 392 -1512 468 -1510
rect 392 -1564 398 -1512
rect 398 -1564 464 -1512
rect 464 -1564 468 -1512
rect 392 -1568 468 -1564
rect 3536 -1512 3612 -1510
rect 3536 -1564 3542 -1512
rect 3542 -1564 3608 -1512
rect 3608 -1564 3612 -1512
rect 3536 -1568 3612 -1564
rect 6668 -1508 6744 -1506
rect 6668 -1560 6674 -1508
rect 6674 -1560 6740 -1508
rect 6740 -1560 6744 -1508
rect 6668 -1564 6744 -1560
rect 9812 -1508 9888 -1506
rect 9812 -1560 9818 -1508
rect 9818 -1560 9884 -1508
rect 9884 -1560 9888 -1508
rect 9812 -1564 9888 -1560
rect 13014 -1512 13090 -1510
rect 13014 -1564 13020 -1512
rect 13020 -1564 13086 -1512
rect 13086 -1564 13090 -1512
rect 13014 -1568 13090 -1564
rect 16158 -1512 16234 -1510
rect 16158 -1564 16164 -1512
rect 16164 -1564 16230 -1512
rect 16230 -1564 16234 -1512
rect 16158 -1568 16234 -1564
rect 19290 -1508 19366 -1506
rect 19290 -1560 19296 -1508
rect 19296 -1560 19362 -1508
rect 19362 -1560 19366 -1508
rect 19290 -1564 19366 -1560
rect 22434 -1508 22510 -1506
rect 22434 -1560 22440 -1508
rect 22440 -1560 22506 -1508
rect 22506 -1560 22510 -1508
rect 22434 -1564 22510 -1560
rect 1781 -1729 1854 -1648
rect 24196 -1720 24260 -1651
<< metal3 >>
rect 362 734 482 739
rect 362 640 372 734
rect 472 640 482 734
rect 362 637 482 640
rect 3506 734 3626 739
rect 3506 640 3516 734
rect 3616 640 3626 734
rect 6638 738 6758 743
rect 6638 644 6648 738
rect 6748 644 6758 738
rect 6638 641 6758 644
rect 9782 738 9902 743
rect 9782 644 9792 738
rect 9892 644 9902 738
rect 9782 641 9902 644
rect 12984 734 13104 739
rect 3506 637 3626 640
rect 12984 640 12994 734
rect 13094 640 13104 734
rect 12984 637 13104 640
rect 16128 734 16248 739
rect 16128 640 16138 734
rect 16238 640 16248 734
rect 19260 738 19380 743
rect 19260 644 19270 738
rect 19370 644 19380 738
rect 19260 641 19380 644
rect 22404 738 22524 743
rect 22404 644 22414 738
rect 22514 644 22524 738
rect 22404 641 22524 644
rect 16128 637 16248 640
rect -1028 -347 -931 -346
rect -1028 -430 -1018 -347
rect -941 -430 -931 -347
rect -1028 -449 -931 -430
rect 21003 -605 21013 -496
rect 21113 -605 21123 -496
rect 17566 -795 24279 -794
rect 17566 -799 24283 -795
rect 17566 -858 17576 -799
rect 17640 -800 24283 -799
rect 17640 -858 24207 -800
rect 17566 -860 24207 -858
rect 24273 -860 24283 -800
rect 17566 -863 24283 -860
rect 24197 -865 24283 -863
rect 14430 -952 14506 -947
rect 14430 -1021 14440 -952
rect 14496 -958 14506 -952
rect 24187 -958 24271 -953
rect 14496 -1021 24197 -958
rect 14430 -1026 24197 -1021
rect 24187 -1027 24197 -1026
rect 24261 -1027 24271 -958
rect 24187 -1032 24271 -1027
rect 11205 -1103 11287 -1098
rect 11205 -1171 11215 -1103
rect 11277 -1104 11287 -1103
rect 24187 -1104 24271 -1099
rect 11277 -1171 24197 -1104
rect 11205 -1172 24197 -1171
rect 11205 -1176 11287 -1172
rect 24187 -1173 24197 -1172
rect 24261 -1173 24271 -1104
rect 24187 -1178 24271 -1173
rect 24187 -1244 24271 -1239
rect 8085 -1246 24197 -1244
rect 8030 -1251 24197 -1246
rect 8030 -1308 8040 -1251
rect 8099 -1308 24197 -1251
rect 8030 -1312 24197 -1308
rect 8030 -1313 8109 -1312
rect 24187 -1313 24197 -1312
rect 24261 -1313 24271 -1244
rect 24187 -1318 24271 -1313
rect 4904 -1368 4983 -1363
rect 4904 -1434 4914 -1368
rect 4973 -1377 4983 -1368
rect 22650 -1377 24059 -1372
rect 4973 -1382 24059 -1377
rect 24126 -1382 24270 -1378
rect 4973 -1383 24270 -1382
rect 4973 -1434 24196 -1383
rect 4904 -1438 24196 -1434
rect 4904 -1439 4983 -1438
rect 22650 -1446 24196 -1438
rect 24094 -1451 24196 -1446
rect 24186 -1452 24196 -1451
rect 24260 -1452 24270 -1383
rect 24186 -1457 24270 -1452
rect 352 -1510 518 -1502
rect 352 -1578 386 -1510
rect 470 -1578 518 -1510
rect 352 -1582 518 -1578
rect 3496 -1510 3662 -1502
rect 3496 -1578 3530 -1510
rect 3614 -1578 3662 -1510
rect 6628 -1506 6794 -1498
rect 6628 -1574 6662 -1506
rect 6746 -1574 6794 -1506
rect 6628 -1578 6794 -1574
rect 9772 -1506 9938 -1498
rect 9772 -1574 9806 -1506
rect 9890 -1574 9938 -1506
rect 9772 -1578 9938 -1574
rect 12974 -1510 13140 -1502
rect 12974 -1578 13008 -1510
rect 13092 -1578 13140 -1510
rect 3496 -1582 3662 -1578
rect 12974 -1582 13140 -1578
rect 16118 -1510 16284 -1502
rect 16118 -1578 16152 -1510
rect 16236 -1578 16284 -1510
rect 19250 -1506 19416 -1498
rect 19250 -1574 19284 -1506
rect 19368 -1574 19416 -1506
rect 19250 -1578 19416 -1574
rect 22394 -1506 22560 -1498
rect 22394 -1574 22428 -1506
rect 22512 -1574 22560 -1506
rect 22394 -1578 22560 -1574
rect 16118 -1582 16284 -1578
rect 1771 -1648 1864 -1643
rect 24103 -1648 24270 -1646
rect 1771 -1729 1781 -1648
rect 1854 -1651 24270 -1648
rect 1854 -1720 24196 -1651
rect 24260 -1720 24270 -1651
rect 1854 -1725 24270 -1720
rect 1854 -1728 24210 -1725
rect 1854 -1729 1864 -1728
rect 1771 -1734 1864 -1729
<< via3 >>
rect 372 642 472 732
rect 372 640 472 642
rect 3516 642 3616 732
rect 3516 640 3616 642
rect 6648 646 6748 736
rect 6648 644 6748 646
rect 9792 646 9892 736
rect 9792 644 9892 646
rect 12994 642 13094 732
rect 12994 640 13094 642
rect 16138 642 16238 732
rect 16138 640 16238 642
rect 19270 646 19370 736
rect 19270 644 19370 646
rect 22414 646 22514 736
rect 22414 644 22514 646
rect -1018 -361 -941 -347
rect -1018 -417 -1008 -361
rect -1008 -417 -952 -361
rect -952 -417 -941 -361
rect -1018 -430 -941 -417
rect 21013 -506 21113 -496
rect 21013 -595 21024 -506
rect 21024 -595 21103 -506
rect 21103 -595 21113 -506
rect 21013 -605 21113 -595
rect 386 -1568 392 -1510
rect 392 -1568 468 -1510
rect 468 -1568 470 -1510
rect 386 -1578 470 -1568
rect 3530 -1568 3536 -1510
rect 3536 -1568 3612 -1510
rect 3612 -1568 3614 -1510
rect 3530 -1578 3614 -1568
rect 6662 -1564 6668 -1506
rect 6668 -1564 6744 -1506
rect 6744 -1564 6746 -1506
rect 6662 -1574 6746 -1564
rect 9806 -1564 9812 -1506
rect 9812 -1564 9888 -1506
rect 9888 -1564 9890 -1506
rect 9806 -1574 9890 -1564
rect 13008 -1568 13014 -1510
rect 13014 -1568 13090 -1510
rect 13090 -1568 13092 -1510
rect 13008 -1578 13092 -1568
rect 16152 -1568 16158 -1510
rect 16158 -1568 16234 -1510
rect 16234 -1568 16236 -1510
rect 16152 -1578 16236 -1568
rect 19284 -1564 19290 -1506
rect 19290 -1564 19366 -1506
rect 19366 -1564 19368 -1506
rect 19284 -1574 19368 -1564
rect 22428 -1564 22434 -1506
rect 22434 -1564 22510 -1506
rect 22510 -1564 22512 -1506
rect 22428 -1574 22512 -1564
<< metal4 >>
rect -484 736 23446 842
rect -484 732 6648 736
rect -484 640 372 732
rect 472 640 3516 732
rect 3616 644 6648 732
rect 6748 644 9792 736
rect 9892 732 19270 736
rect 9892 644 12994 732
rect 3616 640 12994 644
rect 13094 640 16138 732
rect 16238 644 19270 732
rect 19370 644 22414 736
rect 22514 644 23446 736
rect 16238 640 23446 644
rect -484 608 23446 640
rect -1028 -347 -940 -346
rect -1028 -430 -1018 -347
rect -941 -430 -940 -347
rect -1028 -1499 -940 -430
rect 21003 -496 21124 -495
rect 21003 -605 21013 -496
rect 21113 -605 21124 -496
rect 21003 -1498 21124 -605
rect -504 -1499 22870 -1498
rect -1028 -1506 22870 -1499
rect -1028 -1510 6662 -1506
rect -1028 -1578 386 -1510
rect 470 -1578 3530 -1510
rect 3614 -1574 6662 -1510
rect 6746 -1574 9806 -1506
rect 9890 -1510 19284 -1506
rect 9890 -1574 13008 -1510
rect 3614 -1578 13008 -1574
rect 13092 -1578 16152 -1510
rect 16236 -1574 19284 -1510
rect 19368 -1574 22428 -1506
rect 22512 -1574 22870 -1506
rect 16236 -1578 22870 -1574
rect -1028 -1678 22870 -1578
<< labels >>
flabel metal4 11190 624 11552 788 1 FreeSerif 960 0 0 0 VDD
port 1 n
flabel metal4 11162 -1670 11548 -1542 1 FreeSerif 960 0 0 0 VSS
port 2 n
flabel metal1 24275 -373 24351 -293 1 FreeSerif 720 0 0 0 Y[7]
port 20 n
flabel metal1 24303 -734 24345 -666 1 FreeSerif 720 0 0 0 Y[6]
port 21 n
flabel metal1 24301 -863 24346 -803 1 FreeSerif 720 0 0 0 Y[5]
port 22 n
flabel metal1 24294 -1028 24347 -959 1 FreeSerif 720 0 0 0 Y[4]
port 23 n
flabel metal1 24287 -1181 24348 -1105 1 FreeSerif 720 0 0 0 Y[3]
port 15 n
flabel metal1 24279 -1323 24354 -1240 1 FreeSerif 720 0 0 0 Y[2]
port 24 n
flabel metal1 24276 -1455 24349 -1378 1 FreeSerif 720 0 0 0 Y[1]
port 17 n
flabel metal1 24287 -1724 24343 -1657 1 FreeSerif 720 0 0 0 Y[0]
port 25 n
flabel metal1 -1266 -309 -1200 -233 1 FreeSerif 720 0 0 0 dir
port 26 n
flabel metal1 -1263 -591 -1194 -521 1 FreeSerif 720 0 0 0 A[1]
port 27 n
flabel metal1 -1261 -819 -1197 -769 1 FreeSerif 720 0 0 0 A[2]
port 5 n
flabel metal1 -1262 -955 -1200 -903 1 FreeSerif 720 0 0 0 A[3]
port 6 n
flabel metal1 -1262 -1065 -1212 -1015 1 FreeSerif 720 0 0 0 A[4]
port 7 n
flabel metal1 -1255 -1431 -1209 -1383 1 FreeSerif 720 0 0 0 A[6]
port 9 n
flabel metal1 -1265 -1194 -1209 -1138 1 FreeSerif 720 0 0 0 A[5]
port 8 n
flabel metal1 -1253 -1647 -1180 -1612 1 FreeSerif 720 0 0 0 A[7]
port 28 n
flabel metal1 -1266 -148 -1184 -94 1 FreeSerif 720 0 0 0 A[0]
port 29 n
<< end >>
